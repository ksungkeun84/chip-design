%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
Gb6Zn6BAiHXe7F6Sao/7wmvi5u5s2OeXw5452IbS4P7oLtZOwTidAjb8I0gWwlm1oHFwFfyMUDJi
pMXFPpF7AOBNWBFZuy6teKLKDQyl9pBiECl+eVc1TYuK6ks68I2Cz/HXyPC2jyZTtQyBEgxdTo0e
k/iWSscDGyciQCxC9Af7M9MAVPo7I0NnrWvNB+vdCfUg72HLzNN10SxNi+DWyOCOeaKc2y5Pak2i
tJ03gDlssQSf+f0HBNQok2QIOrk8H9m4AvTmLOeAvfJbY5rSljyiEmhS4aLF4ftJOrO9BLW9eL1H
Db+NxR6uVPle5xaE2nijjHNd2Z2pp+BY9taP7Q==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
5+MWLw7LOV0T8SGzeDCMOqPaW3K6o22vszfAkRpxjP5/giw7mGpXReg8JVCmNMzDiVMaRQOmgTEp
a4gwEDdCPipdAjbjSyX4cmv1jy2zSONJTuHYqR4UC6k9QgOSeG07iBCdq4Z2UBfFLD6dwK15XG8q
P45jWOUhZ5HNnYNG4iQ89ygIYClFNzT4kWL8rDbY0MAxQXMUpwzxchnrQmI2Ikl+T1vvzKrzbxS3
FATTkl491KUppxEU1ehLUbRLq8I/Jyr3c+S1m9kI1Pbsh8KDGA1VnNGMbKUzR/rhczTgk86sqxc4
inY6Blz2D2YU2nHLcVEoET5AK4n2B7b0GRs294eyfvDqSMHqUO+uib/NORTPyo/dmiTbKD2gGktH
g2N20az0PHcdobcHV5RKjvkc2xOA9HsM/c2Isc+nxm5t+oRvZGeftV8//Vg0F9qvOTyz+ubUxlOb
BKW00GCNbCyQsx1iApWcwywUBVwncF/fJPJRRGCcuLCUHqqsyks/ViOBJafERyzmNJLw4jP8Kvi0
W/58tStwFReMfVxKwG1647gX8hu5iCpvDOHxzq0cw81YjGFqfv2ahWogls5fLtJ7LYt9uBj5e4qj
GZ9fH1vm4Hb+6jacOxfTtqe4o4y6v5T0iE1jRxpBRdugywTFXD8Wm7kPTYnMQJcNYP8uwQv8i21g
fmjOLpuziWbeunBAdn6deTLHustgxFdMaBrN3PBs+9KDkFqLp3LVFpx/TBrL16NTq3Ye2JecokB1
a/pwXqOW558N7hHgArME3wrzBlcnSXysBW2DeSew80JObafRSceZ2eP0qjqn2qZqcKLlVKQTIiKv
SnOT6/XVuc5u4DxmrT1LTyE8ZuK9uPH3Lnx+LI7E0HU4ciF0qifwqd0Z/mFRZAP0OWD8A/8YCx+g
e8XMoE8MlbePXylilaqlMqk66q9MSe9Zzy3JEjm4gsoDlUu8zBLHMl7IFoWUVoM+qhdwBhLkzevD
SumlBgX1hFQ6KZIaf/49AgRNFD+Zb+5/dLPOrA3v6aAu3LDJqn8gx9kGVK8vVl66EcYu5T2tE1gj
ll5rXD0f/16B52ctDsa2MjIUskpKVy8FyAvenDdGUAHUB3YmjZ+HUU6KGtLEAnWfcLiavl/i7kMc
LmokbNMjmQ0KjQ7aHVeLLo/IFRExdynw4IPbW7CkMohcCvDxTw5GddyJosmB2nBByCyQhsHIR0Kf
xkRPv/VywHLQLsPIf6b9xNp2yMitXC2JODhqYU7ipbaWD6jYVuGVZskUeozy5jKglEDmAFiZmdnl
TEBSXm1+dUReHjJQDHqTPNGg1BpWnVasOQZLDE/LIXlYfbSsOFWpkAkmguiWO7vMFK1gWogORhAU
PKLd1e2Hi1A2Tt4+Jb5pcioj7wXgTvyDNhsS7LNPFhZBInUAD+sonjIuSTJapFRooZDHFjYBBCJh
7v1u3uvC/01UFFHkdMniFeCW6Lbf8aSXOpm6Pt6coHd+QQmRs6ISQaia/ZCmxKS/BUEfa9JpZSLI
HEE+dijHeJwLw11NxpHG5dA3/Iz8oSd6VQ3aHxVaG6i0UHedidkpcgHYA7a/JDqe2PQZMprC7C/7
A3De1RieNQyt05DR1zd/CmNH8D0lxxiDDv5OgNKrUsQ189Dg8fJUsMJb3s6/GEqdpL+Q/lnKVsQx
NMxxa5qKxlUVXDJyn857n5vM0oz9YeT+Bsfm40wwORkX5mThh0X3+7hrhNU3xA5Z8FChOps7sC58
O0+TO8ar5MKr5vwHNNrDQeJrK3JVaP3AtBFn03Ur76c/3Ukb1tvXHZIrGyu8wqSEVI6p16jBmR+0
m4Gu0FLGT8XqjIHPxh/PZ1mGKOEU4lTmiWXprfxgNGppoR+YnFYGjV8YFxadX9XT5v7jGfHV5lI+
xkDKfzED09alu5SnmaP7cpyA7yv3ZCsaAc61XJ7xLl/66jvxzRfkuSWIqfy3HgmpNIzvzeUVYAt0
ZWjt8K6fsxul5SPzjjvrUJLRICKCOMllf9Sbq/TKnGp7MNYfzfpnDnyGXZfQEfdWK4+mVA1x1YbC
V3PHauI7S1BElQHlLq5TsPke59XjD3IdXSRRW2IdtC5BzkCAi0miIyvRR6P34XDfLTUiMjJVWcqV
kCjLPiMNFPeLkQhOaEPsNIg4Q7XL1NNdfW8osS+9rh3AeDy8TG1XTy+PPDcIgy6cu0BKwldOg6qi
mKsBCJ7qaNzqJAOocMmuoZFwSRb3irAmH6I9Bv7oe55tRzQZ4Y3wS+sxuvU3n1DhyMV7pDL+a1zZ
/CHk6R4prUr5X2dQ+jOIcU5SGqnywJlVgfxTXJj+i6rJRjMMBXi55La430OQJfzTFFa1FVT17OvT
7ZiwKfa3HdHo6cKGs4VEmcxhgEAXNNtDYzU9sixhLSSMzDu162cH6AC5aTH2tt+VOEQQZkMROD0m
b9EeIdZISTWRmg1hJ7KTwWAqaTqrmUNFkrWynSJaVyqsIXLNybReJ0C9Z4dO2PNmgq2Gmkd8bfJF
Sy8I2mYoz66T8OwrUbhC7fYhJz1BM5Jo2tO4Ekk00phPcWw71XLHjs37710kyHDXEqes8rGvkAGT
LFGAi2UGCpbf6rGlB+CLEox6bPnUFLHdyYUBrTrxOVP7rbQjhSjnidP/91SK386yYRZNAeHp9xCO
0uECe5PPB78PNUj7/DY4h8+EdO/qr40BzQwNFT3LZoaPEW/1cb/LkC7RB4ZYa8453oUDmBceBn8N
pqdTpM5IXUE4mv1avAN98Mw/YE1R/C6kquvAnTlCFbItuEPdiKXZj3JDZolgLIW81aFa/paK3c9N
OgTkSShWz3buOgtjUQPoR2+Nq0OBREss8KymwH6ILkVJF86hmkbSIlXzQX+UxKqMWmw0bcGyvK3l
ytGeBlcPzM/SlswBuqMAVNzOBgi1jTkP9pvOAT8e3/fjc7kDHb60Yo0uXxtGvbsSOwq1Qo3xP8uG
Gz86lvX5RDrDnIsi28WFEm+xtnpa49ZaIkoz9cA+OPOuUpBqbfoq/dpPbntr1jxasrvx4RhkOlF3
RSAVI6RXjBAJgh/R7jgKq6m924I4IxcqdRrxdH0SvFZNmiJuTTaKqGm3gGH0JRVY6K5YPbkqDZD3
GgMZIFEeLRIQJZOmrk6Qj7DMy2CEDOZP4u2AdsZcvjKagQgAdMvxiErKeJ/e3ujWF8rJCHRaUxVV
+6AQ/+1JbY/fOqj1xkQvUmRwWMkc3/nWvGEPPTTfdf05iQlbagXbs5gWsQqXoiY/tm4Jg4ggUUqe
Sa99IY0dTNeZ3m+WuRKjk+kL8ldwKLX1Oys2NdWBvMNbvoxNnjq13U+RWskv7wQ5IBrBAtpMuhMK
Kiyb/CQfMb6rioIpv4QXRPI3TizNCSgEMqQQtd7IeEAHocp+CARUi3YiD35eyKloMZ4pdXelWcqx
ZuDJ3qSzkEYd2u2iw5fDjPn3s8cIu3JXSZGapIyiTcECGeH2UHfHM3twqMK2VN7D4pUIR9REgWgF
xmo4mtXgilIm+ADfspqol3PxCQ15rIjLUi79By7n5VrrJygZ/KdPtiZk1mRItab9FCQKn2pK86xw
Dztt5Fax3to6XBHpqhlGjyDq2hRGfAHowNIpueiqiFyjf07LcxXjc7378R+VTgVRT43RkmVa9l27
bkXf9HHMXaE/Ntvfx1EWx9kE/bJ2vI8YtoIlFCJkOz+z0Dt/TjXkmMzOdipl/7Vu6EePqoSFohvr
JekYl+ItiCVKxUDhNUzxe9HOxCChsukN2hM+BtTcly2b/C/bVZQR1q2p5mfA/tkt7NTBymn7BAHH
iOL+M2g8PnlcCja8Vs3svbvC3k7oif2fkxGYJOpnBJA+Mp+4XK/F2ZEAgToCMtdyd8YLaW0HiPdn
u7iaduIZGoJ4NICjuL+ATNi/pAFcNeQS27HB1qYUu2S+NX4HD2XdRASZVSkuWUEa2LXq5x2lw8/w
7M/f4eJ0qV4z/Fj79811vUQJd1ds5TjNGchbSM5TGydxH4fEEvu89KaLlPEh+LfWvmVgosycQ5y9
907TQ0cu6iiR6ecKk6KUSxT5qc5y332LQDnsrb+UP96BzotJF5tKg98gQAb7dC8DJSCp4G4vKcbQ
0nKAf42us5NmgX4yP9DlMg+TxlFj8CP4ohhhwufW6INwIysSAMk0AbamH/W3JEGfNtPSgYxyCE6C
EAf9wM4wPvwyPjNjsnN9qnrb0366Adj4adjETLUEw2Ycj88n7rCndIFkPq7IGWdyD6OeCifhioad
g2/JaZHkdqTp/HE2UBRhhggmEtRbKBCOMtw5iashwXJ+t3pGBHIjPzFX8bXCXtYbHwGKroQqh+Li
lmF63KvNB0Af3uhHPAO8IOifXrzNxmxDRCDdIlhC6Wp3oQ+Bs8hflSN1CLaet/JYwJs+MTXvax5s
sRR7/0KOLbYmeh4kcykn0gBkSXXH93qxYC9TOfm9jJubj4qq5DYNdtInEzvV8pRfK8RWqe/D/+Wh
4RBwH/38sgUvutuBs5iCmJdDzW8yRhAaSkMLV1psK1cA1soZc9WIwoC575ssXci5TRw54wgVF0P2
B9riUgJvA2EMR86INCjeMTsYM7k3LQgNCGvEEp9GNhO0neuhO+1ZFpGOIImCdPe42GxI9fjOQqgn
xFoIt27BsC5onog70h0Kj4TPjV1YpFziOjGyoGCslGEjTLyHcU6ckhlLwhPpxDiIOQS04XICvib6
1g5yF6YA6+GV4+XaJ5tFZ94Kn0T28FEDZ7OFvKtaUwGtk1asg6SYgUhGDznwUFvmhNlhDAv4so/a
+T7GGMvrKUviXTcFThqD/+FAHYrgLkUCCWiNC8b3eSL90jx8gdRPckicGUoJDoL7EyFjLnhKyIUh
WFMeoM1YGd2l7PIOIOAEg6hGZ4Qr7Z1V318racyxrIw/wDNS4T63Zd8c+AYvwVqh/Rwt5y2Zs9F7
lsKEBi1hPrPXf3bU/6FtZk+gw5ZLAK9rkczrvv1erwW0S6+h8PGvaIFO9zAE9IG+buoounK14CqD
XQIa7XLtt4OohUdZ8Ifcr9s9YCBxbBiQ3NziQEYUmLk4oaXLDIHEfqMRkGOoajxsk6uje0jkUQrL
g5c59fwUZg9/BUcJL4uvz5u5jaWLJfNVkPaf1wJhmKw+BBXGPgFPFJmVZfVd9wZ7SncnSa+ndX+r
iMpwcmL04hW4fspycRkiz3+2yNhDx43KX3sDmQm3f3dT2wfHPpYb4+baFWAG3ok3UT//DQYudSD0
BwclaWzYjJtzocq2uK/P7Se0gjALcbMtezi7fpTfMYe0ZTf/faT4JyR12nwaTt9AkfNK2inz633n
YM5N4t7hPtWxNrUgCqJmJ4rB6N9/ywgKJJAGS/0pHjxb3O7hQS0x+p4kRoEFJHdHTQKgTYKnj3K4
F0SoPmPLOJYFmpVvIcvkC8//O4hYfGJnW5PXFaII0oGBv4Fxm5W6aFruTm0KKPjG6QADn3Ew1MBt
vi0b2O1f2qIQYudvIDXqz60OjjvEBtO4xaQoCZdTWakvCVyUa748CrtL8eQmT32NqDf7IyKAOIo2
DNl7IcTRn4MeyZkIBH+b0eBPZqZ0UZcg96vk3ojwEokDD6Lxm1inikIa4+0e4ly9k9jtz3ZMrs3k
8kzvlPm8jcMH6HsUIs8i6iDUVOvIstpeZ7H5enP5BsUuFqYKIxt0KWZhVNnaKgARwaxxGY3gN9qc
Q/nY0J/wep5tKhuU1U4YigH/woiL9SeTIhvLCFwLeENA1BbHvYfiQSMIfh1l/OpGqt1u77PDEdyF
C93NybYaYZzO03gT9WjW/I0XLs89iYqxKY+DBaAfxK4U/bYfpSFZwuSjEvKa/QUI5CR3kEOuMj5Y
UUOkeYZmGJ0MHx8DxwrLoXp8SjL+8WwwKIbtVkHlY0Bl+2UNInbbiVE6rauWW4ugkJBApsnJF1mi
tVEjfZ+pCTj6n19YvXvqWxA6QLhHxdy9GzXDPeLc6g0H5mxfZQVDOsZZRSkTNCIJ81kgRDkUPZhE
u0b63RQfyazZpf4LmNJ5fItpXje3w9cX+stSwmOZwYocOmYjtOvaTvR+RywAxcntGzG0CZ4qNU3M
EWD86zsTlSatiehnwS1je6SiQ1JBCt2bOYuxMGkMaFhi77DGyj5sE1nLmEWpCi4rnR3rS9PQZJDs
UolJ7X+3O5imUhsRmGtMiOsKf13TSmE8Muhl4uoO9gsDxOcqd9yN5up0j8R9STuMZQPzAsYoYoBh
DoJ4V7d9lRNTj/LailkTWRWMoe8F8vsrZXJhAockzFsmt29qMda35QSlqOFFsyaKGur+1HXs4eJb
dBc55LlSDDej2tcH3Y2PCUbVDHHq5Pon1oa36wbaq3j35McDm1UaZw+TdsRqsIVd/tgvLrpjT7sG
urYo9XgHvLNxJuc7wr200WWfe1YFJTj9VzKl1JjMpoLRoL/QxG2KU/s4nLb80uGCjHd6s10bNkm0
5nXTKTx4+6fBlfrD4s3Q17Roq+3eBzT9N3HVRROuyj7JmGjsKJ0pnYbbfu8ve2tJAN1f0cOGaxW5
GfHsPko7Ime5wtPHlD3ev0g/5B7h/C4Z/pdNM1wpXOYR87j4n0vFYXuiph5LeXQQesW/r+J3LifL
HXNcdUS8I96P5p6qOCCVfBdYrKxkQO60A19D6mAk774+nQLJGLUFNTeZaXDpo3OqsZL1WRmH+B3p
zklvZWw/DbY6ICzXXvHJ/ZUxWga+Ox3sKUR5oUFUbHXe/OL2JEdCUjAyCnVqOjz95L03mCw0zaxm
GKZrh1H6AIB2/XkU8Hku7gZR2IZnupASY2qfY6tzrhgVUmZIOjRIS3a1PLdSjRctTqXF4Ol3bF9S
vZyS8gk7bnI+TnGrcxs5CbAx5jhIbKH33fzxqJ8xPvagB488z5gK/dfR5jCnJgdWy1k7NiRnnsXp
0RvgR94Je8Ek5QWE4fGtwEQzAYiB+KPLHrhyi72Zuk38ZFPiohWkmWjfQoQhPQEpWGD1OMeAc9tu
rKcx3Yq1jxX/Z/sjf5M+fo8X73JqE/4bROdyEvdsGbgBkPGTdePGiuJqdyA+7tHHaT3raadyvYL6
AmHBmie+QEWVaJPkUu4LVs5Y44mH6fCu2Fq/h31ABSZQvY7u92OklukMuIFKMLZUdhWHETc+qXaD
jDaYAjSAYKK44EjJ5WFOiOoapicIu+jNRg3yUCjUWEDSiTzXfB2snc8wpg+jGCjVwkLG2cqSLtFU
q5rNy2RDw//p1V62BlsR48H+YhddZ+7EoEM3yN8TI0uq8cGrpcGgDy1AQEk8fss8YXZVPM3/piL3
8X3PWNaNuw8U34TicJLq8oaxmGL+SLOyaMzSsscWkPRZkf2pfnxNrEY9Qhek4JCd85KUvw0HsLzI
KaWb+VW9G7m0z4NqOFKkkJjjh0KsxB5f4wxmaymu3w8Yl417K6F6hI4XNYgwO33R5Vrq3wxPH4tN
AO8dKHwpMDX5IS7mx230I7A5csNbJydOC75MdztSCvKS72h0tTEodLxzvFloPGdg4DHBuNPQAWfz
PXy9JR7Zq1Hye12Zb1f/X+wdE6dLhDS/JYpp+8uFziygl5CRYWjiFeNR25JC9Z7hGu813d/obsDw
iMm5ERm6NOFuEWmwq4I96qlS/TO5qLnNCh0dAtEMMqajIurSwQe1Et16U/DVQsIeP0NWss6yPQUX
LWRPOiCR+flRKnKP88LQnuFB2yc6NVFQ09/ANW9tcn4ShV+O0F+r6q0s+LcSy9F+mCC55wHDocUJ
U3Ne3Texy8leVxmPADcldQf44ceIz0a6WcV1lOR9mvVpfRu+tDwqGABPyTQl8VK5vj2mXubyHHvN
ZNDzjRHujXpqJl59LKz1UEm/CIPg5OnJUpERAarKzfxt2Or4KrPqBSv2IVOYHUMU1ZITx8On5kJj
5Z+qRxeXbmCtoJuThagvgesxkCHSiUTFahTNXBoPDh8vKuLBZ4cJoS8qMqdZ+xGtC8CQlWLmeIh6
MEeJUiHVmRsROnGpSkJb9cPcG3PHZoIBhk/DcnH4b8mC9zcaum2iaWgb5zSMF+EUiGNtjhDiWmOC
9KMYBQbFMJP5yaDnkePBnQPKXL3Ait85QjV5jYEXYG1Je7r57R8nM6KaUpx9qk/YL2X8LlAC2C4C
mObTsUPN0C64qPzoRntvU3DTHp0LMoaNaM1w0dc9Nvs+ixYFLe0ejaMTY/nqFWe+D2mEgzXS0PB2
HJchucZcBYUEZJtAOfnLE3bA/4veQVFg1Q6yNgUYZkcA6KBF9PJYrxVFsWiUeYFJ0FbjLi6d+Qlq
pWZVnYrzjczo/RGwuzBB1eewJ5/4bKW+5vc0Y84qD1iFT2Isata9ZvwRtU+Kl5sSds245irCGJdy
l5fVZLGDbLgyR5JbXqRXgPwmLzDTVm5ZxsJZ2jIt8mVWYCmLK8sSz515kmS9ZCD0RO/ILLSSmPmI
7GJkQNyAZqFH3n+Obn2pjGJTphMgN94Q8cNkicyOXMPTBhT4EERYAtGhtLGDYdkdmejptk/fR0SX
UCY5kWYoAyRnzO+ZQ2PgpcZnsm0cCMJruPCKA2cnhI3I5mSVo8a5LzkOa6EMqUsuG2kfy1/8J2cD
JeHk944N7JnY3zl59Br1n4NOOKHXJoEPK0Okgg/w66qGRisbP+BfQF16DSF5rKKuS1ER97KB+HSX
P/zoi7/m3iy3lzU5XZZMgZLWzlRgikyzllJ4dVpqL5uWY53ObcVNerZOByi3qRqHVoTE1JEoAyh8
ypJpfhY3dayeK6SsZASFgjX2dXy3p8QuZrk0590Jv4opK61Eq7oyWywR+5lhB9Hn45SsxtDXaKxw
npfMCZEhw+tA70xBPtnoyVAyMV1L/t3yNGEdpR+1wMTef13APvi85Zai95ulauWC/Yyejlkq2KXO
Lya/lqBO0yd8NkUik8oU4jQgO4y4+IFOLpdxI3Vc6WlaAXpGLU2uDlza0UADvE8LCJySppPv1/tn
2YEWLeRoJd2sDyYle2CbSQcfNA93HQGr5czWJ/qribEJvtOof1Hau9KNyjnLfDhkJ8byeIfNvM3n
15861hp9SbXwA9E3oPSd00VEA6qeby087+aMIoL5jM6EUfgJHJ90nwOtAPvYfJpnO+3ynkuKhQla
SSooSJQaYhJkRrLG9WS7c4RFZFEfF5IMD3avybbxKHWjyLPvc/bRqvaurZv5scj30V7aF50paz8R
3K5KcWsjW55Ihim7TWS5j7PZquGnrrb/5IMugvR7rQe3ElZ9AkMkFR+sV5xZahKl5mqXt5MUSust
+Ig2Li49u/ugJK1Ffh6YudfOqAUuoGvCC3tNJNom/iEs1EJuTs2FfMqmcJZHrGIAeDwdzvgXoUqF
Wp9A00pEafjWDfThU5vVjyhYZiRQZ5L/Oi/3J++DVpn37S5QpltcuhJoZJZsgmyp6Ph59O7rKnry
esdlGaEKIQFaH0fwFyhQX6xCICTXgKYNIfMawQbLCrSNHwD3PBfLFH255dwB22sx4J3CJtqjf07U
x5ul8clXu1LLC/NI7MW75jppC1uzFpjBa1s5/ltXXxpKFG40qOYaprRHjiyLftU1ImTD5fWloKg4
CGL1t0bM6iLhtth5QrGE5KQYtfWBn4v0KpOnbkV5ObgYTemRLUtzYJUp9VZgYeKjsg0DdAm24J5/
NGQTu0lrnax1O8EW20W7+aZtZB6zhJDq2aJuuqWtMh1n+r7AOWWTJ4091JfYKkTx+Mxme6Z6C5rQ
M/0/+h5iNBHXJB+9NxM4Ggk5aum3UPC6iraaEc2z1/t0pzM/Mezcj/ZuOUlDQF7xP9ubzvJ1JKsT
Fhl/DlYufANtGooCCJ14eU1nn9H3OT1dg7fSRHgapXzL5ZozjfCRXksCL0AlxGRykShwbb3rJj6+
Qi6FuQFwGYLBVQMYhBhqltj3wstpSZBGb/5u5kjg5i94Wbt6CRuaOnXshoIcxOrl5gc2C+RSrOJD
NZioE46dwaYSLNp7XL5dVwXcPBSZexDsI9KIIQYbQLY+XbYllSOfIkarU+ck2WStb3PbuZQJcFJZ
pyLy0jjowfnF6gayRmHqbuB9j9+Qb+UqjdxefSpkPySNoHkbpUaiIRldaLZ883g+Z2cDGW1dyLCl
U/BoLJ1JAPjW2BD6rsRErmx86vYaUR+q/BI8mpVxsMJsPdGChwiPW56zNZTK9aUUk3Kx1zXN0o4k
v+wgEzU3svGLOBIpz8FKTQAcU/a3+lHU3paJTJzM/U+uOfoJeDOIVcQ1q61P7ve64a4+5CU/SlFJ
Tu3poMMfRkDsfMsYirTOO6HHRSDhMhlf57aL7/7oDP/67MD3h0fscjukaHuLA7TJzZe6RTZR9tTS
Fp2xsh7IzhMeP9b+/1yJJ6+GIixCJH2deND1fPCZPurqlcSJDeGv2Y2rw8Ijo9PNQXoIzagC0xs0
8HLv7sZCq+B+QEXdpSyZab8DzGFayi84dJYNpcORX2mbPd/rb/Jl39k2FPJyabyHe+9F2bPy329V
rlJB5UaRx6HCXt5Oj4HJXZwUlGmo//UAPO7pO+CjMJpFvUVA34b2zu+QoW/6VbhkS8KacyaNLUJE
qm+kUGG8sY//WWZZw95v44k2ALUjyMJKpQErwuGfEB+x284J9sYvHH2G+fSBO662MRTVSfESFK4U
22YIWbr5vgvmKhO0Ou3mqCRDFUoi3gGUQJDVPkxev0eA0LX9px7odIXAypfAxJVFyhK+Ekm1jl/E
giBUUrmDZor10FZzZIz1FjqOvKkAkxLH/dI/V/OPi0XKQE6TpziL/BfkaQIFzdfxaw0ttBWinSux
UYd2cfPmel1aSsifSKVlTCvtP3CAlU5Jv1xNwi4KT44qTp7XqvWcbxnmKlxnx/6uGafn5gyXyghB
mi1dKvmVznZC/+HxPnQORf17e0BNQxQMWOO2YfZhHOomsG2W2naf7k0PCuTzgRmBBH3qO632dBlY
z0ua/ALWrowQZSnlh+xU6O8yCodVTkIM+/liwi4K05Mf6F5/fNt1pHQ7G/xWpThvzAN6AwJym94Z
Bk7Qb71adUmVszpR6JKDCq83oylm9SsEOrlsddrHpgT2dRgIXSZ1akFEed5/yMjovDLmFTs8QEeA
aUEO3DBvVFoWZCok55qqWBkrHLlFsAl2+4BukloM65uDSnuLTWfcHmKTOP39iGlEWIpcDNQ8AwQZ
iCPakmusFPaAC0G/0F+2+2No3Ra0yGqmoWqAofDySeNrrqnaD9m9LF3+0rPZGjRwAsIu9GTW8WDY
3Q9dzG34xY9TBCF6RmgTSUgBbmCp+izEWbuUdU5jHivhxAJYARQVe/o3Wv6dtqEwiQlUuLZQ45KV
pYTzEXOT8KEmD9q+cq/bywQyEMQkmo70OLqGwmTBLmerLvju5RHzoJ5QCtQghNjzpsnIbhtZ9+WP
ONY+QuWtCWLgZRcfSb1zrq192y//cmaBeYxlRiyHCcCq4XcGElWYpgMsdRwM6ee8yXk8NmxMcYFs
7XtkvEpRexRwy6JirYHe9ViGl/uLOmSUT/Hwz3Y4+PDw2ID0QTiYSKze6+LwgC1KTymlIHeoVaZt
9CH54aix19txaXbJ18iIFpIKTNMZP+9dRBzeodpvj6ZxUhJxP10/CNAw4b4+9hPLuH3KsCRm4r+u
0w+uXscJquJ/AIx7chknupaNB7sJ8W6/haZg4RCxtPSbD/Zi+m7SJ4arQWC3YtZPBnPoi37DIgsi
awPhYbsR8PKU4a1CLh9CT+c8rktG/u0usKbZ/0Poi+wCCrP7EDIuBQ9xFSkk8fsVgqnqCMPM28Eh
TNt7rOe22hkld/udndndfL8jmn3u4UhjEzE5LsHibhXFDIvZXifxhTXeatHOKv2cUBvMxdLNzRJF
cBUpd6YtAy6il3mcHNSFncbcz7Vsgs7yEeVlovMJSZ+Q3kWoa1lv/p4W7LZnttOTTirYQ6s2W17q
nsPUY97o88hehwgXZJjoQ+jxsekM0cxvDQA3iLF9JcesloeE8cPB7nNBab3Zh0A+BPecv6eyqaSK
9YMkGvDtEHNyGOYx0hlLLgQzQ4n4ubEsP3NbmE1wvaXuOqu+Z5haojcyxPuxjZAV7954GthxD1n/
s24qm/EOhWlaGovY4rJ6via9/nL6MGctYCtIS08ZoJLbIb+qxgWeB2HbjsL4LTmS44VeuyXseQne
V30pcwWLmDUR0O7W88dVtAc0jYlkOVwafUlu7Hzb8DdXYav1WghFesMoRlHukylxO50IM069YQ4T
J10RXrfvgzE27jFQEcQ7vceAswca/EkiAO8q6wS6CT249674venSerZjJFpFKJcYvSjYephRrqef
kxNkCmNViX+9549DXoxRuYdfQI34ed/SMJhCOueNU5A/b8ae2iQRnnISvkqUn2udZqI5xEufODHO
bN6BrwpQXAVQEcU5SrRvoRxVV96BWAs0V3etPz8zCufTw0n26rI3ThF5FIx/QJY6hMe3MehL8B/M
29XUf90lJ3dCD7THJrV7t2gDYgyjgtKxE1YeYv6+EtgW7wjlcxOzzxKc9ZFUyTiAFM2GVhFaqlt1
cJCi2/UAQZJ0UooA4BzvWc2xEyGDrW7hLnWXNcAgubUgg/dq6WRzwh5fbwDfHDckAH+SIGj3IDsi
KYeXWTO0XDBwQLnIiscxeO7HC0vqegLaJZ+VjhWqFfG/AolYlagTQhaByrAXthKYaCSc6gYm/SkE
vx/VdrBwKs0KdUiXVcjJNIZqjhEkKZQKFuoqkgMcGOdzmvMuNxhQb/6TaMWOrPzRGOW+f19BWNyb
t3NzexJl8hSSKCwp3k6o0n8yaa9hEIRTVLdmgr7BHIa6tY4M9KQXBZ8//RhL2zSj8jIy5ksQCdpJ
IiWItAhxKUFNHiChwzvXDNj+/qHqdKukwBfMoHgpb/AVk5EFcfmnC40UQLliMPR30P/AGCf6oJQv
rIgORVDrs+ESgcT3yUL0wDAZPI4B/DGgqi7Dg/MPjB+2j6k491GxZc2AhkJvNntTUeRRNxbSBrn/
QD+Dq8GMJdmV3KO1Ds8HJH0enW6OZkaOFFBecFPByU15+LgewXQgIsDS5QxSBb4oxSRgDtMK+bU7
C40Z0KPocEaK7eaItTwaZksDf7EPl57loDmXzm9H9Harphside4UWa072GV60JQmUbA0NbO16m01
EbNljrsA46NI14ZGGgJkTLTI/ctonpGjHG0Okvz+C9tWzyuPsFlwaNdWM+mqnep9qbH/vNAHXJjM
mqO20npa7A0amtmVaaN/4/g9j0WIgG8gth1Imvj03WmH7z03rzR/q27J5yopZk+TiTRwheb+S/R5
tABpUD8J1aJMRXUKhabWumGhYeto2tV2bWz2P62PDUR0yCXDRZsBEqJ/Z0AOIAZ3uFwWT1mUw/M3
wm03I/EN6hynvqPx5vB4aAdDAJsqNQPs7jt0Ik9FFX7IukeXqTQPsGsIWemnb/5wlWE7FJd5AXHN
SK4+UMIV1HTBnDdfpwZFAwAt7Jw9Mr67jp0n1IKpUYp60sV6OLgXFa64I6CjaCCHYxJ8zQoPL0x+
L6qQiY50PdXaD1NGZbAabrEJMX3IaKK9zFGDrpYXY6Gh4Ddw8e89Ud516aZn0Czxi00PFP4AgVan
aBoFQGOu2bmcmQ+mLyKZS7Kl4rG8wS+V+EoCPJBtAxoWypubpuNCAwwWti8osjGdz+IwmPGNNqgX
fq3MBtiPkdlgsYch7/rcd55sVyRuyA8pQpUVEEP0XS1UT5hVIrJuOu1cHq/ePuQ9F3uNsOv5S/ak
RVCuc0onunCIe9dzgCnzbAtJJ5TeGmUw0euZ9nHBK68zbiLEJKVvXKMwldfnBaBSuNyXTYH2lE7J
OOJxnwtb8LSgsbN4kLKSjap9ABcauOtXHwrjoAAsmVN/SgynU9F3Et2/VnYh0CSZt8QQ+ZvWfrnN
8Huu+3X2N3iBqRIEdiZWDEItUcwoYDhJ8YKaqzd/ZQw70RWXSLd0gKqnEBCZNNoK3230QOD5aKJZ
ZUR2LIp0J/zhVdNIdUXodqfNPrP2FeUYSH+KkDzI8x1LaTRF+A5mw2FuIa8v9PjaE1w7OaqtU/Jx
HXIT8JS9didS5YFrGaEuNuetAZig3YCCB9H49flk+54V/yBqq8tXW7J+yXnXNhugKtf0qepRF0HX
9T61qKqxtBOm+PAPwh2bU9uQCPoLZTABmpvY6TGsrbor6gP7fF3uIGhe95kqHUwey/eBgPIZIPyS
5ghqXhJWEfir9SlsficLxJLAI58sQJ/cw6IjItEGZcvNNd8pzVULBdFkAE0WTuSb/qz7f7TIIls/
+mmNvxYtV7StK/O66DJDQk8lmz0bqUxYLjEhUOaC9wVCwidc2JSG50F4qono1jSMibhcGahQ/y+a
GA6dFmyqHmdbS5cByGM4UlT6s3M4jcKyIkNaUO0M3ueYpS+Ge29REr8uc5GE1PKzBY3uJtKAVVa6
BoTiFL7uij1XHNcn+rCxWtcN767jvg50yXhP6m3644BO6x8eLFSzTxN58H0qJcz3XkRQWVzWysO4
mw2TsrbrNytIWxdpS/IWnxFHcH2b1z6hLmA7vgEGEOS45Q6wYwa3nmXyNMfs3HaZYzUSO2V1gm5a
8YxYTB57lbfdAQKSRx819DlzZ2xmGHWp3noyD3ZJ1tbKFwVSBkS61cbj824OcC1yj92dOSGzlxMY
c+Hs2tANi2hluMOgujlBE5UaJzg9Y9oNflYWDz9px7Yjf2+3adQdd2yVWtO0bDjgXcwnwR0IiPh4
ojYUwxOV8dGoassNSlQgFXw1qtJexRu65qHisgbgegdxQcyttVfOg5yPwoOiUZBnH9K7+7kCzuWT
PEJqWQA5QzqqlCJDJQBBypKiPWj5Bm2yMIzAeV6Jx92OzYvnvKj0uLNvelNbx8IQhm1xpBjWlL6u
X2grGRy8bkWPJsdBQm2L4wt9D3tK5CH3zePKkG+UE8b1oCULMk+CY12nVX5irQNW3Xcd4Cv5il2i
47oQkr1lASY88hhCWATADn+aWEqiNRKsvwy9tiKwI4vRvun1QLipSbhGxmarZ5d/3KnB8ZEJTTOR
yDmtRKSnYzCkD6COvY5YisIuA2upJnPzcrs01mclb+zeMtldwQ9/GN/3rj3h8GwHnNNeUufqMxqB
TqTFzMzTSTW9LMgXi9pfq9BAiPuJRWgHAoyDMbDMbRp7bpGuwii9DxpeAdCRKkEh8tJM5sT9pd7v
jKn4JRsv5u1Tee9lzQLno6AzUiFhZPvaqY1AhlLMX3fFywXcwwNPXwWApgaGd2Wc0mIcU1YOpxo5
NRgV4Wr+N6x+p4meH4GESvuik13hBRFuNXsj3oenWJOLLknDOTh2m2pBi70/qcK9LyV/QHaunZzt
3+Gmli5L5EuWTGsy8rXjW1LZIGhdjHLdoAyDhqTbNa8LTZFtfa01Ay5S9SMYm4Te5nc8Xa8EI/mK
DytY6gdAPo2teILhaxUe5omPl3/yPeyJTTWnUFkp4I4a5tbRY++pNmMzDNV9YOBWH/BMGj0knPSj
MYnSjCQgSUYe5vsfj3iF2Qs7FqhMy20TVqvqtNnqaoSOw2Om+TTb84jERqf//ArYQMRbuBptjdLT
m1hKltIqw0PJoRuQtZG4UcVhDe6YFPXfZ/ub+6kgh9y5/k+ssN70zERyTPEaMKRkZ9b9u/yHabLg
UuIsWwHUv4CF/ch/8zjaFgXH7exMtNiO+RhjPN+6Q0CqinmSQQYj+fLdYNP55Ur/qavk8Gizk3JB
aEjkQ4BSQkciPdHk5QS+1Wwqm4n3nB47gkVksniUFZXkbeEYqkPgpyQx7IE0vrySApk6E3LlTm6J
Xcjf4QqQsFZqRso8hsoi3f4dTYCigfYOhGbskpNNv6uUF9xFpWEm4XsAyUTW3i4WcFm274kVr0M9
n4yjTdNvW90LivBpTW8f5PRJBiLK0Tmc9/DNdlFl53o6t3zRcMtnN0y4OHfaRk7CgttO989MELD2
AuREoiCEZ12lcaExV5LyfuSDP17yOCMNoZJTG9Ak06yntv6vhzLqES/SUKH1YgI9FW7+OPtz2MH6
WsEH7uosSVPlFAiiKoEOR+ack4KoA/Dp+m0MFyTwD2DLUtA1iPJT7RZj6u6aqrh5331pbnYU7K48
aC7zoYc0kI4VWRvOr4edTBZdx1c0NRa7sUUcjBAsiL/JpkZhVyqTPjQWTasFiq62dhzEK011/eBX
cqWeTTw0CQcslSP1K2SurHqm+l8HH5mEJo7afFwobqpttjQ4Jjbg/1+45hMeELJjQ4SSDQPWgf5c
2kZwsycK+Gr9uEpIJg9mpgbu6MOm9uUI8ELRsMz9zBUF0tGYvnUOa54CdWtqObVaG2UuRZ8aDLs5
vY8DCeuBxq12iPilch0waEvb813SCyNpzmIs7fRtW7QsBgqHvQoTL0PpD83m8sefS6v5NupS3UD5
ybf2SlXi3eAnb26zJbCL2w3ZSgkHBHb9tkhKgdAhJJEEarQQNxEAUU1dsNcL691z9UMGnIXOEdNs
AfptYUG6F2UihPaFjRsyTnz7pRi3Oi9Gr4fipB2KS/9cEMMtxd+LUAxui8e4BRowSrUOCo34rfNY
IksZg41zXe71GHWbYJ2LYyt8tcOpeLZDtOsveBEC7TAHpsy5d5Vpv/gFS+8pfRKjbBaveZcMuGYl
4L2g7NFF2nTGLObLapqtCjsGW2Jzz6qakQ7QdHHpJ+YlboC3RCC7Qns0d+mKcR6k1jQNesWY9ASu
u4Uc5ItgJVemIwymFe200DlakSqSvP7fRpNwxc92NNc0BLXQfPz79E90kc5+2l23PV4IkDVwk0Vh
e3XF/IUj+rkfIR61GVH629XKwFxl7oB8qYULyY2kxawvjWJU6FkpuCN4PJXf868tjpZugbJ3fFso
8yktzOlTGpORdCSAhyHrrZPZrXpuWi0JMxUegDh+zRfUEqoQFqDU0h4T24firYOcLmMQykVynktu
E+Rrm3rLgchCRfxzUqzlvJ3ww0vhqUoE0YHSZj56gDXM1eWuN+YkWtMOPz7ruwZxJQCrQBFqpdJL
tF+QsGwb/zFAlULk1wpxwMZa5IWqyK/JYO9O3OejTTStouYV2XEDdT2dbVVxuT94YVifGbvarXJP
DqdnwCWRjxI+QXO7Ha8rccDk/GjH+988IaEY0+SE0m1ajgT6VAEpNI7oVtdYphapdxvH8jW9ghHt
5lyUHMNpswZRwu7XxSNQhtQlVY6diLNdewTKg1QeJnL+/GozeEbD3hj12bm8HhJtxBQVQo0FFChF
qV8QiwqE8JJBeqQragl5568T5KFniQgGBS+GnFLozSyOzP4KflvbFLuKmfPYkuE6olLP8XW/wtWi
7uDcLe5nZN2NfLBp+zjXgrDz5QtsgWQh4xAYCsBX+vdf+RJb8CnE2d7/FB1xg/klmbYmwCe0e37z
w6z6raXbja+0mWADfaWzlnBxDGQCZvLFB+4WQqu/6DxTCClg2xifUZ2d+gxS0YInZ3MoShqAUt0r
QuAUpe15N7vLb9YafImEG4KBdZuZK3S699Nru2qNeU9WgvU3q/w5E39q/6rJEj+lDsGpAsSXValc
bmpuIFGWU+SopPP2m0MnX1S8xoO2kbcF1XzGgktdA4SRNvCZtqWQEXmbe6hD+FGoViNLPsbhTvFT
pf1H0m1ASjA6qdHIgAffDz+Jw09t2hMO7u6Yvj/FKnLUcKn87DNt9Qtr+9v9I1sITwBJbGx0X22T
yUwlcU0vLys2GHqXoPzryt7dtnjFpd1p+iQ1gySUGgxVXac55eyyfdEprLi3NwK0TThvsuYO5t9T
v4wQLrIPIw49dXTX1lWI4381kvARKXLLaay9jQ3n4hBZTg5BRAf9U6DQ6mGAlkE9ycmk3gtf03PH
FhV/Ogjjn6l9bDv1o8UwEzvr24Li04d+V+zDTAtgbExh4FvHKogalme8nG/DtwRAjP8wQRnpoP8m
qam5EZTR8MGfT0+ACTcZsGQitATNv/wpx6fe71vlsMRrNxxdxAX1RtUDKAT74pgG9p+WLMrCP5sr
UqqjCQ3Cb6lscRVm7rmkow4sLhif3mczNjI8GES9xXecucqiq0OGZgkBNS3H9IZjwHWgiXRwCQMV
rcoBKZzocxZvnTkxUOUOKFxzj+C96h4S97kNLozwVDkXSMyNO7UYgl2inSr5+RgT4G1HWEEunqUd
VFJH0EhHXU11uOnzl2b0rBpNKZ5/n6Vgc+6+FRmjf2Qz0TwAQSMn6WqaAuucH+syIEUDYM9B5plv
Vvfq1Shqe2iQBuNDcM+zF7GUQlURsQmtd+Z5NDUA+u4ErsE2E9bAD+8mdBwfuIUIOkG+SgDrW71X
KhI9A+GfPjTj8DB8KUOir1DvP72IbDJ4kIFn+4lTxyL3nWeE9YqZ2nk2LhZRU2kROBdDVGTdIE/W
2VSdx8Qc8FF0TPA61kfepOQp5mKK1DFrb3G49/S9tJcfR46lmTG/0m7fJ6dK3DG3AcieY2Luj0X4
RAGE7hrqjjEBeRVXpX3nCLHXUWhLomTfv1fkI1ak36tDisXpwQptf55u2K0JBjNHs3SF8p8Vq+KQ
PBSwh6MAcdToWCKpyAFQERTsCZntVi7Lv/iM8lRwmhrIhXtkQXjL26x07lxA/JvcxGXqP1Nh+pEC
5zonHK1ekJG9w0vBGEYjPJHM1uoXkMLVDsBPdfmqY+QDGUiCHEjj858s6KoIwayMMuEGTbweLmMy
s8JK5Fdr5hyUfb+Yqeukc2jLzJD1VS8EZJ7Ll/669LKv9+GL+MYxqjxNNAwXC/OCXGAb6QjSNwuy
ojotGM83aAZbMfcIpngWlEb+hAHJ48rX0LTZpAZIf8sAWWWYjMxkv2Qrscxh5xcL5+Odtal/pF+4
W39bKs2SsJedhpW86HAI0NYFzON8Rlxf43RwrmYpugKPtRw9kdcwticI8Q048Lrl6CxXklIIn/bE
mJaLiW991wL2hdSZdopJ5tz62mNLzHh8wvqu2A9R1GaEq9AfFyoRAaPJPjJnIVBzIx+zfax6vxdL
wwottqWNsk6P7u5amlPBNHYcfOzqzarMNDFzRlZMjTqoXAatSU8uFr04DLqzH0iw0KTod+s5rR7A
swP02UqvdBfHilDfAhy8sbMv+1AfERterXNRIo2fREY/lmUIgbTCN8o9uRWIQNs4vDHzoKBjXVqE
B6jfGZbcw4uk5fdAOWKRExC2/u+y8USGRBBRcn8DNk1SCDQoq8WAjZKHOpKeta4GaymOOO1SCcnT
MID3rG9p9hRwUS42ljhh4RglCwVBDrXnmV8dOXRj8z/DZbBLhWl5yBe6kEGzFFC3BQLgT9z4h+SN
RHhIsRfzmVhHRHHbyc9eJ0VscuvCdtZQoC5rfDdlICziELQ+7d7UCoh0upy8/v7oSUn6M5xDJ4QM
UV+Wc3ktCRmpVKumGEGEuH1TD1fWHl4y8FworSNku9eaCHbLdqtXeX12eplpPGxCnE7fwZfcHL/C
CltnRfz7j+pnbp+cgmzaogwf85UcZw1W48Nu9EwayoFQpr4fzNlxLwWfs1NXYxwzgAxGJhAY/0ne
KLCltUH/uVpExZbXmJFcWoTLW1btlbnz7BqaSl7GQjU0pA8xBAMB3iylf0Oy0cqrkse8RaoxYaqh
tyJYtjLui4qLonG6EFGFBKgPW746P3UBus01mAdlHXeRQI+A0MPxttJYsXnyx0uTs2S63KJcPwYs
QlSaXn4YeKR9ZXbEGynAG4uS+1kQXFBebGc+oDnyw4JmZ8Duy6lJEJ7R6VFnAydmo7vuUPW3W+87
ud3htbQ8h0FB3kAW6w1lgkefDJ9SBzWSYH17Tp4XhgKRBSMu8DDGBZZ1U4Apu74lPmxiVT4ICpAi
4ptiR/upYKVy33hksuZ+1bPMfr18Pjzd2lo3LTD3Zc4H97nioCn9VBZqWAakD8/rz//0TOIAsRRV
shvaSvnTrdmkvGFhWFFRggd2Uhjy04a5G8Pnq/Mna2dfdXxZmFp8L9PbCKjEXoR+lfVFIK/baWbo
6c7yQve+rZzvaJdw5lD4HbDH1aPpo45YQ23CFoBpGBO2IPWvuE8n9CmqIzD3KPbTCPgVKmBFr3/u
oMD4QWNhvzvNPN/iOaM2bT/1CHRnyEx5j8aeiNx310OypPrCQQgvJ3l5I9YJI5umFEGnRN52hue0
CCukUPpcBDXwl+ATXxqdddq8WPGYUJlcnKamaA1FiqneDqbHuuLJ1YDydMj3lmzDrywz017O6VB/
r45hOo1rbHhbBHGiPWdyKuEChEmwcXgQB7KZ7j6Sg8DCGCFBNmMvb4YqdkHykGaVnZ1CyEJU+Tpz
ujKpadQdJCt28/jfwjp+po7poh1JoLG4je4j7akPexGPHPEyFz2n/9XpiByXpLsCE4I/4X9eS7g6
c+ps+kq+NnS2NnfV2UcJwtSDYNp26JatYy7JXfcwCSB+dKsajK5QC7clg4hQRbK1lT5Dt+ysF5uL
tO4ViZFVhR4XzdgAvSpjcgq0t8ERKui1GngNrqq2z9cA/BE7BnVX/I41xv99VAnUYhgoKRa85Gao
z9yP6WLgjjN2FZYt35ojZZ1+/59EOC2Q4x5xeW7NgMFc/jAutwEnJL399WRecwqL2U3w2MRwDiVJ
VR4dc2v4YOfubF785dOzWUgozSmVGgViZTrDHLJERDnv0/gt2+wGhOfP2qFrTTna85150WgFGBC3
8RBFyqS/P+BlZ28ZPdAltMcGXMl03W+yrNKyiBC+n+1T+nklILvNKm7ycJh4RmMaieHzv6SI25Tc
NlP7QNbOjiKsozbMQ3sFGZ2abQVDoHtzn9upvhmsPgKRB05KM7MEUROU4ElUChTjVOO5woS+QMqe
eTv6v7ifnY9THbebbKj/mqMbYOT147auaYqK8OLqRPSV4CuSQtqTxzVaL6el6qqH1f++Hn/s/9S5
XZbm3qgWnAnVe5gsft9fTvVMOCWmbSSrFrnEnhzvj17ID6qx7CXh7+rowQsPBKBwODqJjWG6Uyvw
pBG94p1qDAv3VhYPuTTylrZfvXgw0sXTr+7jkAIEP6pbkNXAaGp7RfiAJLURkjXVR83EB9HV2hSr
AgioE/Xsq+j1pV8yan/EPKfjPsBxJShEo9LvlTQW7vWsuGi3U5+tcdkSUbKCLKfW/EMw6PS/58Nt
mu+MzcApHLTpbZUvrFj5wXLhIIeLkYHTZ9ZsuhJrBLsHpzcJ3thX1gniRjNbzZmdKyDzAQ9aXU09
fzQpzyoqs8DQYTAU+2tobRBNyrhGFZzg/S5991/wk1c7xU/+aV5CGhBVjSMdkCzsHgHF7FpAGjhy
oYSbqD8qUZFSofB6lMhPlt1xqOXD6bV84yAyQSRd481OMedkrHxOIKtDqQBPO/5NErLptIPyALPZ
Wu3cmwDreXA+OVDs0WprYKjAp13+v8Mp9ZZo+Iy7mhDDWAX2LxQ4/dqgrIaVaKDkxiNjdHfpyXH0
c6OsxTz46SFxb8g05zSUr6m8eJQf4tn0a3kHoyhYK4WIvHn2tQqaec4X6MVgMIV2FPuVDye8j+MT
LqaDKgpDLhWu1JzaZsId0Y63up/XWg3T1TMp76xW5LXvPCEtPkbpYna03Xufp2gqUDw8peUbvrXL
n0v++0cZbbxuzBho8qEc+fN0+v4Uq+yt9uoU9YcK3GCfympY5hhMSkOYZsd0drC4YMxKoDViLH0v
PK3vtSST4WBIqsF8Vo6tawyPmHi4vmYR+2VvmtFnwZVPfdpp288salNeqXhy2bZP5XtemC/LJFxp
xTn9HhHfXdF5vjLUY21d3W6Ntaq/CAPsQb+860fPvMwz358ApmNfR5trFE0ECCeLzNjmWhSRZg+/
t884aA1UUS2V3nEd+n0wqmBK/qIT/lWHgkkGmGmYNfILt7SIQH6oVNcy2tkc3TaciUYGhrjybnnr
m42zegtVz6Ew5Yrcb4idLdIKIgAiC4C5REBvxdRFHlazL5i1GiDGOMJ2Iigfxh1aAQ4iYHga1XLl
f5pPXVAxQRNQhR1Ixa4Utts4BPWmLAkcj467NPv04Tth7EzZ2F5xi1TiME0W5aAcxehcHwE9kw8r
vgqC6dD74rC25j72OoNsh2HpEePxXZuu/M0PEQSRX85YOEGaQ0qpkzERV623wtTTZmVnurYwRVvf
PJU/ImGz2zRcl4ZvvMboqjs4e382gPAVeSXPgNAZY1eRMks+ij7ojlZS/zpLghQm2z1PgwH4R+uS
aaavlbcaH3EzomDir+tVY+nmKHBsxc8bH8nQKUcRCDje9Ry/3oPQjiUNrQjqdY0WDoR2I2i6X8H8
u3LrSAqg0KCrch4iPmKcffGbWR7vwaQONfIiJQubazUtci2nh3Eh9koZS6vdVmz0rPzesCzNiXQz
5jcjC+mXPoEaQ+TVFEwlma0Ob4k6JzcA2fBPfGJxRE0VXar+1oMGdb5kg44/o0t6FD1ChdNWuVXH
qe9Yg0IJjmDtVyg1b13lsCxFV4z4VLhz+WRMeEwmhGYTSbc6/FLWV8krj7ONnPup8aeEzhTXPT7T
fxAsUbnSlWc4vc5ChlUHOxAt2gXzQ2L3IJAFay8lmCo/C59MMfvID9ZCl44yyttZvzZxK2FAGbIM
GW6/MvFhg//4X6nTq9QuAA+lOd/Yq7+BknG4Nor+bYuOBvn66MUfVhf683n9dAWk9sC6vdgwzwAk
3fTkJfdVMdncp7S7io/QyKrpuGQzW9rUsg7FKifvSCitBA6Afo7VceM8PpnteeSd4ke/jLgqYR6Z
cJxSR1ccHEB84Ax9nXmF4L0xb1ZDYBM2N2p8uUmbZYu8tetuJmFrhxtHUfqsaiFDsJRiPr6StSBK
ksXJSuesRciASOf00tLXKv0Q9SVVqk1VXJmUNO3qXjWrqS76Ewv/7XpdTCl8ri/LDsnk86HvBVya
4jaX3YAySwWbj6VfPsq8ybiwUXP5hCeEp+hxo+Zu54S6Sk2dgykm8FsrZmPIuVTQgJWBrfjVhvxc
5ElQ7MP0gkP4TIqAzuHvHd634fJ4H+a7iy+/BrnDG7RIwbnyCGFha6SwUlUK4c8MAyoa9YRB5dJL
WivDR0O4aSZs/WthsidqRNE6mRZT16KUHHU6xe39TGDuu2/YHr3LJv3tK4Dn4nq3FCmdeQqTWBFg
Xb8okMbgpvN74N+vZu4VAz2DPmaIww/VXYOtZic+zsuPQBUzHjV43O/V9ZJ0GRZy7zpThQYA5bGI
xYf1+u/NNw7H7BSGDSu1F1nUeSBIgqMYr90ByiZmnbzEcwyHZL38vKTNXy/dwKnunvBZ4JLhaqaO
2g9BtgoXe2KyviUnWcc7teHzoQWT+D/mwR3aJKdge6B3sgOODBoRc67F/C44dAKa9ZhNQZRpCC6V
qGnkarSi7/UbuUipE5/4SE3AOUlV/Xwc7fpYeklOHYrJtjW6SEz2iX14RbIV2iuLhsu18it6Qp1K
PTjLRCD2T3uz244RV1/L/+7RMYf37F5mgu4hDN1kx5J9LgvYIFIEJCOKPglFyE8Jgn/n87+J7W9q
m512Ri2opNmPA8uMz7HCSBjWn1g2jl8EBkIdDno+dg87bS1/rWK+pOxwld0KpTLZrdI9CReeMSt2
xE/9zaEGR0NRBuh/cYuM9Jnt/M+dYnDCWQHrt0H+rZeiCPuOwLA6aZI/8adUNaow1JdkFIyWSrHG
3WJujDM8bfAHikgyJSn9Cl+nfr1jaWKGod1pTxTB+fNDAF0gG3jP8zMEp98nNdSIhFlkJa+SbQ7r
WcNBFpm91HIcuGYCYtLWY+jRor117SA6MEPKwlgm+srT8npTD55DeSbxpZwRwpvg19BM+ehsUNN6
LqGieAqhrpvmSdZr5cZUIUMIecuP+RheAJJ4VbGkJmoWp1Lwv/bNo4u+gF/+gyOV1RBht8/oXwrv
ucwO2tU1Sp3lzTia1zar0NVKIMqaICArVhJ5Z8ClIZK8chehtbLkogqy2u0UfWNtU6x8ujWIoI9q
LO3hzSFRx93bYhOjtcvumt7SdOPFhBPFmP4kAHJdmzamZSBlQD39LzQ9MeQPwz7dkSPZqT6X6vtj
QLJWpq10aOsLQjuaUQvuUIdo8E3m/tJJPIep4BddQqqp+sv7jfTccCXr3fn/rLBKMNa5ZFA43+AW
qR//Q0MOjYl8YvYmsPrSrpVrve66ugULbcuLflL8xdOSOXkNV4+rqAzgrXYhee8JhI0FkyeV53VP
OYeU9WUUiqsHW8v7glo/hN8/hvxSSNf60d4kuxq+0KQKebbz6peCD9wQ6YXAsIJif6FnyuCKTnJ6
zBlepANWQAwnjQMOSM3PnEh2NHb5VsN+l0RYiix62ehZsCleTEx5NQDgt9V0uRIBgLgrfzQyCp68
qx0N6Yqx8FiNoPAVJei0d7Vcuw4rTL4nohNU9q4xmJFJwhQnEB8XwkJspqY149QFrtS5inFiSQbM
XOwWtJZiteN0w1Yr2iVVI6tRyRv5yMmD8TTOTODoJDq6ORuTvclgd+2nYjAqDAetZDNNRmwfr7f5
ttxV9qBf2UejEFZlYTag1A4tK9V4g4ee3dJ9lssZBlkTKX4brJRvWSXPAvI/pWQZoRL/OkaZLfKJ
Dcc5cX+ly8hwHy8C+cLVw0YqV5wzycWvQQSg1UhNbUYjVkxc5nWPuOxVa7cS9mRo8rJ75k67N+nY
kOLzrZhUDpgBF9q9cFD9BaO97+/S4VLWli8wTFKFAIauNW28Oo/MA4Ap4MswkR3bzAy2gj9EKyN0
ceINAH6RL89yHPC0sNyQbyzujjq2ovzXKg+6wzZYqMEYyPQWAfecz3cXhsgYFTeNJmugXnTcpH4I
Nim+LotGLwwjmri1eiasONTtzWvtRLjIj4mf8sGFsEckpGLsEhvXxOQh+XJokM/Fy3p69PgZCmA/
cl4yBEj/glNqYhsUzO4xosSi2bHBJ7wUMlvSH+qdNcD7Yi6Y1/JxMGb60/jRptz+xEKRboI5FqqA
t8BTRpNIj5sy/hAbao7xipiqp3C5mP0OKAqvt+jsZwb1LlFPbb/H2QZrWi4AptiEA3d2mpgfATzU
gDS9ej0xwyopRFHroOpt3fCLtSDHx31xFPEtWPBhwNMXPlQCOi351w3eYVFNx6iVLxPIOIc6W4qo
dWCMM79wUazCRz8JLbk9t6Oh7ryb6f/DoxlT0xs2JoO8ikd0pH+dLPGXuhLxZd6Vk6i3PMdYF6Px
gP2c2yalvUWn6ycKyci2Uz1RxXANmUv+UyrfrjQjhN6aq3NtlhDVZibKU53+zXPD8/Bba314XKqq
TQ81K4jfiEG+P3P9+w567lJ8oXlZVOVB7zAwuH7SWfia/lwv7+qEKlKIXJDzeUqgOePrYTaN+623
Wb0H3qDBSqssQ52WNZ+TGLfE1AY0ARZwJ6PMLDSNLJniOfz1tYjmjegHjaxfZuQlEsHjJMbzR7Qz
P86EmLe6EoTSC3YSrLhOdVVlyUwBacmhzsJ6H1Of7iUI0HusX/IlKbsmwqYfrkrUzFyJgN3b12AC
Xc6VVHkheiNAX4xFPohqbizAi/qGEa7CvDvJksCz0FegjB8wCMRYPNcigxhZSH8LY2lLz92ilfAd
jpcDqZZBlQ+c4wF9OnbP9jclOUnafZW0Jpj7u3z+nQYDYLepO7+Uu3PnDQmB6FAF7zHDbFuxyUkJ
aoZZu0pGa8kF5eip4sCzsqI+Ofvh2TelLut+oIraombV4+ZCpKd2qhfryE+BjgOWyvuWT/Babh8B
r4wiQgVMEVzqGDTeHRoz0mCA4GbLRkE/slWqwxqQ9jOiubua1wUmOeYST/LhtzPYFk6lvZeyV0vH
YFVLS5J6wcnivsJWrJat6Nefr/YLCh68Yd6qVV9Z2frwEuD1b+D7/SV6jSuirsS4yEOcEIKVrqf4
H5XuTxDWkUAEKQ0x/Mkf3UzfklAn8H9PQ+Z8GTHqa20/h4rrm0uXnd/wtNUllgOylEP2NebDfgLR
MajfwTb7lH8EOGjKEhQFqwzqfgCHrQEulEGPCV1ZrtJkw/MiYADDadzwK1HPPo6SM1F+S2UbHUm5
F8xsUWOKeZh0AVpWVe44ijB8Z0BtGO7VBlntP7cc9baMJkwoEwXXV1qWiQkVOaIq3T/hIEGEbcD/
oUg/rrE1SVpHiqSynB1ZEY+Aan1I9+sfCw0zw+1OExB6WlhKJIomJejl2O1xAjO1eLXjI1r3VN2s
YzoUmZfncbE/xM9puFMLMfutt353pEJTMXc7t1Bj4MAsr2LP1YBwFPBYFzMp4G1UYPzYHKpBJseB
IV5awUIvNWje7RtqItirQT3JBkSALHxDeeM36McwjNdDC7o5TByNliaLEFWrIWLju0JWMNyNpxdL
zdVDRvGC4cLy7MKqWOq1sx1NFJT2Uz/vTgnk2P0RI/RrgO0UXm5cJRORpDfVzAKLxuoIXPKCAj4b
orT495IkJzRKbuPVXtQtVgTEtA77dxrgz71oc0eTjH/CfB9Ea7SNReS5G3r8pRf0ZEveia3ttEtm
+vzpww39fjCK7VDO8dKmDwpDwFqqKJ5+dHN/WuprreCl3EdArzqv55dGfr0C4byikb+gw5kdQFOi
5Vr/R+K6qUEQrIurvCTvJDJ5P2ULoeRshnSLa+XxgCOGIvSJCWTy3OPetBBY5z3IJ4PDrhyCvSRp
cQuDIw1BRNnIzR700Td1Zuh44epsdZ5vzhRZ2inI2YY0VOrIJYkU3i7CaLWBbwKHAMrQJyVtmlvU
S29eP2qUTcSszIGhVa3P5s6O8uR5LB3ztOZk+LVrbtmnC/e0GQr8grd/o6nyJLZhfIocBTIEn9yN
WqvzjZiv/Zqy+DkyIvFiLEOIHoSkRT2etYztfVXDwjZ7t7tBsZKHBiBbCFQ4gsk/VaeF4nx2NVll
Vj4CgW3UY2w340/ghwCVAOoVYGJ469o7fBA3GWMBZ6ZIsdHbIhBZRQL2YSckYFObD+GbdSL7Lj4d
I+hvUAvwIZdXmHl0ecKO14vj0XXq00bbiXoVRCiL5Y8/9ev81JnIcb9MKTGbA667LjKDq8V9it1G
IvIdxl9chY/OWCuatmlmiuzkKaQ+GHFU+io7jcba1CTI/h/nEvwWPbuGb2M/nhi3bS8CUmv/2YsJ
70qDc5hwkl2H275vC2nuQlozsrMLwAvabBPwRIS7AWSqzpladlj5gaShgQa7eXSBcBV71lLbb4hi
aN1y5AZNdtTezBOy59zK/oVfrLhpLS5qVHPUlPuXEuLfrNRHBKEHsTWM/miFakvQl0IjMrwe/V9g
GaDcMRksCWNlUJbc4AfDmBvA4plhmC+rH790DJ9kOzsawjj2QPfDM32HCO07H7yQwk11AImESlT0
LL+knXVXoxz7j+Mdv8Z2bi6w1aqOQxvTk7z/8qzZD+z5ca8fGJ8WD4gGYbB2diA2hSZQXpr6VXAO
VzyNDvVSvvSHe3VOcd4bgB7IEUlaFhAWu4X6hEIf47hVISxIR1gXC6AP3DsicfWVsMDp5mlt3cFB
xct5JUjYlqP2hvKFAtC/DbGm5XNIXHcakX25xLwiy8MkVTdCCM3wpbQAj4+O0kc+jYKfaOydrHoO
5fmAOdtsOyWlRkFCG5GugfoUQKtWtC8X2xVNdGuVhC4ktUSTDHfU/npYAy7LKqQHkXLvb+fiVlMU
6Njgpcup9F0sNzlXmnxK+oa5vI6B4yOrsZBfVtQ6ecj6h9M1cITwTyv6spJUmu/UmAdK7jZHh4q+
N9xozuvNq8DLag+tqBSKseVO/3djtLsE5NNrj07yKAVxXWXFyngDL24IFmTtLcRGexpBmHmaBHqU
uzGvF0z/R9llt7ZrHcI+YUTdOTF2va7mParNg1qz8k0tzWnYC6HTI/QxvwA+S/uyakbxoxjLw92e
ISrix9VWXg2tj9rWGmvTT6hu+s2o29HrPznM97tnMS4q3SKcW+wrip+uilHdO5xu9OSHjV29fjgX
mscIU0MlWdJ5yjG3oNhDeIwSyW/ibuBaQJZEqtihYfI5VGSuGG8/JkyhxdRDFLmFKYFxy5MY5nRq
Wihzo4h+6+JEK5MHgtCQ89iQKVkRHnhbS3o/UBYw/f0js7laHe9uLhCH45M2Eq2sa2qFpM/v+ZZT
O4uMBjgBskH6eqPs/rh3mbmD9aAA4O76v/8AcnEWuxscUA51iCFNkqzxHEIFGXsAQUb1jfO0jsqJ
hPV6BGAItS2VTs3bdWGZ42BtNN/EE7rcDqrDuE0Mv2SPURWOnV+0/9CesGmNvnlEEwynoYNTIgZJ
cWbWkdLkB0+U0Cl/HH3Di/6n9rfanqG4R1fdvqdxt7zvYmZyTRKjeHJzmyW9GCjVMRLYzmLwOqgW
oZE42CS3DoHvOYndqQ3G4GXbBraRzMA4SF4CbdaUcLvm0XzVQs4/1IpW4S0rRivS0j0cLutIwXym
M88JBjWgbHWfWQXPv1CLkK6kv4eizOhMyH5DJ19L4BkObW+GIMd+xHfqT+w2ZnMk+7vuRMeh+pPa
t5n3cOLNeuQwVDaJ1Bb8SbNba9itfkZirNz6LQ+UF77ffmfoYgO1aGvVEHPZxwyBuK5gURe8H6sU
BqPXs37/FtInRZjthI2Y/2GDrm0rmJbla4NnvDdiqgtLQFo19sTI6BSdX4pFQkSJK5wL0vXFoME7
hyA3ZktilPuwi53MA+fsZaJ/zts8ARVt9yF3MeRMpn+Y15sPVX4BuN83Nt2FJI5S9tMPCMeATpXn
UTgxzFAd2dLez7R7HstLyXyFuL7oSDfbMm1yoFDm3ESOgUNtQWPH7xtUIwUtr6Y1EOloyT22HSzO
kuVZlTC9LtxNEEakapllIl5kbSXEp2GB+TM38D+vVtMAhb5qkZ6W5O4LB2k0lVykXYQQBEwxkNOC
sgwdtR0yYH9CwQSOEWzs3XtEgxyi/Mmn0uOlUv0wKIghnpR8EGKYo0FdRsCUEtK2ImokREj/uZX5
v/tII8SYQ0NiIT1UebEMkiseWiEtTUDk9Q3wBA7k4//rWgpmAqivTC322eQecu/oUXkMLaElxWik
RSmZVAqL7zSsLqo3LwCj+3MM1ANlIw1uatHmf5WZ7TFUS+QYYm7QUsgD1eCPM1pK9cnRrvXnDyPB
tO6OWuV2TGaCowRj6HS3HX0W0I/B/zzMbyTmKgbjN9xDUTnfnmoMlNmrSZxNl42ReOCE31lObdhB
YYreVtJA50Ae5cOPL/qmo9b80m+LLUMwHPZ2F48hyViYSX1tnuH5sNUayggyNlmjDmTAbHYim7Kz
0G6f4l0YAEnLLhOZR1W7EUsLSGY6PbKs4E43952j8IuATIKWGobs1zD8iVAXvGOVqJ9JRgDyXP6X
0OfsJVgKKzbcKc062OYAO11mfcZ3VGC5GLPqr/URe3ULynZutaJ3iC1Otui/ycsYlNhLFDkmXTW/
k48e/5HNaHmMjxqHQiEa4rQEtQTK6GnpuNASEvPNEqeFeDSo94z6dw+S9frMVUoJLoQasWzM8cWw
n1qsiPokFD5sFpAIUe2H0GHdPhmgFf65t/Mi9CDp3Q3cAph8yLbubDUkj/iXtwe+rILAdJ6e8wph
kfDAHFPX+bu5CxGb79/UbRLRqniPtmMlKLuQ7IaLd/5RZ1J8FhEsLPYCWAw/fKQ5pjP03+OOVShe
aix9y1g9iCg4TGWE2EbOHF8tQm4yei+8RQtNiwc02fMiv9OqbwrBIwUtAIvRU/devMaEzavsbPwP
3BWhW6zCFw+2UY/PQLGj4sN5jKVlvGkv9V6J9qD1iaeU8plqLrQ3nv+sEHH9tahoeq5N5PgH237x
HiWmTv5e1wVntRparCAZ5KO+uvYTQNuHp47K6/CWgVgA4EQWmiwlPebv4KujduaylU4e0Gv6Lv8C
EHtFgQ2ZSJ+i2y+bu6xPQoKHneRKcE06JTlq5kmxSAp+PGnRF3G4lg8Ku9sRWzv8eaqfudBK6Y6c
3Hy41GLIcixJFXG59jsF1lSQbldeZnnTkmlz0ZDNTB5S7QinFB847hFmTBKWSjCF9B1Io6DsQSAm
5wzi0grYCzanmBnCf+MMys0JHJQjJ/ItnB7lDim0PyPZY4NZU5+6pA/GeOW/r3Qu79Y/P2dBwsGW
hFP/n2uEqt74bLfwKWxUaFxkC4QLBKqdRX/SQno7WAq9OAr/RLmCRMsA6xyEEQSWEcLXgmIb4GSA
ZvDWDmz/WY50Lrg7P0PWH3mLzgL2O3KJ8vVpS/6v9/LZlRTHO1r4y0vpUQlO6MWgkugVm5hTtJyn
B+mq73SvOP3H3DW8aGM81P48rNX6kdu05Q40y0YflsTuTf8RPFGjZ3H7pBF3GlB9B2TOx31N3qtI
iI7JU1gvtTC5Wy+CJ+wqZO9TBmSqcHsRJEmDZRYYd3mtMMZ1NTxzvhmlep3JkBKZ6ClmiURGT6Nu
qhrDYtHrD8iBf4iAyhGhjhCeHJ1cBdWfXmqbU10me1UY5/6gZBXemsgPr7TEIuqEGWvHx8CoHEn8
4+7ra3UzCD5IKKwwxtaxwA640p7ZcMSh2EllQ/t2zsoLp7ilSNbASr0SIqrUc64SG3la/ARIsBmS
x+Je+wUC4njz4F5sqoWvEZWMP8sD+6HQ7guViBD97uPLmqWrf2Zbr4E97g9Z7yCiJs7a95Af90DQ
bp02sNIff1ZR8kGI8xcbj/MzCVWWBwgso37iUTzp5HSviBqq7avxTdVM/BZIR08MvUIPocNvsohP
zMSQS2ijrFa85RouVz7BmXgUuW3UE2Ie1jfLaSSV6kNOu6Q4JdTD5pyKwkfie8xKCme8Qfx9pAOM
c3EsTNQcxyb61AzYy4jFgERJgL67ZWrPMkJ6+KuHCNIlmyFRCMthwtRVEqD6d4ds83vGw0BoIuTs
zLaY17ZwPlUHp9hE16jefmgpbl4hkgmGDzfRezYo24Pju+ufUjLleVUnIwaidZ4zMoJ3/lMKg6ZI
Mw4bkSABNypfX3dBf83OXTQRf2L7imlnuHygCMomFQ70n0wcLNK0iwOZomRYnraTasLugJ7mO41c
u9u2uoSWkG4nWzQq2sAP4HpANUfzQMSdkIICv4WPIpWJltCYDJ9R1G/20ieIpbac9tgdFXtmoRSB
obzX1j4hgA5QLv5KnHz/t9S/1r12QiE5ovQ5wmgpXXnbWETIZ+5JN+Kuayvd12CxuBmkX+ARy0HU
0Fe9fo5M/SLugzpeoDPbO2Txe7US0r4eteGTnzc7M4E1kcS/Fa6Y85gWJHOfxjrbbCpoQbsSpbtY
+SmfsS1WWAkcFdxvCX1Q2n3iijZjyBAoqI15PXYV8hNhy2pZX9Xiwaqrjq7btgPSBq9TKLJPifLR
6ePH23ARMhkR3GLvja+awz7AxCklUaeE6Z4APG7EDmUWiEVEbd4PmjT7on1Z+/westn7NVTx8w+M
2sJy/pmhWmSBuvmzwjD7tqM1UCPQFs7hssdYzzeTp+QdjKaqjQkbhlVSIbNcElt34Qr1FQ8F79RH
sFO7aRna2AEOA0jbG1I7jUC0IPvg68X7cy1wuEfo9QuaiclbfgOAbW0Gqp47PI+XuE5YHWeWEhEU
eG9C7VckdTvPqKzVtbZx2ORlaT5KFPiACUS4z+0tKQDOvgZlspypfE6pHvndR0lylBE3ndjc7Oqe
RpiH3x8IgsTFYp/8prv/DkQC0NtbN03wyWa3TEpzL+2kbcvrbDR2XwssQkR4OIOSzz1Ldwn4Ut2/
cjM8pfB+ZFkBMYuPSL9NCAx6WkHR+yZhTRTgtNNv0AEE0qrXxOsrw+cy7hlAmu/qLipqwu6PZAg5
lAn7nu/XyiIQwVahmGfWrZK8vA/dTLh0jHeqG2hQ/sTSNN2uW69q3r8QUXqeTyqouJ2IMn0QCqX3
ytgRxqC+3MLsCMC++lBq4VPASz6LMj65HAE8FYE7BfgAiVOOVuDqVIrhV2HE1RMyaPLRAkL8Y9V0
yt8VVya756OvolidxNnWS61FTCyt5lICG5y833WWOK/3EmZvjJL5ax6FqbjltvismASq7I2GAoiz
bEoqDMd52G/zUjOf0s0+asdUg2ilkmJQv2o6SFKTxpRSKCHoTyF40uWKa4gvb3YjVN5le/phcjPR
9TnUlyuA2seEMsWgQPXpNQDfruj+30ZO59WgzNt3MWpUOHKZJ4AKxtD6q3CY5ELl9SlQfwbpOjYC
+4ApHBSHg2aoBtdP5h3Juy9XGMQWVgAuGp6DyJCN7nSH/TxPu2O1voLETZdDgsx7ipYCjpTeDGeV
qaTHRaPLt+0S3Iif7VPP3i9EkUBvIsvdHa2lKi3ShIAM3Sp7SqAbgO9RVDG7tOg9waNxkwjH2U16
lwa8ezpdmlHvWe9CEBHOqwVkGtyOX6yEHCLyrOMK/fYvsWdL8IobafDcHiO319GpQ8SPGKd+4GU7
9pVUa0+vbmEhmuDQptOVTG1ZEcy2fdNchBNZaf0UeV1DqWmSQ48ExE/YbsxfwhuXqUca04Usti5V
TNemnBaO9VgjorD4f/kq32mqFWnkotoorp/D0B5xiOdiitBGCt0xczMGw2ffuCU5XX8jC1+41Vs4
5344ZqWTTfGklyVakAcu8oqGla6gEhsKRVcsH1qOUIZSAhDLBYk0ntAYIglDfQdjWY+kwbG7xwM9
B+fKlegX9sF8MmGeFs6um4O6PQm74Y9ekbXCaWrzLshsIhxni4BbJ+l2J7Mkd3a5jwd2/M5+4Oqz
sfUn1p6kAE97RKhkWc7TJKrs9mOSjAgUXnB96Y/+dW9zUiNpKonqQjtGidQEPddPkAK0Z39gMHCG
gT0sLtxpu3pPl3eeQnh65/xjq17MS2SfM1Cxhdm7X3jpvOLsFgkOh+Oz5j7mryilo+/bzxmCVPHJ
8YAEVUFPZ3HevTa337Q3P2RyWUECLtkg25sOvB0/1t/6UNvliid67DpPjynoZptS6T6gKciTRiE3
kF44B18y6Lk5VmUZbaG30VViJBQjdRxYqM/fXkpM71m7UFB9u+XcZAiSrMCTBUHTy30xxfHeXCq7
X7MoSZYy9K/T+3kDuBB4fHfKgHGB2NwhwEkH6bDTew5VEqS0Jn+TyDWmr/ZwbH8Eg7hB6gw/uyDe
IjU7zhn0Oe3az4bP1FWAjN8DHjRwBWY84F2oUR2wcJOjn0q2yodCvzEP38Vanvl1p5m4oLB972rO
OthP3mof/CWE6c7Xiu7Q0k/GDsg+oV11ph25fPgdVn2+cssXfaSSkkdDwSBnWwe5k+snz29oCG5m
oxdABDphqAfsfJPNC0OJQJSqVjAMHV0wiosumlGvXaF+tReWPFTeOuHBs9m0DD7TRm8b+YwN/Mhk
hTXA8CH9MInkqCLqkjD8Ng5tb3586cFwM+MTKTNoHG6n2Y7uprkwI2bYstGpt7AF+V+4X81Vg9tJ
9c5lxlEehw0zZTdX8s7rKTCy7tldWZz3yVDdXl9Dtr5ucksoSF2uDkA9lxzjJQAn7ByWfYS1Wjab
xVNpsHLB9IvAnxqlIhTHe71riEK/qWKHqUscF2LWjYDEf3dLmL+UtufKp30/Cur6tQ36VJMRAI7S
XrIs/6UAPdtajEyjqE4jRnFSPRsW8QWI0BI5XgeUrk9uOymWpa9nDv9QvXs7QT4AiXmc3H5qb1UL
zDWsIqJCNZce1D3F79txDhnxBAL8ktsMwBPOEbkkW8HCKFJKWydvQ1aBMXuPzjdGZ5wmAPwNyOlt
YQXGbUtsosAwT/rzEvQuU4bv/NZCofHqfAF1ndut1UNplxzCPwzEMNeelBIozFys3tNQHqPZKVcm
Vn5Zr80i+mJGsWUFg71IzTi5cjvJPOaLYMVoFNhquBYAKtlf2fKoGJIgf3zY+WzNBkWFK86PhjWz
2+iJlA44UPq/BDOYeHc+NEV0dr19e39EjNs9CW/ucjI1nBoI3EkjNSF4hmhP8BolQ9khdjSTCmw1
aLf1jMsAECkOGnffbgKlra7Mb2Cd5PrilrzoLlaKYFquh7gA0A5GPFqM3nrh4/hb0ierZAlNq7f8
KO3KH47htLmyj+ljOmTQdXHWdqteP4JfzzVYzk58/krpDBm5ym8ZF6yJUt8H4GuK74crcZPKoWLF
jeWpafYngW4xgvMujL/m+dxEzuSAPNqZzcoNXVcQEzTl0rivaBUCIyOrHsGTuz05JLXwoewMHZh4
nRXiraQNcwewF7glsW43L880GX4dAac0pHckWVna0/5nGIs1TMOFbp8mZ9QRsZ64k2K9qM/B3kx2
dXWR8aHxRqUpSgIH1DloYRUfj66Hez88NWsl4D+V2ty0bkXtKdMC/VaCnzFT8MW94FdTdmA2ELEk
qVMVPKdIZBSzjQO4wZbIa+GYvexhjDIxqAqtFeOCXsaE7Wl70lvps1AsXOGEpxRzZoeKB5QVTMXt
YfblsBp1JqvubGRxVV4SjjMPHiRJ/eLbkEP0neZiCK8jG6BAza7aEn9W+4O1JFqN895YCEuhkTca
pPplhOoKFUVARsZkwBFvFjQEKv21yaiABPOrb8QBhyOjWnfdqRWTNo4gQnwUYMN0eWk9PQalaIkj
sB0cF8CDENK/29RYqdVZ5wuH8BoFXu7IioCbLL/RTAtH/W9tfs4F0mfM9crH1dSwhpMGkAALt9KQ
tnGRolrq1M8wawCllh1oFnoxMX5nM1nS2D9eeXBvfKepqInvZqN0iPJSPIP/Y0Yl0tFJAF2FEsFr
MgN0ij0VB5Sf4+NDsa4/bSLeeA0yVrjGjSvVv35iAf4bldybCxlriMazOotrEAClFe1m4Pllc++Q
3H71OT9DwWf6fg/1IkusYaF7rAlhTO3OPzeeVoNabbTlBPMM0YJADDEYVgPl3dU+PVxyyeNowJ6B
COrsXrWLkIWNMa5EfawhC6pWOpf+2mRv1CFQJacmJLs3cZC5Sg+fTekKQ2mcxkeLnRByvcIDmVA9
DGAoHGRTZZJmFHT2NDVTKe+20bwbraGNwGex6P/3C10m6eKkBYR4lSqc8LmlW7L2xhYSjNtSRxHY
DfNkYz0658Ybq3OT+WZix78kbBXBDK/aBMDbtPmwkP2ybjy3fJJs6+C5IcNhsk4/c6O1GgqVdjB4
S2K/e6bq/kTeoJXrPmsnUPp21L2wIPf1vab4mkOviVp8cXlxZRlvV2x2KwuiH9x709YF1vGZ6L0a
fC8BjdMBOdh1eG3nHrYUjObiDUm0azeaRA406pZOwJYbCfbOc61BQpGsj1sfokUuMZPzdZvl0sqs
WhV9RVMrbcNNWcXq1iBc04xo+2KhQiRQO3D0BY3JGwboZ7zd7qrgK6uMugCxXnRjtyUW0IfIAF3e
9cvSucuqzaWYfJpAQqEvKxYGyKKUDP3IG6fWXQKkMPLv1Cm9vi3D9PtlW8Be3eVYHrPhwazYy1VC
LClRmKocr8coX/r9QAmD9iL1Ums2lxN82inw9sNnbkzywXdl53Ipa13QstEjulMUhrN9mw4WAc4u
SEOQ6B/2JpIYPgLvVY82ywW7HhFaXTfurx1b9/YFh7EDtk1WM+7R7f1wDnCvlPLBds66M9HMOYvp
+ubMFKDGuOTXTuve9Q+Hj5hZWzljuO7BwJbdFqAuhj4YXmBt86LvgOGP2BbBbLnhC7ZoItrUJpvv
SEdLXtaQijTg/czmxwqVDeS3bL2ZvgCmDUYgh99q3CmIdgA6B1UnfEUag9m4BuTIXTeegJvsIy66
QYnDrtikWwfzWMVGpGj8x5mSkJPcX+7J63VtZoJsLXJRRNB8xFnyP7RxaFmSkCP+ol+y+Ybo4I4Q
Y3ZnlfinAD571UPs8bwLTM7iFqms9qAnL8lvS/0lMT2govTb3oZNfghtTPlK4/LnxJ6anfkHR0Wz
1WxrDJQtMMcegc3VfYykE2YpxsxPJSze3HAfn+ccEefCeaZtBS6gLj9WYQ+ymhwOYhYq+ag7bx+x
Css5TVfkuZ8ptZwChC7josa7/jXmhnXGGpHIqqsS5nbo1RdnJbIuYLw+LjQyxf2K1E5KHw7FFpgL
kD1bCO0eJA6StS7hGOgoppbOD+cuSqdMt+mJFVkBzV4hfVTA4NUkRd/PWW0xbcm7rPJln1v8av9z
GsCsCShHYF7jJ3gsIO1m5vljcZHg77z0iw9xFTDaqpG+EeKWRyoPgeaCjYeeE4SIqpC+v/7+SyRe
E1qTyIljpCFPPPbSPTHZRcOP6dUTM6tieLjhgo/ga6YVXpCgMtrworvOtdB5MGnu9okuWODk6K+T
It6DT4R0jPyIdP5kW5R9KFhtB3iW1sR/3QFqa9w8dBuSr8DfnvFz8JfQAbM6mrYiUngO+3r8hPTb
EQkv0W87ouH5qj06kK06cnsOSVofymkGYb0j1RSMZ4Pe3oaqd2IQoCk2sQGD3uqJqBs8ItdAFRp7
1G3+tmEPnJIVuwVyYpTY/0TbV4MBf/RF5h4t305IATe++DKXDq5dlLDhMM31QfEIWU/K4cK/zUn8
S3eQJHtHh3cHSV5c49gpuUHMNF7CpXnVRJiXGJVCZMCrs/AgY9ddiu1dXK+7lHQn0bWuM6zUT3HO
rN24ZlSVlNhEUdgWCTIwlEhKVvjQorL6H/zlfIqCQVwTrB8l4HTJa5Pb8Uf6+pmio2L+GoiJC3+c
2ZpHodvb3vPGokjEJbcjy4zfz4eGA4+8iZPBZkRto2XRmHznuALFs5mUFMb5ybuVVLthL3qCTEmq
jWwbfC7BjnDPFurTjY46hqjkFXGbCFu80b2cKlEukqJQNDGou6H5tQPz64cnkimUYmKPf5q7cZfW
GxdYGtDFxG37Kw6M117vBgv/gR1dV4g8J4o0eY++F0q0MP8NoEOVQ5LPFKRdfMJO0z4H0u/SZRt0
95uCLuSaX8ULtw52nXwtGtoDU3s6unPffZc4bEtdvupYvoTcHkROhoPZIO1OFM7H7IrEt2JQ9l7f
LcxWFlgdDPGbkmpNCq0UPRIhWfECyPrBzNKGKBXXA1DW1t9DIuGK7hHk8BPCjVMs9Ez507JTmoQC
wEJV1bcDHFfK/s7mx9F8WuY+4RUhg5qT87BhbZESjACnlC7Jd3kWBFCGaEVQCS+n5mQ28+bZ0B49
DCmrznI4W24FO1HyyBtczuUWU5zWtuG7OE03A2/mSOwM9ovi9Gb5Cb97tQIbfn92lsLQEAbTSp8r
bRfr4/pzEXmt4nuY7xYYB027mp0DPbkFJ/Tf2hQnWFtuXbOMouIdGKFMXxEXCr1dibLs+E4QOrux
8Las1VPuf2uCLRvdelHhTqfq/bq/B6mSGfc31kyYshTRn+CrTshEXjS3lfV0S6B1K6a9Kj6mEOWr
a74fU1nKOC0eg/2hPkEyUqItxpbYHkFxiOangKsPJEI4rb+29EHng0smg+JeKeZzvAZ9+Ak1uiNy
QtB1QLYqBhNIHidAAVvrZYax2mIzrBGzTW26q0mpffeB3ekF+iqViX3VIbO8Ii3J8CHgqQIZh5wF
7NWoNhuZkNQop36bvxqRBonpICqH9SAaNLj/9lkKw2SWXYz4mDkzMWVVb09wSm8rw+XHoceBWTd6
mey0I2E2p0/n6Xdx6ou3aeTjK72xeV/y0cMLcvQDTdAZmKVn1eiw+FNhVAOu2Fy4MG7tq6Y4EtOk
vcCkggZGthhgW4boAQLpXVQkz7Q4K02gVJTvPuFBvacSOPggJ4/H1xVzhm2Dre6IRf5BHhULvgr/
ohzWQtjWQQLAmiCuBeHNbOjQl4AaeHhZ8i/vqnHbiIUc83cKW9ly8DZG9GTqV0Gl+LG3tciqe82I
mT398YyaJ0XNfHemE3Q6QMBnFUq3n+uCRCoDsHN+BjImX2tQS984msohdPAIRR7gRtszCDETCqpz
mOe0laxTzCBWWsIxKlDoaOasyu5Y6FkRibMMkouFYXiArsr793eVoETUZb0YYV6LipY8tglSpGe7
rypfkF+DZ8cxGuGC+AJGfkcPnaIVyvvdftxSGIpI4TBB9kyVHZFzm9gx/DrBVKPP1hTZzfVzcxI6
0RDOqBxY+fUmEFiKuh6ybfJxDuLnbkP+7zSGozV3U5lFzVlYlz8RbUQWTLrmU1sz6MaFofdC6oxM
Y8JdVVeWowZgk4JuNW9CX1UotMOCgbSd64QGj6U24Daz3iT7LWCNf4lV5iDShNM/B/CWsy/o7I6D
9S1H+GcIALm5iwQ1ljL4MtOv9r64GZl4/WL7bJKlDI0OL7Aj6In2hsXLiha8NddoFuKaeGOqkyno
tsr8nzx4W8CZuvTDO/cwzA+yNv2GDD6GJiOJDgtrOV2kYC5LtRz4AfO3uFWtIsyuR4IRFjceYD4W
KPuulrQV/yi+b0LPfxN3TwPIpFNHHP0t4Ddn/CNL5HirQapaE/7ty8MDlLVFuzaXcbRkQBLLCcFq
kdFQX++N+B1T//pwWDAraPX1tHp/c9uB+ItPBEWBxcEGCsgDSUek5RtzFdF/KB5gMkYdJkuZBm6J
aqIkBeu1/oJu00SUC/jEqZotQ21FGTrKgpSO8jUawNwwPJh/+s5bG4rqO56cTZ7fcvml+hzYq0YN
gw4ISPoipqj0AvdXY7FHH3x/Dics9AWQGrYYS+KHU0YINGP1QCg0Yj8KVSLg4vKCV/kdboUgPVW7
0Lz2f4NZrtHan0i0iyeugJnvrZMV7K7XwZhlk/Ks/Pu5hhY1hwKy9ggogtrKvm6sxoO3+ciV15SD
WbFvTZmIq2izfB3BBWpfGum42Ts18WZqjDMEixbvTNUlFj2DPj2hazstaV0nIdlEea9Z/lQTd1Zk
gTgDFCbzbTjj4/AuhWZRV5OZ5WBrzOJpjFFQkgUMr7GJnL4ZsZ6VtMtR/bfc+ao63FHwZ80/akCY
b3AIJFkLHuCDwd0iwFpzRgMRp4IzMs0Ax9l36+l1serGOg0/puDYSzGFQlmNBmxsOexnd/B+XJMy
KYi/Cp2JPO8bT/erDRgE+jU8HGCdXR9Yg07dsSKxDNObdS1n8CCn4NsEFEb1sOcJlThW1IHUmv+J
WRY+XbRpCGaiYcSHFdTwpmysTbzY7VJGJT9LQ251Lpf1gWqES4rBbKf1q9UzZXVEB7JudibPymcs
SPnd4bop7mp7E6u4c1PpmWtD85bblh5Bs69gSikTGOJsSjC6Aws+t8uI9ARy9WBbr8H3eOsfjxGO
o67RoD/ClBtMISMzX++ddxGKHgJD7fUouTXoh0rkUDZ9cLwpgyjYbymRTEK/wCpkbSIwYBoXMdJY
eM3Fb0xzUTIPDi+h/R9P8X1iq66IFRshXyToGmOAt8FVF7XVgj6pHpFWLGqgnOkNiVRpDeX/YZx5
7/iZ3/+iZtys0k1+v1Vr6lQYu0Zp95YDFsNB/1z7X51Lhv1JT06F8zSyMqVK5xjBTvR+gVM5k3EG
VxFNneHcCgydHU/86m6piZPT4uxhkeLuysOnGqvpm7X9ozFdticn1w3bN+Sh8UMFNbHh0/3cP7fa
xTH5vAWbPrHdIx3gSNgqmy3ReoV6t90CjzfDunsPCjtBd0dhhUdqnsuQqwaj6rk/kGp7/oHT7WC7
uZU4j98I7FoOo2TBLsReTmvB5LNkkj2YZkCeYtuWoX6zl7biGLosiXQLDNNdr9gRAq9F7yLJj48m
FHL8Wf5i5atD7QCvpaY8TSoDpvqmoNxVP4fyu59lFZv6p+JyxbIHQjC5OHwURL+I824XsfwnExeT
zau6FAJlL+BsKHp3T7sUhtfMBhv0HUuAHodHprm0kXCNtRnKvCf/EJ+p5SYtLQdEvLLd8VBxQfnU
CzbzDCVLTrqCU6+hop9ER4rqsSEmv+d9oDrfnMyrK+6yJnczsakUBSSBwdSqLd307U52aNK7cuMg
A/DhxnJiYNXI6MQCBBKwaJZQjwKVUXy+Z3dWXS0MiCnZBKfntfbitcjVHnmXhqu5Gdc/f5qO1ezs
cEedWj0uys0pJxucajXSLH1Z02zVbf7QR3ADeOXodjVfxLdCjeiTD/LlOitFLX2D/mKlSkTii6XI
G4cGXSFMthWE5Lk42G3K73PT+z3coyng3BcMoqqQ54aL7m3jLSdq7oMEq+1uKviIUrw+sDeFaKs+
DS9yXVXmQgwBU1ONfusIHg//EyLm0QCUiuJ7+NajwgG31HUfweh6qGCAZmX2l57XpTx//lKEsXQ9
u54MuO+z1OnEu5kp+SwAyUrq/dZ+wbgvjtozJaVdkkQac1I+vLWRksJoYYS5AeKUxIlDJctY4bbS
OOTCdhr7roRx8CgOo26cjvcB4RifGUvKr+aKUkE2JuF7AOZHcvHpY3z2+LDYZs0gPcTF4kunEwhh
53gLhL0Oo7F4uO30ws8q6b0hYqvwNwRdQPZ7spsw7fugYAZdJiZSPnRkvz2CG2dF91Z8FaTKbvuO
02j+mODRiegh4bqc0owReFjV/mW8nqk0KYJD/qzSVQBHX86pDQtbM915a43OJ5xQnX7BJ810pzCe
rTs9p9+PFu/rwMvE27EXNGFnT/cctUvC+nG1y0BjnyiczqueBoUUiWe/vs+DI6CYGWw+rNyqjDAt
XtkwcXia1WaW/dBVnCUWR1FQCjn5D1cJsspsRqqqnEJqvV3JaPEJWQCLwMqneqSyPaUFX/OhBP2h
86JjbzttRPPYVmMllMNP0dE3uo1TVFbZIzEFsalZMQ3lYO1UdTupKr26QG+qCC7p2XwNkEdPn8vl
NhEUATcIkd6tonBIB69k+JQRecy7mh36sz9JBUbv5WDneNqNYi+nNFlwPP74gqRkqQNI2zW2s5e2
YNweQQ8RzAcs6Lz1KP6XfPwL2DUd88rJBmpBUa1qsqUiFFeiJUEZK7IZmK60wLe01DNVO0Y1vWbN
9Iy3s0MRSoy1LXSKCQQLeB83EyyPlshCcrCIfscNQsGcNpSiNtdsiuJhoO4a9KqjqkFjt5N8Ps98
E31qmISPCk5iMzAkhdt00tASZ1UpkuY72VSHTmg4nBS3CfIVariyWUF5lY3CSZ3tWfPuOTEEq/Hd
Y+mQyHVADaqRswbCX6GkVFaf7+WgZI99Yoe5E9sI2US+gXJctfxURVwAdD/PJEZxhMIXXxsDX3cu
JBXTntGHkONWWzHQY6vE1miiiPAZkNhqy3BedNA4qD02G/1v/yWzKSTm0rOh1FPjJIxSh+GcpGte
hiVANu6uRKZlJRJyPxYEvy/QIq1q7z5eJb+KCr0SgDDKu5oZuLP1vdSVIMydGeWahPb8dMqAk1h4
eMHKqbZOPkwgaWEDC4n2AyyFkUutUOi3dLK6phT1SOCtQYRONA6d+0zlyd62dcJ32KpI8o7kaxbL
Y0jnpYQJS7MnNFmAkXYVoLSe8qWnwIIgSwJLlhuXnY/ryXI/9uEnCYEo1d6aZd7jokOZtrCZbGjY
FlQXA44XeT5LGnVGvoreYqq4WeI7KHgjsOnVjoKegKLQJe/4eq6UWWVfuZXQFe6Q7NGfCP5RGFgr
hfqkRyIBXK6WTaMcKbDwHul8esJxKFan6KXb5D5oAZGuqgepyxHyL0Xsf6WN07/B5cwhCVxhTjDd
cb/kvkm/7iX+6kqEYf3OLPqHmX9dyvh75w0lhPDq7ArbyhIlwZT6VYx8nmo9JjsXZA88qR7JIIoV
U+8tDj263KEIy+FGdLHgvUJ2pUKfPUCaEnbMZdTcN8Lrj+fRqvrFiM4/NQN0An8w7wuzsksVLaXZ
dXg1z5ilj7Ad9QaR5VJArLsPwHYp7FPM586HYq71E4jCwDfaaVqGmAPWE4BH51QLlaCwUmAXdJfR
WIcC5FR5n6zrG15aA3hrd2JGA1jT3pnqZG9uRYdHZMc48ZiyuBnthVCQGqmdCPoNQa67q9NQ+6yV
XBo/KAQKmyCvXxLl2eTSrVLvN3NOhlGi+Fe67Y82dcDTCG8ikkdavutg4JDzRg9WmcJ7aguJlGHJ
+X2WV0YL97l2KSvG9SnUKu1S5hdbts7+FjxoHoHSE1GUHa/AMlP/Q80jT5mAxp+8ruiCHqRA0Zke
2J6KOhzg12vs9rUIpWPS1+/qVhQEHkewt2upEJkukwmHbb7zvThdoLNXEvLDNwc19pQXpBpBXSzE
3jU7VXH0zqoORGgYQE1lMhbK80riszuo5nbUMvJpp7m929L4NHXOk50ARcoZxwCIOcZN4GPO4QEO
UPvqrQYJRJzOc9QfeTka6qmkIFNFTwWYMRIwN0Yc1VY4wGPD5s5v97uiMO2tZjzk505J3a/1FvAM
O7ZyoVez6eeWZWRxzaMFa/XomGDHEwrwbOGkBcJQAYZtZz0eDjgFIoQFP/9GZRhTFngw5/VciXht
YazgXOGYEA9NuaP8DTpWGTyB6GdB1Fb1qcwGxwFsqzvtvhe+9AjShrqQLy2H/XyS4s3EIbP4aaME
YUL6SJG2+kns/sAvShwy5DypTKq1KJpT39CtVSdUAs3Sk9CC7qUcyMe2YGb/aMMog8WtbY/Wuq8P
YbAbBgvpUn075oa/fBIJIQub0/K1nj/TUQFrI6UojGKvO6O99nJjN6Y5dp67N8uXaJGMGdNcXHrD
BXSp2ZpjQ89CPU72QH4cUDthQmBBA4XgD60+bj7P1utl9J0Z0gTD4TexuloC0gq8bFSFlq8tx3S8
jbKWB1NWaL2UpY3FwLT+v11xj+ekpU1IFGfiNNtRH0nfM4zhZuXnpht/5TzbmBLryGLpUY5R75H3
zO65xOk85UhWME79JAFgQk9pl+MiMavY0ak0xEjOOnDxYsnduRnIdp7dzYVl52gjQqO3DJb0bBgO
RMUvl50AuK8VUKeLOm9QwVY+6VqLsdKRJV+ZH+RYXIFtBDPJb1Vr3tCHmUmg7IEL0WZgqJIajkG5
1yHEDkS8d1mOncLG8QP4TJ8caJ9Fr5PjjiYHeP7Y90LiGcZiqqNSHv2zYa8McG+195hcDUK94jaI
PlaqG/nMVGL2aVok1HPSjA+8zQkAMJeFtyhQxJmZD1xyrlqocTdXowIMcOm7QNDdqNjpLFdsKbYR
Zc5SLd808/dPvQzOugdBaEtfVpVuDlvc0z5sEj/2sc76osrejxREZIPQ5dALjXQtJ6z/J7/ucqeg
O+jUDRdIxcEyv5c1euFicQZ+rKYM9WmOfXca2v7eNR1/4C4VOqkst1HyDxYkSoIgCV9NUS3dbf74
2AbRCDQsEuOq7JtfbW1bWwqSFYXRQos8WCBD30/jn3YenTNHK85qCBI/wu2bUnfjkUmRiQtvimzm
AehlMkWu28dbHn56HaueOgBkgFuQxJjw0m3tTqawjiMBYpyPZS8Q6JEsB8XvgVyB1KVXnbkh5C1V
R0QmEfeUJbDoqRA0qcX2ABmaC/TshORR8hG6eDi02ovFq/QF+hj9P4k9gj2Z2CZ/GPeTpiXrZFYg
s5zoO99c6i0GgrvNua7IFJeNUCnV5n89A7aDIV5qw6zz017csSwQm1Hq2DegawbKxCuy2HrZf+/y
cvKuhE/yPgRHyvTMolgs99i+ri5ZxbngmJVN0/Wze60Cwlk+0GbeQeCnEm5gPuip9otw9eHZu+CG
IZwTRucwSbeDxZD7IYBMneQxpvQfcPaeTasLfil5WQ9Pd8MDQMGhg+zMGWl1H8UzXvA26oeXFXgb
RemdNTJrvi7BSgBHSqTvFa2TpOfYzy2qmkTH4mi6xiy9HkPu5XIcquJ+F0Mzh8+z3diqku6skRXW
cDJsMD1G1VoqP0R1LJPOovQuqfQG8cF6Ju6khdnmhAnhx9xJ1mGvO3aeL9Pkezj+W+Gk7XYE7y2y
FPWZw95iDEhH9gVmsgte2DjPfaHZ0dPhcbIlnqwoFDGwykGKzAgFamUFQQWFFdJmk9MFNTC+3crn
ap1e4r6cYk7Ha46aW0ExZpwgvMIlEn5Vb3r/ORhdtGmq/St+MDVJVjwbS4mKgnn3qZsLcExGDWne
zkoZUcZvza2zyuZ4TE0FIsdSLuyDqcOotWB1RFuWY4mIRonLJbCHB6GIdrTM0Nh0M28A9Wi3wRvO
sgBcpBY8uF4kOqy9ERTqISAtMGfhBRR1j9xDqJeWrXCsSlPeK9FyHbJE9fsLmQPGzqUpCTsyZAdP
IaJuXbudLh7ysmCrco6sVgzE3LY22aRriPddAxp3WjROVW6ckcC5gm2B/HOXhL8hDgpL7F5Q85fr
yCpyBXtNc4DzJPXnltgAhf+zcS54TYBWPnx4SD9Evq8du8iod7Cjp84U1SfdBDUCwFv5wOALZdxJ
nZ7uISaO+1PR8FzK/aYs0wDPB6QYGjz7ALS0cTuohA1FkpH45ReY97aeMwb2/sGIqWXNMpVauRLB
udr4OQsxN5AYUAVolUVyL9QHTl0LcnSSJjahjus1Ufk3mRMtZAPKL+zhVAFeRX4QFy2Dx6G/P6Ql
m/T2pfDfLnnzUMW7FZWhwog/Typj6sG5wYKR3KSRRN1EiUwFUhw7AG8afqTlIG2LL7c5ZSjkzpSy
PstYeCTf20qJ4Dhmt1RBCC3ql7Gi0rF+/1mJNDgEBRzNWKmJhyqvYNr8BWc8JgxMU7EZxdkAa7+Q
a+GBA5WGPLPebXrFWhT/e5NqZ1Ijt9GgI057L4g67rVDQbIxOVo5F4DvAWsex431txMOb1ojqtlw
xS1nxzWS0bWvsFJ/sJlBzFBxi1hirnFlKXR00oRjkhywPOPVzfwcw9f4x4Uum1GKOEdCUAhJQPus
EGVYSdOoE/tdwSua1aFT+LtK8R4D2QYSmxDbAa+218Yt8P6yJtFffFbt0+8jw1ea/JHjZ+JK07fY
YzoAnGl41VsQetreLK4UXQZqP3cUA/tiBr16KjrnuaQ+fv/vxfVNnH40ENXWkOWaQIjLtz56JMJ8
dAm6x+aGULXKGvdvrAtu03Jochl52GWiUeBKbBcgvaFLv+Peo2EwNANPEE1q48og9CgLjiTPcTdh
ysYz1pCg+buoLoRiSFnpf5sptBr4gMbvXJhmxFBhEn93jpU9CvSxzlDKxm8HECQ0eAcixBh7VYCX
VDq/4A+xFZSIas7YUV2A3DgS87CGvVS1vBt3nbcIKCheDfEa6Tq0ipla6RSkDAKd8OSXU3N220zU
UHYghK0sq9wPBxVJshewE/zGoAhKDqS01LaSKEVwbakCstrhRhCvYHdRKbpdqiepI2FVXRH1Kjv5
KlaJiu8BecWq/k7B6iFezFoh6PTkxXc7k8D5UgQi0OtSwa++KlfzR1yxe0PaJj2bctv9UdqSTwTQ
8om0EELzmGcxkzfZdlA+DpkwZ2uAJvzN9mULRhSaBgogn9ryj+oUycO2sCaA2UwUgZtYUwRXepAU
OCOh3SBBgIxZ+l1+x3/h4hZT8UiyX/UCvhXlWjykRQjnK/ppuNPID0Fmu+3FDtfJac1CP1V3mIRx
z8OG3mTN5rw67rXaduns5JxBjZ1XAjR/C3CwtBrqkbT5U0EYAwx7FCy/31Ll8Z3Eg11C1+zXwpIU
ubwMbvhuqYhAPscWoXb3z5ZQjgD0h0KbudojZ36x06tQUKtWgX99P7DPlIQaKnVng4Smle+7BC2X
p7X7h5I6c9xmOY1eDhyHbb4p2hissaz8wUHjpQ8opI25sTozX0tEcSNgRzz1oMsHTFjC7EYbIuj3
pOS4ZGOYPhQjec0usQUyjM73B0BI4/NZo7ulqxl1mnAZghDLpMrD4kquyKkRvJr4wL9AmZj9Q6h8
yrRpJtZlMKLdmUYjXwPKmdCqMNS+/guJOP7hfssUk1pYVM6bye6F7WZTtuQ5nvIefhf0VR9K9d8+
+eOjME08yK6jW7UaOCxTxrVa2jp97bWrcj+YgqXSC+2dgRAqOH2C+g01jw7zQTUzsJCE6kU9grXt
1rWHYofVXMALvF7i1+uzUM3pO2KZRBgEEbNSRwaooGJTCszcfGMeeZsXD58TqCa9bS3kml3lWCYk
NLcBAQxoOwgmnPh1y+J8TkJrEYESRltz2KsncjzzDxdGVzBOj49eOrlfR/2fsvThlHR8Zdw+gYxn
zjskiKUjFuBKwTmCjvR73aOmmY1jluNbrqboI1lIJb4x52lY/PvW1Dg64f5W2l9a+SFc5RQnFj8C
6nRwB0PCpI5TmgDcqJpK8LSeynucDZMYlwSU3Z4t1pBoZs4DcFYpgB2KJnWyGrCx1bHSltc/f8pa
DF8ERIo50rzNzpzX5pxIJTbwltDWIL4dOV9EhqPUrkUxnRL3C2DJWQuag7X6KIOqDXY+5sdxXFlQ
4WinO6cU4gPLpYo5vR/UZ44oo0zTNG8IOjRi9deRDEYEOnO6o/8EgaOlbw1j237RYsizc1AXwF/i
gD7P/GWhr9m6Ltx+6BHNeWTKjJcldfbvnOrETUCv2LZAY86ZobTBc9040c77mhwJu9eRFDQZ1ga3
Gc1yx+Cb1a56GZh1gFDxtg9TT1XbyO2LoXEL7nq1knX3xCKAtGSz7BlojmPjedjYkosHmhY1psKI
s/C6X+5lmhrpOQYzJKDojyU95Vg8dnMDgCzNtcaQdXgJ395jbVcij3OgKQb0ygTOO42rWh+7TF8Z
OtdtIXdyqUWVi91ZGcu5wqv5iWvzZzjjuoqb8RDElAhq/KGOArQNaIY2vTWMG8Hy3BkzXO51SGCo
x1iFKRlGHXEBYDONRY82Qkquly4oTFdyUwqBWIJ5PQuHV20z5d4hjARKH4/9cfojuhYVJdZDP7N3
cFpdNgi2I5q/euXEjE3cC4kqM9OXO/NsBPMPYmn4GsvC4wHMAX94BuozaKM5pjqds8xQzDTBWoLE
BoSTC28jXhXnZ5/VuLfnCOO310yl+pqNFK0SBPdL5x8jCN3VBN0iGrRMTRnVKRYQ/I+BUH1H3vFN
VzwyYuEO8zNVxWVExF3h18TA5U4vzEPRGLdOiwFgNGmijV5DZk3bSGsuJ0eP/149T44+pSYTVhnF
32n4+2PMVH77tB/nXj/LQ++DtjJjpiqN5dO25kmm2a0DFwQA393EfLcZl+/hYVT9vqxJnwilBivT
TO/r48JhxM0m1vRKr7xkzzUzrJ92J+Flax5acVl4J2BIfvsKNGWJsmI4iMvTNrJqj86IcGOFncyj
vlRV2R4c86XjvhtjB5ZL8EzRbar6tmsDnBys8d/arlnUsim01VQZ2KNsjA0SuvU2fVMZuWq11Fhg
2x0mhHF3W/SQBg/edNrt83t5ChMlMDfQPDxCgVmC6gF+5DNSWnVi+rw+OzLsj2UWsTybO9J5YdZi
M6jbwKGaCsvMwldfNvT1Pr/nRJTeZnQa9JH0lpKWRFirRzNDu8S0+WI6RZ7DYscaV9Icvzpwx0BR
OefmbtCZLjJ3nIWxVq31mbFqVwm3cNna2CLQ1o0DzUDD3yQnt4aj/Y35QOi91q5Mk13tAPgkpC6b
o3E1kdjFqZORxxMMfVDsPgf+u+ZjLbJFGPqUX+UkGosQa4J6hD7W5f5jMuDTbbn2hapF+HcUdjKd
H3iRynm2PFgB2dwq/d3JrHS1Gtw89tulPc3fYof1bIwrykxbBtnamqSRf+7gNagDXaoskyBBTf0/
9vfc3ow4jsmR05MulzjGUrjAerVv+RkCgykhFo+jQa1F3ydg4JlzoYIZJmz9WgFC3dwBhdlY8iVo
Odi9wzymurYaFEMVC1/Fc15i5b4ydmCAdOWF3a1zGwnGZdfpNaSZcCHB29Jn+XwZ0rSD+SdZLDJ5
n/emrZE66e6NUfg4WZDF8KqgREE/19KdscndoPss5XIdi+Lx2O4z1yS0bf69QaA4ZomV/9GQJJkt
/1epAQbv3lTLFr6CluEW6rNBKX8ml9lXOvcC7PnUurPhMvKfWhc34plTERO0BHo0in2yYzo2+CzP
JNzaJWbR5nILOMvjpZjXzRMIa3shFFQhA7nrnzQ+BSonNGtuA9BYHyg6jC5hXmaz8Ofj9c34BHnv
VPnNEKyCv85iJEG7qVYa2YtonJM5K8wq9ZM+2nzxbL1BjiboZBpi+nElEygd3lOVctF4r5Indpxh
31B0z/TCaYNejDOvNQ+aLIkbQkm+MwbKc89txPUoHvMqoMAzI0I2qadYxIZjll83Hc78TR1VnoQh
ABdCsiyDqfjXF8lLjyb1c2PJiZr6A11ilWQUyY7gwRqc5Xo6P0C5D1d+6ZkC5Srd3gMJ+SoHaTPN
dmK6MbLD1OOhBIooHEBy3P/PiyqXClwekUieqh1N3RFidPyopXTz9V2piNyiA+FcZR7Tkt9vRGr0
DSkaM4Quh1oYvZwJvPDe44BYZfMDTrajoqkCV7cy46xme0Zs8KzBInODuLO6gdGaiE7nHhtg6K93
tbOh4iAKcsMUvbqxIOqLsMmYJDRlKLZmXwPel8nX09aGwq5S2tehr1wUy0a5HhxnamI3PMo/Z5uM
bY18fY02rsgQYuclJPQdyfVgTCbPNY8qEHZqhtfVtxhunO6a1b2vhq9ro9igGq/OeVwC4Dc57fjq
l2Pbvw0Sgi7soHLrlkaCH3SVB2E5lQ58wFbziqWVh+08xL3o+FvUxM1H9wMhd4uJlXP15tFT2L+X
VUMopG6MLu7MyBav85bLcS6Nlhk3Opb9lQPl5WIqfUv0xBS37ecqhYByKvbnwfmKsWJ1tGK4V5tn
bMgtCeikL1cB5cB58CmCJQ3Jq2AorQdiUzq9H2HJoNBk/fdOWyWIyxqkp0z0zRNf9UFQcp4R7YdK
aBB/a7bv61vW+FyGXhbqtydNndiTPwEb+nmK8ojpN4/oudS4AzRfZgPQ1jchiPt+HpMJRjF9+SOB
ZNphwr8X7qFzh1l0EDvhXBVnttDLp08YfYIXZrZW9GI+76oeQTDVUldyDY23hEJFqBUeD18VGodl
IoiSYuTVmNG2GTMBcg+a84KWxiV8VsKg4BLlgR+6wV8ehohTegNd3laYO2XlSZk05cybQEW5vBNe
rBXt4Ir4Pvq8gfrUlTgNz4qmEMCYWliWAazSvtuB+Ob2LMcZ4V6NRu4lIAdoEEhIoEpUqYZC8yW0
2IF7CHctul8QTXqK9Aj6NrkqsvoBgsUhHk6J0C4SP3vbBq4Fcv7fthEUnzFMFCjoF0hlD8iMMp7B
E/KLNi1Y7uELdlE/WO4SQDF/V800LdSQZLISRphTFnu0r6mOFP1aZrNIHdqgLHLTOWROYcMKuwpB
SvxVwtkvfxq/mSrg6XnwDpOALZE96gAm7uvmTWsR/Zs02X0ZleRgrCw8ut8g7ka2sQHDuFgxq8hQ
vgpU22+k+hZb+hKy56Psqmt5IVDvZCstQbcEhZhSK3YNRr4XRuSbyg6ukZhVhPdUGLTodS04PecQ
PYpRy7yFqNdmWVQ42X3YML9gqu2hfISXw8sFK/zqucS6JfGov1ZwzewSN4y84+cyj27cTPHNCK9e
rn/YfNng2Oot4JjmZ1pIdO41ad+ss3dU3ucz1ZkTVrctFYO78jMHpYsE1jo77+2FHvywgDdp3gnq
ZEkBpJsAL+MqzkI845gMBJXRShB/wDBhGZ9hrSgP+rueKJdRJxypdFrGEwx1Q/pbeXQJZeT4IbKt
qRVXCZSVddUmf2jOK5UECPArJjEjCmJST3YIZnrj71S1g5bxsbe6510yFQz/okAck3wnC3iCkgzX
nf1TVnf83oQ4xy9ULtAb978msHgJyf78b4hEozIVxYytiZYZl0wsqRzzMzAK3gUZTEZt5f6v6MF9
Pp49pyANRlGFR1TcohjmjiOemDhOb1nAEgRBj5j+CsJqH6tz2Qz6JXECkYYhNntxBzIj77Syxb01
ZsrBtr/Xeh3r1bud/A2U8HEGeOBR0iRl2o3fCbW9MD9IRdeZq6xJGjw8YUsdi+mkS+KjPPDmyCdi
O0qdVUsEonETnIra9f4Rvgc+f6EzlBK+c5wPGOP9LOEtGcIqKitZxGA21k9gRwINmBNd8AhohehF
1yyHC16DnYnc9QdSnAqo8cQ2d595IJ8sfra32yUsskZaxpLIrx57EuEnovr+yR1yPORBxLmxOP4c
yRVCFACJctWosn6W8RZqilt+OqCh9ob42HzuQsEaKXAlrNrYpSa2btTtIV40SoiBud6qLk6Dwj2I
8uyRBlcC+3a6OBZR8jDW8rJQI/Qp8I028kFiZG2NfTjkSbiPeFUHa3pW2G7WE7eUtPxlSOmBMqNX
PsrwXdxdkwuK6m5Gr08DCjXwvZ3pm00olwCOWyg7PH3n/nxQmLGN4T1nqx/BGJCsXG8rQEncACdf
x8IWcBOdgVH21FsGGOT7xeqj1tW8pfKWfr/jQLTJ4+9oSLTLyONfJEL9TaHfMHAOW7GsMqQOQ0YX
d0/aYK6BL9Bi88+WPam6hF1QqDlBH3ILAxNSdP1d4b3kO1b/Q/ZUAtTANxSxOs9bvf3mbEoioQrO
rv+igIjuacFAEcZJwaHBzxCtndmFmPpgTueZTG62x5nKdHyWEL3CCB+AMjINQd1bVYGynZyEIU1O
diDdc7TgeZ3q8piE4pQDusp75JK4Ee/tpAHCB2yXR5Ni2G7JNDRXoleFcQeD5OClOspPmwAXh+7S
ZsakkcXddJnuus9v9W5drNAU3/N9sps9vmYXfqStBzTR9giJT9ZIobHFAGIUjQqWZgH5+HnLlEU0
XQuTqmE3HfH5GsjshypS4hPVhmPGEpVKcuTqNfO1cxrM3PhFqyw35XhgFRz4Z5867MncgQAk1gDX
NAHmRKkZcERdevKf4XM76MvOB/V8Wr8qZUrkwnUesylMdxFgqWQXlL5lo/+jY52t4ayv4sy7jari
tZWbqJcXaw0JviiZ2WP7EAaxF/oWJjmhOIh8yfwI4nkN0KeZ6y7g01kiaKkYPUFURKq9TQYjLxuR
nIaFfdqWzPzfCd2TT5hEZW3d0C3QE+0yV0Nn595OsUIubqrCU4S5v4E3FfXzDmf0lTgVgeIlL53z
cwVn0+okHHVuKhb7fHocLMi/Hqj2H+uo8bAQe7rntiHng6ewPcp9PmOgTxEhb7fyXWLDKPWbERxA
Bd59b/uZ6iWVVm1pFKsAfuzyaiToxuLNzEqV7tPX5FGVWFElctUTlhTSqRrGk4MkpiXq1uMnsZ39
k5B6eHzosLSZm4JR5k4sPFIS62DuVXDL8eYt5DCm40OngSpkrUNB7Lt9yfCQNtrbOhhP3Q8MnHZt
Vq5+GgRZnR2IraFNA1+D3FZC9yG86jOOhTmKpKcJJ4MzViKLAqO5j+flr1jyfVQYkQobS+dcv60j
rRlUjyBKW6ISrNi7HnLnU/75MtiCKSADVEeUK4zlNgoW4tRXvNxQNou2QMVDfvnGHfn/3YVAB3kQ
j5//drp7zafHDX8yqhO4cccWv4Ce8RiQ/i1Lahj6masOo1fJb5qusAmseAojygZyHcLISGTiP3gz
zogdqLw0z8kqy3VetsNOHoNf99LjfKYH/nzJEOZ7DBfE2JsKTV8oHdmn2dCmoVTeHf9oJQJbKceL
TvXikk51xUkD/6dN3TYv9sTu8bDxFnPnUP+l2NJusy6Ezrwej+IyVSTU5HCNFwHjYHreoSJjM19S
qDzAr1AASc6jGy1fiozIv1Ms+gtIgoLCLJyJ0AyDo9G9UnEHUy+Xty8GVJz4MppAfNJlP92d2QSb
469sUhZ6ee1w3HbHyCbRoD2uMFP4wZYI/wt8of4M5EVGqjRuiklKsQTNdq3NKZJyFjo5qjp0oVUD
nnFZu9BwWSbXZt00SdJXW2PJb6P46kHkVyBtcRlqXkCl3v66Vsd140EwdUNPLmf8ey7VQbCgcOCh
YdjdiG2HMi0oTjedzh9H+OTt54V/RV4ox/s4RqBzbPy0y3SWqwzFD89MAs2aIBhC/RbnGYwSDRbU
vGvy02nBYOsNp1xv1OqewanFqVPT3x9xI5CzAXrpgAA2AGm8U17shCfPxYYHQCfZOVhN1RFvTfY2
isBuMFEnVHPAqalxeqOnf/ErTz7pvP5QfYHgKBzdJjVZk6sbPF5YGBWw1QH8o5xqQCnb9Fk6fLpt
9ehwL4wKNY4PtoiQeUW9sYs8mqdphht2MsuC7ZT6GdURcj9vji3fvEwEwV/dHF0jBx8qfuvItxc6
XLvzJWekN3SCdSKjfH5vHy5Epq9ab6ApcG0sB/5BQwOGsaR0zcsWapNGj7t7fdra/mVeZeuc5qeX
qfpSJqg18YLBWTUYrNNw57N9KcOCDEGuj5EAL404Kd/OH2nuebU8oICJHSOXf5+a7hWplKn0sllg
T+uE58QNsfaOz135lEgaOrzkcTHlnUfo01mCwe48vZBIr3SLeBEXDiXFF+hWNgePY78Laoo6Q2Kd
uEBx3pRTTjAL9ufNP4z0QF+nVQXnTaPYd7RdBQLn4GVAoFhD8738zP4Uzw8P+ddCTMJBGAz1ha0Z
Wo6OJQXkAxw5lzmulO8e053Hy7Zl+/8ENVdhyXi82pyxEgpUrSgKf4cVSeuSBRS34SrTCD5PBV+j
nXkUkqSVDCRwIQGmlKqi8/r6IoyIlMikgQiqO1r6fFsFqjR5O5qlKXYq6h6I3X590xvPsLvu2C+2
uLf9oWmUcv7K14vk5qqSAet0a6120QdBeAyh0IBns+eIauUOHYL1M9McaNMpMzV5mBpTox5BjeV1
pvBkD8+tEMFHBqlk2AevsLKbBK6TBoJgBxvZc1RJ6j4A4wcsqqbQlC6YS3RJ+CUQqLczDpCmFvKb
SxVEVHS1HwFlGUtgWZsma0oVFOO11NZLyuPidpuidwGAZZM8PxY4lofzQHYp/qtE8npQErsJ+9FC
U8KD8Ii+litvWpImsikuOqS0VYlaj76ycqoy6sKW88gPSYg6OM4Z4Kno1/AcGnSpF3+Mounnj/Bb
Bl/04pq6SjLDiC6BK18M2Ehk/vNOysYcIJPrJxLtEj/KCn8BgIalKbKlxV05g5gcUzD9BIpJThW/
Od6ZIGkR7GuFhA0S5RIrMsiNw+CM/xu2lTUKQMuMQ67tijnL/3IyTYAp6B6/N3Jg/ygZxZUSdVVC
Npjt344jIDbJgnZMIlqZyqGzwuUsJ4cSnTgCYzlbg2w2sTecDi6S0HoQnUHvoclyqfKkQV1PflfB
3F1ie8AesYDx5sApOQj2IlEekwMzmH6eVEUjhrDReIy8X0jNQP+LUlf/Xj/zLDAznxkPjaUteyE3
mTTeVMzC2+mNLAPXdKZYZiqOM/uBgIsw/v7ls3kUhuoewWTJyqwmzWqKRFD9Cuir6ljYt2MO45ly
8W+3vZzoVeSAhhWH96yeuDOy+5Pz5XRpVZQZ95xb+gP/7njfo9hcKuS6YaXXbfAEOCrSfcQofJjp
E10imxX0zl4EO05kUmh46fL9vP/KSAAw8ORh43esVKSfmvQHu1nAQCHtS/U/K3YVxs9YwaNVSpT6
5bwykSJBdmj6agIJTNk4OQ5iNWLbiabvPsOTWvsO4UvJ5WyDnUW2Dzqci6avkKlxVmnoRut0rO/9
AdKtypfMmyg3ZK0fNlgfxlPESLS29wMpfqawGXY9skrCOIwRTNPFmdJvGLS5RL1J5ZOBcZ/ILIO3
bOEKu0JnoPYJvWzhLR8OyrTw1sXeiQt6H3YxDLwoZdta02xROWRr4eITkyoK21RQRgi9l4STcOlm
59PpQwAHtRf7nO9cNsIdXY7LB8uwQx1oVVXEk+2RGO8imPCPHndClV0Swu2tlEcLkQ1pBHNo6Lte
k4fJ61BIwvT4s4B1Aim5Mr4fScCvWkAUc+r5XrwksE0HgmrPAmJYjSD4R64ymS/bWAkd+asCxbIw
+syEQnZMTYOgY2SVxR89x1sD6lMrfm3Dx6Nfu6mp8tc2Nub/EhC6xCX3rr0ty/F7nt7JK042xgSU
FYepACNHFoUqvYWslLmi0XrOHkHcER0hHNndCyt7pUCJC2Sc0jwanmYaeuDHMsoalez6x4bbh+B+
yxMpkff2A5CDBIg3Nuefxkk3gzXA97XDumjuYlb3+7B5o2DkeMgFVYtfExDyAvznZodRCMxXKpkM
6mDHIep32FvBNKgy6k/MNrM93M9dIakrAV03mxyIW86Tsq4pIfltBV+n7fBMqGT/OFN8Fl1/Tcoo
b/VlvXMPr+efK1yUcULaX0JszP3fnnSdyL9hgOthJH8yHkFG0g+VIHQqMQz9caaJZtRB2G92OLOZ
H1cZybGOjB9Sl3qVCzUYjlvBMnqVIYee2DqgjbxaMVBd+MX9oooRmBB/TJBo9MLiKjxZg5djRhN+
T5Evs3MDKESKd8UTQwRQlWK39Y71uTt+9I5IKdj32BcWMurVxhiP9exWLtDo8iFawqW5RRpmZVh3
tUH5NAOwe/d8/WlPGWEim0jt3CPKYjwezcsDOb502bf/Z8QhrOkRblaE3o9p6OvQKg7GZBNQIU+5
N4bUPIehdf3G71xD6Te9jsD+bp939JjEojJfaG0uaDPtIHv+q6MyhZzcL7mIWUlh0FmSn8i9mFuF
8bEKZ7EY43OQKl4ClVMMNkFS4Wg4233VCX2McpsOg4PHd7V7jk1NIT+Q7YhK+9WaJJb4QG8VzCj5
d6fe6A3OfN3EGlNR7TRSjAXeQ/4jb+6CDk0z3EOP/VVo4rEFifF5cIbUoEk9+ONj9gdjY0okwawM
jIIwQ/wS8Db7lHPGou322yiFBTPJ1Q4FqW2xuoVuGQEWFBGpVX4ErZc7JR3eQj0bet/nb452GP6f
B4Shf+Abg4fpOdHViwRWcWKTOkxJiJ2KqPZgaH5jC+aCje1k+yH+nirHs35jCO9zgplF5xs0QdkU
hpfX2hqGmiVplx645rIwyfXvMNdnVKkx6+dYzfKf3SL9vAhYMz0L44rxaW2wOGRwbN6ANOUQT3Vz
9rm0XhK9mkTFmJ+JuNzenNuMKMep+Dk1jESxZjO3VFSfVn5in+7Rci+mNMsioCN/aI12wkaqgxjj
wBttxOdsicDut68XsKhzlinQnEjZVRtmPxdDB6/KwGy2nnVxPPAFrZmSwYf9+wKx7BIcWf++HoZO
bEF71ubav/C6NJ9pv60E4G0Xv2sIUNnHKc39XWQear6EHwwNnRABpSRfWXNzQz+QEFpWz+utFdnv
QRjVfvLau5pOOH9Zf15r3RM5Xi3oGbO5COSWPsqsQ4Dl8EXKtY02Sv6Ld9OdDWdDPq+viCgf/TTJ
+zic6vH3VNF0R/swPMRj3Nk2LeeaL21vvrZsxpwR/EjHFnPUfpHO6RE0UsHbH70SjJh8MTT8tbgH
Pya+FIDBbRDmVRQpHKInH2LYhi6KaQwDzhEihiXN3K4QuOfc5Dyf7PFZodNOO14teF7gcg83XuIV
cW5nuT5jkdfLdTSS3tFFlCMH747XiCiGE4b6yjcfQpWyb9lIk1RMWDTNFjBHAQv9uGIG1+eM6qk8
57/efx1TZaQS+D5A8WvUFSqiKFEr5eSdVfG055fIYHYaz++uJqkSLXQN8TxTAr0RfLgEBE2YXt5P
CzxaUH4x9ojSVHcoiXfA+yrnENsdH00/mJJDmB3NzWVLEJf35QIAf4TPIdSlZnYLY7Kg25VCXAvj
WvdyRjMC8hMotFNHHwnHE+A/ufRJJ9fc/XZXfRWt0XJr6aUMf5upA/ERNEy4uUM9M7iEenSXFh00
SeUmZFhVhsNcrSaYUy2xr9Db0guCrUn9WNbTlB2but6p8N42lZqdM/8jWwXyKjiNwohcCWLUhFic
Tdnk17p0rTaS6B5FvBH3v3UVhkyXEXzPi8UCyM00JI1ZobQapFrFOE0wbQ5+30NrAD/pC+EenBvU
Raf+QxtK7JI+C8ur2x2R4VJfK/GftBqQo1VDYsugmDDY5cBrOZ83g6lRpvk8Pnn19KMDPg3dfZnG
IFniKzWDMV6iDZs0g5TfBekNX0I8+M6t090LRKmfeJlhjqRBp5wqzLXSyLe3hALDdqEZd5k5U9JA
/zwFj2AThAF+7RDZNsH0vPWy2A1rX09Euv6FdoFioIpHJ7kvhX/LTxVEDF/DCFt+OrYHjcO1rEXQ
KWZJW8FdJRsgxfezZmbSy8ZaEB+b/WXPSKcbXn16g9bVtoQSZYCxLGin1TKdNkpWbTDLa/EQZUpS
eL/6EMpuiMNMUwVCehEY+4Bu3zd3kb1My4azV3Bc3QwHMIAwSih+QbIbX3ZfLbRaiszxY4g2gowO
gD1estUXS88QY1Yhr61LK+qhWyyy/S/XBD/ekyReXZgXWG82tmsZWbWlm4F+l5milO5/z+LZ67MJ
VpRIGq/Bp3rVgkhwYYebwkvDJyrecjL2FaTzMUq0t5lwEw6Q7zTZhr0dLkAaBEv9oSHuNHS4HMgM
zBZnHEummSODGEzXzDrLOZaZbknUQPdHSdfuUT+NScpzN5xbTTlSUnLBM2weENDnQPQjf71K3FL4
5+W6xmye93wwWybevL0Ifn8ImHv7cGOcuTXgPU/fZs6Zm9MSNVmJDKX1gVfPABQpOmPotKdarX2O
GM5MP7SFl9y1fAUsW53HU3gbro7uyF/5k03igoGK+cL5qhKlW7NROJIUoxQUOslf62xKj+wKEj5h
TMsBwsFx8F+rCXorKAIHIuGZF2kPpgrwzP74yWLCzTcFznR3PHLlIz7OblAqgos/L1/WOlPMe9TI
8X3zQkDP39dozfXXVmUqRhAwj3ON8VDJp+D5lfMo65R7kN9g6PyFMcAFp64SqCI3uMnXwouWHiZn
11rAW/JYb8b7u9aMsT7X9G8xgUgDQ8x5B/9PB3pYK2KFgFcO+M9F5I0K5ZZLc3V4ERV+bo39JbUb
cHUV9Pxj9779IXSbjaS7Epc6U7pwDw89CYSoNPNvL1zwDBFc0weNQE4dhZhp0J8Xu5wTJaZJV3JL
NQ0gFq6N4hMFm7zQWmOYXlCh3Ki00SeTjQM5gyYxi0IZmAJ7EiNPGm3YJr4hsW6yPYucFdea4DYC
nr3Tu9TKiqvR7QNODLHS3bd3/XRfV8+V1n0nqbnvIkyghT5lYJUUhfu4CKU9oS7AzIepb48ektMO
Y8snCM4alLqcAV9xVY2tFXvBBOw47MdYxYI/wwnjJCbWTwNhltIiTXFeANp1xAqGUliY2WCayCqy
w7zDoouTX5ebR7OaWQFhAKRgDGz9AvQPBdzmGuK7gNdL7qCw6NYG7P+z5I8y8wdRSQ3cQpQAe2gz
INcN9WFXNYT6U5wbWaM4ymVeaSntfS+WyZBoEgGxRSK/Of/aPvqwLSVzvGmfd5ZLRIths6CSDOQP
2F4fbe/3B+iBBh8oGQINNyDeEL/4X2O96dwJb2UPXRQRDP9CvYWg6oCaiUUnTAnBJp0iMsMgj73M
3Hz8sooFEHuiCLkJHw77paZy3RWtFfhwswt6gKI1lfnpTH29F7mVhaK6reB2FETjSYpbxIqSrXAa
lon6sykGYQxVnPlkfP91m327r8GLR8I7f8Fvggebv6CdMYoknEOlj+XTEwHE90dmczi7BgNagEOj
lWsV2SrYBKgr8ZdOoFEcEkiPe+aSh5I5yMuFdzR88sgGh4QApIVCVd/er2SArYLPB69l/jeDaEu3
7Xx000aPdkbWE5AJXSq0w/OzvPNBQWz41ja/x8gPDIlB2THGtsenGTH8lCk9+Htt7wpAEANsl6aR
wOQSssA0k5KWpTquKuNPGgFRr+zoB0N1mCQgvsNhIDB2M/Yo5H1np4BkvdldtKCnanGMtTYdOJFb
dTgy+ekzlu/ljeNlTeOCApqX9351SNhdadtkFYBY519YKY0KnIjF2mAO/VXj1q9oUeXbpqUUSi5V
UwYItVU+md/VjJUVnz0Bp2pLdc6xVIsR5fFp7qPhkVM7lZDvcP3DCNtnwaeB1Hg06LZ/cQInvLEr
HXxQAlsWsaAwQGd3oEQ/7kMcoujDiV4hg30UiMp1aaiJVv0NzmzlXC9pI0RNbOSMjLlBW+YNZCnB
c46dQX6oBkPgV2AqTV7oEprLfQPCKz/duVqxOWlhKE9Ou1ZBwoWt1b0Ahe90lmijx6MA2hHh+adr
GJzZLrvgpuftBPxaZ9bJJFBmriidrWHLparlpP+d3gVhBrnqCvKIHz+38xn3Rb7UGr2NgIPSGwxg
wK7O9KkjwtJysNwuI0kKf2n8ne3Pt8ID6jj8kNHqC3O00e1Gqd+7gSz/2HII++gy+etE91p40XmD
Zds3nWh6M3E45O8kn7Wp7ctKFUMS8rkjMbRKJJ+tpdVKKdvT6nhwK4ZfLw+FSxuVNhrTVHHZa+1n
4G/4wOjHXZhotA2i5gz8HTku42z5VVRJLig1FdxjiUc82FxYZWBdw7f8qJboqxYla2qWR+bQ7+0E
AHyxY+/qxiBkGd1Sot0LzvdiwXncV7GtsJWL6zWxZcdg66NiaWQ16i9MwGeDmnmfC/oZP/qIvJT4
l8i9OluWFxbYl2oSZspU319GCm+b2uJbELtisn7rFrmMHIAlw2jnb+ygrQmov9d8MQ92sAb8siND
75SPuRg2lS6OLXtBoIJrtd0DzrRYGt4FbPYxHkNdDLbwbxzteWHpsCKiGe0WpykfRJgxUGeB29P8
4Qx1OvZxdQW1joGiI8EoqM2YM7BWqNtJLZpEIGTdBPpP+vvPPqu/Pc0JPvB0dH0cB2FF5TMRGpML
gbQj7fDsaSAOPpWLPpUDSEk1pt53mMLd0HiCivnmxOpy1Vk1PR8x6Af0mnHzroP/Sffu+nooQLDT
E1JQh4bJ5LwfWRMTuhD2snB9oENcnuyEyhEwlee+C58fFb/g6zenSHe/kg4XBMVIMrvrhuzi3hv4
UA1xGo/oBD3xjkDUO37NAT+xbzkcrXlZVUogEFc+f8yZ+cSJR+n7hW4nq+kP/3b+l/WpOJxH3Lx8
1dRK6Bg4yfKgk2T8FuGJS0PIN60azuXOx81yFtYmiWueAZr8rvEbAmi58WROrRx8N3NF2oZ0Gr3g
IWq3hSnwYIS3m+gTsdqbnYJcfhuPzOUYSf+eThe9UsPS9o/QUWoDMB9b/YyU19qHyKGFBPpV9JXQ
e8wOvDGYL8eYtSdrnaQf/9kYMmGi2xhScudTq+XxcbZCbqIFfue194/e/TOxGU3Q0fW344x7Oxa9
ArXF6vpZniAIRuppUgZN/urdRLO7PILnZbetdndtKOqpWu/y0KaGdcmd5N71yCSnv/KG8f4hENCZ
dqffpj6rnSVTq8JqdWDPTgLgU2FKU9YFvtLVqHaKMNLdF3IYAeVcFno2Le1m0FBuvVA0R6BFBSS4
78e3xUromqZZRVSFQGZuRkkgYjpvYrW68RFS43WX6s1rLTZ7PpJL9O312WRHsAomHznViOobAgKb
MN7wnTLCxlYzEDCaqstu/5C5+LAfMXfOdKOuzqQ6gyN5bNm6Lzne6ao97eHQlLbSpCSj3oj35Nog
9KAohjNCaFEgq8r8/z9iVmi82bgX7kntlIKRt0+a3DclKe4nL9tKwvTJxSrQCUs11gmwOE7BUQQC
M66OOD4DwK2Xem/NlLFAPKj8FQuZYc4SgTJeR/27mB/aRRp6bbUPxgEyKCQjTpNZykS7jyJuUh6z
xlylfsPX6GUDRsKp8nul24x95C/qnmVnm2jBa4GRPuC5GyjVrtlrmxptHbpmibMrzUYODrBC9jD7
rt++xcmxFZR8L5szEWxF0myVlwfEDyUZHl4vnY8kPoys+Z+GFG0s/3tXNbURgNQe4xIUXjSZGe2Y
2g/XM4IvqFs0NvY38HuTmTqvFJvBepZ3nM9g1BW729Ngbm94HiOUE8ktMD9aILrrrwwAUdKMg7bz
RZ0lAeF1hx7odP+dle4Ca0rbV0DcyUPNMeM+9hplINZaIS/T4eB081m6mHQWgJq9ZpyFOJ4YUOjo
NAq+KFXlRHCwjWcQu9uTQuVGGcXzinvuibL/VPgMxUTK32+5v06+14u2wC6ExNnZjA+iNdHZs2Cd
FVV2lTWaQiUMb9E3B9hXoPkUWph/x30LohP3XNyZD5wYfz58HUSnuUw93bUP7MLfWKWJcDAyFg2/
Yckw6eC6/m+FeVanGBZZv93NdQ4dnblmsClBRj9aoGp3Lo06fFkAu9HMgwkbDKPYEdKkcZcA7d/Z
nxkSWg+oUZcjWfmC64bXKJ6kksMlmD/jAyKxcxKipk+Ar2xxmXc+0ZVnoUGmyldZz70lAWqw/185
3ohMByK8TscwoE2AS/98s0El1QfdFXR/gT2vJYJ55KD9D+glhxugB+5TdBFPZ+IbABRPvSvHH5vr
wml5Ae7LhLkSdAaDHfis9wVJwB9RP7mSJSRE43/nawUVs9D4Xz04I09/6SWEpWbqDoP3SVzVdbvJ
2KlDeZlCZ5J+Zq0g71TBu5fW7/2It4f7esupvO4yLxTttgO3heqShbUzpS7+AlVFJzkXg8otVftj
SH8ZuagrXVq3EUq0+2OFVNcQ7zWvex6PWW13xGvxuUi6/7zMLDipr3UoRGvMYh2UGIvnrtXwSM29
ODkUW7zDAWjqwmgTtXtMUtXDdQ6wdmUNR1nIW0eiQDkbP70ucEEyP4e0oZFc5nFkYtwA3EJ8aSCz
dlzhHa4227OcJvc5+vxiL2zBUVhvXVtqJn/OgNPt2LWMlQ8j0S5xgwZ5u29uqcVYw6JOYDwcspwu
3SAJoBZfqDElzeF1aUUO7c19VZmCHLouTK+pB0kjNJG2WHEcZxz9RinRtlOfnVkT0BX4rXLqlguF
2Veo7OeysuOvP32usBFIMuV4noP+b4rEjx9KBaj6cwb+d8rCAnTl+7SXSyknY1tJpYnF/+aRj2lH
I8FJnntCXhu/eJvHgZjIzlTL0lVfFF+3N0VOCnxaYPJB6D+3iCN/BS+vpcsJf+Qt7nfyt6sqiPLN
wxoWk/0klIvWsNdghHpcUi5FTCM2dOyKpJhwouTXdOIoe5VwECmCZamSv056oASK/WDa0v9WTjri
kwnE0xHGofrRUGH6yPmBmef+hoIcCvbXW9X74DEWPPh9GiZ0c7oVfTnON3xJKw6tsgbfUphxdQBY
D+JnRhQH0UQaTSY19gWw6aM9ojm4ZCIi3FYJ5jvOIc2K/60ZcvRiuTu7TFK1DhtiQ2J5F4hJaIi4
ztz5YOMZtudPND1Sc++bBmw0HPEOHZ3z9lawt15RPTlduHBzdxJ+mSZtUrVaILKRqyFR2ja7WpOy
0jO9BpseAgYAu7U/dL7FLOnR9h5l7LVTjh2jB3vmHeRIUBJGRq+z+C15Edm69G4oNumX9pW4M5rY
s+S16UVXcEJ7TcKYNxdrGfihMwLn3esKJiKfxG5v8Bl0j/4+yNjwSIF5054BBJN5yDOlkLnRUmTG
EHKHcvzXv8AwWynp6+LoUXEvj2U/5TnukSjinUq2025jr6c1R8UnODI+7Uk2cWPDZhL/rELnAgny
GjGObVh/q3/IZ+kVwpgyUTxkWGGWJYtu89n6IyWXlZ/+x4WuO3XG2wEUvj3nR2zsg+v8hAbvUM1J
/frJoF1emSZLNqsTBiFHF+5ctcZ5bgneOHiRaxyMf/J9tzZrhAy0xk59KMpH7cSO6uwNyHVOh9qC
FaV7i2H3J++KP6vPOYH0eXGUD31gDkYnwqz9SqUWU2DlcPSNNZXsOZuAwx3qJFYxWm8CElDdZoDn
HDf7ensHC4c9VY9ZcTsuFAsSPUB4RHfA6FsSxi9RBFt6k6w2R+oSM4YSJGHwHHhBmlhVM5SJ+dVC
chvd9BdUG8XJU03yNzgGs3bZw1E3rhopMrHkL53rSSvmU1+DfhBMVWHvcy62LG9d9taSY5OBcKme
ub2hGhHad5QoGubfaUEhVPnUOyX7rowuDVJ7lyAGYxu1mieZDYTXQeZNbVO8Fc+vTuhyf7zttCxQ
+Jygis7ifMBmAqLFPRNq+Lk7DMxlY93pIpRrKe3EOCaPR73EEaT7Hj8m/BBb+y8zUtKyQbwo7bDO
VNj5K/TAHSRWvqnEkUT6iUCAc/ratcuPZcvHEtPOXU8+9jWjiV4YPhiq0TPPPMyCDrr0AGwjkX69
eSCcBqCL7Ed2nI07uG+fdYL6P2w/wVtj+VSOgN/K5TuvfmxMBwpw2jrSVyEz2bE4izxS0RU3QDhz
tZ9iAcqEFdLvVwP7ftYleHWHyhblfkkQZgCdTXzFWqdtxrlODj3xuZ8ljn0qZF9/Cqq7Q0ed4Sss
IHvTVN/iORFzOsOzL3Z24PKUhlwswbTv4rJCkNAV2YZhICmrL5OtNQ4A3Mk3YgOO2u25dNRj7xDf
pzS+VT+rOvPXIARJ9QxghjC+1fFrzuF10lENnsiJhERMcWUNTeXLa6SLG9Tdz91nsRS3ZnbDrBPq
qG1R3F2onxSuJhYwZSp2Fa+tJXikVONZE8s1czyYI5a/iTdq1xG5LnKqkoPEKsUTKLSnsDATaA9W
F3DEienwMO7xmzRwx8EXZoRyRk1pudGF3GS9Jcfrp7YD02eC3F9UGjGJQuKbPovY1FHmSE/cNPLV
SL4fq3Rp10OoA1YTO7Hda+QGwqeiBGSjL3h/Qh/0ErMbLO9rGw73FUrAEPCm6sFjHAE6hknNus2m
974ine9oDTT5jaekc8bgaaqvEVIppU6XZLff02fTMmq7CRxuBlEry65u2uXHLToZs8XYlV4xJnzk
yhABk9/62x/DNAWLcgm9I3sC0vvM+9XpEcqLmL+jCk0sFhUnAJqHEpVJJWJq+zrg8GwkEEXnoj9r
uHMiRRtLZoAwJxdg9bEjVtqmgXAwwEmM2Ods9QgM7mlmO5nG6ULnTgInpa1vHCDtIRYy4c/66mj1
t4FaQsca9ovW4PsLIQeYPFgzmkBIb8lfwGZEaZut8RjzKnz/Rr5E/YkMErprsS2gGVj7UJ8XRcSt
0MQfPRJ2Y4KY4VFdUEcLDTyT4mXEwIeYP/1rGoS6ZTZXsbhPUbJ9OuwirUuJgeaq9Fz5PZBk9GmT
99EDZ/YesezeLWIisbvjtZuM3NKs5JOTFSrM4P1Ccz4U7KaQXbDYVfKNg1A2BTGytSZ92wGusv3e
L2fw9NinzhZh+vnAUvHW6dCTT5X6SJEDO8GF2lDzuYxdes1p1n/OOTcJExUvn3HGKfGh/i9yqLBr
VJOkM/zEgIel4EoMlegblIVZKULFKabGMvZ/bG0909iCAyjbQ8f578zYpwhHS2AWB2YiY7z5sSrb
7EDblphdZtn2jB9dSNnfsbtTZtg/Lp2lb66isnF7F5X/aNXvE0eMuizFnuqv2xihd7tcR9Urim+r
aUwbxJv9HqlVGb9B7Fz63eVLZKVKXHvnJa8wTJ/6udDeHECptskCTjbDDoz4lDpwF4DoSXbbowNY
aPadJ+C9QoucgI0U8Q9jSqDfXYjcN1oSIKF6ZTLcgigbgX2K9JRuQ4NT1bsuNyF03iX0Oeh6uXEJ
/9qTl9zTA0xKNZvia7qhXSpEBcBWDhI43W14QVflvlZiFZzA/AJRV0hnIPXTsv8JCBXq5e/Hz5Ws
mBe3IvjqrGNk9o4o2JZOvqt4tXgJ9gT50PJkU5X7ReJW7irwtct4r+Dan9yBl1df21vC5MGxIPz6
ac8Z/ixbSOQtVoiA9hVv3B5dlQmxoQ70NnuCjNgb+80W1jONggL3dyqgdPgcWUfIaR4guZx8pjqe
YKzwJwsbrEZ/lUjiLdWjdPMqd19TBtr1X/6bD3gMDl1UnspyX7eKUQTVghOKpKlMb6QsJdK6jQ7G
LQ6Pg6DRiIt0nxCNEgseuY1pARv2xQGC11Wx4Go6uB2dn+AfviuzZpctR0+gfVi53Qah+eNKpBiT
pmap/AWNdtnnnsb2VPr+Oak3XOi0nWMCABJkgh2ENiELroy2ZGABUNIDC95qNc4ZGKFfQw+O3WrZ
snED7xFCkFO9PIoVDk2f/F3IACtSHctCwlbB13eHNXyzP6XY6lMf92AxnuRuNMPeMFGFDEC4NFY8
lbKB6QBl2CrByoL/LXP76CzbDHcQUivgVn1SWi9CIYFLk0m92bMtVSgqE8ZnivifNokgOkZcnYPC
JNFlqL++KM4ufuWWvTl53sGpUvGdLIHLI6Mo3klLGf9mfjqysLSjgO9diSRLb+XtM1SBWAe49A0H
FDs6tDd9CJeIbKftELjK3sM1IwHr3WgfIQiun/NFjihzrMsrU7kXrdYdlVvFXB7OhIX25UmA5M/s
+G2l2GTu9BQVaX1d78ShZDN9TM1emHlX8OUyAnwlSIoo5gN/U8qaFUKeO4dT+3wI5TyonQ6CWCO0
jEDF7Juv1hKdi45c57Up1Ai0XVUGssfUH7yCduYhNCLjyPlrQvwc6cX1XrFa5j9tQAXezEXMqyKe
B52uDzgGVUSSH2B55diS52QXlPQtb0zej2NOAdi0jwSELqllMiXAxI85FxnQLeztA+AbsstD/FkU
At6kB3bwCETDF0eEommBYty19d5AGyAGSbv72ygudhiQMK5sxjkdRkW5ua1UsK3RCoWDXIXEXHfZ
kWCs0FBOIPSMvF6OTr11Mut+PJfAoKqbF2vCQzbj2f67AnMyZ27GYc7cpbAOvXEjGz+xYiWLRQIC
H09RNYGJ0SF3Ent7J5AUfUnq+Tf3D3vCOoqJ1NCiXrRJbWAPsVKTg/5to4EJlXT2Ox0ke2HKmALO
ZNjKPeUjM4hUvUTh+YGH//CfCdQgH91gYoCrCcpMm3+ysm+y3Soj5SPvq4Lkm4TgaKXjXV3ChNNg
+m51LGs6MINxns67IPPIbedlzS6l4jfL+cWRPvUmUwOgNsZYUc4mVGUzuCBPDLwUd9WA3ntO8QS3
LxTmlgvWsy26DU9HaRtypYHURuLFCbk/lJsd7BH7gQy/Ll2XNQ/FInIp/mJ57RPpYCQ86HW/vRsk
uxjqYlCnFiQvY7Jk7KC4Pb/mEeAyHApdVEL7CAmLFCMQWMsH76OUq8dlJSbLMivz7DYQRgGCs397
pld+yrI0HQ49uxT+WKhsvO70T1GLCGIXeP0+cxsZuNodzF1Ix3K44wIDtLFmX23/M5I36yGGJ2C7
REJS3IINNjokX3dFYTO9ohUU7b9dydiTrUWPu/0D/bLsLcybPUYYk4gLbAElP2LQ65IWcbReK55O
ksrx9WPLy9TDZpXCQCKjFI8ZifurwqClO9y3yqjsHo8OWerI4lcZ2+s+Xcp9c8a1DDYJk9k9K28D
UZ2KL6WwVwG6JOtvaGq2+sDNuEhvlZ8J1u8ZRHerhsCTakC9aYIexxZy/blzhdbnnWE3SimKo2Gp
6qSGwy9dorDHqUwq7fwuBDoRcN0U301EQrVzyRARv82R+D3RIaN2BMOgzL9XIReDbGEf70UNSb82
64BKI6gh28FRjViTZ3R0FrzmY9qO1WXxSdBvalnzufF1m9GUPn6J81ScLeuJNKPPQHhwPmax6TRV
vSfZSiJ0AR2DCsd9mlVTgVYAhDDW5bRNsp475XZVP1wonnBlD3e77Y5tdC2JRQAlbKMxZ+4we6w6
OGTdGPh5hr7OLgCeb7pvgtd0sx1vUcxNf+icZaDBcgwxRKNAAPVP/PtIc5zWm70KcGav+FxrNqru
xEuzX9DKt6r1/mGCGczEGrA9+ZYuYXjFtV7i/Fj/G77w7ZSsSm/QS9jk4hZeqn4Z7A4NgjxHui8h
ktFRuPSQWJhKDgy07DhW05F6k4OepHzTiaAwNSiHyvXttUFOgXLQmbX5XteHRKktEAayYO7BlTyw
zA9VsvyMAv6+zKMWdr9H3FWw5h1McojeVbPJaSKsYrWHxGyUZtZ4yxLbz3Eznc+JaEffelQcGf7n
s2wofpxjoiJJgTpGmWVcg37L/rntufo221Mhe9nm5sFJgQ48XuFfTNw8ZQydWV5+6NpCk1QFNTMv
PE7nMreGbAtCGzNW9RimMyujKOVu9PPZg+VfGTtF2pvFXgVWAflRRyrmBPiblA/j/gKHOItevU8l
r8n8UNoCr41fsW6Nm6MGG6ascuDM2ycO5+jBEwGAVUO7+dcPSc2rw82QriZibQvMv1LRrWAlRjH5
xonSySFe8CS9TzFDbI3/MKaNiZF0JsAGX6Bz9SvykPsfulxkfbjmS7Kqb5HTQ10B8STieYwJnfZz
VnqU/sAXIGEX8aYTFr+j0G4YXyYfcq63UczYtHg1x3GG6ivKCm+xRvDFEe/HnQNtv31iuo0cMCrO
T2UFghBR8RQYksgINoR86WbRD6c4hEqoaPc0sGQcgtPp+IAi4JBRhhYbS/9z+Ve9WKGfQW2snxYC
0sxDvr63bjOfe9/Z5MWBmz4pe0ArmGviK/K6Jgu12/pM/qxJDhthWcKHG5o/o95w4oP6dbQh1qp1
9fZhf/6qwhVdh70eh/m8agFjtsrROOC1sxPeM3Q6mhB/JVkxi/nD5+WJwQp2tyQK+F69TUukxCyi
4oyKb8//v3VVlb34TPfG/o8Zn1mtRiF7fEbBK1o2ebOVF954qBh4h6e6YmA1iH5bBqcvlflZjIyT
v0B19HHw0bSHgky5I82XccPtotqUtZrruYRlhK5TIITdSIoBCXsP79EePjFAR3fmE88ToOQXDR9f
cav9eqGfxppg319WKuvJtYbQBRJ5mZO0Tcbfkz4cywL+O+8WYdx28LIQ/+grcg4cWx5J9OFHMzpX
6sAjEmd0QcpW8HuaMyjOAywC6m5gOBTayaMp6b3y0m6M7aZ7+1Bm6gpDniv8jhPQVQAE7O3F/h/F
C6DwImqD96JlrDchuomtbfyHGn4j3yYVEhnFH1neLaEboogs9fl7vY51o8mr2I0VFqQsYULseA3+
o6gD1kFVjwe2+pzne3N9AurcYAD2xH8CFj4cu6PcO++mqgXhpbTpbqTjRQLtYNsT02G8+X+WV8mt
kKJ0XrKSpuW5bOlcShoV/DehdNACyDJNazL7kDENJBYF9IJfmhP0OT6WblUP2k4WXfLh43Cm5Xn6
EuD5v902+iZwzFPh7mIs9ic3NUr4m7uS/D06nqAgzPr/azoKNvY15nXFcdxYjCHPWpF4lwmR16xe
X9XyJIuABmVZdZZw4GwlMTd3VA5p/bkx0rm+6lX7hKutb32pmwFP3ZyQ2IWjJ/R6572ynerdlaiy
PBmSZEi8Z84gMSPGOSI2xxescXLfvd3zug4UdoL4/TwA9Ir6eRvSb2I2voKW4/FnXtWnHDXeMGTt
/XSBR5+ZTbU29Rp2xQzAW7N696H8Q5YCkr+ftGVddb0U+JFhSAcrFG5UShTEvdnRZRAmJR8EKZeB
VNCdUuR/UEOiY6R9w3qj1Jme4vkwMtzxGvSNRl66+mcE4RJToKxB4WIjyzKGJY5+OOqc4MiFZ87l
CghOq6Cg1h/+xNFLjSmKTsxc3VwNKBEj503/MCmq2YUsAKwiL/LDUp08pr32+dMNwm3NbnuH3jEg
snwWZPjuuguBhpBLRVZGrnkoe7VDXeRbM6GO+AXc+OGbABz8SzLWaxkZKz1YwSXpkbEmm8ZdhACc
7ekpbRQNUSh1jGOJtfPz37yrWYwxwmtnIVy0szZA3SJ2pfZ9EH0WKiXsfS73ML9Q5wJeGdWyzVq7
QwdZjOCRS+EBnUPAd6JTsYQ+1NhAwf4ay05BWFa7lgViH7PJlvbExGOOT9/9XIkd987zn6JfssuP
ghW42ydbz7zAQ3USEZnhzyEwZLrKSH2STg6jumABRnuJJSQdbowR0pSenydWx8xpJSRMaZ3jzyLc
SgyX4POG+wa1aCiMe7ITLGG+0aCvBQ1iM6GwW5Rtui4DAYIR05dguG6zZwt+K68E6elHhvK9LE4g
0/W2slWW3fXT85lxYFwS3awtePguYAUGNMJ69xDyiNQjakrnIInP2tcTnwaIRU6U+gkgs19KNANN
mBQDScjDMug4iJUcU+qopUyHYXurysx2WOm9Zs8LJ56njcalD3aicFzDHWL0GDrjOd6f1PJjnfra
mUuFPcV7pcwN+AbQp2hHHkKcAIifgQQDs7d/hgWyM06Q/8EynhhppoJgtdQ3+yuU+8ZOnfSHCYAF
5TOMwil7f5P3HRqnP9JEvjT6ArPef3P42K1pXIBVEu+dXWs2Hr7eILThSVTrm39o+uG+5SeXJtZr
jYlZkSurxo3IIKTVSE4Q2BQZUId8U/vUT1o7PFAJ+JcO90w/jpS0kBIFPFzbXif1R75mKCn+Qeny
ez+h9WHN3Yy/Ug2SoOnZOgaRK9QkpZnT2vaBg7cy+xt6Ox78txYbF/gYqKaBX49+rYTywkP2j97X
vXlWiy5ssdqx8ezisNDvoromZ2liAocCaEuYxOqWBFM9QlhM1cBEn3vjJUKw4Je0WH+Ct8G/JZas
o5MBiiiSg0FutT9cFMQWCFRY5YLpacKi4F8fKvBplt3hbH0aVvZe3F5KlRYiwGXIb03CHS6uG+3W
Nis6urJjcq2cGf5kMGa052hrie6PAyUYOqjg5eB5IHKrr+44tZ9xbtejH2QTd91emshEXf7aTbX9
zwIPXs8PymbCys2JrHwaM5zGClaWEWRfPP1rq2wGMRNXWCc/Z0CuYNBRx4SUn6wmNr8wRlqoUKt1
O4wuWSZX4IjjOosJKt1ZMx0YtHRAuaec7WcLdDB+8JSnSF8uc7sacoUCnh4Xk/qcoS5b2+UDuC8Y
6gT6sszYLaLMCbnBbUKyqPDnsWugMlOdqaGmfOOst2f/eVAvgL2YMhmSxatp9tQeWZ0O/j87u57I
nusfj2R65RRTnFM978OEanDJKSBMQ6TWNWzKeOiR4+dSvC8IisHoGiBcThjlssKpBgEuy8/B/qGo
LXhpXHq7lRrYYW6T8tVPvMmrl4u8/gGzE8RDku5KCI8c8b6w/8lX3J8TTdcJ29p81djPbwZd81NK
EckdeU3GE3jKNbHoLHXKKgXU+coY7NpwzzshxTK2KB4e01qlJNOusQKr0u8nP6CBAogoNRYhSvS3
DRtkHD6ByklxkK4lfCAkmeCD+VXh5TL0woefx3LYyzSjiaCPmaFckEXQWitIvG63vSQWNr+iAy8v
r/gmeZ7aW60W51HBKCb80DkFSe+3YmYVjND1SdlG/BqD7koJW/rMBC36IA0sFKxGgCnwGS7aAOLU
hVZkVaGBgMltLAXXXnf20HmXRlv93ukr5jJwcefhY8wcwpPbpRfBa9OEK1nUDIVQDnmHB8js8455
2ViJ0siG2dSN6bwErlfnUX33zja1bm8aKOcdVpzkdTsxfQK3woOOfRuLnn4IXYt34IWTmYlSwgYD
dzvwmUtNSjupknlBB1tdMldsXgU+BHmSHQAN9iL6vaPGfzntMj9TURGXLImsGfWZUwLU5pxgJLA2
kLQemBd1NcwNBesUqiTGBignC2UgwKCTmU9a/+lP6hZsodwi9b06jZdyqx6YWyuC7k/WMde5wlgZ
48hJZ5QbicJtJ+C4f8ZNCHil2upMw8LyOdAiYEorQcj7dQW1RVNzY7SGuP6Ad7Jeb/zS99rdl0kr
OTDKvE3rBGI3W776topH6G/7sDjgFy2lAhA7ophx715uaTx17c9o+qK2r6HnAPAlkeOpW9lx0WXy
OCSyMWI+l1podm4UeygeobrftCAwVncs/8UrjcsW11gaVdC7JY2FKc90K5xCXS55QKyOZKlNQZVw
DS+ajr3OUAkbD8LN8qX5NqAbKSyi5R+nKpgxXmxVIPjet9+us4t04kHkEkmupZUiUnWcb5uFyFzG
LZNxHLinBn5+1CQaGVoS65Z0lBDjE3Wppfo1SKCtHraWSNbvcUiGRKqoKY2wrbR9qiM/Lf2N7iGa
XNWKzYccC0peRW3noVazHYPKZwZIT29SM2FPAC0ZBVYA5mEtAfNqRdpDwxFSlkULJXVHWKGp+09r
5FtZyEqyuqAVAN0R/qvRKCYhnAs2nFf1c2bnGwJ438AUlnFGaKjiMosCokY+4b2AbYEEuYpNwFW5
RniEi3sFoXRXxWjpYkWCEqPwW1rAOYSJBLWAbXMlZBxwVn9QtwKgvw1BSb9K8pvoTeigJeJBxuYZ
QLGoscVc59Re+w5zq6pV0vdXQSDSgWIxaQpOf2MDfqDo0cfdho4Sn15TohPn2rgaOR65S9mKqCuF
c/uvh7P7QHPWtVaGc88iWUFM1MlIXK++1bDnXEGuxPoVIbLCbcPYSkLNPzuimRhrPUEZhZFLouEg
odEDRio7r5/PL7eEP4Mj89SVQd0yLgl67Bl4zsfi8srxfmFTIn0ScSf6qdsIN0P/s5FqrJlUhFDY
i3l1bJUEK0BeAQ+2ZRDkDmddwDkRXp2nDVYIEJofKBXELgkaWUS2q7cF/HEzUe+T/38EOZvxVA6C
v6H65tWzMzuiEEDhdUNoCnZCID/BefVYhMeE9C+y5PpLJXb5HijfpAnHINnvihwSk+I+x87xgOZ0
G2pFudw5tXmXQJtHOfzMaOkrTHMJpWG/nOVEdgMEeliFL+Ib8HjN+AtYHDywtUySX8E8HWBb43Wu
oh3EaEZCFcT54iYLsKtThjl7OkaV+HxLYo4vOEEntpO3qybyva2s/22D7LcCKJlAAO2fpBN+TBJw
QuIf6WQqKWIZ6NQbKlaC/HuNiyq0VMEe26VahGSytbKhS+DIMIdLFWA4q6EUKUgyxWmjCAQNiHOM
fHgmnpeBcjB3CUWu83hVVpsEd9qwPGdyNakU0lSOQ5UZfMlCy+XyMT4oxpJduidqDtequgIg8AJQ
D1vjhTLvqw6xIi74gsCBTgmTFbYvRwXUxLFFqmiwXrYUCQVxsxVePvX5bYNipH4TxTAP/sjP5WZV
sL1GAikz6A2KIGtaW9boS0ViY1AnaHOnCWbjauHxMDUfI1TGK19BVlQb3l/IPyLHdmma/zlxNJlX
M1L4Dc6HJTVGt6h/uUjnhDOEmCvuwsghfhZgQwvQMukSLPaZJQjO++QWJBkdSr3Q9QyklEWtr4OH
pOkc0Sk3j15qh65+ZQkIMepur5Z3fRijg1qC8yQquTBSqig+h0bs5mW7+KoRL5pEwoawTe4NFSdt
t6DyH3Paf4zI4Bl+p+EqO+CVGSz9EowC/i87J+lYIIPqegD7U++O3qKIuqppq36H3bUMxramq0FA
GznEecM4wU1UwUK027GCnjppTI5DH/++TmpTx9/lfZ4uifmYxlTkw0kvdcfj+qDIBwxjuac4k8Gg
Wof1OWIgN1ayMS//d8MEzr8fx25OeE5pnr0N7cpo2Bxk1oP1xyxSJxAHwFw0++ymtdHeFutsn/Mw
upbVRpGldUDllNarnuvzhh/W+gFMqdQjxzKS00rucIpebDCTFRU8rvhsYB42ZQ25XLqUPpaz6+KO
zeapV2KTVhED8qJjGKGas56yDP9lBK65ohZh2qHTBva/oTKujpGONgDoXiYIYX8QJb25Isf8UFEf
PA4uR2IqmZ463Gklgl5uKZjFhJSnOdgsnrTeqQqBT28kN6cufpf1lCLsWXkabJ1rjeCVHLPI7oj7
uF5i4qkYDRv1TixhGXCzTOYdgYh9D8W7R2zexAZVDxHhYBA9EQoeigLs4RaV0xvcI46R4w1pbajU
TSrL5e0haRgtP7mxe2V4Bz9U8Q4lyeanmAN9aedgHwnCMW1ADtN/vHQ6k/+HyiVT+lwCBc8Y6Wyk
oyMlxkpwKxj69ob/M40qWS9VwNrDWqI4nyy2lcgdT42OuqU48qeF6a1nPvKSA2+c66wePFWaWwvQ
XJijVRZ13t+VQpbHZdpKVFbS6q41zzCjhkd+gBP/2x5Syu3WzjTNGF6NY/BVkV33Yc2jWd4FlSPj
eabkEhG8XJW7AyYASuUBgr3lAIl4ESZtiS2RcJfcCIbtqRqrITPPYSdaB3Qe20WxHJr9tQMya9LH
eildFuX1orzXlyrzWMfsNP6cT552wrNHvROqq2dokhnBGQbNFDg8q4oqGOVNz1EmHMYhn4cgDltn
xDxAw5+KjYN6+XyBHLqzrMpiPdPFPvDm4H909w5W1FbmCQwN0KTPMUkiHb1ZJWkFUgM+TpHaW9y4
XIOpoG9YVd7wM0TbRkxY3zsvg6jjOiIIgfwcsn+9Lmc6M/bwJOy8ty3Z0eP+dNpz6zaSZ7fN7vqo
cd/ch1s0muy++jfRHScbpfLQMz8NtrN4XP9d0kTBgPBaACqddZ63LmUHF0GPQnrpe4vVzTdiE1gk
RxkRosa9vOYBvLg2rKJLlSMfrg9BHKouSaA9aOBODp51f9hFCNllY+fKnSCIF5Aqcoyx6mcVRa3u
C9wMVHHsPPTbUPI1EqSroUTsKqCrGhPyt8bUFP+6Qz0Dmv1BKw20btOKCOFbf7J36uiuCOqfPXaV
7/wJ/qF3PsHocX7tOOk4eFt/mJGQujDg5W6BkmGLIIuGQ+xQEeOTyvcYZv5ijH8vZbEhYDj361Va
yRwJwwsAIpzb58Y9e0c73S+ph42LhG6LFZsM4vgSnRpdGvgES84rfqzEhzT7EBwD7PD0fgq5PKhz
EmPgS2SYvPCSFGK1gi719EWFoA7m3DKwEioH13jEkKaxiZW1ZrtWEKqi2sHd1DxBEaeVyuGy6ySe
z3MSUmM3pJ5XGzUyi0FJMzuxK0LfybJq3il+5YYd6ftpUPsKEBuk9/Kp5HUoW3J6ii61t50cpMKJ
YSYU/M0hzewAtjJGYl4c0jdR20uWlg/tdddLYmGEoAg0mgxJrTCMbi9dlKjlo+svVfRSry21FHrk
UR97a2cQSHxigJXwaSuSbiX58LRxLwlvarhHTNGRAWBlkdyWMMSl2/1ZvYTmP4I+V1hk71g+YzW5
/WaQ4lp4c3ZIVJmOmcJT+vPH7VStKzCfMlh4htnc4Ks81OMxX1R1Mdv6EZQcKFDF6WISCI/PeeyN
byVeRNbM0n64BZjqvkiW/QF8Sc+j4lUfbczX7EkOIYxq4ikktEi/foc2j7DzMpBLbGViz7uZB8gC
ZC1ulJZER3LeVo84M0gmHtuOsorm75Xfr/OKOkjSFhFP6w9fjD03E3JysCL1rKYJKLbk9Jtnli3T
rJWc/4gh/GcacvytDxxV1BRgoZuIuWb0Z39g/D8ewcfCG+RNbmHUQWMtMIGpo5aF0IyV46DnHZ7h
C1SSmNvgcgI+TPe2llTC6DnnII3DKTDhu0HBr78ve260F/KzY46sh/C9cbGyIuijcI+aDnMuInIn
HVH+EY1oxECQaZ99YZBGPklaMnV+fNF/DVoSqmnd4kRbi8wgI5juY7gzgJQR8GhALIC734uO+02Z
Cz72RDTJw38SEaSfbUS4ZglrJVSZORGvOlb/hxjILM7o0bVGYwfC+tIeEw8fLIvI7jrj2mF+ogp6
HCcygWwvp2njWchGkzqFKgsJD163v59ksgUyXdgwuiI6e/LLeD/gXpg/VIIiSn9MgxpNqOBnRqYr
HsD6TPUBXvGzLebwr/x7GNNzd4bhhbDpLNHETaqOJg+Eq6t7uN+TAZ0ePBBTu+Ur+OPdkS/AvP0h
YuSRadSkPqm8dLC9IBACNYvRwhHwpLK7QfDx6e6ThLMWS+Fs9viQCcyZMQAXgQePvRMwWpI2CBc0
8eFSTsJ1r4VxXMgEsGlJNyK5ixYXdtP7EDremLR3ssM9ioRpIwWCcWs0yZOm1LTesjBy26j4an/S
Ts1BlmXiCjqVJfTC7OtBGdEoBQp+eFjdNbxvB5m1KyuWWtd0qyd9PJigspODfkXa55ACcK+MTVkt
607eBtRqmC6pRjcf3tZEnyAkO8/DhZ3mK23H9wZsBLeIsm3t/9uwuE682i4tHE71ytvP9nrHghxk
zqD6wQOl4LZQ+Ea+kErigLNSstjRg96inqaV3/ueevtJ7bhMyh2fAdSED81A0dzDxX7MjOcfJ+si
y2bI9k0Hq1VfMKbzo95SCA4OpCiZJfJCRuBKccJWJjNT5RMH5jLxNZk6r9yKQL31C8oKCMORuok+
4QfTMA0xx9s9eLhq24OiRlEhsaXMzdUUahodhnQ7yBlppFm6bkcS578aLG3A1tsELIPjXte+kL7o
uFhqB36LnKRiW8ADdD9XQzaF10yDSG9xRUo1hMuGAuk6oMW/17LCYwrGTxIeDLfTUx12yWLTVllJ
BKyB+j+SDPWfdm1AKy+NS5hnpRcylWc5dHIqSdw0rw/CLLe5EtphGtZbEqdja88qwxtVRy475ByO
jp8goGNQkS3JEvHvmBTjlSZoKbWiTlwCS6QH3EtlB6L8wTOU2BMHOHMCcGmpOin2aCqf+lgYlxam
Gtf5CyNdLq+NbZO427gOJ+n5l7KILyqQ1VXz6IqJeOByAbvWiDJ0VyRVXec2Tcv7c5YbwAiz24m4
6rUYN7taYXob9hfMq/Keve/1jlyKUru3UbJDUXAvkyGO+TKqqpjvAqGdaHYx82xD82xIvNsG1VKU
qcR9Ns2B9kE7wl80/YmBWq3FVUqSFU0Jl93cFNcb9R9CzXqsIX+/b6s4Ddz4fqqAogcP9RXXdic6
M905iCvR0LJyvioJCEofyl47aBNhTuZ6Neotu363YBrM7QDBbnNrKBfLZEJprCe8WtaIoopJkCtK
l3nqUBV4Z5pxqCt04mMIuRNi3sPxWYRtNYvFu/SgcaOTWjV7NKKrUyBMYVUF/vBrKKWMP/01kovA
7V3TvB4/0XcWL1DnxVmCacz4YDSbcPslIDynQV8fy2+n8kis2geh5y5K8WCOR2vs5kYRC6ud1aVk
xcuTPbvRUQk+DwUllStKhwdIu7B+AygGkw3SxetpXIfgBNC4dhOEWiOtiQPAXLKQ6yOCdeEKC9zN
FKSV3Hb3olvcAZgcuLMhHc7O+dssah5xAHDJgugVgx0dOPmf1Nsp69BTNzxQ0B5OGNKAv8eQ+7VW
RbDfWU4iyyXCrLQta+Pft2Z/Of7zicOTt7CXDGneGTKOVcOYf6yX/0t9ZaoI5ocPnUmVuLpk3c0K
4AITSHjntGa/Wxt2oRk13x9PHzJvGcEfM9V2qWQ0U6qe7z2Z/FbEVpzzLGh3tQXKbxWZmhq4Rf05
an7BfoTBqm1Rb6Q5in6VsgLhMMyeGVbe7zmkMScUIER9ILfmaN+yDkJk3kn4jDseFnjQkByWX5X7
ngwMkRFypZVD4uguWt3m1qoQ7ImQAWbzn1XAjtMsdENoENSr2p2uKI20jPrhnMwItShpdmWl+/FU
cEe6JsJU4sutmrQfr18Skamw4+frVsdewv663xXTxIJkY76z3HYICXgIx5uOsE1NttPaed4DJwNM
7RO3YVCD0S3gbp/htMdI4xWlVExaB2d0+X9PWPC7vRy59xaIJBp7dDTh6AL2UUGs/Vp6gH4+iX4M
MSEsJKnorV6o6eE5SwSm17NcLN4z+EKchXMciXZCnyDt9n1R7jnpjh3rja/U4VZH5naleIUqeJ0X
fZK7cKGq8x8Az2vWQvL3w9yGOawQfNPDb+9/xyBPGpll//gYMtrXd8UWJW21oQG4a/cJ4d01RXVC
SGT6tAGvOx3t3XhkXZU48OUgBWa/bu30Vuyn85noDYlXYkiRYhf4csZ3tTY92gZ59T/JSvPBf2e8
mY+ZFcPhXCfR/IEHEfw/b8tP5wsoPJ87g7WXNPQuSv9MGf47Ko9LTYyyOdBapz4kh/2WA4F3P7tb
6ibUtA47PgChzOV13LZE+pazDRtcUmKJclG1u8LcJICzdyvhRJTOCvy2ibLFbuPG+l1wdZNtfDVL
IpzuR41jDl3wGTGDIYmrX874I9OXUKP9Pc1BDBE5pIDmCVptBXG1sJNNgLdi5WymEQQmVQeUQZfC
m3NUiHtcSGZQZlJeozGNrMtj7bnyGnMAWnIVgFDbwrskQUVtR5DUzNin2NJEMJL1tAshzll1XVwk
uGj/y10SG62RRSmLUQQ2JD5+/6uyra+vvyzGOBD35177rrdSBJDrCHZCi9gT+L3100uDhUbxjuYz
49RZvi4lO+NIYkBFZkwVKdNUkWJGOEsLDG0ejDVXXy8wLNKD8BsKLoBJEnDz8Sl1uFdAQoMblV6y
Uzx/asWM1IHfIKoZEYfs+9/ndJma2Olcxsyi6r46kjZtZsVkjqMk9inUv1oOk5hZkV8nmcImA2mB
kUWxD0YmSIb1kQD1eYZGI3WSsePYs/qnM3sx7KzlXHpbQsUfMexBA1pSsEM508xKTOmI2F+Yu0kM
sP6WZSijuk5kS/ly/L9liCpg5/0s+ioMSZdpJpuH9IFImztjoWXtXrBwfUFmC3894TIDrh1K7ptX
bVVYI4VOUF0gHHlvYs9SiJtURTzI3xVlQEGMCQ/oM1dBUl+/jAYowBBXbVEKqYmjBgh9oOxPiDv6
oLPgb/EJcIOzOipgvtaDkyIu9XYGKBkEw1u4YICmU69QHG0ixvgsJaHHsHzj8lwtJhr+XMzP5p89
XhBF9lk4GvFK8B+Cs75LIXTkp6JU0r3HrmAFxNbI7EUkrjtE7JXOI1hrislOJ9A6O/bWh2Cc5q7e
hVR1MHM4ieLfbSmO6ClFiGYAHugtwZI+d3lf/vUFALmsC4qmwYbkITq3GcJMsz3WF6JrSkoO3yKd
SDAVj7L8Usf3G9oNy6cUZV6wit4SZKSzAc8KMNIQhhgkQ982ufrXpyM6xaG3c8PjJP/5wL9lOcYm
NPZMUfv2vu8z34z7YG8r87ZIG57obGulmpgOh+RKm+clyOz5gzeczJyZmEWbMCAF+IZv1PQYH+ZY
KpnCH3MC2cXKZr/ef2Y6hAh/tv73VMvKwYRJQvuc0r3a/uHq3FNXVjgcpTzPgIydAS53EzUv90eF
U7Pg2adZIxaO6Uy1hiYUS4xPzrM/3UT4IsDWbaEDb0wcVnrd6D4G4qB2ItJ1BFaW0L/S7MVRRCWJ
2lYGkArmC6te+wwqMhmi1mYZrMnq5daM8URlJfldKE1f4lcHJ9Zu8xwab+g0f7UBAKzV43MWZPDQ
WlGaihQyFE5nzy/d6Ftkaz9jpnL5Bdtd0QtVpvOraRiUXFY2kUtrAXpwitRaKthnHJKz6rwADL3G
YVom0g78qyOmy37xPFsZ32nvqFWj3jGrOi/MgH9MtGL3I2nVTooat0tphq4N9PirqDze3AfeXJ/D
f7LWc+vZ8mC2c9jfRFa8wYYtkJOE+LlynBpaqzSyaKYmzL8gEAJxbwzv/2xWScn7ytHf87Wdh4BJ
JSaASXkJAEQsAOK3eekNR7O0C4Rz8p5Fy+F2URTBM6rxrhHM1wQaNYVybdbojpj3aeFYHUf5xqfY
iVLjXqHCmscLtEUAwy5e73lLCdokT6fgtXddNOILbJHXEgW66aM4He25rGGoUfYF0CevIuC3d+KQ
1hOH7iFeZ5YMhtyKhgLkKzNY2IXCVj1vnPo8f1bA8Ol7goAJAa8N1fl5TM9Y1rJ1iow2X+HVSPQT
LjNfmevo0V/ts0g4YadDtC84v+zzdAC4EFwS6qnP306V15lFWTbNZ6cHTKIVyclUXmtp0VmpTGe+
ftrRWvj+Ay/SejkQon/nC9T76aWgq2AnJ5M/FGcqSVzFCeZsOMAuhDT9iRB06H72OFfdFFQzbG2R
CMRRgCjDdVc/m+GkIbh7Sz8x/2NpUtU/VykOKZ+XXYXtWUEi0MPZme6gfK78WHDBCIcAkiOnWsw7
3gIkmnxa4znD2Z/kyWscW3QuwxakE/sRU34EX/2ICEuX+8hBbKkZ1QxSyWJ1dZPYApAyqw3oXzBh
v1Dxy2CRV/EOuXWIbTmJ3ePVWBxHtsLVLujhtVD0XvGu7WdWG/+PhUpdngKtPJJ2nRtUbniVjkl+
wyJSxq5gSSn1+bKe8tn4FYS5/4zLlwVHC292VYGV6/0o3Sdr5tehlDbK14KNrqSg2yBQFSfDBzfw
m/UM9STXPeCEF11+c1f2WFhc7Cm62/FiZi6ExcVfqZx0NmOxFnO3sSS++zbPtr1JyVFieHZah0ds
diNtl2Hh+sM/fCRWYEPTkf70kse1/q4zrEolLIPL158yRR+Ga6IGj0RmWdUYun/DG4CiSCdJLntp
6YErIPu6ac7X7Ps8LlBp/RpKn4nXxCbGt5Jzww9XvXb5ixNNenKjG1F1AMTfGciDk0tu0bHdaAhT
WeZzZW1zpgMskmN5/sKmBkv0xcCx3fCT+F/IES5FQqtEbTWQ+n8iEwZZNQPlThMSJxkIEJq1qRjU
ttB7QDp0fAIlUx0X27GhOv9uZEY2w53vVZdL6sneXOtaJCZCrEsDQ+WlbqeQmGoO4XrI1DrC+VaK
UzKZRIvsr3RNhlslY3e79xnkA5+ksElHAgRVwq7h9/FWE/5CIg0Ckf/ITH2bmpCFI/WaABfOh1K9
zn2XZd4u3BhAjT/tS2z+BjHxrghb8w5WjdqpaL+ABxEzxssfztjdaXZJRnMIXkX87xAN76Sr9B+I
64Wq6yGzBXOARXig/W9se+aXza9SENuynK76l8OQ21GsbqW6GdIjaXuk+q0kmgWnG+/xvL+99NhX
aROIDE3KHDVQkIxekF91RPa/cQmG/NbrFqsbwnYTcoUv3l/1FqnwGr8DKApuqn9rZMMozFbljI5/
4EeLkU0Tn83UNimCL7WMuZ1hrNmloyP3BQMPeUYAsNyT8Z/n4ACigb1Y8gGYIIZGqrgv+a27dZEg
kBLpJYB7nDCRC534jGpu0/VbX/G9xXdEi4Yz0l1eptaguDw+dYO6Lztxoh0woV0vtl+uZflEQJaf
fLa2dRvOPwIEUtlINHAaRMDMBMgxTBsJBcLbkABvRgwzQIxVHEizE7mm9Qvguux2Orgrh4mP+a0A
XEhg2qKexBeNmLmJD04UlKJUSuKFjzqydPDvrC5UIEMdztF42pT6aOWDxaEo6P2mGisYJp5im+/q
9VLYAc/4xJJTCF+Bw+DF+3itQ/NuD9KviKmEZYXWV3QQgENVrxyNp0GMl6wvDj6ZHrWq0UqHZzob
Vacd+HsA2yaGKqb0EBeIlDHOpESZY1GoaMxFyibU+bF7O2Hf8yYkICJ6Owk7OhYcHyQLEyxKLMJZ
nGSz0um3TFPwLtlZgw4m16jtPveLxv+oAOoX5Fb0o2c/j0eKkV8e1V5kJKGdPLrnbnjoX4r818Ir
4/kZbZGMBEBMci8/slFmSb8Z6RAM4VILcTdgoLCJVJb+ZMDkSMIOgtGXDPFp/SauUw92x7wPOqVS
HCVOIZkw7Uj+ke5NMRsUiml7TnW9YLdgOEDzMdOokP2nmwqrnK6QeymM5+yMbON+ZiBSJ9ti2Hq/
ojT2HHwxJWYavOm6FMjkrPklmEo23zjEgBa9jfQOOMkIGuElhSNc413q855kiQQheewf8//C38zS
lz8CrKNU8ZEJs/m46jLITisLy5LvszaCKfu1dz3+RJ8i0hJXs8aJFYQgoUF6qgG/CHWevvnSKtPf
IQwp0uaGKMquM62u7J7YH7cUd6m0nUl8pE8mTSkJ7lptTXurMXdfjrH3Myw6RUHedkX7+ZyDs8vb
3Lwa2WO8dnq94yXUfNA6ISt9Xw+TUUy7THECZ7zdoPoXWXIs3tf1fCchouqxhjOqrSs7K4g/pvRW
0472a2SaRpLRnU/dbHWRkZHI6n5dz31HTKfKbxan88ttuqUfXpLHEwZUQ7EQy3Ejj4+iM3yOAx7K
mW7Akv/0wpk1iG+e7XrtN7Q8wE61PYIP7a2RsHRYI27U6sL23qG9cH/1leNY81bjjRz55VhVZ05T
ZOlgQ1P3Rl4suHPzHAj9Fk3x/CFVVO1AKK+D8m+oxmsaQfqg51bYczEOOYXeLQGYFRVgg4aMEPqq
6S7E4KajdKxS/xBOI6oUS9aO2oNRYde32NP1ZgEAgmMw6TvkxcSJTQSft87HcfIy8ql+W1it/E3B
p4z7d7tMh2VnvQ4m1J4xbwtGYKg1mKtH8/tg+fViLKGx71z+GGny4tHV6ZRB3GenAhkRpbsMUgVp
zVscSuTSWL0CP4F/pco+7pYBAeLMSR8MynqvH95l8WJLgGjilfxas/vg9HDueVCJP4vhK5q0/6YG
MfRwCm9X6hD9szUw/5GyOZkfnRlqmvbYqhmJ66flcAwQEZd+KcoNmu12HtSmM6Ff9jqc+l03DU0B
EU1sQc/RvyiHX/1WGA7xgxpl3ppWXVHiCnM+mfk2pmkpMO3H8gvwjh7oActAeMGGD686kcDdQldj
Mi3CogiKS9OjdKnn7O2KOGDv9PeT+zQxatGCjFo9hqB9nr1zTvNjhZ/Nk7TV5A4YM8Ze27Z1gh/7
vWjknteo+D4V031OnQ/Vrdw9Q0GEEMvbA0iiakhMHMiHAKMIsnQr3LqNbR0fLaSYd7SiiXxOzmPJ
3WWV858e6pbcWrWru//uFH29Vew3M666ePJ2bVEL7wbuqDKIuQbBn+bC1AgSH0O1uEUzgK2sNkkD
ArBRb2uiCrn8tjHs6VUcNuGKMK9Nc9p0S8JCnPEIhBd+G9EftD9aMKfarDO0sTD3aamYVEM7Dh1o
HTlV7JAAl79tirbN/q+n9AAc97XRL3vvI6boNSxAp1GQzcIm7tdkhSGA16ti91HhREZscqnf9KRl
DJc6bEZ7EXAjOncZR6+YXxc3tQCC4kx6KcRgH8hEhVykm1vwiAzueHxBVAuZAJM2BsiSTK4sXLVq
6mEleHf0bTHIzA7stbOGb6Qu6X/5cQcwNZpVVG3aQE5ssJZSNToNdPxXmg4aetFl2gFWaVTBwJAk
Duieuu4qi8S13OUSdwBBtKksnJxIHImj95TOTP1kZ6g7o4hitDDriul1B+DH89dr5SzR0QtvI+UG
5+Vlk7QmMK+sJfl6VgFi1rN8EclPJOAHYKlv0XS+Fsiek1yHuTk+jdvf89RtxIvG6tqOlIYxcnxI
RhCZ08VW/4BQ3H3OwAh2+5dY9pRiNOXBlgIXz7O/wUlcj6v4WDjaLBJyqIeTcR7R1GkqCn2Tp0Rb
bFNjGZ3xKSRaA8ZGyfn+hCcvj66ToJgu11aR+05UJaRBujsrF0vHBwB4mgPmLp0+ou9iYSFy6jHf
VE0KKXLus1O1UlHQH0pk6FtD568KtEKLwVuclI/jHN+Y6RKdOsCuyGUKsvbCTy3iCpaqQN1++I4K
kdD5LpEWkQ3Cw87EQRa0pJHzuj9uXpA6yST0aCxMOoMTK5Xit1DMDGCUU4ELcd7QSxR2xab8TdWe
80esvH3K1kC60OpMKLhWOJWmuMy6VtC1kSnS3nTeOXHyenRsDF8t4U23SgCj8c995C+pCk5QF5Uh
XD0IBd06VyQky9GXckYgDCQJfNhkQd+LEjQKw2AQJbEILpGaiOWfdtowYhdvRBpPzvkKt9mITSAg
gnB3SS86cikW39afU/J/o2UzY2pg/FAkwZLdaWrYHmnmLLFdTzVqeHqc1qrlMs4RmTML9j5XeFJD
y8OggcONi4/4xFPdVxD2zpNG5ACxxroFzzXsOg3BHuehvPIIbKQvav+HkZlaaCECdqNJEKmioMNZ
1c3Yn8sWNAVOi5WZ/jm0Quo5UJGgnkFH73mpJiExwJ8GSC5Kp8AuO9vY54Tomr3O15/GhxPf54Ek
cooK1mIo+Z+2LP49KJtvjvGQbT99NZSrNERJzmDjRpnE7Yu+79+QEjTRRcB+GDyNfBEeR0q1DwXh
vHpkIMbF5ud6An6B9YDHe3nwoHHgSKKiN3cyq+ucSHTuyszDj1Dhq/1zXuGOMHSZC37FI9B7kQ0D
uuUpChYeNsBZ9n/b0cRVK1PQX4IelEBI8+bYE3xKhh4g22KVmBsFC1lMYuCs+s2rm/wk5IS/XWW5
dCHOvj0YrXbg5cGqY429BoGJTsFSybFmZ2gosBIUCySTKVMKGoJIGoIwbqaNdhjUtR+rsy1vaWjv
wbWN2hi/V/OLKdho8YVrxhpj7YFipn+9KNPlS3iRSC09nvFy+csLBb6bDrpS27bdijz0t5rn5iyD
MOOCKB+9JFcKTvj0w12nhNxhPkMDGNsCf6YnRBmIhYC4orinOpf2Ho9u3WnTbTZqlz5QRAlMxkUl
pk94OWijE6/zcsPrMcgs0ucjHtgBZyaXqZGX/aFYu7m+P2nJPRfhOcGxo2jCy60qN8LncZsnOoHL
4iqGn2YfkU7NDqHHIoo+CqGaJ6WH/JzplTj5kGNtNIgMDqASC6THtINxOKNVjoy0UQlpAzv3erEP
r58lzUoS5415KEHIFM52llrnI6E73ybM9riAbeHkDPmu8k5EZLrpOX/dhRFSug5ElGmHmyvnAwkd
BRx2oxAWONBGSNAU0sh8JcBKq86K/avO74z9Uwh78u9YlixhxJCSAnvKQN9IpgsDQNCcpM//kqgh
k5Z67zJKXpy5jrNlC2tyPSJo3Iv18gtPu4X6gTskYrZCduRuA5YiIynrwanagiRPZ8dwvD/VC5Ly
poRKP41sGXYPx1DTD03iQpsw4nJh9eGP3o7a9tLRvwZh4kJ2cgJiMm08QOOWiWJRXa1nSH1k7fj3
nQYCSISvueZO2MfrNef69mhouFK3VjAarJ5W9JhxL1DN6NSXujq6fqxyx7sk90qZiGycSzIYR7hS
CH3Q0igFxL80pZDnF2+D04Cl8DL2ssBppLUa139YpGyHBXme7VoNUE1E1nYq88i2PkRw2s0qUijr
4o9ksWTWcuYnzipZ5yO4gkfgwYpxuDAXKTN5oduikhaNN5vLL2Oze+eV1XRWPAnZUaqnrQqjhkjm
E7+rZaCUsiASWo8HR5P/ZXixv3UXud4eBiMzXmBWWPrwk+pvlJip5DmrMZ0hRH/6kS8PBwipuumf
v9TZc3gZCTM+447axqgcBFLiRryKanl6+tYqQ+DRmHh+9ynE7AMDchSiCBVaupWbjqfF+0ZdGM9c
oNZuYPT4BLlrw2BWb0QjWMAcdsM4kRADETbwBtZ8Vpr7xCdj9sX2Hx8obEHL7YS7qrVVI1FzAGh0
zlm8UmqhkpTXaM9MeHSJitn0ypm4PaEpU/iCSG0t6WdYEEA0twrJsupqzjwPLUABxY1Dykn03zyr
GYseJT43j6ADbmXlnDnmnGhjCkDNN2OYucjjEFfGLiZdk2SxPPhuT11iB4COzgDsbadtdwo4/vyJ
U8nxmmjQrEinKQ8QeG/Pj+Sy0W7DPY3J+aXk24J/cmy4yF71DwATZyA8ARBPwqC2OHhQSKf32QWh
9LW7iAPPLix7AalV1xr+Yw5b1bpJVKftvmUl9c4mUsEVX2lJJcsNMVAw+/mCYELv4IewFnJgJpfd
WZvvYaKFexFXkclw8+kntkG0Yeb83u6G2T/2ALe79EOd4Vp0BRrvPb+rPjEpSCThe4QQUMwBX+z2
SCNxI9/PJgvWY2rHCqXrBetEl46sPxkcEg8zJnT0EeSfxu3+SwWSjYJF8g+OxIa9Tcix/NTT/M/O
fbuDYwSyMAxug0HrdpEo4u0CBR4BmBRiUT3pc/vUjy4I0dDorrl9e8BfvxTnZMo3PDDnZDZPmQ6M
x+xNOOtkHI+jdMwNIPAgoNDyZAC3Qi5Q4WKloGcBtrTUiYkzGa0MxDLBO+8IjO+O4on4ATDC0F+x
GD4Tp0mcNK0GQJHRhkitEu1mFUx1agPIOwNMhZMKJqpvr9jfqCm4QAYoiGODFi3GgGiFOahicmId
nGY5XVt3zCRq0biqIR+AEuE36gQWXPZIqZJru4UC3vZUdjMDnW/v9N0KSWZdsUw8dLnZ7LIMSUKW
/rsPlJLnezeWjg1q0OWXsr17zoCKkzJ1YHqcGPm5L516TXMUnwrpVafwz/W5unG00u31KepU4+o1
kDdqhJNuv8r9yLEmtbEjwbmqNAvHhKVzGox4i91p534TurCMD4rulaWXrphjmDYUN+vcWgVKzspN
i1OSZeVrqQ7JzpdL9txySfK8oQoV6I4r0OlGnYr2Qg31OfOxBPJcghTz9tz1+rIkSdu825UalT7w
aP4Vb4TiRjAKqJV9uXePOEIQEJMe2WztyCWy2zakQWhxvjlu6LAg4r4SrbUYtglO90q8rmo6zi8n
djXChkN9MJ/mllVeuhE+s0fcYiO3j0n7Q2oZFkK5lMw46Vuk46RWb5dKqXt2avrFq9lGalNlT8yj
3Zjtwt3su5ixdblYlOBHNIa4zaNs0Si7tulrmosdRBCPXE2LUL4ZzK1tC1cNorjlqs1oE88nmurC
h/Dv25ndgAabeXmnon1q2ZlgOoy1PzIoaJs3tPDFfzfe+fdRhQ4cIRmDxEPaEz/iFco6vVqhBNOh
AGse4IKC+wRV5MkJF7SiUxagBZea1WkWR66nkQ/X0yE6oBMW3p+Pal8TBO56wIBLGLU8xk1FEceR
PhfN0xVrvtf8Ud2dzIQ1P2wjlvB/67QUiG60UqYQsxkpA/6LihxBodgghmSC7/oQiWfr+8emJd3m
JToombddviZr4KpXbvxDDGmpNHfnXgiVFb1o//NAat6tSpgM9lSwKZaK9U6dzERe9A9126lrxQFM
V/Uz5Sk1iwqjZRYqgaKjDn0lErzwv7cddQ7+4QIeBRBdDgDHEkGMEnfHOssoxpf8RwwMKpRc94KO
a1BqziSjBcdi7bz+kcE7qPlinWvtMM+esUudWWrDVH2CzbBd/JzDRVg40L91M2S81gXp/LQstt/A
LMvQjgoeogiXEA8j1D22i1smfGGV7d52q65I/JltTP68gaWnDR6moXYDoLEtFCfnXEXbwfd745Da
ouBVf/ux55SRsTPBsRNpROTleICtBhomLS4PjfzhuqKGKK3GfD5h0v/Nt3YEC3x/VhyFirjTyS9P
r9jA9jfm02j6HKKV2EksjuYEmSXcA/mLskBbYrGXTTIXrWaeA7Q0F3EFffvR8pqrgO58SpJZHiIa
Z7sYKv/K19tmEqnPHDVFPKXIjK4tOcBeCvmaQwlAXnmbDYVo016QLhKfAjv668n9w+ngWmCkFXJm
gcCfo0WeewHFVkKxEpVK85z0tBogv8+kjSBYDrbpkZKAw8CC7ZD2v520XjJQgNomv2scTftcO+1U
RRlWFkC8GKNisHq4GtPHRsLEdYU8PaP1UtJq5lYsvvjFPeY5JX2n284ElAQecK1Rh0i1StDdvzG5
GHPntV+ayxJ0HURmG5UpyrTPoMvMr/UP/aLcifxpxH4unRuky6y68OCO1mqnqa9L4EbLBQR4kxIp
ucX9fTKrqT4o1cmBvlhxOFYmwuUBBeSOSEsRNWifd4voeeEWQMjRHJQZTqaC4A3qHTUrZlKhAb+0
H3LDz9/p+izhaVk+khf/HpDqOMusSxd17JNExPc6wbn6acqZBu1YygHBwQN9/nX75MPXbF1guhhH
+n23ziDvyq/xPttQFI47udwWUzImyLnB94K7YDo+yPNsNOBesacqI64CP80e6Hgr7fdc0sA58AqM
od3v5uuSWGTgMmIfsr6FX1AeGYfF42y2uHhSgbKhtaar7f2dd/2nJ2XkJZ1IK9kAsw5TxHBKhu3b
2QQl11TOkLAq/asjr1c+WmMaUWb9ax/yCKbHUgbE/NNPB1AQy2VJI6ciLggoA0CRdjyaI9cm7JgR
M+/DQybFKD0nzZOYAsSiIxHhqc+UUF56NSxDp1sNsKBeEXn2RvpH3G10Fa3w+0yJAFzSM3R6ticT
EkPWKCbKqrfPeF2ufnXM3W7lZqQ7cvWzxVt7at3uSmuPPTJlkuy408D7MlU7Sx9uKVGxsR26XYAy
DJFE1uuh2+KkXbflLSZCwKQpDf9M8QLTkqEpLOcpYcjmBdopNt6VCR6KpUuiDclrJPHTokPzLgPl
Sp8dqV5rjM0NMLfwJ9yyaMvk/DSrU3yWYZ6COpvdRZJOXMsjFIlgNutzMj8e8gH63kcDw8gyYx3+
VeeYEjEk7ESkMm1Sqo/zxv9Ir/SGIvYojofTMGouA8oLDdxE/w3UowltaKiNzg9a38HvrUd4eKOM
G3Fm2NWS3VK2CzZdLkW69ueZuxbrHqnXvur6x5LvOuOsryvMZ9EK1A1Ij8mKjVRezn/0cRpgiWry
TwO0spv3EslLMorCQcWvYpTFgHrgCxirQrwtOb43Nh4yop3jARL14UguX0TYWLoz/V6bCULZser9
Lws3PHmMYBAbVaFyOwBWBIhH5vgNpzLcI495sFQ+Fo866qiEb97zUSYNf5Q5mGUZAdivYN4WpDT5
26SxhoMeGnb9whCNJ72q6chgaZ+v1RNX7BzV8mftwXZMUUolYT+DYPvFuxGlSlH79fx1snacDiWW
XwfIu6fWWjI2Lsa6A2GYtgI+PR+u3kvaGl5cVxPsDvZnjvWnnVpXo/OlIY0JwV2v/O1OPFUaLCZ3
BRWJG7d8hTEhHPbga2p1k25hKx4Po9dvp2Hugko0kynQFLXmtM9qOqJmNVtDD2LMlDQ7mBCj6lq9
rWbj+nr97Zrf/+uuUQXXwBb10jAmQj9W78pr0M0hXt8c6IgQZSSW0idYGuTJpxuWHfq0HGw6XEEC
Bw3z3c/a1ZMdg6Gpnua3hdgEjQLDzE1+8u1JbzElQCSzWEJ4Ada7aKWRGT5kMEIe+owmf4meu5nx
ADLfVyR2zkgq3lqv2F2Prz0LvVkgXOABkn3IrVXrR85EfLY/p/jCTfy6fCDtlfTSly+vEVjqVca7
f+jv4a5ev0JeKlLIwx2MsQequLFv2xlI8a4WVuwf24HFKIQ7PGUPrCrXrcCmwlQhD5GbMCa309rb
5Sxh6vmnIh+6iCgZTf2sdCnw2nAXRJVqVSkxz+LUaZR+bLrRYmn5Oni86OE1orMwsZRMrRdwzO5z
4PUE/zXIq3CGaobvko7E3cV32DCIY3nyJXi82OK9oypZHxiUANUCCbuYqvekznT75e0FZNt+vHrr
Wl/Xkf7/5lWWW7Zg6QawWV5CnrkH3KIXG0p8uBkobMHYD12VHAo7iHaAeMKcJBtQ4yk3bgz1xLLv
GAjiuVqlzDFn9g3f+MtiddsUFZ8f/z4n/ksXsZHleCkO11oy8vTXWhTXy7ADV3dK5KPQkgmEJSni
l4iIcZHC4r2Jyypv5tSkolhZabtbQsd19aEvwRedcmJFmrdYWSyVw6P5o9TmNeyNr9nyas0ordGf
ukaExAh0n3SF3IDX3AoXp51sGnkNIrPaia5OnwVooT8zaNwLkLNWZan7ScoTVNJHgGIRWwueMUgD
yPDhT+rZ89b9nmNwccVwvA/f4Tdp1MR51fuM2i4ck7XgvMZHIp/5yzTtl6CGeKpqNh3qx1AJVljY
NBN2RmMHqkm3knA1Tg7cu19whh6Q4uI0p9ltSZMUi/V1tJqO5/CEIkHhITTuJdoj5bGk5V+de0LG
cjZpnKJPznhr7i1Uhxe2DZJ3dt5MEX/T3gGE1NasKkq2KaHcmkEv5P/f1iFyFs5d5QqhLsdNHSHn
cdKfaHUmM81X6LgC7FC5nF5NusMSoNubD32ynutVkCbA/eGaaR1zgOrv6brU6QTvdVVRz9Sw46iX
b9jlOzDMXTJysKo2VZUQvOAMqciVwPGrQY6oICxlaNPno+zrWhzO9fq2KifUhs12vlW4pb8GzuTu
udZVH9gkTslDxxg5zrmsTxTQG3bkFr2nOB1ojGO5JOZ2WzEoX9rVRhJ6BmsEX4JOL8N7ObnzNCCY
bNdaVatn7kX2LxsW0+cCEytFu6Dii2owqnod4A4W84z7wNoIi+Ca7E6aSok6fe4zPtk5Z8lsnp2V
acnY/JsO9Dl9HxByFvxGOMFmL6k9QmdWdfIL05dqMLAfVhOkY/cwmQ0esBsEHCyNONRn5zj9RvCV
N0QqACXfooJmICPnjCdAhYAWc/ggd5Cr5FRJ1FTz0e9O2V06Vy0AX78CgCJUT3x18+gHT9or5smN
Ba3uJWExNPOyXDAzVuCX20ihPf3gfbcmNCZ86i2TrCmYbqNM16/yqXgyKDhbH2AiRANPTKFLQ05Z
gbaB/wpBQf2wOXZByaen8Vf+31LQHUzT830xytqo3kfi/i8P0YYYuJPANopy6g+d7j780nrPMBsE
uPj9HXE0KsXhizYNCe0pcX3wxquBT3UQTvPjAVHN/gdMWqYfpanSU0/+39dmANYpkFB4tTCd9e0j
dxNTqBqMTsA4LPr8Yb/ZSIVj4am9KoZBlNUs36WfjutZk2ldmnVZkCoQJlW6SmLgJY48LtLoKug/
9gkdLc7JDjG2jJgKoA9NDV7I8vD3T+VN3eBQcxI+Toi5n0OI4VbxAt+M67Z9pQdCaD/fmKnsvJ3E
k3Z1JcdUkgNGctLcJ2a9KTJiDDat+FaFOQLIcMx7n1GiLEiLGuRABo5iPBxNT1bynrpaPCQfNvhR
HxzWWNS/IdY72XIvPOdypSlbeZBlQZ1PxtiqfiOymRowlNIVtfdLulGG/827ngY3yG2bjzi5tPFB
dBHWqzCO2152IQJEoGQt4VnIm2Nz2HpmAGgC30bwa4/7aVPmLZ+pJ0Sl5gy6PTB3YojuHJXuanC0
i7J8hGLsHuT6+2kjuZkX3KZlIymffuZsHSl0JdB33qlxc665C71UYuGjVyl7mzKQokJDn9AxWu9c
k4dea4rmxoMDIECkknTWCfvoVrGgHXU9QlxMzH2FroATDYz2B9fnVZJQDivxzb+bT7VYRKh0fB1k
jaEOxLl3Xh8nsChunLLlvdBMcn/luoba3Araxo7c/zeR+utyONP1lPg1CMXguEegYhu03pP9WKWG
CbZvkSpfItXLF7Amigocrca6Z0Oywk6/vLcvjMNFBv+KE/IhxG/8E3b8FWigM9Q+8hO/OWiANfvd
foMt0DlbMpx5lx9yQYbI5U7S3TYGxQpOT2mN9WNA5xAX9Er82LkI9ks6gposLWat8nnD+VQxHdxp
//nSEBB5Zf+uFK0m2YnCgbgYV8eox9m7omzZZ4O6URDvsDKUV76PIKvH65A+UmGQaaTBzcAe85l3
KCUa0YhgYNQl13sG5HRmMidu0Qu/BR0XO3uqtDxbiRHY4PA5JMkGgdvd/0Fx1LqEixcRooep3JP6
oGPxeZ9MnXElF7iuxDgYOfEGHsoLszqBJlV05LtbJ32TbM5moxlYOIZzYBdcGE1mVWRsLOsAegy7
Vap/loSUevLtZRdlzrkGtK4MByAoYBr/2fR6MgRBQKcgedC53O0Ms1HH9oNAZk6KrP+8LIKAUB01
01jh3UC/YzCbXI+qG0nuxTdEOHUUJSLLZ1nc6WJi7rbfA3mI3VRiaqNlMnlGxvL83Z/3R8824ncU
dZ/nXNiZ+6iZaJ8O3pU60UNzoPem1TqU3n8UAJAS36QWCSNS3Ls+qmjkFg7Zay1ODx47DNcRKOI2
RrS0mEX/+t6pt6XlL4T31nJwG9ntxScX0kpUqkJ06rqa3s7C3mrLNi9FzYuh/ft+x8bkfPO0XiF2
iYpcJaC+dddS129ZO4xknKHq6I8/iqC+QLAUImCvtLSHqEGeDA1ijnmGZ9DzqlbQj7qsPWvT53CI
XUxSnB2aCf0DoVpK7O24WOkMNpWm+kEUzzF1MbA+JZcTolrkKLy3bebzQsgSQ7M4H1OkW+aIcnEd
6OWgu6hlPzp0yfVDX+dLV9QMGR6535JucboWNin1q03CUs1nqqMVpeMV5qBFyEVMIl/fwnisvFbg
dkxXZVzTMjkhJIIbvlRHsd0d96OSxuARUiztY62p/XGcDZzOLPzDMQMeobIlNcxg0NBpDXUNr8U3
Aa+sXN5Hpz8WJ6afcvSdrpZB5nD+yVRmxNqlCADBvNJidGj5jyyfL+5hkIzmDO05sZFhfyGmLxbC
8YAhxbQicVKwOk5abl4nv0QMPEMcFcCC/mkf6s9YCpd/AHV8LLWrjbCEcHgpDx0f0GFsF6XN9IjH
a8uCyiIfmYg4EPsBbKH/g4hMYV6ygDCPfzCu3ngfhb9qoV2WPFxE6v8/2QPjAEDBGWJitwYD2/sE
NjbyMb+PDCF7KAj3lVXvxJaeVv56vRjfYhS4JdxZq0CiSqhMiSxY723LZN6UIl2+zVrEtJH5mUzS
N/yOh4lkNbOyYfBTocI6VRJPXn15iBeVOk6CklaO7Q6AQ3vV377L3mnxYP6d5S8Whk+g0gCYZ6gy
mqHMq+KQMc3VEV1VwMu5e/FZqHJvb/FJTso07nk53TsveCcNCua8wrh6u+XpUs5Lc1ctGss3mQBm
+RkilhKpCGr0hlNUDawf8GScPs5WL4vl1f6eypJbNG4XTvsgZbfFyPgsD72q3qWINLlQmfveXG2f
NqS2JIhEzfzOgtVacFSrDvWFt+8GmnEQAj3Ffn8Z5kmXjUYxLx06YhEkJ4uu82K7sUb820MOj6Xm
oAmZBbpiCBDjPmxAozg4UVRmKcMoDqBwY8v+FXA+tzP2512xtTz98x6ucMymdcMqTqDmPIIbQtkD
RRvr9HsuY33hXLdskSI8OeEmjEHJWQr5XSSuvLwGh3gCvmM9uUODhEFJ1a7MU3TZAY90NzKBAHbp
TQ4N3nzNYGuzJOTrWGgEEgRPvwTYfCCcGBNSZyk3NeCxyNi0hWq8NVErMA1RBb1l2hMMFo8nMtQc
J1GyFAP/nTHPQU87HAapkmAwurSA4omMydj3WZhm092FpdpWzXOfTgLl8pG/NTnz7G0NYiY74Bdc
HiNQPrE2Z1YfmJxQ0WyG1wp7zBYrJ7CcrMzUa4xOOuk5lbwXDIcNeMFrf3iQ0fPhdl9t6LJpksuZ
z3f0M0Vkhf7qUW6KKYDkecShnFqCaeQIpA+SBXPll99Nu85GXGwcLc6CsdMJ5enFAdb7FVB1Z6av
W1xgN4sji+HEvbOTpxcC0alTERCtXtjJb4JHm0TJC5+zO7tKANIbh3QnLRNbZ1ssnX6foWkzhNmG
d6S6skNn5XNlYkQpkvut0ocNU8b/GpUI1QRXCDs1SXbfRXkYRkHr3eRqaIIvwYnUSSCe0n9inic+
J9ai6ag7pXqLwa4LJv02dGR20tCZajMxrvcgi34a8oA8zoBLnWuKm/ST5Glt3NBIsEl3/4Pp4EpL
1Fd+Cxd7Eb56I9gqOVzkSza2F0zzD7TqpWol/2Ewqe1GZ5uZB2YaFCyn0jw+Y/DTbU+nxPGZq9Vn
7sRTWO8Ltqbvq2VJB+eADJY8sVBXQimwiQFXr3x05z/UBbz+buwFhbDaNQ4Xq2cQ0eSh7tNFWjx3
iQ2i5qCX//nzx11ZpfRov7m51Bam4c7ybTB+KXKUldu1kYa0OtgyXrgrOBe0bUm1ZkRbr3bir3zW
/SBKMwNjtbS85MVKi6Ze1keQHMSxhs1uHjFUNRTfQhRXqnW/jUxLCn/62NeczSM9L4cj8H4H+Fop
NCd8SqyaN5IHPEsBDWvIJtTJ7R4TxcGzHPjc3TH3dZDLIpP+4kU33hpbKbVrT1d8D8g58jwEgoeA
oStylMMluOBMMf7kyXD6DwBkoVXqyYHNpQ05Q1Z7gF/CCB56OABh0oiOrFpvi0D4MlqKXf6rYsmk
8PCz7c0Qpxk1Eo1naF9zfAwqZ9nv5+5/WEfjg7Ny61aEr0txC/UFphaIF/xtwVkjPFRR+y0f4Wjq
xAavLvjvG03hFMdXISkm0/raqftACBhcA0I7Pi95ctt0MiucFYTkIGQBtYd054Ijma9904RN1OlM
pHF0ka4LwISUPOYvl5bQ8dq4vRBqVHxJu5G4RGdfXeslKki6VuGf1OWGs8dRHYJCyy6eAa6uiQl/
oSPYWRUmLkeBLWGl31QdXEB96OGu9PXvfNncsn6pQDgx9u+toxJLY0cFAyhRwsvhY3T1YvXdSctf
xw/YJSHHaX21go2onNHvl6SGQf0i7Oaiix1H9IDG8MS1GP9Lv8/R6h0ovb8BDzgDDae7J2eEVk4i
wi5WjkgbOmXA/1dLLvlcT0e7o3vOGrs05KX2GEXKghhmd0X7YvWOR49NmeC5pOcoT2m1jlOLtIJF
23gYueudd1C1X7AtWO8QrhFKi/HSDQtmxETNRKs0bzPgoB4Jk1/YauI8Fop9ahyZh42INFrQaYPo
gTXJrY+HF2+jX+LPkyZklyhgzilmN+FvU6tvmxtDEyJ4qL1Pi/Aw5ri8ndC30irEP1Q/JyWSEHe4
6hR4FsEMGS4ttimll2e+llCQlcNBmz2Q2AyPCHF2Dsd8ulDDPplI6+wJP2dukJ19PU0jhZgLcwqA
YOnlKYfzr9/+UOliZeG+x0N2Si7ABWczPrs2oB73vAMtIQrxQcB8F0AdNpWAHNYiJqrV8O+Goug6
7RxRtSFuAvQFYelEeGFpNifok33Kc5tq2IklHdt/MugyVpQQ5dk0T2Lkla3r25mrNxh3B6GoEcIG
6j6/P0Fc0W2shq0VUXHOPJduHdtp6nprfrdqb8O7BkRaxZcmyJPe5yQKYTeZc31VXUBJTN62a/O1
cbL6Q8OX+jII2rB2xj90ITCeNq5UdCfUYJ4XU6KSOkQpApDTNngwvBhnGxO9jptLg1B/fbhx0bex
mIulke5ATjiFfH7YjXoNgEjtH/sudrLcSTXgsaKRjhF2I8STmt8W//o0ThoZuT7Ia0MHyF1wkM5U
mpTjGVSvbUuAhYETltKaIAJTqu9XEe3YM4Z6RP68oF9tY7XrT1J2DWrf57aqKvVLj+Tjw7Stj9ru
9K1cfm6dgNtTx9jUucPA+cdrpIhCTrg65w9x8xgGYc7aFUNcJKO0OZC1hcYZVJ2RFSbch0/xJUVq
SDsybZTotG4tHyEsHUIB6QvSsI3oxSX6u7/8pNUODWqw/aZjwPmlEyYCUQYN+02oqRJnZcNg2Iwo
HLJC60x5g8XHoGhFpJg6mtzp6Q8PV6CPRECU3RGUSSrX/wETUMKNysaQp0S3TdKH97YJVq76ey6c
hWA1MxqPaNkGo83MZBJf9KhCuN4ZeP2eCApZn12P16usZmWqEEQRIXi8XxA7qysbq/kfupEfBoM7
E56g/4HY4Z/PLIvrGBwv90hUmJPDrcZtrWY8kNexRAiBmc/ElmDQlJ4qhdZUtGZEptK7w+sN41un
MahvsulRRA2831H6lr5kWNZA4MiLOvFFYk6N2Yj6igutnA9udLhrp/lbpdsv3yHc9R/MT4ehcu6O
ztNh1z1JaSGyyPvaLkziPWJecpPLWpokFNoKw6EEsxbUHCEOTadSTSrggW6jKx2s8RXzrrC6CDfd
6DZ5GBnaQVipXItXzKTp31w5wenxRRXZXTLeHb7oeKezwPbrMzattqkLcO0/YOgndbX4fksecPTr
xokxLq0S1RcWkgt9+rZ5DVbLRBQL5bb09IzdKtValRhz/XEcNcaLQSRMixerd8cmOscfe2dkMQbR
JzVXfzn1SCb/EGTHDkoo5DVwnjsyQo8TQx3Rb6hRy05zMq/ML09X5mhrQqEkHckHb8Um/KERsSsZ
MW/XqQM5c4jTZK5Z9yRoEIC3iqFh/eErHdo6u1c2/hSyzyG+nimgCv/EhdqxFZqOVbIb6TEdpsr3
oFD0sdvs7aOKEsj0pVajHb0x4x/MQK94rfeX+La8CQwMDpbLYKgidWBCBta54ebyvKGLfi2iC0QU
tOXzmS5Jykd4337/FxjHY8PnpOYVjHV521XFjZSCmx6y7s0iCjvU5P93cr35ATjxzfes2wyIoA0g
EZznMcUe2x5c1SPmEaNP+mFixiPITXdKGpkcDxOwTKlSNVDCs3FwFoLoVZcRF/YYKJ30y9oRFhQU
VrAOqxdTYLORJOgG2P7Q/xULGJk3JJGKXWBNg1kDb8mhU5hqfbr/nC2xhddY8spNYEaGzncT5jz2
PdOUWeneGjeE/axjBfx0FNShEv0ajhNfVqznVfePFsfeq9jgghVLft4a+2dda+ONTFcLQeN+md6n
8gXrMsCjERd7808/poGUmdLq79IPasb4meIlcbUJje9tynU0XoHJIG0GjqBIp3qhgr5NxXekcBau
0R7pqGh7H+xNyHtnnOKgASR+sCc+khGNG5sljmVtFP6PiA59yeiA//stigV55ZlU7GiuRTuEr59O
QL7EDGrSviG9iOiSrDD1OwAulb0KsMo7Yn1/A/nbTHCeWxeS9rSxeAmoolqTKeC3fiZqePznwddq
Iqxiub+Sk7oTeJfYCVVjuzB7tSJbYYokESUlG1/y7BjAYfiD9F404LPBN4YZXMQSTrZ9P3UDGBAI
EuzwQ9pNaNswFiT8YVksmD7IVQxd9JPDnYL38GvuyIDj/TsfWmcPLiNjyNHnSfqBgerOzEZUF0UE
rsXZB2K29sr+3hOPxgw6MvRUqeIWZLaiVA3wPexpjtHUBVLocuJyYu/4cf+rqKJOIQFgMYmChQ3Q
D5mS0kft2v3YyDn96gazVowmNtk8DsiXKUg7HSjpkwyTZrv6mgNXgvZhnul3U14jsPgk9MisnPRa
Gc6/jWrWZanoMHMpAvzF0RwD8zaQqm3TVr1WzJ+id50WqY1D05cNKnYNjb7hQ8DUlz+FUMPwct3a
hpAKVfFEQsYys9r1Kjk0CfeQPUsRyGEvRbszkvuq5EPKkbp40+Hs7SrmDqt5hatmAj60Eld0WeXl
XbXr/DULtOrLNGfi+qf7gBujxmoPNPx9ANeIvyYBXapKT1HyIUE3zyz0aC71n2XuuEKzr5nmIVSi
ad7X3cYFLaqBKxAALN6sf+Np29lTNiyUJum6YfLZjqFf1/ozUOvA7gv43cbgN4Psgbu0CTLHa18T
p+sXBMoB9N7mDmkJk4BhrxodJQimcT3/enUEbvWqG2ISyqAm4fNPeLR+2WFH+8YOsiwwnwBLn2o7
IlwqYTUMqZ2gk9TYRghPxEZ60xJnhf0ULPK68PZX+Yqi8mFXHeq4LB8fMg/K7sqXUICPwQC20d4Y
3f0ejdXW/845UlnYlnh6nr2OITy8IRBoRw90ogRw+kjUe2BB7OstI+3sykP1yIB0q5s96cef9W2J
2ZVtca5JQOeTVhrkcb8wiShocxuJGMSKlyaqCr+0/A34ktMdP9onogYVlrFmMHvrf2UiyIvZZN0A
Yug8UTtvuGE4wq6W43xszLKcybCZZoXkjiP+8cedEIrwoaioMvL2RqdW0SnOkL3flnqfbHJap9VL
3/TUoEyhmxudxzyfZWVA246gfrJ+bhTdvniPYhLSifygQO4WUrIx7TxzphbHFOTLJNLq+yPrPtnM
V0NN3q8UUeJQNXb3swDqLozikv0bDuSEafnasA6ssaFiWmuimc3J05MoXiVwU+1XUvCLjkTXEebd
YPbTAe91gvc94PQ/X1AuSUhJxyflO123zEfGI+WorY7DCb8yCgU4739LYpQD2vl+CxBE+e7KyLtM
8tR1fEDg/eBywexmcS4lV3i/TcATvTihTCmLRmoNCWWDzDG2nAHySmlV10mEaB2AqpxF8pdUIjXI
tMkUs3ZgVUnRuU0uOynReSAVB5kNLjPFkrQ86yQ4p882rYLUKhEVL1YvkAklZK5k4Tbe0a9rJ9Db
O0L+9/Ecik9uSOzcQSVG4LGrNBKBrNwTuT6bXe44GRqhq65luBF43Op38ByiAI+ZfWeBVchlFsfm
1Vd9mLcErJ8J8iLR8guuayjrialiHLdz7OktRXcqdi5d0C9bNv6Oo+2uY/tl+aCOKCJBalgMVCq9
vpTzkI+MQFXQAIyqCh2HNH4P8bUC98Qi0FgvEzPucq6Nu/rMKzBZERYWvKh2L/Ii9kPW9JyFFKMc
d5yOmcz7rxEp59r33sWu3D3ZILCXQQ9V2QBDfNXTQqgmr/H//G1DgqDnGWLttTZzs9GZ2oRalSB/
gD4UQZ4MieI9gscq8sOw2xrrwWdWrDh5dzyWemZu981FIL1Iu/a63BQuNIzgnXQuiN4rTNFg6nHm
JXzbRHzVvD2Yxbg8uq5Czsuv+l5k42Upp9cAWFf0Ji7oLe5BZ/obRY7nxIjBMXDwmbDY002F3wp3
KzXQnL5EAuG8L7ZQAHwAg3v0a97QyLg/KVAc7GqcFvrOWbSgF5lzMeMPVA8dy0algaKNOAGieTZY
IqdOvsfiVM4Am05Vto1MR5M82x19lqDtG0mGTAFiqgGjxGP6mGM3uqmXiCLelKE00BqRjkHKJgUM
SeuOnm5nAKmxVMBWOaJ9tDYUvpwt39bR0ixGOK9CkBVIXLorKd9SodIaygTfpaq6ARw+VUbXgHHH
7kwKAPMUvTLVmPt7B6/sO9LW1/0ytpZyDmUwVYMlNzPCYvL0meBpm43if3+8jsYNrSN+LXYBf0nl
iM6z1nbpD2aMZ7YaPDO8D29auSXGNeSZjVrerJvFXp4/vUYUIhzC9Tbs1iP7pNrdouoDcEK0pqyt
CtqeKH689+WZVEiv7h4gICeDo+NLQTJ4JRfTPhV7I9c/j2dHBuMTxFefHfaFYQLaHOzPg2mOc22G
9fwbX22kMMG0KPdHQq8dR6sOqwjyCVo3KmI/DCx/T8ES1uubVflGMgUnR5n7qwwe4fflsHwbbkuH
VkdTPqnykIPt4CH/sUeLXXOQo624UzA5i6BtvUOmTQAXqQOtK1i8+Q5Uhk2Ly0UjUTxwUloTtgS6
j1ihmXOE2zJ/itWfb9PDJO04EdA0fKJzRVtSdz/Vi7F2dl1FIREGEWxz0xFDV7ErPiASt/Vai6sL
DZvj2Ol07+jw+erEBxxxtRgTD7l4qABQmSMTFjNsd1PF0JO6uzvoMLc7dXXDlh3XwshXTMZr9v4s
0Ku5K1fpUqIB2kKSUO6L38AEnyeJJzq3OpY6WBjkK6Ib0UrBvhfV7x0rvs+tlWVzhEXFjyNyIRaC
yVSRPjabW/Yor3ZyWpCPOaNT2eKPdHI2GMagU0Ju/c3WOB/lUfVazXgcyyZc6sHDWK/LOb9z7zz9
kDNUOy8H5HKha4+XZaM3oXWA2Fw1u+7NHaZHISPDXNFQLTegbnq81/dmHyCp0WQOGaCc3h7vnZ8+
j/hXmaX/cGhGug1g0oFsdTaRmuULtuVWX3ExC7uL0xmXYGahVWe+FITJJsWIBBPBi+BYArAavxfv
q3VkH5ia9uAhApHWQ2Gg8capvr9KeG5F4hGPUe1666dzBAlND5gSzyu+WJf6KppXu4sKwJj+Cou7
zBe7QQOd/1B1ThOFjmfOWHBR8a7qaV3KfH9Lxdwh529dWeUU+xunEEQg+kg0jxBZiG09IyejxOyQ
dS8pYfOvvTbHrBD/zWla2UUSGCktgh3myydnHQf4qvD/wpoTKblXh3YaCkWgvFnXJuHKy6davheh
UrjlnAQugX2FffUJFz18yARQC6oXVfCpLZRdRkqn26SDUHn7vPHDDsao2dqaUsl8TdMPPKQESt1i
Wz7q3Pu7b1ryiWyHxUZTAwfBHtEcSg1pIenfOqdJD18NldwwypyUc4e2FzyK2d2Ga39Gac91UQ7R
FPbWO0nDeE1KS0L+8VDx84V16n+GJ+srv9pJxpfRp5bYHUABU7ejlUi0OE9dmRUIxCBu3SEqRkIQ
Oe7KRame/+FWkrTWwysEWsVFelBQ+A473ljwq1odGmrdoHiuu8zVVj2QdLLhEal2HQHg815KRqGt
bD8PuNFH5hD0Z+vDrqS9Bp9WbMyZ15ojY86exYVddnSFnvRaHbQdS7WdIkCwn9z0D6EeWZ8v7oCx
1u/TsR3Ux9MUuYM/RsvxUx1v+XDs0UMz+Xg0ix+NWqIbqXqG+RUJFM/8MdK8Ho0tuChs7lT+bfVh
Ih4c6pxMwrBO3QQFBBa9yN+38ss7o5ke/+I12g+QPXN0OdI3hP/nREkLYoHPXV7UcfiRjDHNBGr7
WYgM36NJMMGJnFPtja5r4ij6JAYKKkImcF/7qjs/oT3z2eM9jLxAOuwlJjJPL1DRCJOsokpkMdfQ
qh8Ql4m4m0BfcEer3cP4k4plAVJ4q3IAfQHMZVr1X5Sq046HtQGXmKR/fABkvzTTDM/evHD+M/Y3
FneR2Hju0Ufi36yDUYQKGcLtIPrpalpjuqivmvTZ6cdK5CgnT/YO4serxx+ppmP2U5Fx4pgMWyUD
WoGS9vaCC25q8k1BWy+thz47fOwwcQnCVwRhannboJ6Q08sTFPrB5MCK/ulQcZR6hW0KSLnxovuG
Uc+Y0kUKr0JO4+qqy2AkTSHbjC7BDUP5OkekBvIDHykFwrj057IYBimpHc5R8OvbfK35UsFbWWTl
zzQbDWzN+L2wnLkSPhEwStH6fpXwLmfdlt22Kxl6l8d8ndWQ2qxkUL0CVIld/gEtaHekrzOFK3Qo
+dxZSvA5oK2ejJG2IwYEz860ZxeDt5d54vrWXjnxYoHs9BVk84B2agvITu+CE8QfQjOLvRaFk59U
eCui+y7XPeimSxqQOVf7474TCdJw6uUPieATMoPxc/c9dJbjmHXCx1wB3rsBvGxwv0cJfpzSCv5J
R++vcKIm8xc4/KGz+5c7i1114QLEEJDeCuWs4UB+cZPbYs+3H2CrRc9fEQrazGCpedeUNINAIJU2
rFGnnhhAzvuKu0fUTCuCxmCQLM9FvNoVURWX3CkPZC1L5hm7GCgYnfTG5CHTFcAil07bqS5NVQHR
7Hh7KnWfsn87B1d2R6aF75UZNobS7ulofJXYv4WCsKZSy9uSfB/P9rPBgIkLoLNA186vcQEJMpbW
pnrARniiljDS7Snsp8xRDgPBOmOPEZdC1Ws78Vm3U6DBQ3Bc8GY4q4wWgXuq92gy22XK0uaozCl9
1cXz8N/el0e80IHncZ8YnMY729W4thLefdL6gdjlXYzG0LaeTsn4lfy0dDHqQY1gcXI3yBazYanA
Mq+CN4QWXEh+lm/T9oqMVvbVpRRpQWEDkAuxT4VPjmqrlx4iGYJAPajwCWLiDhPhdwI/j0tLMDsB
+LZ7qS2dO+hw6tTtkHIqRN3eDrKjTYH9/RnBett53r7fmMDp8rjcVDDCeD3C9wezeYXirfMv2smb
OurP1QqihR0Buf066XcaDRDSOve1+0JG1uOatbRsTiBOUxol5YSxPeigJhaezwZZvNBXdrKI852j
rYhUrSsZBFB90Bc5ANv66HcvYJqxwBSnK0lU2DF4nCi3IdcGLC9/aTsdtnpOSZ368iCtIVlMXA12
LAmP3uxpbcGgz5UxrISMXVOYe3kzyS6ukN8xoRFPZ1hNjW5rCZFOMCow/CNBaZmArXjT5Q0Yig65
Nb6qXi6TNg12HwlOjI+EOj7+he4/PBt/1SXiJKxEbA1Kud3EZNy4D0NZwCF5/HmghYFgqC+MYebI
Ql/TGNUEY4cYHdakowMqBaBBti5AwtNqwTVwey8AMML/BQTev8To09h7zR0b7/hHTNAalXbpCXto
ibnotAud63pAtGxpejY0ZhMb9efkh/EJyj6ri50jbxLfcRaI+/Z0X0ZiV4Z5Msnau4/RfOsVr3/7
n/hAdJQX4yCZ71mXWwMcd3jJHrVY3fqF19TiPLSY6ptZeQYDFCUwZo3XLD/TZIUdUPfs4QTlUDER
sG1gLQIOgUp9rAHWdsNrKrOyKZwryxVlLQ2cnnsNJijwWp2LEZZp80DAoGWZWDJs+E6VLl2S+TJw
jLgYDfeVDSPvd1Ks8au8sXCzs8jSFJ6Te4Ync/0mcyStNccH4evZ2scuO1A7lz6xqr6lt6FlXWQp
Ehbvr0gC935+E66dPUo7jQdZ7eDQDT4V02gdPUjR9ss+xmgXsXJ022fTaWG4bdcQccKjxywCxQVO
06EDssLkjBWrz18go/b+3i9B2gIu4DcDGZCjM+LupTd4VhZznvBW7NphHY21qEqPIkOF2M0IjlfZ
ZE0r2kjMY0mr1z77vX+DffnzRX+a27vjlZX9qVYsdZmksjwtGLljI+Edxe7d7SeTpfyN09Vm7EWv
NbYu5pZ1HSejhBzWhm3/GHCdXfCyu9ySHlWs/egQ49wwEIxSaFD5D/F2aWqbGr5FvGDFxSrOAgRL
Hnu4rjYRiC1BQAoAg5kZeZMszi9IH3zus32eFGyEB/ivM/y/5kn6NaDV0WgdVl0tmTWcPZzj43Z9
PW0M4Oeu/nGnw12z8C79qFMbT1Yh4S9kfRCFtLEecyQiAZcLzCTgofVW6XR9EuxZcNzpGT7Z0amU
CKz0WjKGSwSwLlbLl8J9Li6AUUXz9bYCZ7HL6mmQZMiGZC2rELLI2ZVJKU16WXfueA83m4xO9s2Q
AkUjZk7AE3wVkQGV0MTz/AcCL5O//zW7UMGCWw3kwxBX4Of3g77KTLTlN8Ettd7XKmgoLshjW6ju
9IsLaHjQHkn5kmcymyEYOHzHR1vp2uEoq49du4IhiRu+gd4pQWCjg168nZDs3y4qbFTnN83ptOO3
O15ChT4S0e31HixpAiPwWl5Ah6qDx2DIBC2fcDVmUTID/5QP++iXfMeJq99IAaLI3d1ofAz6aD4M
7i4UyXY8pYtyUutg1NQk7X6ImrSScT3aswYsKYDxF9Wq7DOwUM0mBWDTZZ58QzgegRNfWZnzUeUZ
xo+GBLLypiIiowVhC53x3kssWZd9ZLXePsQ2WThgpmiZ8o95IDTq1nGp9ANjXNxbCgjN9uokWqT2
+/IhszZprFX081pd05EzOpW1F1jn5fNXaFsJwqsrcignI9B94dI4Ul330ODctnj+HJ6iCc93gDAD
Ej1wk1Jb46mcTmC58smcOIfvf3GC031v+o1DYy3mrj1Rlq4BkOp/9Cf1bIsiMDap8OEe2ai+6v94
c0V7MI4cceIKZw9VnGNFeP19MlJ1G6odmb0KVQdQhbDQ0bBztQmkqdpIr+3zQVwFZ43Aod/kQcyd
yXfAYqH1Yz68X0004rc3nZXdu8Lpf+7b5x1pxV3Jh4vvRmxb2F0hEA9GED6BU1VPkdr5JD3l7rbb
3flPjBXA7ho7cqfHeLeCbMbVeCw9lov1OgxgqKdzgWOfKUxSjzDiUP7hlBgaP/Ul6OJvB973JIOX
1myHRXfPJ8dT0UqqOwlR4G7ASnUm8QVNl+egkF/ghWeZfzJyPkjOCj8QuoUp9NLO3ZUTSnAmG5b6
UuulF7CmYWZlF3CrRSkVpC2ZqCSLAef9yr02Ss3HjntgT32eSWZ+5/y0/dxgDcrtZ2LkNcIk/iTL
VATRDBFgQOxob9+GvawnMk6GMIUAEUw9YpSMBfAKboqKlyNZoHve0F96ezMKbWWypgvvFLB19ZCZ
ZnlNna2GQ7aZGgMYpAWXKnUTRbDumnmrQgcuEOM4RUqsZyjdr2LRrzq40uohdUoc/KYETUqzNnTr
EnuOoDn9xYYAwOBIG4hJSUhyLJ3+LZMqDGBHtN3ox447xJS4zuK1Siut5FCnzZo/V+eD0VJ1j1dY
CvlT3Ks7BhssuWgevadtO5d4mQuKef/xOWoTdi1oiGipDunYPgWmDo9IJlGEHxDPKehk1dIpiX2y
1lso0Yg9/ew9uZFEkwXUn/haZfhIuMuHN/e1VD7aMzU0gALCvFrrHwR4raCuGjGJbWmaAgYz43vG
5J2xuGodox9kMKePT4mPFiMGHNbfCpsAP7W1qvJuavSEsJ+kWruzANiroYx3Er+YLjYK+LsKHqTE
+E/34JbGudDc7fdwO4OcDFg1TUVjwMagt0q3C3MbORsQuGZpxZPgolXzsSaZs5XOEIRJMpLrbVpE
S73A/kH0bakCkKg0JXwCo3k7JsRE4W9z7yb+VtsOYrvHB6YS0UBe45OTmpz8QX5I/32T449IeHnQ
efltwYf7H1sXx8MrVYEDij8GPwlvXr8R6IFjK4+oTq2KaGiSPLrHnUQLMvxF3KZEa+zyM8s0eiM9
50hg6Ibq2EOywmHf2gItmZdLyk8qWoYj0wzA6BN8q6ultxa/SFo7CKV42PUDBR9yNdlfbgRd2Fbm
dm6t3R9zoF9IFGEWKx7Zm49uNGaR6D4gxXwRlECWzQn7eNVUaeUqzp/vnsNwPUDk7Eo3E9I8H6Ze
OYnyaiEvIXfzmLS1Nx9lCXdwdwQzQNoYxDpD6tmfYdXHhPVVmPTervbRYLyqj65KBFMy4tf0mNXJ
wAu6bImHUanFMcjkpgYhXZrXHlkmt56OqxbPTsSB7urYBBSC58Bb0BfCVTv66FRdr6B0Bd5fvYWI
HT55qtXwaOusRbOMmdG25n3rIhfpEaO+AEKIYiHSfAebqkFgmWpxYPl9JqBJmJlvCQkb/x0+3RDV
RAX1CAzmgeVHnchxSM271Ey7P4LhYUlnETR+GdmJ7RZQAbIBwaA3PJFXie7TqQtn7+/NlpaUWlAL
unxjE2Fglk+dp1ku/+4dKT6T8g4kDjGCPZ9+Unch/jGdkLkUOyvM4bW7vmwnmvZfgLbJVyaZDgIJ
lD3vjqCeX2/oQqU1sMArm6UntQqcVMxaFNJdx9BMt51/U5Q3jJG0cZsRqovfjdkKKX5hKAcMXBHJ
tWbhEXF1V5py567Z0EFOwG2d2oRe7Xcn2+8YZ32Rs8mXvIVt3ROukNyOtMKLMNVQinhEC5maJHRE
2tScWhgSYWYcGT7bPjZxhJMRvGEkzN0haGWDJjR5moAT+cyuRbS9koPpxLEIey1lGET6xUeljbZi
dw7LNE5SyAQ2ZgkHPkV1kUnXOz1xBtsBNzu31HNPGbOAF4aTN0cKiEqSj4PJoJ4nbYoXnBV/0PIP
3cEAJ500/b0QzXUXyhNDogRH4thmS92uUw/z15jcL5r2RyI2H+KyfZBIg3xvn5bqTpXQBMUo1Eyk
dQxCz77h3PgHvY9RWC6zpvyufwECaioljOgyj1bEQC0VT7bm8U+R0x1I/MT7V29O1Ju4QbC8SdaE
X6SC257KbXol4h6dW6CEApm+tneDJmV6mIbXhKypYSxCWr/OvhGy24GP3qVwtKXpMkT7xKDNieKG
r1rigwHNLjEWvc+JQimja89j86vvTTvb+mrMEkAx9dGrzZYTB7ndrt863R4E/KxWpkHtoRaV5OTr
CrtpPs5Ia6igjlzr1oLoOKaTY9HvYCa5/chTChgs9U9/PruXOIthBtK7FGk4r81Ep6PVxs713+Vh
vB7Ji1UuzcKpqbdn5ytzNu94U8/6VzyZ5susWtnYXen70S/60zI3ftuyJa5PLuWKLRcRgi3+z5zP
+3KyBlVkvPWHlS2R1O4sPWPVIiugS0dVIZ/0FZLYKz36kOxf7UFOfIaii7GeWnYMBHjfsn18gE0p
KuPZOI3A2kMI+woxJbGV39HYjrEtkomsRj1bnW/mQKtDNN0wFKPv5108I/NEGW6OVh3mp3zFA+qZ
amdKC3d6V1A+KLXbP4JWzRd7XAkKcbK4oivcQ+U4mcNuNXBS/YejBffn+YHDg1uBTAcl0lzvUOVa
hFXXkYoJLVrpMED/fyAPt1sTcStCsLtX5MZddEl6k94FpypSQGkWXNmdbeFPz50jXE2/MvKWbm3D
eQw17AzUeNEv4/RzCEv7RjQl1rOvURUfrmhnzD93i35OdoxX7B4LE9GLbqEJzUW7kT8ZSTbkZhTD
9PLjo8MupBS+ESrT948DL53geR0YLIXXE4w0awbSMFL0NYhbxutuYpKUlf8M3dvdOm8UdZZksDhs
4qrd2pGVZnXnjp2ryTXBG/SvunKktzqkdzt/dshGu6/B85ym5MEsD+FLF5VCtkKN+VPcY7H4X6HO
6KfU87CFwFI4c4oV96/TrbT84hu3iOmAEnog4P8gRIUQ77okrlOBgVuBK198Ore/Bn/Q5B6KMSOm
+sAol7uO7DpWETRysy82j4RrkvoS/M3ClCluNPDao+gfdVcysbqRVO4HopjRnNVNBmfaMOcJAgx0
MrUBY/F2YhhMZ+p6qo2n5+kIzDqcdO8kCkldCnSBMNwuxJzFkQYhluPFg2IIYBTnYa2zzBl0Wd4J
pItB8zA69j71/saC9VsTZLu8+9oOhRXJ4I4p2RUsYvBH2D0l4ZnFnkuJsxuFDllUyNhM9H/6UQqA
f/HPfD71eyjUk9HXZ2ZTkcGavVVdZMkW3xb8V2spnPKn79GSp1toyvba505GCULrdHXD87oH7B4F
2ZQF70mtqqJzRIq5ph/BKOuNX/5iWV0TQrKfOl2XpeOjZk1Tri0RBSSC8AG7Uc6coTlZlx/xUJDx
I6oteltjD+xHPHdvBZMorQBhURFq6Q2rjt8G2ohIcWREuTdurLlI9h/b3k+GCSCWGfnFJ/oNQtsZ
FpgyUBRpdPrqSDmnFlXnZSUh0pgvb+eyGz1MZ6DE0REW5iEY61lXAWJY4j+0aD/ivsLvjRd+H2aF
IMru1qaNY/MODuOHOCUb95ekSgzQhWLSwEzyA57dC5NbvieYw0KR8av3cNvT+s2ie9FbckvbspX5
OAzpoeiZYI/ckex5mN9KT2NthPzm5/bmcmFebETQ64VKy4PaZey0F2ZEucQ2V8+SChV31iU/aYLm
q/EYaSsjfaW5fsT/cNUkcQAoW4F6zusWCvHWvFsj6Zp2OA3ruPIfZMwQgbvtXnOXjXRPEvOV/4fJ
sZfhGFWgyP9hVL/vJlGZ02J1qFlThb7RLlIMjLci5NJv2UIfWPfOEGNtP6cSK5d9BwoehSPPWg55
3U713iCg8QXTvpHxtMD1XzEAjiC89zKc+27N5MD48OpxPcWl/gsdgOl7DYs6CNo+Ao+gIIJ9bhMg
Dnqg+Oe6buWqoK/62IaR2G8lxXa1juFYomxkN6txa/pDhe6SI8jUPCwx7rZgwb4R/akeb6IZZpIe
fEN+cPVicmcSQn9TOVGR4XAmYuV7DDD5XDWklq2bXaqZ57a2mR7i9Oi0ASnJg5/uw5Z8JA9WMjXJ
QtGX2tPrd34LfFOP7JTS0dBHOOHhtUkeE6e+RmSqqbZMrdAUvlUIEqa1eBbwB6phoXS6DEL1NSKa
csgwW8uMsbQ6fFWvTxCyzqmmLWTDWzSRzaCvJ1RX+mKkvl45CLfVsvNcBvIfG2QpnE6vrHB8ogbK
mIWbJi0QNCjDjuoI/dR5+hIy8odkLJMc0O6qwBWgfiK7YMe0Ez0nnc6CB+oThwb0c2+aJf2THtn6
w+iZ9Pi3pPLep1Bd+X0+TmAEJXA2UmFYRkG4jjK0I8szzCHyZM3pu9hrxnioB6yHHz6fTCtMJSBd
7Z32WQiEsyd2yiBu+InIMPSqlQfu76HBfB4EJWs20TqFTIDeTwK9Cdt+3LBKSLdluxFZ7c2jyJZD
wmZPUlwBcqb27rq6HZdpeo48N52b83q/8sODiZYFMn7JZTalB3SXYTeiwOwborqiih5uC6tXdTOy
lF897pe1gIk0JJ6RaYTO52cVpDa5QjOd7uzXDn1ugzLgsjtkHeEFjpp5xpw5UfiYX4iYrRMcrPAe
u96zTgQGVdhjXoZJRfUiZ+ihABzs+P0voig8VV16MrpBurmaiJSroX75Vh37bj10qoH444NeZHl8
HReXD8ACTEGS4EmdOo+9OsB4zmXOKzanJH0UP2XXUZZPQ/3qjggiujaMRxdfg/H7/SsgYm0bs4YU
EtRHwjQ0VQoEwDOczKxMEbWztXa0n4HELDIdsyTfNIPOMrOmtMFeUh1VqzShq+ppmU41IcJXFeMa
l+GuPJdGacACctJGl/iPbJjV8zYpwA6ej/0vxd9hurQi4rBA0Yp1ckG2zTHOKG2fN1SR+0WlF4p6
zhlJpEfsv/VqDIQZzMz5EwNLVPTDk9GEhU+f6rVJ2QgCuvPgIUUsKQn68V70NjfoPNircl3bHF3Y
zV4S6LBwTXNgTCWCg6J2cIW4qrn5nQZLRw6VdZSNeeXYs9zzp1m1SQBZl6tQNejjxRbKAZ6EF829
NmxOrimbJPBPFLef4KJpYa7rLgpOiRfcOeVgvoP94keZPZiWob9cte8yJk/8ZqKlQJc7iu5s8Z7f
gNeg+vKv9UrsjRYddjnjv6XWfhgXzpmBsr2paQg4DL12NgLGj4E7rALz4+gkd6Hv1fW1bjM93kJT
c1zIoBlXGi+WAVebxELnOcEN0rhstSiN1fGVkknYG+zQcs3JxxxW6r3Y8moxlV0TDgV9AOEfPN1B
2aj1nf5OEUREMpX8m7bYN9kqhRWbB6EW32Ds5aqypz63/BLicdzf1BUV6/OpdxvDkilYaSGO+cEQ
8ZvbG4fLqis7eDQ8v0yxgRYMDfZ0gtfd830VVj8RvxVBJjcNHsSik/+clVFwdD0erae5xXGVpByC
Hpkw+CRP7oZrDaV7trhuK091afESTIfnxwKr7iwlZ42IZdSQKPWIn06EqNGOg8gaOdHle+gEO6Dr
s9K0PpvXKNEl4hFOdy7tDrK4KzQQ3RAnJSZDymwvg2n/TodykhML/gBYetmq8ObZgovonxrPrEz+
fImruIGl8ECxzNHiY5t1kL1irJ+O4h7kDJA4SMakyA3b6zPTAd5yiBwHIdEtSVqfs/mkkKb3/CRK
l9DSSwQtb9LsYzanwTrU+KZ1IQiWo7EAvLnUbs1mnqQbPvlZhiS5oMp9MLmdJvbrB2cc+lLNU5q3
TBB2wrv/lnehnv/9GdV15Qf+9Eq/xgH2wUgwva1v611C5X1Iq4IWYh7SNCqShfAJ4sS+NVY9FcJu
c/rq7yPfV/ZiUDnCw0LmxrN0EdlT/etyC3mtKD+bGYYxSj0QyLYtNDBKnulwYjYM5NcSgkW+VNne
tuiFCkAzARGxCJt4PRw11UEhRxzvJdJPwY4Li1bj4eicfujjBf6T3xXh1LSquuCwkQv+BNSPcoMi
PmpXYQ+qc18XHYNLTWB6k3bQrc1eE17KCVuStEbmZQEhE1VfKSVKGwoo0cuoUx627cYtc4Vn6w1h
LP+QtvGRTEK3ucood+h+HinbbB9PclYghL28NNRpw6oP2rsOOMXNr1UaTrzz02h/f1bRwXSUuLmR
yinpRxbCdjXRDC0g2eOVHtd1JXuPh6/OVik+4UdfQ0UhI2XteQ3J1R6p/Aja2yRY+bkVNGg7ahoM
hY/KC8u2RMgGVgT+3roFGahkfBUGpqX0wmEPbrSzAhjYt+l0E8VSo1WKo/3mi/GrkFV+DLbl0zbS
ZEjJScZjqa/hDanBo2IaZ9+FDOMb+MdVZjBGcpaMPrD3iiandQ9OIEPOlQYNZeGPmMEIPQ8EaPUM
MZe3No3olceYoXyCu+bec0xjzfgo5/RgXmw/3MAr8j8jRxgg0iJuyuZgLq6DFP4CnfhV/+CzUQgK
DeACeKyYn0PCXIc3WZTwDPnmR+xuqy5txBoOrRR39BCCZYl/Ts1dvz+IXqm8XNpHe3io+uRX4jHZ
sok+8A3z7hywIjRHiHAJQHUT1SoR/U9hQoNKW3ZmW0zBTpAvdp3v8mCoXE2ithxtIPBEk4IBlZtt
GVYR9s6GIh5JsXetGiIVDncmRceIxDtqmNSRqg6+00ASwGDqtTvZbYJQs9FxdpkDo0ZmdSWSXqui
N4VMRFbs1YCVHH5b1bh2HCG1pWUboH87Vypwd9a05JtARmVabnb8OwTJktfuhCb2+z4u2NhhAmdi
MvfHw3GWrXJQ7R4lA/8gnifK2BFWbRGpMwMU/emPRIJD3wxVP4mSO0+UzpYnomcMVxGEPMxak4iu
sBk8PWFR5e7DRps9Zq7gTe1op0TTdE53ghNYUJh+zhOARSTsZ8PPj0c3OfFhDivHjzovzqXDlXQJ
2FjfS2wyR9SOw7lrpgAJRNwQ41RD231Ymw+btnRG5908T0diqULFv6MV0LSSDihPyxr+zZhAWOhE
exnv0iKY8zjHS5KAOe1g+GStQn99myRKwYC4gUtVlKnZlEMZzzaw7NvKNYO5PYmDL3qiOhWgMvJ5
MRwi0sLy1Chva99hFNAk0E3RmofAd2aGW3uKY8eaIENYiRTLpAWFPC25GiRyRSaKNvV3pT7AVZ3l
7OUYcUJuIpkoFDJBqRwzXWsB5/beDlCIXQztuGWu6kaGBEFqfog4+sT4yPsQF3JzQ+NI5El/gGwp
wD9QDVvEc5uRgNa6Dw5ONhSFjBFJoCjHLBYIpGIw5D19gn3m4NN8o9yZwYADuQs0b+EnK3vrW5WY
5R/9pmnzZpZ8vnuAH9sLkHHOMvAtxo31MlS0Zx8TCkiSZY+aemPWRJNLJoH1mqPtVasfkicWbuKB
6Mpuu98ELgQPzKu/YFuKjXmB6N7mGdLOuViJ6dMkYQeT0CjwRfW1/6nm2yWBxBARinDpZhhK2Zag
pKOTiheIqln5lz74yXdWddNXNuedFNAHCv9TRZx8I4y4h+P2ANhKR0PeyUn3Goyp1LqoHiKHJY2D
XkXT1Z23rk0rfp4y3X1LVmFHsIrz5G5yDUgXRtslB0HM2Jdr4qddtrzwyIdMtgmwYiR1Ee7JwkFL
It4MT112roZBvmKcaBAtYXaI7OTMynSMq17wTaaD9cPGhnGZyUed+kmn+ndIeyDAaxPNRjR8Hfv6
O26ISUFQyh8HsJoVTuKDjDDTLWDhvR4QyUnb3RQU+X+H+5WL9tDcesFALhoSeMkwoGE1zftn1wNF
oYtd5G4FGZCbob1UBUwMMSsbBOu7ANHw4O/WKFwG81A45BhipIpmSzdtlYU9oZnZMqGr4NbYsKyW
R/GSLauRaNU3MaxZw1G3NtZnzbVds2SCZwj05kpH1z4f1ATwSiW1U/6SGgP/lxJyY75L+fRJ5eMS
2y/hCxGRWuNfz9GnKgCf5mEPGqofDbr/+0wRcWVA1y90yLkXpCVHN0mKI1RizTvzVYY88E524W8U
0y5YatuP2/YUu0iLQx6jytOJPCFAV9UoUZCuQwKDbW1uBYB3Mb98CZ4Rz94c+uyUqo5bd0VY+dh5
gwV6FK5nwCps7gEp4DVrxKhZOxYWcbx3kptDMNO+uiGnlYIwnlsJ+BAAc55m21gPvROjQtrzE4Yz
7XXMZHQ5/h4XF5sYHx9dL2SWR5Gu6fHgZdzCOEKzFx7H/Sj1GzaeLLKjQWURzVcnVbT9FqRKqAay
1oXmT8Hv6nkZkpSsAh/f0KYTFKlGLVC6f63XR+A/NB+n+GH9IYVKiO3I2m2brRB+iS2FuZ/df5j2
ARGfFDhZD1EXpQMOJLvTYlKSagFthMrRrGUbBsWBAMHsnQfyRhM/hGhO6WXdSIuf0B+wERE+OEbh
+6oWaWG9hRHWp8o1u3Z5G6s3IJbFPC/TlVZZZVe/Rru+iei18LB/1qphspAhACqog0uXs9daFOl2
HvoT1HEkSRhOqoW75RqLHnQjZxuY7IdcgYzz+MWpWx/wx2J6uT3GVMlxeqm0xBFrDy7OxJR6M1Co
FZg/aTO0OyoQGS/fZdSi2EJSpF58FmCOGgWuc9CEQNTtc0GbiSbB0HNSwwZLs+F7PJ2L7EYfBm9c
qtnsFyv7fFuoD4yjmUuUgQRoCyTBwtY1tz3j8RZak2p74f5G6Cp6jXn9z0MYHPYVmuW/9/Uskkoc
b4kypjUowzNmSdwVPoe1h1LSMsheno/qDQfnCY6+ixpzD+hlhGKupX8R1wLPG0rmV+qbdGYBXizm
pe7zMVW3xD6cd+5NZBn06CccsZOOfv7Vp/jmR/gItmziaKDREnWGXJdBnXtXj7K7dhp1PsK25ng2
3+ivgyXnYnX0//NJeTKf6V2mVs5g8H7mjK+lQv42zkd95dyMhyQigJ0C132V9gbOr1cYcqcgU53U
OVdoo7iBSWtORwcRAqwIayCydQb9CcRKHArVOc/fWVPGL5qFPaGnu0PiM09MUPfGZga/8VSsgjQZ
vTzHb1kf2gt+nDdSeRBgB1Agl22UI38j/j4Kq2GSrTROIR1tPTsJ0HsxN3TqhKgbps1+BIIl++8+
8YPfSMOY0VuiVXSwFYNo2bZRnlzzu2n9bQ1iUB2TX99Z5ZkQqp2WYNoTd2OI8bvSWl9DytYZV2G0
DhIYaikgAVLT6YLuicgCv+yhLQ7MyCbHXr7KDFy4jzo5y2akko1M4zT4S6f0xBFmTuaSAC7Y12cV
/Es/Thwn4h5tX77q6B/tXHEilvLTfVORaw6nYFlqY5loXdlqqkCJqhT6M3MTmbbs3uJzDb4hufT3
vSddWUlUcfdmOga06ZLBMM/pnKTaifWYMWEgtie4lgZlKn3yCjoOw+Hm+edslDiXYifNvZf/wxGs
itSRN9lGMdEDVdhvpx4C7un6Y4ySzK7LoHXcbT3WIm7d8McxK+yVwaC+RbCIw4aSRHePfShlid30
sReSc5pNZqdoCMYWjIkkwg1YXHH8KgR5TMgOz7sJ39+J2txpiZvfiI35+c2rom8iDTqQaiN9QYNW
soQAqPIUb/rcWCD96XNJ6mjSR2kHzYUWTLcc/tOzy6n5096bBlZeKzoAlkCvEDyAylfTam7gIbgL
eOtvYj3Obct1tFPMYrquFqbxe8fViDDWxgKxuO21Ncqr0l4ujgOuIBnbJCmKxAD+dfYlzcH2OWqU
0EG1VGGmXDsSxeyGYyp4KxLuclUYCD42vaCtfvpMXQW4sSwaahC55NN7RiDOpauOL5TY+GHf95LZ
QvWet4rK0cHlqbK3opxAxhaLsyAJONSuH+1GhcUrdKzVFu8aS7jyTWAEtxakvyRHRwT17hux/mSw
IkFagKz1NITbNcolm0PH/xq/RGVifJhhjMr9Cj80UEaycyaNPFziP/jOtHxygvfIQHobyIV1dMkm
1PD8HUeBjDhQzTz7iSqbyH8erhAxsLd+ByQAJsiaaqpuAGv9qbCHuNGnfg7XQtxf8eRHf3ieY97+
1K9axLtI4axdJZZhmHS+m2Ue43nAtOSntmwfKaa+lCGjFXXMwKQ+Yew5lSRT4DgDEQAXfXwS43lx
ZGy6UzCd2Vi6tfq9XjEGkjKRBRaD7gu7OHl7UiUdlQo+xy24QVjGO73uRRs0eo67RZ312WqsVR15
LIzzsggASFwtAdmy9t1UnBV7zrFr41sS6DzI3o88U8dgBIB+Hm66g2vgLmWtCi02V+K/CHuLTqB6
d50GLREziywBa+gjLDmG+V/i9I/zPHMJQhcMFE5CtMANYbJDYvKyj7wydM363GTrHJxN3YAemrR8
Txb2zGYOuF5Z38Omf2qF6s18eQXqziS4flPzoB3UqHDGzBrU6WgnG5FYj/DvJji7WEigaA9kq3yk
wZeIPGMgY79uLTyN+u4JaUr7DFSDBObYwBNQUlS9b6AV94K8+6GGbuGVDDGsj4sYFylX5UfKtJH2
0RxjUcFWxarOZYV3UWju0MtjPze4VpTG+tBw2hKvRfBvxLgUGEn97T2FJK8nVzmP4Ck4yfNJ7WaV
Me8jXPnQe8P+CUZMuK/mxy3axqNcGiUHWT/szhmGxCnITIXqyMnLmmm7B71+NExS+0BcB+bQqazO
p8fsq/wwf0e3Lsj4xQ65YgfbGbYZIAHnJD6fCGZ+OFSMa4JDF+m5lZmFRMQZNDdtE7aogkc1FSgO
cp1aonZvhyvJoluFkXcE/6qOYKqAXJLk9Cf8POhUo2zGeO4CjVCEvO0hYXkWvTiITLWZN5UjknLT
uC/qawpbpY/t78lPyt7IpkTQhd4i2lnqs3U7eChvGQ+MgTC0GMyLbRt8wo+EpunX5swMEHX2Ykm2
Yli2vQmpxCMMiDDZLZgb7Vpa4j/AzGy4YYnfr6EjT8vzjplZUk9SHcQnLBLlXGVx9AnQpC9n4uL9
hm8lfoskuEPhlRGgepw1Q8BLH56kTcKniriq1uMvrfoEpc425iGV7PPn8iC5McyUKeM5gJYYX5Zb
tPgRe+TmKNHXoBoAkfLrQH4ziLAS8CVJASEb8ylEsF5W3y5Iz7YzRsULbaEV4hOprT9FCkU9E/iA
CTCXVsE+zy3ZFxODlROt1kKAfh3vbWAH6Q57ca4OpdWLtbVelsiRvEC24M0KShNSCEpcTES5dcMB
3xDMiXcjqun7xFMpiNv8Qyu+TEVbhGB/gvf+OGluvH+9PvofFx2vRBxUpmwcRpvTrblxMkxuf+25
/bh5P/iRW76iy3ddyx9rNk3H9UGcHeCeLgr7EQlV1w6vgmcOIm86riymVa9STCEFwy7DauLOkgfl
R5PZ5G4wAaao7KNc5YLULMZU7DNZEFY8+yA4ewa9RaBw92pE5Mqet7bskfwYvLwDOTgHXnv5MBix
BdfygFjMoI/lf3nT+fu9/hI9pPSwK7YYkIsHOqiDKV5soTRlT/TLP6cptRJ7oewBQR8S9RXpOkGo
cahWjw4Y1nxJsON0f2Dwi7D71JSljAoARCb8CdE9EU+b+FtztWO3u43SzsfWkD06K3OMBBdbUbmd
QcWaNk3PHU4F1mVAysWolejSlvLUKc7uCH7g6ZBUKjdWTJeejQS1Sjf2Fwq+q0iP5u8aUwKhDqVe
+VuW4fsyi3fZ+Bq24zw45w334z7KH3RC58RkzandZD54fXgkLvv6hhIyGc9wx1UgZFDFLTAoZukF
GwP/sWVzyYK0czP/f6QrszJwxV2JBQDMN2GLXLxwgvySeP/E9PKd351D60LWJKsVfCy8uLAekqAp
P049Zm10RWeER8093JRlYSSC/ULELduUUXZrDmkudul73UU9iC04DoumDOT1Hy9EYun5287Z+mdE
YGHMrnPfE/wMAK5bpG/prnQMicnvlty9LGks8l5Y7VMwGzg1F4C88xGD7RkQiIuqIqxiby3eZ/8B
SNt8ixEl3BZRR3iyJimZzFcXnQ8VHWgHIMIbZ5uDBCWIvZII+6REEKI5wvW8D3Ab5lZppvBqiQ/K
uhKkaQWEiJBbK3S+2Ii8IlqIib2ns3yYz59xO87Nkr0EanicRAIQlUf6hpRvEm2ehW29B5vo+uhA
PSNbHSkMOedoj6sVcxtGMmn+Z70Cae4/UTcApl3dSaSw30+svNiKHIZx2AQIn0hhLRBsWchqmqPQ
SochT9Ibvk6w5HxbWvNu7FzpYC2xuxSUHS6p4WeugsewQmVcHbBOZBOss8apqL9JF/bxknZQHJej
akoEPethrJ69kp2aQN7sCoY8ttoJTmtYsOrOMa2CoUzpsD1/2EI3Cj2DxH4f+actD2REtM2k/A49
C9l8fQ5Kk2oQSkQfocy55qER5+TPw5ZIzGlW5zUVENlro+7fbe1sar9UIKMBoW3vGNVQ5+4+Vylk
iKkFGYV3pyrAv6VK9WDmYGpzjAUS28n+DHgdMJdNWeKfhxXqpkV1lzS9tTBzxAqLwRQcXLgdnGNz
RCfeHlJDwi1PZeH39LMkIcR5+qz380WWPj0WXJHAJySf2qW0wMdb/uwD7HSVzIENFB3zgyK2QxaF
xUQqBCnFuMUx0T+g8ESGxZueMpFM8gb048LAvodLizotPIRLBnPiVAHheCNXTXmvfBDYyUkZursb
2zTBMjinIV/BW4oqlBiJkxg0tT0kCvJnnWXyOzd1vhqzv/94m5tBhNlkp35N70WJxhAzUiwiVD0W
Acek7enQYxkYZs0Yc9Xy1WeVj7HdslYg218qDJp48rI+N/tvza1oqN3ghce4ErPTVZJuCwXHL2+h
oCSOIc6TXDb6rWpBZ/iJKOEOEmLvMjm+zwCzsaEXAHvH7+QXK/v67kYxK1TeW+CZFKTyXLzUGUxW
UZjJNs/lJF4WSGiAeSCUAxZ9fZI1xWO5IkqYMrc2kCj6dP+df3yjFzwYxdNgQG+v6dSOoKbOajBI
mfbU2lxxdGz86xeWpcUL6RDzUjsM7PyX1fsbBI7IAgNjK4mk6+g1qxk0REmV+ADKqi++PlH0pN4z
aWstEy5sqJEi0ImX5/rT44ZeymM7FgAzj31XaAUkLO0AM9gAg1Z/3vvMki1+hOkXvU/1V+OlDFsx
DrS5cGmOedN20xF0TU5IY3R0xyz1gR+dirmI2KxqOfIZsIPLU3xU8U33xl0iEOweH55+e0XZsNaf
elR6g0yHRfc6bKjAwhLJySTXOvq5ADXYeU3o8Yw04iW+v3TPV2zzffJQD/8Ua6Ukeb+oSjVcdYxv
hfHTMS7WI1BVImrTuGBXn/15eLKexwZHp5Lt3Pp+2C90dEhrmjjTaLLLdNxihZ79zkzlO9DjmmnB
JCdkL9qt4o5R7obr5Je94G7xS1OUKM50x+o2s9dbGh2EcjHlVJnampMnp9+zU4KcjQ41fmqxQVZP
HSsfwfeUG6ejwKZxrj+0jgbYZSJ9IUaWRZLX+vGSQLE88pKiT6IuEPPjCbFAVpH0VchSdzfm/kDt
NkEtsAJjR32R1cnMG+WEODnL29C50sCZrwhJKwr3QZ9DyPVXc68N8MaH+6KuNfUhDc4GywRu1khP
mNOUPMNrQ+YkpfjAtjkIS/39y5ZagSYGsEJGRZhy+jx5Up4Bk6PQ3SBSGObG1ymiXteSTr5HOJrM
UdokkFCsJw6ilo9QmmUvt5SW4XnRoE9MMomexZRNdn15iAKjISRtqZ8RN+7m4t8at6LbUWRlFfoB
gzT1V9BQwZ3Te7aWXutD8ZhtyfpApHpIMn+fk6S0d5pX1jyA/jaUkGoYuYo8Q7J3ob7TBexpXEyG
5kEfnzHAFX5DE8Kk99LD8zk2wMQZgLSDLo8gHPWai2sb7SOskoE7wDcIAHSQXfk+UQLlKvgPCUlM
SgJTlbOa8NGGYXu+WVEAeU4EmjGk0emK3HPAnxRMJBZNXIudxXQpILqlD7Mj0hzvivNx/rdMEFrJ
EK3E852oFpjfMMn+CeAMWWEepia0MKnhwtA5ym7ZHjFdhRNg9whBGavB08fkosufSnFJ1j1Z1Lo4
FWYTasXoZgpz068WutSObIkqDpACehz7DiwCPgWzBZnYH2KmHLasHwBXgDTEL1AF7g/owahplSCp
7740Ewb9Z+YOIpI1aVjYEl1qAdzCdTDQFbqK68tcp3fG9HW32+hOaVYQkMQGf0JnnwG2+Z0XQ3G+
nZ4yALwzNZrFJP5Dyurgf75M2SIuceYHXhOvxkc38wu7TR6JMg1aRQ6iqQAIbYIF0TdGu64K4jv6
GFe0MqkrxQmpuztUK/1CP9njkQ/5Ar1cB14KVulI4vvL5riwnrHz7cEmkhN+Pgi8O00Uoo1oDAt6
qNi2be9xUVDn7b8yuw/bXXjr+UxJI85K2FR/rG6pA0vRdOIZztxP88WM6XcV8z7muGczUUMtKvLE
b70YtFII2WCqrrqwt59Isc51qn9CC0pHdUvEH/Z8EPZ1HH+eVVOYdfV+ePJAg+m6x7fdCBQ4UL/g
CbzD6rJiM9u1etSaYo+grwx/Uafg68fpX9fGV9BZLdY/OrnsYklzOLI/KsJyiYja3Egwv4DYB49p
zIRSKuuEraJj1iQ2xSwyDKxb6I4hssdqF/tanB/uVg1e/8KruT2h4cU+hojQow/09MJPfDi5ceK2
WdE9sTJou530BDf9XNHyfBJ3zikNxaVNugeshd41FhgV29uykZojBlK8aeQdKRi/ZBGZcZdd7cgE
5sjbbuOhWnucNoiSb4ohbEoTGr69aPdwTfTBUV0GBMBjdtY1pUfhELRJpG8wOBxiIfZa7rPO9bF3
WUrTraLo4VDvhWykUnpoL8Oih2N4cc75Zvmv/8KYLRJgN9og31XOwDYeJFiXPit6cFKaRWW5d3gc
nzxLzNdGaPZEff52FRRmb6tdr03CO+PRmD/sFlcLuBLcXO3gp3I0d7bUywy/l0mRtUFZLPKF3iRk
F0G3+g0ZD6fhd2wZV3YjB5qBZ35vGGEZrThQpCmssIdZ7WIVThmFPV51CvyHXdrAoNk3OxDeKMxZ
tkmziw9Z9Spa45/WDA/bc3AJ7zXciIjTbl/op+MiOCiThPtp8Uskd4lPoCbVAAJ6oybijAfZsMaZ
7ZUQSl8IoBKyyJzJtB5bpk67J5LZFGJ7dEJKPVIoDPmqCarSNPDthbMVreyRCvOZ3+fhHHIMx4Ai
xTqV58SIJpniVAFezx94BLuKuc0Eso7Xa9Ag8w0xShrNNyvS0pKBzAg7/3GBVJw7YGHXGL60CRRo
548pOeAnKk5Tx4x814byglN53YkZgcaq87INWe5RpbOAaPZToiehhb4whkhkx24GmCkSxYcPtBcb
5xRqMcN7gZO4vN0w0OOoK7n3lMWUTvSi5bhHWAPDKQCZhaPeuSjEfRnwzp2QA5PFZiQhwFsXa6G9
KEIEVZ/5wYiSnQ4LGdGX9KteS2xcVCOMa7KK2dV6TkbttBRVZxLRtC+7yoYPn/hD6hojSch3uea8
YqONzLt+z2eyKRM6blkgnGVb7ZYVZXWWI5RGQnpMpVzVvxvDSTGEFhIu/PF1vTAOVMYNU0ehHDCm
KLbgHN0YN1+kdrnuih9ddBXlfNQT9egayRBAo+fuQgNzVfx8fSKA2tYbIVPBuKTVrquvJQHWahNK
ADhkf+2sYv2Ivbn8xltd5MtyNxg11BqK4ONJvucBGQQwl6lUjI61hdvf8Bc7pvIAf8LqnX0UWiYt
WON1Z7OpYuccB7TwasMSAELvQMCKlkSc4F1ZMcuQxrA8jNIVrGAZfcPVy+gmREIcwzyoLuid+YUz
j2FBXgMfjJjwtt9DAxTrgm6+JvMAqTjX3HZOB6yIwpQdm8Si8+J+vg1zeG/JmS60bPeIJiCGg5NY
/W/+FNMIz0Q7F4WheJwuA8bSpK+7R1WCt/6oUxNl8eBoVUygIi+YbNdkAIyFDPIFv6QEVSCfiihh
W8Gh5HL7Cp+8P8jZi6BQ8UcbQUpUAW++rmGTQ/n0hOee809BwM4Vi4M3jPLQnkkCbL32xNZHtama
U10+L3ZWs5kTg8Zm7CFw8C9Tcrup17YZYOfsgDAmsLLl1tWRv461ILbN3jTf8r1QL7hDbMJVJ5J0
pw0ogdpKMtUq25zp6F6k4UDe6KNuK0N+NU+B5gp7dA2YqyOAoDsn4+Qb1fjM5MpCKs8yKQnIaSFt
dOYTudAxML4KGj8a77Agz57aK4tZvjmfYXDX/MkXu+PzJWAyg5eV6BU2ilSngpHWtGYaTCBsXw2h
LoptPYL3XXe1vSo49a8rRV+fGGtIL/jLvM+0NBQ4NfTr5tLeHd1B4KQANVXWOQQTZHrIRo+LOqAM
fIBT+lrvtqWFgM0rZJJE69AIyNprUeByU7omKA2ZLIdLlBWSg2b0SiYvmY02963CQjw8yUoBnBHG
90xVdy0MpbDzsj0rMfbA07gUDdUHxP3mOFkkuBycw67DItCOvtyQL0CJ4sTMte/6u0/NN2HzO6Ly
O9/rAr/2xPExLpWvjQar0GPuIcdJQU1RQ3E6mrF1UjYMkYvLglWi3TJAQrC7gaNveKsce57IThzB
wAL3OidEmpG8uvd0XVaOR/Ef21/UDrdxLSbaJ8krHkjv4yMLCp+X39KkAn2Vv8+PPjZNKydZbphM
2MueEO7199aI17H3SbnSLdF/ekiCai3IK5+6/BQgwyjJtpJXLU/wOkvqb0sSXa6HzEHm8yuZsmGz
xbXcINzi0ZpgM/lGwTzw5FAnJMzItB7D9IF3ErY9TV1dmiiCXcLEwRzWty1i+FDROO3UffhXjyuQ
OpP+YX+tOXTT/oRb/aD2jcex/4bRUw8gjmCHtiJi1SLMGdtl1AC1YpFceOv9QfkAaqeMFHMmdsR3
X0j8ARFpieLTx6J6QJ/Ir2SgqIIh1FLo1sYm9pPdOJz5FZl5ESsxED/eaCOV8n3piDMOaQkTvK94
M7+4rV/P1FSeB9N6hLayLN9Es1gtnQdypoRC0AkNGKGxuC6oRoy5J2QEfcSKFfQQqPAdA1Ei3bgG
56GSJlMxNqFuK81bDESulfWlZP7BR2hPdeaBTK0/l+0t1xwofgPUE80p9OSs0ojD4pG4bTwFfZh4
iKhx9Nj38QTTP5iI9w/whhQocZY+4J3H81WaLGynrRezoLXIHJAZKCfUZ8KcxTjVfpCdTsjQ8JQK
Nxau6MIahBG2vBSLWZP29Mm0WV+RgTdRjcr2EdRtohzHOQJcjGXTBSU2lZ3xeolvRSdKXjSxOxlx
24hNYeoOvZB5TX6GXNyrG8X4RjeWGLPzb9zy8FtUsnLFsjM1VtxVSDlE42TaCu4cDBFZSlkgZQ01
wEWH/6KBt35xRtDdNz/TlDdokOooMLQ7XzOOEcoMLH7pZfS8TO6nFY5pCNyB6t/Puuh+wRMjwj4w
uWeA+LVgh/Njz7E5o8ChU9B3qpPE5W2Fa5lIrOPEV11RXrvp9ad3Q66KISW1zXczqsXxDodREZuS
AbSrma7N/ZBaBOmsqLuvb4djFnSP/QdiWwzZ3/MiteqHwMvqVEA41etmEO1khstAXaocXnkH1aAi
Fbei5caLIhOaJJ8u3D8OnNBSiiyhgRHyqwOcbZ/r8GOrK6E/yo35R5KOcfjeTbbavNWVLPonSpw8
cE7kharsiiTsnqs/XSUw6k+fVUuzVFLFmBnFRNwJ6OIl8lLwPdAtpqYBUgRlJrOx8u56JRu+oyi8
uP9w/b/BpNsnKLKrP4ztHgatJPo5X1kQ4bV72/f3SD2ErFOKG7i8YDlCnHRy+aIfJdaDmSYH9aws
A/6kXCxWUChWkC5JNcjb6NtvHtfsv21fkasmYs0LQM38fayD6YwS6W3fxmnQbkJpAY3vxBTOZp36
6yctfWvhUXZe5EryghxWP/SZC/D0AEAeZc4SYdg7//Fb1OjHdlRUSIXxuHiDmtjTUyvTF2M+pnmi
Cr0szJ9sgbnk+7cQ9iBP558vGDkFZDD9DbHMeZamyzdDBMwkBxzzAEDV/jJvPJEDmr6b530UKKxH
RCUIB6CStY9fPMJXCTn5CTQM2XdnSmB4I3mjzOhksi/tjcoEgxgwLt+bKjp5R92kHAjRYPYZx+GL
BsWAVWmKa8yXfK5pHToX1MhCcCh0DZeJta1tvmuDiQbVEAKNyrHisEWu5tWaF1ZdYz8i5MTL0KLY
7ucspyfvyC/DmKhP8DXxW/x6UDU2UCvxNwfqL/bEt+PwgnkWWdEb7ElHe1C0vd9JD88C4TvWU7+s
nb8cS6yk/MxEql6l7XS5JSNaLbyvOoJAYd4L85s9z/fH0Qopl8EiCtBwh+O404yfZSyVNQ3cO8Rq
Ju1OM+OvUCb6x4n/m6rth6Gy4BvBz/AexEUY0ZeNVQxo/PCSdZaGf9EhikzyLdCPVyHU5KigtiI+
Gl8uXBm+cvJgSaJ4PduEzgwZ4tKaGaqWj/KubBC7gCyR6hDF20vJeHbFzauwI5kOXkGs4a7tGjEf
OY6GqhdAcMmm+Lz48SgEDdUeS3IakUKu0bMrIvi12Slr+mWE6yDNsh8lYrlEKzWJu+Fs+SeokmrZ
ZNgnPE/1vYdYrcxRUuoeIaPhOCKBVBOVg+TInzy60ZOaywO4HgXbd+IMmASrLbqB51B9e/yBgFJZ
Tcu9lzAc17pFTc6p59rdaDOUTkgFyarmffgC4YxiTg3UVaGISGq52oGIExyw8Ykp55SecT8QzpEG
UOfyTiaT5blSMKebuKEDraRbD9FTDPFqkFgJb+BpcboLi+ZzZpkZ1Ypu6hdGhxijHLRq/fkePZ0X
lKX8VWysav5EJKQpu26UUKenjw5CS48VtKXSLZheeFx5yOqDFn92gipH/pi3VWtAbjdJG8sqO25W
UR2BT02RovsnNZWtMnonxlSie+/xcNSjqSkJ/S/qJlWcRq20d6O2DBCg4O0p1B4p39PVCR6DDua8
onRtwTYQErhiIa/MCehnOIAjNXwxffbRz/tBRaM3rn31wzmFcuqTzC8Zrx0itKUpYnJ2SrEnH9eb
erikDnIRWb5e90hVAnpOF8YqwD1989aE1kOi3YHfaSys9D9bEj18O/YdzAQERYfOE1pvTOJSpKWB
XA38iGSH6iFCKHvBxK2u+SSE6s7FBJqRdgtgWvxxZyyN8AhzhjTsL0O6mlGlx0WntK2hGpTa0kKm
V6lCVgTahPH5C2h+zu7JncoSgZDUua5eOx9ggTptORP1vl1TEgHTMow+VrvsFf0cnIuLpqvxLYhw
PvN0bHkrjLDP6RIFb7ePjKm+TYTwemHSnR/G8x6VjG2IVGihd45PFuxY5Sx1G8fCOZzo6EW1n3aI
v6/CrictL3m4u29IWHnRuKjLY/GBKye5lPfrk1WrrZv4LLI8Ov7X0fHyXDteyjeaNcTeq60mqauY
fFqjgtN3y0BQ6UC5y7EHayH5YqA8s7asxmGcWG21ZpRzfsJM31/d3+8TmwC4uriwB/VjvSmObzMh
LM+VfUAUfJja5uzKz6CZ7LsXk7gjjztsNWB9IUCsL6XTBhZcoXO5yiYOIQT71K1cZV4De5tUgPF+
ufrCcml2/EQRlk2q5pNAP6D9FpyQr983TmmgiYFripsFU0WSvDUS5u2mT/4LdXAIZgcnJbpdhGxi
7LrRNS4CsoOxvkuVbjZQAYnAg6JB0CezRRWCb7ihWxXlWOUE4HdFbt6gV9UdD9ySpP2qzwozF7lx
fyslusKQXeYudxIoOysjabWIOIZbLp1PBkJ8JZLhNP+rVVhitQ9llT8Qe7AGAE/vQN2VoHEvXvrO
A7CH4t3XZzJpdP3goL/KlC7rebN3PE79Q5iNWK8yUicEIOUEcx8RQdNaHbsU86bpnZgIipeBjwCp
qDYTDQQ/75y75EiVti3TX+JHHxb7cQcvbdKqvNcO+NoHNzh8GblxCH3MQA7WtSOV1MTh8Vk5K9+Z
P3ftZ2giCfSt/+BKDv18zEuYVFxecFRm9M32Fz/yDD98lR2AzZ5+CdBkIo/vPupzHkwL9tmu1iBY
khK1D9M9FVoI0f3umpptKxAmMzsJfHl09GVRTw4HJyVv9374skUx8+qB1UZyhtdoppg9HHUelu34
Y4T13XyNLkqO62XeBP11f71DZVdm8CmfBZotGtgP/rOTP+8fL2TMYup/O8lnVn0rhAJdaKVh/AMd
ccP13sPOwk3ceti+sx39TdnDEGTlUYVzD36BuZCVip5HZNnjr+WJ3THFJRar2aCvjpRbTYL5//Im
M9ljfZjgm7ZpkX2EbLk8GzfHaIqZ2KITXlRZWon2fliN/QupxE6xGybFCZxjq8yBK8DCXHE4Ilfj
VAQmTpjVoyWnKyWUkeaf7d/SRlDwuMXHcxDTJ4MUXM7jFwteSp0amRuhciI71U8VVULPSzhmcWm5
cu95uws361BO78NbzF+1AHCtNfLslH39QlIIY2XnkOiDwGDrRAS/tIN21lrnFUmb2M3zuflgjA4s
vhDJC2nRMbqT1OJhMa0Ccc53/U6UVwliP5AzjIPn4KMgdLi047dIybzCYrkAD+nBeAa+YkTCI0/x
+k1sF+7CrytU2yTYwWyzBQwXQvxTfrf3i3vkJWB1KpUxJRXTQWP0iVOuEY7VL2knkHVFFAuptiAS
CJxPYMqqBh70+n+mw2BiGIZI4yophNN2L5OWCelYqTp0V/zmSgTl0GkbqIfD8Plkr8/8lwOs+IPd
OB8LJqBPaLlyfXIvUHyia1a39GDXTU0rDT0lAEetspQ7vn81/Mi1Qj2BQyWI6rxyKG+M764vN+hh
LYkv0x3xOQ9+a5mMz2I3J5fN2cIYHz0F6K/AGhLw1p04OiMAFHTVL/6EHNyg8zNsX3eUFqiPnmJP
T1HXvAdGNLF+BhuwXGnaEeT5ECqvAm6CK0XCTLopQP5qRoqoXC+2Ek8qjuMOR5yIVcvzetjnmxB0
JqWp/75U8l28BW3u6XCA+Kj/0nJ2KaDBQhoNeSYhDh5vcK5obf3rM0UfdxXc/OCktgOo0Y6A2cp9
mB/gjv1Ji54xa2D1qiOlXxCZWdGS+IzKwV7SA1ZUKWh8cf8Ib6tFWTV8TwZXdcc5RJLeWvxoU/qN
wrOmT+EARwwTTCeNfSCEfZB3wi1VjSD9aqf9V39mJC6mV79Kh/4WukouuZaKAOFhbEeRRiPkvBWL
dZxiNZIIB6WZNfTdslf5HdAqxPQLbHd5RqAi4aVE7KqOaeDTsjY2hpow+B/k/Uely5EiNGQj1cwc
z9EmzuLulSw40ikb9LIqB+CGz+OW3wVmu+16cWlVsBMIdOfk5ByrFsHYaTWSI88fWcSE8O/sofgg
ZEM4S2GGDT3EQq0kdz538BgMKfCtPwOxyqjWqnUS2gvDFCbp0iLGuEp5Vhtx5VX2OP26h16OnI8v
hCve2uzP2fuBRTj3LLYkgIUetyAuvkPicPo3RuoqVSOlaWlU/gHu0QamPSpUOV9+ov4F/ZomKHCb
hTdieb3OrCy8vxNb5IwbU5L4jh7eVKU/wqq02Q3Fkp+UJy14NIzxE+G98Wxc8H1nMUWdAg/q1f4E
tGgPU0e1lEVezgyjfFXk5Bp1l23/jcuaFu3Uv+lcrUy7iLsSaQCdIKPQMqSt4f+HqKbGuVAzHEBN
8tz3nYlBfPa3pvgL2nA5f7gD/TrzdwssEHFfyhFcQxyA0CvpvdX2uMki9lRrmV5GRxKeOk7AO8Ts
bIKg/2quB0/XYtngrvneipC/KZKAN3eynSVPpkXZdx/P6m65i4kVhNYSNKnTv2wyT+EvYEZBJgk9
CuleAnjXGPyK81Q2v8eEL1bSJnIAsFOTzotI/cjR7mQalmine9ng+eOkV+kF/txk3sDoW9xwouHa
WseuKXHVVGr8UgfSJzuET9DCNLYVsw5fvqmTSyEpt1edMGdrJUFxT0th/z58meW6+sHU/tdDvJby
u8XkfDh3bJsEnaXNpQza5i0vlmMCENVk6m5AKR+WIPdRTTl3CktsNoRv4OiNFIstm4W/fch0a2jN
2aKDiG2KWa/6t3RhbS2QhaDJusPPOTZKAvEil0A74MUQRVoyqz5RXhOl73fq/9yqQxlPnFDV/Vd2
K8hex7WYlF7/1GJBbZhH5H6qu4h8lOdfe8OZT3mGnWkKTmbF7V8HE7no7GsMFpZ/0gm5ulSe23NV
M5qBMLe98VCqD0AwSNtP3tkv1wPYwVoFYMix70aYNtL/d3d49gXhVGKFqeiI72xHlJfYFz9h45/P
91quSUornC+W6EMt0h5/ZaFIxIOH1dXwPSbfrpH4/tmMAx70X8ZH/BafqCFwdHWLYF2HsTPw93wZ
Sl63AaxIzgmEneJB9k4bniezGlj+DGKuIm96XaeVJtPYPma15xCQTNfIK/MSxrnUKBCDRr2kn0+N
KHHX3q3X/J+nX2V8Qoeuozx5BKACd3OAXSPlk3At+RXf+thisUxVDmRUs6o0KybwO9LN6boTg7cM
Zv0mpdRT8KzfcN/0CvDhNyatfF5WL891g3EryE6cWQubxdbFw24PdE5BVNBOSRVijh7gP4K0FBjK
tKpIaYezo1sghSVoS/uWFDetWuJSYcpZtrLX+S/+5ofKS+YR4XxMUz7GjWuYcKJDsKb/VJdN4NUU
n0C6IjvZRyDjobUh/D3zNkNPpOO1lLz+O15DKsnqqe5Awkq4xPiNjFPKL5T6OaCD64JCF9xsHKOM
LVD+bFiLfx/WrJSxn0RIvcDFqPZuenCgLGL+VETPUfLrzPQCgC2UH5ehfq8vPJIcxiEhstDvHmP6
x11iA9PwsaT3hw3f9ooznGJVf3SzJDIaavB//mLJ7LiSBB6ydpoKSLeW4Kr4NwCDR1AU1fp7UvNC
BYtm7Qn7J26y9X9cPoi7OudNypBHG1IWXO98AKgz5GZGfvpsdOU2fJUgDGu0sdk5h05gG5iN132l
o4VGhMpnj8WdtinhIJowqQT0/XcxXiPkctvRLhmbICNDTWzOZxG7TEZJl8xlpq84xf2nhIdMme7W
bDge714k7Kmspyce4vwWlmoJL1LqqfpvSqrwsVKDrC3Ua0x0cIjHE8jnUWvDck54iL5ZBFq4Yg63
HfudEtxGQ73kLYKVvS21CCX+nA3dk7SYtteXcUPqS8KMLb4wFNg6TwvQVTIzqAsodhnyeqfmEIkD
ZQIFntzP2bri7bBxp3qOW0sDaFQQkHVQvJtIhELZ/58Aw0z1mZeNJ9eqUDGJLASmt1Udf1PU68Ui
/3Zts18/56KDygmwyYMYXHt1n7YfNohv0+qB3yxiS6RVAHbHPVLOb2+cXG2u859pO0s5KzR7XoQg
nOexaSTPZm0SwRThpabwjHiZnU2c68uBl/hzaHY1qYBAFpWoA8J7y/umZHoiUWxCSgPoGkGNHSQr
kNrlXYUzuSTIoH10NLYBF9Ecpnb5WCuw3RiUsIk8mKHaGXKMHJJAKyXazv28Hvm3YwmunOqnwfaS
VID3OCiPL2MNhlTHEs15Aj3lE+WQNzkYFLAkUz9MNqbI0bS+FPc/XNoiDIacibZExZSumk82H6g1
xjf1zREnw57oASwqi6DNtgZS4WwVUI72tZH/Ubhljatj8nj5dc++pTyN2KW36SYe5ZWtGKjmziEI
KQ9sSSXlbaAjCZq47w3v6PCT8uuU6Yru3fEPUsdePbo/ghtqvxdR5cmpLJmQxtzBhc3o9uUjpu0Y
Zk138rVp//N1YPUmJ/1BnfaYraikuk/39ZrEtBwyvaOdGc+WiqcmyD+qWIAWKoiiTEy/fsfavxEr
vL161KrEs1fNfohgyB2JNhTUEpxBttKhdsPbmm7GTOANaX17rWcTgfF7gCm1wrxorUQ9eqqce2M8
0DMnEWGUXNqy5cp+6zgfyphR1UEcgi/6FW9NytQb1QVYy1a8358MVsjwdudUWLUonPEYhuAoO/aR
EhVhJBKqvB+BGKv367gSxh2FpT8IY/UMVVKmQ00EBDq1s5OlJQFWuCtOM3FZWN5gJwMigNVF4041
EukYpvs5KTzRZ+R0wSdXhOfwbhUVqJtE/LoN30IGC8x8HhfOQn9ZkJCievG5ACCACSwjC4AK3GJH
MyhJWjeFrGaZwGVRbwo8IZ36Aate6wxIFghn/cHki2cM3IGndhKUl4HqrU3BIvigiuFgb6yj3gSu
Y9RMhkLJMBCyZ3VcE3P6kLWMOo/HBjC8+gR+rQnSVXpVhm9v7YvGFHeAond1EeDPglf0nzu9FUNv
WjoIz+trZuJR244rx7IBKV3fxbbF2hbJGx6o1oCj2zUBq+axtNxnelEN+U3cHl4oH6hWVgL29RoD
RDe0DrZD96EbcjEXFtn/vpy2GbCjO48hRw6IOenBImbXU3IqojbyFqwa1VZmUGamA2oxiGG616gZ
y1HM8nm9ddoJyK+Rfqrsw7ds5b8v8RTpOGKe2o0Bm2zkif3+mmlxVWvgVLp7GlE/867WpKbEjSNi
KSG1MGmQI1J5HjHlTbD9xWwloYaMKfQyo+xf1wBEXdRApZyL5vQ05EZrItElTWmALcCt5bt7yynw
d079KihxEXJyHI4XKxkMFjpCAqS2Xg7w3BbVDt4CQVSSNY2lJPQUiAhGbh7Yat8MhRcbfuiVWqiI
gNWE2pcwF+bBI1Cxs3ElJLRE1OKscgqQ8OPiLdeL6oWXsDaOWoJ+/Xk/s6h19zTBJVzCJgqK6sE2
WN153FLx341Ws+cHHApYef2h5Lk6xiPVRyAR4JJEKUOvqKyTsyLRsMXclWlguQWNqMRuit4gf4pV
QCE1alhXrL9wu+mefIvtklr93wOxUmcuEGyPuzmBPlbF0oP1RxQmTIOKxTJP5LwA4ZZGl7yj+1kH
qqrzdKgCXaNoKvn3/z02L8E4g2BfkAHaxb/++/oNKFFJv/UvZAy9mJwOchU9GtT5W/kJEeOMai5o
DY4HiuGc6dT6irF1wpD6qhNeYE0iB1bTRXIUnS4glhHeCUwzltQCiqO3FrKskZ/op0i7YIK/LOpF
gssvU6FHOaohMq79jllFoEYjpzVRpd9v/TPrN1e74oLWs35VNWk74L3OUDpmKrCyrmfoT2cOIQ7Z
OEKxTU7WQnSkB1b/C7VWSNh4YtkAv/MTtDoP9GZrkfQXeStnGppt12/z0jqd4whwd4oaPvvDAUgz
PPThXOw5QapsBoKGd9YcyaHKnEtjU4Oud7KWrDqTvijbp+fyDeo7TYfKFSMeVie0s+bbEHQoHnOY
BIXHnooJYA4IqEXz082xT58aukQgu1e5LAHYVuSgO9dIH2J6W8bkCIgcf0UsAaLC+ofJzYGNWdGd
ahQOdaDb2BTTUbAos8AdxTjL9c85XkAw8S20lZFXIku25ibOz8urFEDlbIxr2Dlq+n7hkjYle4cS
glx9hNDSZPjCyE0bxj3qGtDhjjMXXNAPKGmvhEvOPgP+7Dg0EkNAZu1q8ijpwOhmBVkKtxuPicdk
LMmMc52DmZrkKLRYSO4X6jY2QilmufRfrWHwRahaD3J6c+gzegdHbq32kP74ITZWlaEShIQnnkFg
hdy7fiCG5qHwjGbpg/29sFdsgXqOm9SRMtTbaS0hXaH3oJ8mt18z6KN+P0gLtq2tK2/iZ4i2X12y
ybD/u9WUSueZc5o4rZjQ1v9taJ+rnk0pU4yuffbp6PN5qR/WNs/luS2eH5MhFkaw8fmDOpZnxjG6
5+gnqvpdN3x8lPhYKRVPbzi0lV7zee/ZVQar0AmoLrwhF+UJja+uuBoxi3aNGcohRgrCYoN+Q3LU
PAGDlmVo9pggK0kuGa1KmimVUBIU2L/9tG3Q3OvRuqq0jxu3QIve0Z+T2kYAcw3LuDRdRTDa8hw7
UuzWZQZne2NkwHR/22PbNzssn7uUbXUO1FEeZyv/gBWaJG5XppDX0gE5/xmx2bRrBJZ1WizOIRNx
fm36FRF/dOUvX2/HxxGCLcb3mOZtopxeOF35f48ri4dzRrYZpFZ4b2ls/lM0MaCMmWoqxUDstzZk
kHXNMl+//BMeIfnUU22H78ZJRN1k9jPYwYZkZrXQAsyPdVcx6jPu8aEGFBosXRgpt4QRiJoeEXRC
l5+01k5ibd/UIGX4/CIOjlRTCBBOlij6FdFUhOS0f6h0a3cSF3cQOaV+5JfzfbFUSuBTvJQ/ZftN
l4cxYGKDX9/dCAdKxBTrBH0JPuhmua4Gx+AvbwQhnyOfepK+A6qTmgp2AFmK5zEGoPBxzm0wLsj9
4zAxsqDbNiwaW1n2YSHR2B4A2VUAgXzf+2YsqTYHm3fDQ2RX5KTzZvfWQ3v7D/MR9wFnGS37HJKi
ly/bvTBR7K0WeqjNWUBSvU9wUdTV2DTJTCXXiNqBxOxwJSUZU8+XAACRE8hKhJimhpM5oZCSXHtG
qty55/6pbD+H/GTHIE4DSu1kSH+C/OxSIrzIzLDVyo+pM+/qbERuXM2I3Pm6V19Cbbun3hpr4WHZ
zY/QteCiL5y2A5Jjmep+ddAvoP6AXl4JfCggXNs745lgYI72weZNFok56T5/1WqtIZ3MLBEc/4Ms
Q4s+q0ZmkkYzkDTwC51Wj5Yss7NXv3ayZ+7tbfgl83DOLnohqKeYwymV8VJrRyTGZC5lZwH7Kcce
8Co/1QJ/0X6OI/jImzZ5tqZiQ/UJmZ7hIrqhn7GPEVu+L9eswcT94GlF8yhjgCvruopuGzJIABZ4
QFglDCahWEuzey+1O7FqotU6wI8KFPCRGoGE5ztbDxWaFEuqWIi4/iew267MF2nAAqsVr/1SBS/A
07L4WUbyUH19sxT4SCzG2Tbm7F3So64/SDNR16a47SmHd69ueo80cYjDbpfrkGW9bKzSlAxQGigW
2f5VIcxTBa78ROlezB994Zks+z/8FvKlnoCKT/oZSVC+5Qla8GhS4JoVkoFAm2KPHsBPmidihgU7
48vFtqOibOjqBdIeOIJg4CKmN5B0rcux/AdFuR+taP4v5m7JcxVz613jC4u2wWqqvZQkBhAG8l7Z
hYPPEShbNk8hqAsEqdV2FU0DEX3fjwJ0miQizHN4SxW6WdqLbv0G7rqO5PfYTW3a4Ql1rrvMsKmd
LN56QaabhbybsEVua+xx5srxh8vVHW9J1uoancQhVam6jp5leDMIBlmSE1Z9aBo0tk0hhLXy7JQU
HJpSa558qscg6HivjuAfLLEfmzCZ2rfGT4Yb9UNVIw7cLsFAjF+MwUV7lU+yrUTu7qVNQQLuLbvx
Ma0U4kuLTKrrv/As3NueXIyWbu0Fb4jzRBWTLIGoHFaSfuZpdodbvbqXZFsz1xsIL3vE6mlu5gkR
9Z535Dgis6SvWn8v2drWBQ7+nh4Ax+fK4ZKCiGyO5G1xYw53hLwOPRmi7waSjS69zpqEbz/zApGw
Xl1I+q2SMPqdvLjSK10O/Ret/k3P6MmsgM2eNxTNHedQxEF2NuKtZ0NCy4UhuY57lr3fOTufaox5
mXvd80Ct4FEqGcWJItJSloYRrcr0ObxuBG9PIalNEi2LrRVZdbNAtsFMhslMEkGCUmpsfJUOi+yy
hl75oloa8KhBy3wBc2+KlJvNsgFaPaFCJNNXaxfEk4lmvRdB+6MWebwkv/3bDfv3tihc066+29eN
Og9uH/gIg2Xlog4yfTq7z8yi9IYOKufBUsfu78WXvO7Su3cxrYWUOEdwfTDesB+oXpMgjBmAf31t
/KMbwhDWZ/bnda0p+DJ9ouijLr78Y4olFkkVu0UyK5qrmSywKeDb+MvC4b4FXKlO+nCtEHM24j/V
ReijPNZinov+mmWSau1n8+TU6o/xcSXDIDgjbqaiYUJCQiiSlzvCLEobxUqjM4afoKEDGDrhF7xD
Pk9XYPgYmNqizzyTgOngwwM6wquLdpiFC6voGHhXJARrZVIfv0xP8cURiYHRiariD/PnCDrlwnlE
YXUjZTPhOnKmonPrvUKaj7LMZqECSFOhZU1vVOiFoavBMT3QJSd9969Obw5r7ki9QOISdCIf3EIy
IeqFsPxox94MgbwIF2jRldbgHhn2ASWtdRWkcIiV34KA0XX86KDjXwSy6O3KOHBsRejcTmo1GuW1
TzUMoXUo8iN6HrcS8J0N8ZS7wusAoWVpIczGr2P57FFrQ/qO2ji7DyMtstO5FNlJaNto4paoiRD1
eLG1FwRmup7QHH9bnsneHnpAWbXNUJIS2pYw5dnnoz8GqvzyuGgyOAjNc1GL8SD9ZNm4pW4QOe17
Jgv/uitNtMqKMT/G6ry54vufGYiGwuDZlLHrurtkeoBKU2xoUlbYHc/Rk7ENGz4ib5GJNXhEqw/H
Q7TT6p+J/flBBoTTNzvyzTUHvQS6LSGM7lGSlIKSVxc1sWgeTA+w9tVClCsWVW57oYns9yhc/EET
pY+2wLFEiVypNIsqFcZAQzt4EUQs294Rn5rDQn4XzZHj1Y4Inl2xob2oYZv0+vFHR/J6HHuThT/h
j/UzPuNJryiPxT0/VgHKapMZm05yB2g0PLfjAaLT8no3vNR82642/7EVP6JybWSU+XoAO0t5zdRW
9Z78b95jJjlSNDGOO/kqTFVLWqRjeDdZVhBGGckm4fYxrnwSPjbwmjXYOGMCUBcbYPRLGvL+oUZF
VhoMidR67eHYT45/ACrSBFgfku05mJLhRZLw8hyqHijgM+pkgV0WAB4QMkHzyqP3hUXUznXX1xuN
XwOYBhfVaGQLcbBcxEzhUvkUO7GBXc84N7L9CgXSUmdJdHe0zHND9dUeBxE8cJ5KOnzSuWn+ngC7
4jtgYntftmkgmUBtFijIl33zGG/qSrRK5Fk76bQrufqOaMsH43H5n9CIS2frSK1U6zuT/YEUento
wiuaRvGKoqNU37/TO9h8/txXR/MT6wKx9NJSXgjPra3MrwQCr1O4EBXHvzSM52lMMwD7G93yiLF7
6QA/4Co/PnUFeHTdyrVQH2ULJR85SbBPwuu+us75fBr1GFTmFexvfvoCflgDjPj2o/2SfGDcLB0Z
0LPojGXQo9vnIPb8v2P5RsSlL5XuD5yqqzhZjoJORV6PGOorltHe7gH/vW4hCT7r1D47r91eJ/Sn
hdBdVawiaZaWkPzQzSUTAyBMe6X4Lxfn9Q6jE+nX/81BRV1PAEFYUSB906YEDiQiOQH+Gl+BOxfv
bwFarXJ2iXySfBHUtP1MfizB/Ai0hEL7F0pd2B3WSKDcx1AmAzhMqGnE9skJDdd8n4Rb9pFpmX2E
J6B6ekRkDrhdxnfGDbLZAq6kOY48OFNtoN7bhJrFWY2e+tvXrOgaHxl8v5hcoXQ0RSTMf8mtsWse
bPoMVDSVi/KiI7tXvtOimXa5WTGY+vQWqplT3yXxAcGrAr7UunW3uX3mFCuQngQB2BdTHhXdl0Af
hXeFmcyivzQDDp9N51rrTtHKa0w81A2yYxcVhATKBgLOrfXqS8lW3IbwUvJmhYkKAJQGDo/cQ+LD
XLP3i3yyk/t3YpBIrzv+weX6ccj2ftsTDQgbIDuL7saDChszz1ou5bA27IfDY7ND1fLxdlRy9wlB
EIXc7LwooarL8w62CZCd38l8NxWNrtueckJEmf5MeHbrUyiurAmvY9n6FuroekxpZLu/9LwuiNhp
el+wtCCalKIxfQKs+aoaaBMfn4YQqfj+CkdRCcP902b74FSI9GJVVNo8A0ipuIZgvlZWhsjsdHfP
wOBLLETGZKS/nKgD29DZGZGv815s5JwvUlejA8Mu6MlUGiwd25lWlJP6TDmfO7Nwn7UMMFUT+7DO
qzLL7sa3nhXV4SRSDZZPPnxz59qVNXg8jx9EXVRpdCRlQdiW+l4YJuwr3bSkc9uLoMKBw43bIJ8S
lSA4ODDz193g1aOlI/wi05cgpr2eL0Qamjy0Cs6prRIKflTJiafMa8geHUZVm4yvUFL8VkVz6PZ0
oAuWwAECcdXO89sljVPfEQS+tFjjrBO3fKYcT5EDB4cj5JXQJr8YTVE3oMz4KCrp5LRYlGhvp3Yb
+0/f+UUX6mrMNJ+bGlJatQEXsJ65aR5Mku6Aj0m9Xazc9NQaA2xCvqhWFzlHXhRcrlxsH2s0xos/
r7Ni/zjrpzrlb32eHnax0zpsmOrIsa4Dq5OY9gU3TTKesanJRbtbRYwKyBKKL1nuav5ZpT5Oy0LP
is2M7X4fIoVq7DLztILDhbx4iI78yl4JEtMW7HeXzZHxJapaF0C7p0Zgp6oReNA9r3ECNUVc4D4x
mKqELi2iS8P+HksY9poM+Dk0Ck8C7EE3P+0hIXVJ7Ab6ZtDpII+S6DF+vKY8wfkyHs7KbqCFmIsu
bo9uGrSzyMUDxXLsRN2pN7kT+Z2t61CXzSo57wAg9wgUz/3Xc8gh2bSOpNwDGyBFbtXsSAsl6HPh
rDo1FfK8YmlDs0h8L1syQ/9z1pHcWDOmeNrxfJ2iNCCRwYv8igwWz0U5tXWJoOt4JAm1cNqdxRpp
TXm5EmIfuiu8UmSqLMiyLrVxOjGvRMjjkmYO4DovHvxa7B2s+wZsIXbUgcLHV1Gk7+6RKpFMocBs
8A5eQHZsL7VKh79km59FFLf6LH6pva6GR26k26Tqhxfl6Gnv3K8/T1xHIdemZKS88dz2E5LmBtH6
b6fZonnIsu3/DkYnJIv23VHH6xBRtKY6gVb9JY7I8n3SJfRT20QpO/SX67VeaA4nHEJwvQS6btW8
262VS7cB1pqNiThfJclOstMiU5mKX9mOp6XYUEa2br2Qzw0auKGnoC29HMBlcPgpl1Q+bH22dBEE
GxJoI7+PXpGz6xrOWKIgRlAUxK5wAXszi2cyxbkCMFmrRIOEYys2vAKxMInNIUstGsL8iIoNf9cX
/2pX1uWDke7lQPlSldgdnF3GVJ1rqwoIkMlGHqRFZMGVltpVvE87pCtAD6TsBTtYsnk8EEy8oPqI
Q3hS9+2l4Fcx/QoA+83dk8iL7l5EALIGVJduPuOieMtGoXt1V+ZurHT8H2KRMma754Faul9EQaYe
PpxG1HY60AjhEvtxQ2eQMYE5u0jyd5t9Jo+uPL7D5p7iEZj5YtM+MMD6+meJBaeTq0iha9XuE8FI
6QO6K5D4a1+B/kKMsEiESE62KO7ZR52flMAaxdgTjZOU8TJ4lb3RNGYPk4tlJLuPkqwKY/XoAy+w
HCThJCrCsnclzL/hEyJ/AKl8B6Yrib7w0OXALbzwIbQET255UH4aiR7M5eSuZWRZc1w+FFWq065C
ITtrG8HJH+xhjJavqGX3ZBe8iuxCdFz0+gm73qQkVMORbB4qaxd1vlMLh8eBqrMmnPbqGRWAmOSx
rLID/v+9WdzgDGXRfMtAXlw0RvI+9mH7HvH2nK6zaoAUG3IjkvJ076BSeP60OxEtyze8u8Ei8Sc6
CUFH2yNKDA0DuGob42TuCd6hHOj2oTRCTF+tfbgpufu40+r6c6fnj7u2HGAacv7/J9Ba8r1nDQR5
xuIVW9GqENPMyL5WQqpZxEz8GOoJbW0Jns/WZIiTJ3HSMbq4IcnXxmVVGBl674mg7POY/sBMbbZT
s5/f9AfKTw6bUhj3vUgmtPLNI6NBMxo+dS78QHU7CoeA9WyF2zJTuHFDsX75/4Oxmiei2/YNmIrR
ZXqRWLwRxNcE8NPQzSldcecjJAPLnoTaFgo2+iFvM46ACH5ce6Wy2/e0dkGw+KmPaBRiv+J3YUtR
J+D7LF1yBLdukDNmnx4qctEdqwFyCVMOMo7UkM+PDunUO86YBjxjsgyp/0ANvsOLBT+llLwdx8t1
SpxhntOkux+Ln/rqwYRX8sauxtpCWjyo4LKvV5w7FNKBk9jklYbv2sM5uG0bCwN/i+5ppDQRlwlQ
QhV/0lwadCawUHpXaDB38/gkthrqXcM8jITsVbXr+u1H/Vvv+Hkz7Q/a0c/ofFO981sz5Uiw9eaq
TRiK3CvVl/Mn5JwMlCgVo8sjv1+zsEm/imbLCo61fnUZBjVUtQuJLl/Jz1LWKheZFcyoNAH27nwK
2warEu1x6/1bpVYqbL5Vw5HQmQ8aRMQKAITwukCYo+cpyzNv+l5pBY1TVGQkF2nbNjajwi7qkGFE
9IKuCHY706T59fIsORhLSjCH9y50gm+7YzNrGIre1AYHdcPKzlBAsMo4P+ARNsy9c9632u+1Bl6y
ZhJ6j2DULjONHyJ4OJ3lZOyhH3itkt7/SfyDyLDL6AQN0s7WQaLgsP3T7oxrB5lXDx6KAUWSfoI7
fSf7HFG2895dI9iNQO8IsEKwuJ/6xcT05KC8R53gFPYxbHNIGGekaeqKY98NqCCFO20oZKWT3ILo
q5YJwCIQjRKNSc3npKXTo/BakjMOzrOj3w81lIzsjtPaaxHXMOd83WZwGscVGhVZ2LkKDZJPIyVi
ZgPFEqNzM4BIbQGDlBKJJJfD/vw2FmAr1kEgrWgUZN27Yjf68NGkXGDVtka7iuAQ8uF6mlNhSr4i
d92z3ly2vTUa8wyfOH9Q8ZUt5asEYqMRv1v7Ac8re4VA32ezDYBH3+/TqC7pCtoxFf5MvgftB8fz
q3THbqSWOSgKsb1UTN/k63YRm9AUwchmhdJTqFD5+hgVf4e+bccd2e27lS18vNcux/0D2g+YHRin
2M13pPac6mKpa4nCKkYp56l8c+qPAaJ6PQAU/XN0AUjQvDxtj8xyJQAmKy5QZiWSX21zSM1/9CRm
m49UH/wd0G72MWZZmmW9qHLFINUBcZXftHC8/6DznIQbAHipv8t7q1CrrAV+plF3RZty0ZDZapfu
cR09YywhefEqNAT1JlRsvjlqI/jaTSByV+kTo3CA36YZ30HtpQf/PGVEi2OePvLZeOd5rC4tPdNd
D7hOqWsAakl5oe7zdA6v1fTlt0Qp04hTXAPogTAzVrtdpCU0/Ni9W+r1a+5yx+7Jzc4jbejeAFhK
G9WNqAhFqsqeZ1qOF7lh3QbXzbK+2Z8Ahep9M95ndTqrO4M0+curgntFHWUyWAqPA07EKFhettcr
Ny6CXvrwMxbdkLuAVFd42qbn8tcaBVtSQPCOJD/71q6HiF42sN1UCJ7q+gH2N7AhhOm9Hhr5Ooj+
/QscruBuYgzJB+VA5eqjFkMmLO1F7YLZOUgyHL+6JU3L9c+dIi0h48BVc7lCx6g4y6fnmmPyYXAx
TgHyAoESAXLoAolx+Vl44dhfDfIUu76ORcCBo6W81Lkdo18ZFVEXFNxwkxSCKhrZ0r37SXywTKIl
AZMqtMCugxKfj7Z19d5u4JUqOkS+O/ycxXZAtx4BBMOWXroG4Tl8BtJOTfr76bq8lAb59YLT28Fq
7HtikbQa11x/dycgY3dMb9WpCsO9UOIdCiy04LHX+ssO425oXzm2CVDuj5zDjVCm4JdbplPN8VhT
7LWvhzMOkiwKARDMERbyTIRCMI53RTeH1hNaWS7MQZE64BVWtfbxILEXnDrvkpR4uhxquEiNhceS
KuvGMTouIzGGBATua9WvCcmArECQ8WySAilSuTEdHJY7f4KZqOKdGp7zAPfkliwKnMGoUPiFTcyQ
P1jvuasUh7P81U96nHlCOHe3heiSM1RX30O0d5G9wJCKjDVFJGgfDuGZwLS23yi1zB3q/bu5x9ki
dUW+qHrKDHuxuiyuXBZnzFlzWuYDZg1JpBsA0kepW15uczWFJctBMcpDiuR3q609Ve4eQeqmQcGA
sIcNlhYkSIxELq3oIjygnC793yGRIlLE69kT4iHeLe/DDUkwem3hEoSgZrx1OKdVBPyMvgcpPb7P
IwWHfnZ6hDchEkMfqjvxAr0pxw8DzIfmfdhMi/zWlhw0+4NDAN2lxP8V3awAxc/E39p6OFIEu6Fq
76tArlYQA4B4feYA8wG/LVj4RNhaQi1iB7pYInZgS9MYnhbL4OtFVIXL6V41m7KRSy9tT26rJk2x
4PK42Ri+jMVPcYJFElndeHMwjaWJGoCp1w8ijWfg0DiG6lq9UT/8ePllHbZvtn2R3gzKj74fdZSc
PNbMrsQKN6BBTo6zFOpO3zb+9zoW7viqEM5d4ie7rPJprq6ImAVyQNp8geXmQ6RO6XhPG3bVQANh
TOpCQHK0yBVF3XnGRk2B4DQyiyxKSRbzOcdQ7p89mgU5yYNatuTKfmvIocHGbdKyR5x8B0d6hfZc
vDPSv4WzQHymH6uab4AZwHAtbxJdxsTgxRxQ/+IuzsxJCJ1INR2jVTPvrxUihfnQDkpmxmaodtPh
VZPmII2X8ilZ/B3eLxtSNX4ZT2zWAXfm8pDwPnWv80lukiBARp9LvX6SMogygNjjPXvV94EXwewt
Yepu6s97hNXuBHcRDju+9c9Pkyohq0c+ZsmgLysCgxjA2r0Yt6r8VZRDZ4lDxn6eVWKNTUCLMuru
9fsIlqfWM215iLLgpZp9fNSd/xt+v1kr6wu3uV4Fzz1SteA3ySrY91I/d15z8qE/V5PmFyttmV+L
ReQMSvfvb4tmWZD+0x62Kh98kaTKPTlNE8xcOZbqy5jzoFyICVZ+vcFbb+ykCFgws5b+gAsMwXjZ
R3g48rxme8O2BLCDYVnWZqE29lsV4HipPS/fdRHk6rqHFiN2PYSCbUBsAb8eAmD9FbeOzaD6Px7w
NT5hErq72nUI8FJnPM2WWHDnISZA2QgFveIMq5F8GjM9Tv2Lx1tRzxZjHaYN5PwlAfSQBSW5SHOG
FtNUD2mkt4Fnti+5iSacdgs99xMODYF5wu53Y+1TOStviZ8LlzM9erHGeuG8KS+YpIqZnXrPdH89
C0u5HNrr4syIDi3NLv8QYGm+Ed2zmHHLQE1OUxc3dNDyID+NC3l2+IMgaK0siRBnyoV6kBh0wY/J
n6FpgN8Tq+RtnOvNIUS93X0VKFBaHEa52+6szR+5H/oju6ky39P8DqNmQgCsRg0oGHhp47JYXcYI
3kqXL2vZo94Xr7AwD7Wexiur/K7zE/u/XuaodCuP8ltjgsKrnpJrVfBMLQYgFwI11C+y7vCQbh6Z
40j18tzu9VzEesRKcyO6nyXUJw0L6TEoEejVbCRbi8deWn0nougEnSFm277efGxaVD0hVVqs9vGS
A3SOBluYFK4D+Y8ChjL9xsP7kcXdOjwiy64Dlb5laxW8UMOzqMuqcC6u8QHdGDg5z2+Ucq2nt8Fp
PWkQrQxCPnbiFk4gZpbzdOsaLE2+2UBVesXU8jHcsE7zGFueTJy9fR8oy+baHiGg17Q/fpGG11Pe
IrpfbP0oNoVCDgYszuHTMH/Dlv4V3CnTjFzgxHBvxya8ymqgwY4X5s96o6NI6BsMaovq2/mdjFrJ
QpYpjRdV2HmVV4M4PZckSF4zVQUiXXdX5UmQjfsmNy0dwqhK2ketpjhFCoSaFHaQioE+nn4AdEsd
MIsWwlGHCbMgfHQ+r43CV67TPDPlHeazSk/L6L/y13t+vyX9LNrpQ5Pfpabl4vI5LSiGImsVscOw
8D47dBPWFVX2NdL+5f2kWAhKymxtAnx49a56c1uIA6zWrKkCUK+DQENbu8oDELGhQEmGQo/ZYahR
c84URmmD5B9OSuVkqTJOhz8NgWGK7lVqR+mmkVUvatZ6wzOtQ5RryuY7T/KLZ3plNwnrRa5cYs/J
yeG1Aju7R7+YDAxjltc9nVOd/vSLxNsj3DVqiRkeBCDEgt2p5HnRov6s1b56Xx0tp5jICPwSeBWu
iE527YWa9v4SDzihFsjYaWhPOhBDn1KqI4hEQyvbUGNjQPj3uOK8zlATQ3ay0cFMwyQJ/n/snb93
dWkZKdUB+euPKqmJIqvKgYPh6tgA/e/ojoNJUh0o0MIWKSFbEga15dzS7/ZIObxdLFDgvQlrWKka
JrMEjcG09cNWEJpqS5vVTHyIWST0NPtzmotYE3wZ+XAWS6hzJq4qXmtA97qIovVG9+PsJHvFtejq
Zh6fZ8KQTLOoPG2S4Rw2F9+bFrkFMny8zV7/IidrKRENJaEhymgaNpU2dZRc06O/lZdNzb9z9YwZ
g47IjxB+XAJ9atMW3jiBTlUX6QplmjPI88AWEoQ8/AiMp2bX8xinpcCPjUaBCryusHym+9NmrH1S
A2mBSFx7WHkKAmbrvBzla2JH/cx7TY9U2gb2azY75Bd2c1Ik7fODhx+ixBNFvohbAmtKPlmFQvX+
HYt4EyezYWpipkSlbzzyJnvcg8q4PxkLaSl2rRDCKBlhkuFfvBxYQc464v4ZbAOMziNjahMLkCrA
BOk1hh6Dei/7eEX8I4KYXCRMZy4844R2KSb+W3oeTeA1Rb+hWs3BZuqSxfP8U6HYSYXAegcP1+d4
Z5Yilv+0ofcNdiAadNDCOHWZH8hIKcZcKF+2+oW08jz7ujBANWOrrEmpOP4LfWg83x3QmcXw+jvx
+Rh4FN11v2SkUgbNbR+EHfYhPmZiumIDlUqKB9w2bsmZDHtWKjDVm6bR3VC8/1+zQkZNMIArfyel
iNEpcFSmvmeGqDz22agW68X3rYl7A0FQUfNwamrUHtHLOml79J6rtdvvrDrkXTIO/FUU1J2wtyhQ
lyKuruFIGy/NwpIxha2Rw579D+7setVq5sOD/bRSKg78gNDPqDLaVrDOSKAMF3iI7Z+wcVjan05q
GrOdLmga2qdvuD0P/Usni1rxft9YuA5YuNPUMagOkIBH3lieDKhKUYxyKQA8hP/4vhPMjV2qDaQ5
J4T+HEJic9iUB8L1Ih/9czUwtGLs0BHBsYtJ9tAQoHUYTU2n0FsiyEdDBfHi5oPfRdKbHnDqNJrl
dShNQQ9owzl11Pq0w8v/iMXTIa32Z9TNp47WWrham93ROwmScG9KFuGQkixOBMJ0PCrPRnChFqDB
P8GWNWQGj4gtlNqD/kS0TLC417GMavNDr0hUmktyOfqPr2OI7oDgdV5cfawlS0psCNyygyIeBSlT
MEoprkWTaT3+Kzk7FDkLUFm1M3LG/padiUg95CZo4RtIXNoH1n94SpY80+b4H44NyCQD/65hzwVo
C8YnSFAbVCuKwf3xF/QB4Ko3CN7wbEF99kiPJoT26p4QnXhsT2PJaZeG3DMB5qws0hJctHQzJ9+G
MGjXQIEitS9kHLm6f+v4hi1cpl1M8dG9cBcDiH2ertHv/+lUImRZ408JPFU9A5O6VeXWMuOCHHhh
pPbRQZzQH9BugRPoMZReWQaPg/EEq1cugQwY3Jg1ZyphC6K/ppmGRQ6T58FBfl4fNd1lvatxdVKK
lRm2HNwV41v4dEzM99R4X+9SyXI6rUx37CS9Pakc6LQ4fbuJKVszUV++hwxF3cNopIGTh+AcoQbs
RT8qH9UYiWfTXM8R6Si6MGZUzZdjmsJthiyb16kQZG7s9ReaJyqu+y+GxfFcWckBJCVxyjBd6XlH
StazoI48Enuq64CqAbYDMqX1VpdKu9QgrErlKZXZRi0bub1uv5OC9YSR3SZ5x7SThY5XQjsw6TkX
3tMqfBIt6xc3lRNXrtvuafz7XuJUXEHqwEjt1VDQK0+vPbwK1HnuqJQKwOEACzHl/sHU9YDwdV+o
0hLs6oxjkjBkdoa0J5K4jsIHcfZ98NlYUhxkGP9SBu5xfZRoMiQ4/sv5y0GxUKQom/19N7cP2yrY
Ti5LAhuHtzEqva+AJEmC0jrEjlnLWMjFpWLK66m9elkaQpSykyNb+2tDtiXxhZ8zcLO15YEhjlpk
1OL6jw44Pvz8lqcGsC1LBfm7vP1xh/W8zVUAtzt577DviOem1s7F//Xu2JpqKJLkltO1JmR8Wbck
4sA4FCb4d5vjipInneT3JxBsSamkkHni5dkARHDPEyGZklMA28q8REgvNONVQJy9mRFZbCAtL1iy
vSIFZfhCsbAc/oYyLnqbyif9qbwFBypQSGtm/yLBIbjmoQxQzE/3MIgnHZECcKADea2YCvyopFaM
JPy7NEbclX43E5atlSdwgl1mvLizUF3lBXdvjFTEKJKTZQMiTfHXCJ0Iw4uRc6F1XVMluH05IzS1
7GGHewKTgVp0jydYrCdV7SuH7dsICo8I4EKaJ2/0BD2EzMHzNTD7ZMYXk0aL/fgaCIGxyJgBItU6
cGu7z/kTVLH0sClpHrcz2/8GEO8DMpwtWy/9NRV1DYRaqr2/HgQd2WlXXl4wh6VPErj1s6akXt3p
h6yQ3yApPW19p7vmYddswwUwA/udKIlFYZqdeveX2gx5c1AYfETk/6zxu6HBX2P+VTR66rEGmWug
UfVazogaTxymt3JzVIMfQlE5ooZs6pyWM9BvXdb0OlVMhwIkFnoY79WshSlhHBm8Xaww+V7E9115
KvBxv4ZNVX6tBdJRdPjJ8+uf7aE0fdIT1OrGKZ4YSf5A3vHoI0+G/Ki1leSIB4l6a1dRil3neEyt
FcTzKaXPg0BznckEkh+vD0tUwjyNYlypUMEEpKsjfPBDTul5vLBW+hubNdbFfkKIzpArmRhhYiHV
sDl9HbOe8OWdJA2wMZf/jKYXMMM/qSA5g4M9UiRtNQj64XzHM/x8ySOA3rAJXWhRUPnEdGUlBATq
5ACEIEfAcJSgzq3cH9Qa2D+EdYHFwT6lo0tXF14bqInno00AIry5KublWPjnamhF5RK6JcK+HYh8
a21DUnBvPEPgmYvL9+61lsqOaY/zpcnCoVQOI9kJY3dwiLRxwZpwvAD1RjZE9YMmClR3+Xsv5NJH
If02zuijbI1LnMhBaanPZeIavGcZl6WardxC+Y34vLEqvTkueQFghfbAEHAWKbLu/lDVhp0honf0
Sns36UhpN0agrLMJ3jZ9icYQ1dm00yslzIrhRJZyz33N8yIQHiJXeeQXl07nlE5Q++C2+BZ1cOH9
kseOQHmz/1hVllSlQIopN5Bm6lXZqQYc70BJnV6FbUPReTVOe+u1kxS+/tZ+sZ5QMSxjKuDOtDc9
GXazS04ST5jjZMJkQJETciZ9Xnuvydey4/CyA/MOPQC9g7HymcGjzPAD4Zb91ifVuZWxbX2b9zgv
VRwww302hawcmpb+veqagvYwpGGr+k1O7HJPD8MhVecAQDcYQpxkwHIVT3B4n+ck6dOCTWlpegLO
JANDECHnUD3VctZty7wbpdwJVbBq2UM30OutXGXIJ2xg9ieJ5vzRj2LtjER7IhOOqmwYD8pYmGF4
HTnKOeNawTXwBSksgaHnuAPBGdJzbhcEY+u+6AG3xnto1QUq6Yx5KSHuWKQ2JHwX6n6bq0rNV0ni
gCO/ZmTpyKBTIEks8VSbpZg+wE08i2LI9Yfg5coB5lfxwonMvb1Ir9+2NbYEwbkwh4HLKXlviC1a
mX88WnMR7cU/2U7P6s1vahSJx4L2KysKzsodYlGdhVD8hojp5n6ubO7Kriw2LCfpSGHljmj/F11I
L6alR5DVbbTcykCTQzNPwteNUXhPS5soHaiuUk7iry0BewBQWnZzgYxFX8wWiERT9xIVQEYAtkyb
Gwv/TLmR7oCrcGOTYmCp1Lytov/3Ib6/Szw44Q26Jgm2bORpxF8rL7DiMNBDzn4Fi5AVrKj/HUW+
IVsk2uUo93Qd8XFSYYxBzC8ZouQFClfJiE/Bv6FS8l3wTx2t3u/+iTeKJ+jjdX6pnqvMNCbpOdQm
Eq8MUI7f9FJcK0pOkWPl02MuNE5FT4nbA818m+XgcDOOmVPfXDg9FVUg++9+y1LzuewXIVQEFYIR
ROcqqVJxfxQfxdNE4367qVU9Tqms8YataP2JjxNRZFnox1+GrvpyMmpci7bHSu9CBt0RtCbdYEeA
QWAOn8waVqyJ8pEJ7SZ01txSQKnpqLXDMgFWbMSBUEqepUnseBWXMt9Yq1FVoQelSDJODRlq7/Oi
rmeEoq2R/0kybi9kC7yb5LQbvH4UXFvrUtM64KeNWSwU5FXGx5FvEIrMtNG86QZxiR47N7j/ATbL
9ljmGeRceRRgyiz8QwtGAneFtum//VF93+zI032QN17uEzk7owqOFQB99IbBQIOftdxriJcZkB0/
BjMFZg3V/JXNSHggjMUu9auz1l9VC6mzaGn5MCQMR8bFqq5fV/BiuCpl0AbgXjdsg4rxkSk3Anz6
pK/DHlWHdAqrmJgP3/ssA4hfhI9kRNf9jThkgz8zU1SvTYxJEF9duJGY9w6roCfaIp22Z/bjI3qD
33csoJmyV5yDlqBoLrb0P+VPop6otNBxOdI6eGGbdn3ccaRGwMI67z5VzztzyTf2ON3WPbUxe2ko
rGAsuFL0i1sjyEYdjshWoAJO4KKXwo/QyujU1XWFI1OUBn4ehG8iEwZkdrcjjOBT39ps7pz/Oghn
z0L2laFf4ylyQdPO//OEdpVjzMELhXNlYDjtigV332Tb9EjXwtxnPu3bWaPesv39CN2zBn/wFRQU
g5m8Q84M9f62ba8n2gWgQSpxpELpX3WCrRkVTKadWUT+DOJJnsDvjWA3X2SErVxZt3oU6cSgDZqA
V1jLGG+RZHlQaVK+sf4zYICt0NDZZ5slZKor2Ra9aYDLbYrgV0DWYx+RbX1Sbzve0DG4/JQ/dQBD
nlNoHwdfViFDXpTsE1pRAdBZhcji/zWEusbUFjx+lGBJVJTFNqjHAirud48fA9nl2baensgB733e
pVnpeY2gJzqGAB6VYui+xOoe/s0ZKDY2FImwl2hvlK4JObAZxFEcenM9Zqlv6aKAGv/3+uKeX1lc
a6C+xWNW/1whukuhnojD2fW5Wy/qM8VZ9YbTk0FiLN1mDEIwkugBhN3wKuLbbFpIBzf7U977dCr6
lR55vdgFx677hj2/WV6BFTust5Hu7LyTZJa+8u5ohxwVWua48l7CxIAvs3pXWOyPGLTcsL9rcoNS
cNDtLyrRaFXBw5nyFZNj2kQduOfs/eEos54/kDA/LTnRXd4Mv8c1u+DS12ihGsSXMKfOtbVuwSE3
ffEKArGz5wGYO47X/24vftiqUfzzYtKoMFRlHfUxeDExc6vIGBJaUY5xxrLI4sxPTvEQ/fqdLElV
UDiOFt0E/MG/nH0aXz6/2OD746yvVv2Ydq5w9Re9PSw3xYeD+8zwoN8UYudl8mgqU7jBHKczQQVy
pcNxn0SIxSaizx4zedYTe5FZW7b5j9Nezt5vCstqBPFR7PksD+GzNQh64/7yTM6lbLqjdsa+Xfr2
xpXP7suTxy6tM8uq5z+TyLOcce18U/IMMYS3I+cIqij8ETzQiXzLmRJ3thRMHcNXLsa+/JLfjyY8
ycnJOcwS33XVd3hSkl5QUND+sx899h9ZiG5qfaO3aOuq0QPwvgWefRPup/B5y/+WmGUBdXirnkMf
qAskzKZxeTGZNfNd1hh/1tCOlJz20cmT/JTHhq078LqKFFJt84BM22aTEcS31AX7wZ05fOkc7cdh
Prxq64mwgsAq2ELWPKrunXLK976Fu7i54KmVNGxYmCWpR/Mx7qZOhuiUTz0zhbydXvB6L/dMM+yW
sPIB3KdFrYX8OHePAHb0FL79tkdwS8Ia0f/0viSBseUXdrZ1+Wmu+cyUSx4xqjWQ6f2b3VB3D8H4
cXGrmfDuX9gtHLwphaLG35Jjtc/8cmpMYDLYrCBiNcqYcQxzEHC7xS/ya8bN6+9Ikhj3D9A7Cani
9XwyOJltxSr/jSKnkU3cNczR07niU6JE3YVibYwW+BhwzXghAybNm1218ZXZOY1Vl6mMBaCEaQoH
gfkqJHIi9NWfjRXf/eY6pVgcNVJxWPkhs0cNco/TfKEEW2bAR6ADvJKB3444HGDoXomAivg8f++4
PqtYNh5ZSdMr5IBBWQHCCS9/e2P2gMvs7eKpwpyMsBKRhP+Xhl/mEwdHndk3I8jSB8vcrF20ihRv
RpgaZt7CYOr02jmMda3e5vp02qMbInu0jFF/xOfjfdQ20qD5FZ/E1MmsUi+2Hshay4aGdtkKm7x2
0kfBJZgNbmtWZT+eeER8jQwbI1Y/9qAvG/uawH2mqUa1QVXhQ5en7mgcqGSUnK+5PzczQz7qR6pa
hom/1UgRS28WE/0nuOSuzQH4lP0yi8iF7gmYHxp1BxHwQFNZjOL6kebUYVfvlACDnskposMMxUo/
I2wqn2WTWK5gZCEeqLnAZOIs1LSRfYxZ/RXL9oQsx9dxCCToSQJDzsJzDEnBfnDUlg1B43t4zgiA
KQN2h36K8V6TZK/Fm9m+q9du3OQZn/sotG3zR/9kwff5zCL/zou7Jk277Rnii6X75oesW+0DEUkB
GampOkaEXfZYZk6UuWjmFUDaQJDtm8t3jRDJnLyG5Vu05tziL0LzhJYZvIupu5E97oJO1egrJHUR
8RzvHpD0oiAzozSOLgQYzBD0PsNJ3w4lEEGTdNo2n3crl13pSppp10MFDMKfcC00YPN/vzo8PeQe
38CBwIdUceLKMfVlErDWdSd/epqChTgmisG36evI3oLiNPVE/CgBr8xOTsN8N9mWXY6UXIIpYMRa
6j0V2aOH28xshY94WmsQVJIkmzl3GrDVktJVny4OocHcceibHuEvJH/f7QwTbCUUIvuunQj1DcUT
VaRhCcoN3I+9rqckJqMyjqzNsMrQDnBo3o9bgoeE8FZXuryQHzfTJs4EAlc8Q8AnOQrZDxabTuiS
1SpcZ9MQpXOa33Ady3Gez3AXJIIck1YMe9qJZaEVfW1+AU/gVRI+ovw4i8lO3XMEMBiMk0JRsxTR
8E7rfVtHv3zVh/yMPARYsZ37sXfBWUDvmLH7gT8Dkf0f9P2F9YGSNsca47omrXl5yxuc8v7TcIW3
HqE48WEinWSfqqk0g5xT0EwdolVbXDyVU7xxRN4/F2rjQFp8xXugrdkmUAvqeKiUdUY56hmCPvUY
IaC/yoBi/LJnGarP2OCvb45Z2NiTlxKWoz7PRWQdRczIzjRljkBrJ5Wk0sekSknSpUPQrMWYV9z+
o0+FLEr1WJ5bKgYT3ehVE5Fj5eOQx025r3mcdSPHGf6OxXiMR1ktCFiqvY5RcWVgl97VO/HT4FOk
vhmx86eoCVnEsA5tq31F2Lsn8DMlUNClUSPk6CkJ7TcDV+OgsEJ706puCJ30inixeDHpLTnksrha
u+kToMgtCiq8dbqK4NWm2+3fKbUf7K/DbAKP8LrMemkEB+btUk9B9QgSHNzwsbOEeh5At3ir1r21
/fMPMPz6bTs9TXX3JVo15ChDl+DPdyU3crPINi4vgbrRhYgKhk8+Ms4Ws9ZwAx1e8Z00lg8uhIBy
I5EKOdQ/KQpvfefGy5gKTOYGkHPa9PLE06Zktanu+7NN9Wrk9vvhvZOnjSbXnL7xhE5duzsJzzXn
Xb/Un8vT+r2DGyYqoAstGi5x543UqslL+W6RVH/OWpRswelYdm2iAJDVFPj27qesnB+1pLL/YCNR
mSbS6+CVBroZ+b9nGm2X+JmgYEzE1EuDPE3wDL8o0lbkYdcVw3n+H6jv+3EvUcyeDMwq7OX35aPW
lutYQBNFSd70tFs7aWzEFODxY2XAe0IAOQDv+DMkUwnED5zTCcHYt3Pet2XUebnvCsD7XhElKT7G
kDFrvQgpa1j05QeYCf/aSem1gLQBw6dh4cNKuRxQKTTVq0jL65XZ+Gi/k9tEU+0mhLruNOVtf/V+
hbTwnyY+iimpJt64+2ybAUdGPKG+YoAYvwHLAMK3ZfuKPAD6p5n9hIrmsSesjvjNG59vTWYv4jxC
fkzRNPAAjMO1QYpW8M7T/8kjE+saGeHN1zE8fcJSfxgsIEE4TosQ1UJAx+JB1LsqZEVTmHcTs8kh
H6eHm25QpUR5ietFzeqFHlRl8q370ekpnZQBZhyJd1imCKYwRwUnCL5W/b0SokKvgZ2LQaVt7IR2
Bok9jsiZV8tPcR5xJoM+0Olt4waFBnjGbGgk96IWOycN1uXPVVGewBpaoe3nauxdkziOtospDql8
TOLVpvWinLXahEyi4xbnziPLuXe08crNnO1dIKkgnxqBF5GuTW64V9MZobvmwJEpDgQZXec1NNpq
++i56teob67WnmN9rKnAusbh2K7R50YKsFUCaCzFu1vzigxRd/XX74yeGHSIc/FQOyLOynxsd4T2
xSK+SAnMhPSvLKPsbss/ZYJnMdULAW/UG09vA+FNqI9siT9Sb/44NTe1H75D1u0lzaRlpKwOGO1u
vi6EnkEizH4re0CzKPHs08DwMfvDPXjLthPJVClr3fKaNpGybx3+UOSRmUGyXqC44RqEklKjmu7m
WmYl9TDyfd/euSANyroQpYiWSktUmlm8P/hiuR3cwE5BWU/6mhT8aaC0GmSUK3/L2ZirDqjh5W+6
ghsAUHJsoGPwPwBWhw1DV/nJ51CWUC5zO63rknTWmcajQUb1qHcmAefAe+Z/I+rF71mClBU6AVh5
xu4bMs+qMny7CX6u66MxD+642KCjV7anm527lQkXFhYI7pGQlI2Z3EUwcLBZNsYTMRzbXRgelD86
2+i/Xr2Zzg32HSii+v0tLMT2B3GMGtjv/iY+jetNdJau7BZ0g9/FbwwupHd+1AZBxlahJIaZ3VqA
dhZBVfaOHq3JFt3GveMZ/IBbuUiiyR/ogw32PCeQm3gvuDpQPrMAs6paeSvqGQJA6K59LMv5zZFq
WpPFXGpG2ULFZvC1mIkk0C73/tosXvnVei/ZpRUJrd3YKQfjBMxfFSuYRZ7R9MJt0fXhi3RoVYiy
hHSxD/YZe/peu4ksyw57SitZhtAEOKL5ocRGyB1Y/VLBQ+M8Zh+u3+jILi4/3JsFVpdMLMZ3i0JT
4pMQLfCtcO35Z0aNasQzKls+ELG3quSsYVYCP88ETOZSDqs4ZMzWRmbTmvyzV5bM+/jSzTujuNab
qHFD+/3gL0vJHmhha8YdTrF8Kg3exNPpp73kYN7GewmkjRyPq89nXK3bZc5DFCaoVTJBofLtR8pf
GzYpKUJIofCYspzQdKl3g2QIJxNIhGJlhuFa1B4G9hbYMtJ1PKWDuCJTJ55isy9Grrml2FagsYq4
/6DIsmk0FPcj3V4t2bLSRYoqEfMhf0s5hF7n9F2Lq6CLs1KoBvBkAbqROL8gGM7Y8f2k8G+ZGAm2
atBUmpR2bj0AEsN40CuaLo5sqTKr1AK76LQHS9UQu89pVG6yKqtO8uyX94wlbPpNZbldXpirztUC
6jmA9VMQSgJnWcf1cIdOr1QgfZfdjShUPsm91+lR/dogfTC7e3VwwanSA0KtOl6iWV7DWPHmRKIN
t8aIMC4NRiQP5+VJpucQlSQ+tSs4Fcu4tW81++wzv7HA4WFwSksPwNA6tMhxGml56uMmwTAjCiQl
5YSgbI5LyFBb8noif3rw7czAnWySwsoGncE1gLl1D9tt/QA3/Jq5CsCNghyInQoHLyXVwXBfWtd2
c46IKfQ9/HMA1Re6H1NOhWuXX1zBT/60JYg8kWjWptMA/4dwzsJAhWjHxIvFeE56kFB5la4ARcvw
IWDa8r37C1z6OZYjhq2oSKu/d+REI7Ig7Lzatx0UPSGL4E4OW84kK9gA0EAhv3It7gqzNy3SLRrp
K0PB2t2X4v24pAkIN0Iw/I/B/8QDCfHY+zWcyVFuPIIFvGiflQXNXYoUg1e7AJNAh61zb22i+lGD
yk1hEfqNjBWgYpe5ClSAzs3W80nNjEW89uu/xvikp6z9CbrlBmxc/XpkcQDzQbyjjWunK2LrNLqz
mts8k5YHp2HcSTqu/WI2X4nO9NbR6Kyq/+xhhhLOVLz6Zj1WVwO4EH7IZlJlM51I82SjL4gw30U+
JRW3iZPNdssjCQsbKQeXV86kv9hVnQ9HXTLW8wETzeLiqP6OJuGEz9l9yJuai+6XB8ik77MclpxK
gjPVCQSWWJbMRJCQnBbbpu8RlMbJlcJAtaRA2/4/8JQt8o9JLb1PO0j1pJHsen45o7iboCOB4TqV
nghGfuxCHLUU7M0n+uWiWu7RIFVEJ/D/e9f6x3Dv0w/Vk8JKL3VZPorNlT+W3ZKdzx5dqWLAufNE
UVhuycc+wKrMd7O52OyuthOTtSOtb8SxPsABtjoMT2rh+3SNqhmgARakXazY4PS/7hh+83o8jYT7
5GLlsmWdnd2w4Mk99yoKicw42GAQuXE2R3xtL7fMIBoc3xf86AI8AIIV5VUuNymm4IqGYoCWb8Eq
JXZaxbPLlMpPcY0EcveUFyO9V6YaJlXAOa5OXqbWbRiY1eZdtZYnjj+Qmp1BiZKFMnGYXqzRYmtr
LOPI0IDdDPs6dfS33pCP7ro1Iq6GuKdmone7nGi8OQYScgtuVZ5uLIdXKNvDCKpZLZM5vUA8a+RX
JqrFKS7r3wTgn/0UhsRwgLa8QHq+ON19NcF9GOJ8I8G4YQ59OmRVx5mUHO8u88FIk3cz53mL6rwr
zT9MALjIXl5ThWRKeE97okaqzI5LUKUEYKa48v/bZjuqf9tIai4FpiPZUgb49de2qzsJ6x5TJXjb
J3FCT5EQhUyoHG+fXrX5MZQso+egScB3hDmLj/2UYl/4M3keiGHjSDkGV4ZxfVio0If8WqzEbuBZ
hgqAL4qD7xP9gLyH0DUTWf51FrL5ZLJ2tA6FOlQgSCC412KEsjsvpeTBelRlDfKg1cjk+E9C0CQX
fBfDd9nWWnmY6JZhTyp2BVYVsk3UvR3/LNaG3yIQjrEhnhnv1O5d+1RjhV8kMEMTTmIlhlj3DinE
PmnJ6n0IQ8lqG4G+98U19iPS9lATwsHwmSkaGk+cUVjwgQxb2l57+ZqS2XvtGp/Jcxzqi7PFeOOg
uooZuBhwbDZzOHUyiPjYpDG27hQn2DoHs7/Yxe2xJqM5yhajVgECl56xsS4musDp9nHYLG+2aJyA
/N9GzV8qfrkyX4btpuB7O+pKaNf3+Lv28+GeScGTjhK/wbkkxOjQeBLMGttBZgLoYpxVDqEADyEo
xFpFmp6vy+TFJzp08P1+6k/6MxJOjb3KEOnzBzZYhK5ESQ2fN+slgzNRnMd2jrwt204UCOzFRLNL
WZS5FOIFJA2fKREgfnhlKQNyoHaVWWinm9hZpuaE852aOUvTlWaqAlWipU093H5hUuh5BQby8UnG
+txhmCjVcSq8PPPhBsfjGgRKvhXQxGLRnuNexWraX3pGXoah0nXFIaOWRx/P4JTv6VCtkgGx/O0w
krK4u8PAKleCHx49OBkbnhjHaTyHf3b72qc+UQk97NSnNuoxCn1TXU9MLGv0VZyAEH0Qheivp0+M
iYTtm2TrMQg+Xci9uv5dxD1+eYzCEAKq/nw28swF0rG2Ifn+vhPOxYR6gkiNlSfXva0d+ZZvOvZ5
CvNKw1dwdCkDixB3Di16o452DIgGjpdFZywYkn/3UdK2G2UFs//yLAzAX+F4ftv17EZtCg4eSUAv
i1nWy09AWppAgRIIngTbsR5S3yyLjipuWJOglEun4rSiwWUgHay7xbVJab4Ip95KnJk3fjwT2PAm
mWQc19ZkG7fLOBn734yLyGdJ7DfmwIQ8FdwAqD904hCAKHrt3aNm5RArtvgz0W9BB1jxnzaCGrW6
PNt9PZRyVQOLCDIsFFIZNyyyH5sjeI0Y9Jm1L1VLRFV8fsiArUzxT2mZZCQHP8Geold7CzC7r0CF
6NG82UWxO1t0BtUxFaaAyzUU1Z4/dlJ7Qq0p4T79QW+G/PgswKK15Hk5AG/3mBmJIe6CAgsBFCMD
twdiikn6STQwGns+x0i+MO2ZXydsQgxJRmeSuHA9w2IhU5MK+xAAnWENfSHQMr4RrfOiNcYNBGGU
AkDSX/7Q5ysUc/716fCHTtadieJ0f+zapL1eVT/lI/8ue+eyHEdIX9OKA3YbPilMeNrA64W54/ey
RX/pN6LRalHpH6xObcuhzNeWXHX++tWGUvOB2ELb9IWF+1uuLYX73xGdfqGppd4oM3vn2DijmAAg
kGjID4DQvUktnbn7sbYHEUQCMcoAc3oFa31loMzcE/802hDf+LK43JmUsTs3nvaHrpikzHkAmges
Xsg3w+pp5g3i6xuQ0HYL+ScZ+hZZT0mZdJsSaDcFVyyD5L2IbH8zyxg3Ppbn07gAruD50uTvnGrM
2FUxqE2YwAKSWYnJVZPi0geNe6SRY7+FRCAk6NKacatVyE4kqPwZMngl+L4K+TRjlE0dDS8qrHtE
TzTvFuEAjUT1NdgDIkzeU55g7a7Kwr5uorneW82cH8bh4oeVLurwgRs9qYDbMPuXc7JKUHg15ghY
0bL08MZWCUoxF/V2BKaCZ9AhSC6A7ZOVzHGbTP1oco+WohZpCQ+MEzncxd/nAnOG2nckK4eY/Oav
mSuNMlOatRPjw+OdOCU8gSIELEi7SFEAM6cP8TFivtzs+M3uOouaPuqbAZZYDMA4xQM7qNGfyjUf
ox4J7/FnYVtyy/L6i7LAW7Rd8wwtcOsLGLoUDLtQCivDVRSrhgfkhzaGAjOty1wH59V7O6ADG6o6
/aajiqsx3bDPkxRRzy1IxaG60eMT/6+KRPAKWvanKBHami/cNvz0y3jPeFcczZ7iA55vRZBp/O7F
5Nhyi2lanQbXiAZWqFnmk8w8vzi4Z/zNGUST7jG4PpkLCmVT4HEjKJnT6HuZCwMKQR4vlXeB4QWM
9FZgdEqXqK00KNhK4VoieoU4pIqnMkx+tCuo8tXJPtUmPC9jx/EuQ3NkAEQnDMVUoEi406E3pqCd
DiR4GwZy0EoVzNajBQDPz/EUnia4WIeq3QyWgHJHibqo8sauLO9e7D3JxSLp3gPvOwA5KQupEYxd
lr0dFKYydLdvZ1XHZBxHTEBT68ZT7usy5A68D3K6deiN5ERi6mSqvEGzxrDyL/vLkJoolb4eivmd
EZ/R/Bq6yED0g4DKhymNCURnr9Kk1z0Qhd/i1eFTH4+2jLzc3a4NOUevnpCAY1T7DQEt7EvuUzh+
U8/TEd/W6zNHaTGk2wY+/OmznAycLhRpTB0lymzVCrCn+AsdJWrEiyvYRfUgkLAmtszSqZZeH8/T
wyNViOAwpBhbsIAOxPTj582sxIw/0/WxJG/3nbzwQW/76m+IDbu0HPLwr6RrW0gxzUMTAfm78mzl
sR90h7HkmbrcAD3XoK1WRrNl4Jt1q0rGkGAKPIwXxxmt3Vo6mVBKcVTCKwjN+JN33U9qPANtaZBG
yBB3zj/SfNclbLjCwtz/6kBALz1stTguZC9eotHJP5wunQBnu72txt8VGzQRdm2WvWcEsa8rwD27
nZsJluUHvMvlwgLe4Q4w9Im/HtIO3obZDBhD9euU95+idovm4cCTkijIdhqGHTfc5gUdTBj8PILr
Z5AIYNWcnmRlY/La1nQKqCbITMIWjGO3ZfBrHqoaNRwBZda2dD40uE4dxA19pPW/wAe98GdkPvKj
rNUAzli9cutFwDSn35NgZqknThYKQFFAG9CHe8SHr902TU6ouAIPSf9LXe/4Eolsp+u5YiQEDs6Z
XWyYbWGnXNvW+I4LlSRr070a3sPuJ/MODGSkcuMVRG5t/N8XMqPhl3Ee57JYRywzPEhlsVQTo8Zq
SwzWH/Rbuj/3uEsPLc2LRf4OXUI6wLR5O+7s3RTS2vUqfT64e9SxqSpx3HhD1Id5W2SUhjB7WDGe
OSt/o8aFp4A9RakvZQSwLv5hKZjOyyiAX8aOaRTguw3UzbyJgt2JLDhVwndnkz+vFGyrS49EigL+
GefotvkTqP7L0b/1jFpvXa42KUn9nS4U1NKSwfH6le+u8TS/BOc50Xobfcz/bJQyrSHgKh/iAi+v
KA04It5vYn8AZYV6rjPc0Lr0TlrPv9t3+TPjzMevObtxPgCf1C1H9LnvS+oSoGvzc2GyqpMZ8VZM
QvBH02KoyRBU61OqUnAs1y6NawG/s/pWm6iCkoyWq5IGdPl4Dg+oRoDBBedfl8txi4RYD2EHelJH
AtesdoTqauewxMa+uL8bq/FIr8COKIjN/g8Q/nBigzblrCYt5Yzvr6EovZPSxtX4C6ZUyaQ1voDa
pjHD7/iQ8m+30a4dVlaozOd8w3x++wYDzD2ywpg4y1maVkt0yJzFgq6sOpsTT4pi2CUksCUhqLJu
z8cIcnty/u5zj6mOn3lgi2At6ePGYHSO4MACknaY28GTTUdzip5hy7kAYIBjFUAmECI8zEo1KJi+
OsormMFoGVgvhD4zc7oqTyZDpHcq1DW9QfCgy3TB8QvpmY8VSKsu4RkrLeSTzvzib/AAt13xdY7F
DVAQTWKLIcGf2Ib7sIgQyM4LtdaZ8a7PB58PM+Nq+cyTksKHWXi365We05MpdZxshmJu6egIFTdk
WYvSqedT46ul4KpKFexdgTRRVWaQJPW8HwQFDKVya6q9BQCLBY4Gb++I/4VCVFbHNFlb3dLOqmRZ
t51O2NP/JlQrKwdWfv0q55QCT83baSaLb9UaKuiESR7PfOih9iA6OvRnyIdYzFv6ybnzHggd4iV5
/bj13x7ebBi/DICTzT/SGET9IK1DhNwaNpG/o+tvbmUoLT/ec/0do0+qS5A7n0dnpFTtAswzRGa7
uwDkYRB3vPEuVsqs8sYDFoPDxkgaa0OfRaxIAaljzbi9XJJm7DTeKnQx6fuKyzt8nNVSh0AX8AS6
+0Vd6pMEnY9t1qVFtatGc+GSg6rpU/U3qzeiofwxHJV9DS+yfCvlrawj9iaqoV3fjKzNT36lVZeb
IqsmMa/3CC2f+EOSBgVrCFKdf+tGgpQQqlqooTXNWLPis+aXNDmkMJAB1nFlnLsQrE9OoNUC5p/k
7Z9XWTXVCeOgJXneBPNjwBbduqQIc796OtGMPdFWyitIpw1dvbNO/tPMXOAznoFjH0rNJUvIWRoJ
wFxYdnzW1traqh+QV1ekIYOg/WQxFD9uOMV/WLTZbbo+RBw+zBXivDzir4Ep18Qz3L9gP1VnmLKr
0jW23AzLZtlfKxqlhm85Dq5hprQY6Qr8bRcxls1y11Vk7ZpHi/hNxokxyS7P60cwKnrBy06MnYpK
bT5xu5ik63Loq2EXNSggqaLze3NJTnYLGthLC+j9SOxH7IsyDLjGyv4A5h2SilDLhqIsyfUFGTeK
GPb+fatEN1gH/SLvZzd/f3RRc0LYG2kBktZ4QcV55Yb3JG1T31vd4u+5Peu8Pr/nCn65kCBgyqi3
7OoGuNWH10WAwILaM5x1c2mclAU61Nz4f/5aPQ0JS+8UIoIn7Mz+hW1QNivBaSV+J8FpewM445dW
97RXB606ggGaFznw1r4ixTWZ+XAeymH/Fi6ClOql5ec/wAHpmWvCEC3jLxZivs+RzIAD9hnK6yd0
b1KnKxUgKSd3KEUIdKRsKMLT7WU1pqITNAatS+nupPb1sJpKaoWbeaH5oK9p+5iBA3g09HvXuopE
EkxNzYmrZDpiEy1p6/j7Y9U8+D0BaeoKs69QfCa5Hdy1pFIOTnjzQTdKQqgu0lJeGPBvzeAjQss5
rldAInh0pl3MzSKE7nf0aDQHnFvmHxGvTdh+cvoGnWyKsaO6zVXo88ENR2fLv7smwxcqInEKMc5+
f3BGzCmb+HFqWkdHTH1s0hWzU+TRjAJfyK5Q4t4brIxU1koVbF1YDJc+SaKVU0lH4VnZNQ3oPFzY
uNovkP80N77OAF57myJ28YI6Wae70QYTDa4GQpabV63sK+5adNMaoBFGQ8wwlgCxvUOnXds4E3vT
RfVmiWl6JcKP4vicJtfiJHThAYpEJW4JYygiDfTOHh9EhVp5AX4/QgOU+t3/V1mKEtMQY7R2s4t+
2cgZ0NBvUb0GJBRVWeNyg9MMgsVle6haB4mZBOtg2zsYstvR3TtJ5oh/yBKl0oo7OuN+ICUsysTV
VaGc5YOFPwo/+kR3PnGPTm02rmQFlCItUvHP1F64uK+mKkveG5JwxgRxixwNLuE4/o3uw78Z+H7a
dSyiT1YlnG1afswoU/DfilIJe72Hld4IhClrpUV9pwf6SXTBuJxQbcqpRD6CGeSkiBQRoRS2kS0/
JeR+nEobAaucOlxAfW/NCz27nznOCBwBIavtUVS71aOMr/GuMNeBrfll3YO6H2TKPD/MwfhZfNGJ
WUQq2cprbDNP/kSFYKRT9KQ23WjNzVN2abZAiiSnjHwwHOU92K0ITOXawtVgqmlYT2X/Z/RUCR9n
VmuvI3Rv6x+wDD5MrMLYjTIJz1Dt30qVX1uAyI0cCU+y7itLunhkjn8D6r8idUaYxEZDq9Kio1xF
vCBogLGXNmcs7PLu/FjXKVVs9s6ent/5vf+j4wkrqJ0z2JLYb9DCkA+HS+x0jHeA9oMLOb+G0GTX
UWzy5UA1/hZTw0d/wBggx79e8yKEddATCk+gdo9IO/iOXN36rkNMf6xQNjEfuYdb66itDnvQx1gC
bmUJdUR6qZo5qBb3RyKMV616wfM2mw5KesvmxkYfI3GGVCHFs0OtqjLTvQ3PR9GnAhnEVZKJrnyT
KHEE8zuZw2qyv1QdVQju0x8NNpwRk94XRoh9HZ4HmAj7CfPiUmbuRTyC69yZwGjL/BlB+6qaDccW
p7Axiv0o3zF9LrD5kMOtZEKatTtnR2exrlLxm6WhrC7s7ZsaDW4wl68bkjCSnLvfODGoErwkuppE
JA/QiNDVG44YGDSMx6p6LC9qarJ6K2b9SkBEpL4HY0m4ACwfmNufdbOFemqvFCe/hHuy4zID8e/I
BD7L8q78D1zCVexyxPYlHMseJ55fMxUapyRAt/6R1BeHHnJxIoTVAPrqTLtPUhmai/uyQKpBQEQa
negN/Jq8mJPfKuvKSOwebMu26Pcm34xSIDiJaDMgsVV+cqJFqAFLe5yZdQ2e54eQYWt92PW9tmrt
N5j2VBAItF/NhO8cayWoMk0HX3JWic+bRoDXCAD91bZoYyMg/qAwluNYbK85JOORiWX8ojQ29oJC
hipNScGD6lhzMZUSgL2hNILRFwCJg6BE722iHOVnWTlQy0Q4Pjp3OPovd2ocI650nqnZw7ytgny1
XbRoBv4lxT/U47pBY27xiksSuhzxMmlzsTDfChg7Fevuftn21R8b3EZuLOTh2hvmj23dM5pDjqOn
Y5tKzMgASesQSP4qZJZHvpzQHZjK0VnDnJ2bf6bSBViAtACZiPVIAp6//2HNYI5RcY/xoyad9Vln
uqmoFq/itWKrUnGgqimWjAVgZNjF3FbfmjjrV6L4ANiKuw1czGf1O5b+zn6JBL9zVp0gQggv33vf
W7zqRHAsuGexM6WghzgKhGYkeD2LgY000lWnoxkMXY936Z438mJEUJxMX1fpU14Lg/IRnyZowN1S
vfBlxwbZLxbv46BME3joY1OO31bWkLBLKzgZCRmhdZD2DQBrSQx3BR5KZt/YItjna3MeAq1kjxAN
sJp9/uFO6rrv7fzNY3xYJtmV7PR0iG9QARLngqrVqdx+EU13d4XfB6+AzXUD5hlLD1f1P8o5B7xT
68E/HqSwR8OKKjXdFebZ4fOi7qDQt/Wf/rQHLXg3AJ52UYyGTBcY98oG2bal5ia9tirdSXR3R8OF
dMw6hVpJ6WddA2J/ayf25TKCNg+VInARsxht6ATgxRGzmYVMHxIu6STTDv4DujEIhBDBVRmTfdtJ
AN82JVFU0xxJ6wUuTm4oJ6ydu/CAgJs/1+jLvlX7A1uuVn8Q4yx0mMa4cNIHVtTe8asFAZXxU5gP
pFNkOyO0ZaSagX0Hz5a3OJ7lykVlSv5YCw8jPFdnNsK2AL/zMONuoTFKN4SK80TuP1G5GJr48hbU
NYM7fEJSqD8ehmh8o5SKM6bm2qb6Kxr2g4PezGa2DmCeArHPWpAPVx0HCmDYY9ND7JEHOcrZCGm7
po77REvV3pkwKxISLroSKqpMvMv2OkxIhaC9L/bNPsXdgdpYNqlCD8nBIbAJOKk0crA6PJ/h6jhf
E5MORN+Yo876lC0wZEytBpRDOBSohTzwFQodmCKJbF3Dc+9tTv0GJ8FAspGRkVJZ5z92xWTqgWsH
rDLjslojflRvjX+wNFqpQyVYQ342CvXC+88zwLi8EOOv1EA3rCmAe1wjYrViek7JYfULd30g92xB
mHYuQTGU+hUGdl1YGZi6j55R3H4Y3pY5MOFVqLt69n49wDlPN0nsUyJmuKDtB7auPufcR97JmOWo
LfhIoQRLM9B+/lj5XQmROl0rmvzE2RRDuz38wKoB1A9u/B+6vR7T17sADcwYFUt12R8DAFQlu8AK
g3UdHzy1x5H3awM1aUpDhpfWmT2P0FozY8FFXA9W9WFj/s6J7KOKnX43j331heQtOLGhfts8VT4j
0LJKHELN+pT579W79Es67MDvD1rtxL3v0lkeDEYJJo1JBgzRonGqngle8RH4mkoSukbltEK+rb1w
h6cg5LRGK6nU5JSp6kcqvn5+uykyd8oTY507V/iq3t/7vXTjiBPMZkC6bOuAd33d/85o5tkbRRvW
ir13vQ3gkAQDlXhDoPosdVgzKr/Pze/oISLIRWlynmy2KMYQNmK9rAdBUhxeUrxNzg7h9PKgVPr8
373dxiVF7itWa9P6m3G1V4kWcixByxE6piVzWVR29hUhqEOQ/mkt68ureGtSg9jfVLvo3J1yOI7J
yz2f1MSRx/r069hFjUCA/0tKUPQS60lCY/Mge94PQfi+GryZ3kbL7kwkYhNRbjnbYa8Ow/VZD7uR
tL44Hz/eLWVfCWhKWcaBFmBJOThetpo6I0NpQRj5nKY4/ilUWUSDiZnU/R3GB5ayg3FfRBMs9Ye3
sO2LI0zhYZ34g0OsbJdtKdM3H5myzLw4nlnuffUixwNELoUacreLe0rW3bxmsnTU81EO9u1zg3Wc
Rk2HK2wrpV3emscdKClu3T3N3JSRkBnKTWuwtMhard18XYNflAfYHLNqMyWhk040Wzk62N6YrHqS
/pSIfJNEVw2gEj6/wXPSBUb6H/rn/b8YSUHf8b9/bklBvpebLji3ZLqxi6stax5Z/GWfmfj1EUX6
7QePW3taYROV4wHAMUoiWr7Jt5qddnw2Nh5qWCXjUstNsm8ETzsGZuNnJVapM8TCBN2emAz1vevd
Qzqq7hklznnU94gos4/JiI1AaSeAUvB2uHXE/+3tkfS/ZSzNpfyBhMlA8FW5n4HVeEV4dCWVXY98
WieQ/vT7LIC2AGVBaqBlyF+GGa99qys78nOX6ph3ZCcdRT53T6XaqlXsOz2Ps6c3JBsNcEqTQ8MQ
JmKCnbvHPeJgt6r1dPWj29T80lSTCwsTkflto5wUd/spOvGCrid+IIV1NtMN3yM/6ud5IBT2/JOF
Si65miHc8wIPFzWZDCafJ+CjQgZPSjOokX4LLPp55ZEXHKaw4ikX3ybricAbG0qO+CfKP2ZAOsbU
ltuhwDVuw0lOCki3EmRFOk6oN88xgCioiSeO0JZNU63/r2nvKdvRCnJBgjbyghwMq2VhAqflw8eP
crYpAsAkkPHtI4ewoVQBXjl0qa/jkcrCgwhm8/uhsvA4RsUukUxha1GbMnMMafA/ZmEA2t5Axe/M
u8lT1LHvSMjY38AS7noRjNbyUorKZ2WsxdhB7INiRu1fo20Dy9tduUjRwv6fx4JpxOtZK87WPMLd
1tibdLgBlt0umLLuuFaDIRFPPXITprS6k1349wPMXnTGwmTxFGTStFYaBvhHwMuVyUeH2HcPdvx3
vL42aPvouYLdPs+5MPgRuVZzXD4pDLpsi9gCNIrZhvpyzZ3ZlxWvNSFyXp893MLScgGnFE29wB/h
8cuB2hG7xmTQBLZ1Poe3DrhS3rDoHZl5gTd1OmPy96ZWx0DtLQTtcZ7d/myV6+D+nFExAf87/DRn
YB73ZDIASxQ7Nr5VCbbzspsxFLZ3x3WPecqRR22KNuBFFSJQr+7SVkyNWqszw7aRv9YLCZvp4FWu
Z0pf1P5zN+iKGbvU8Qyusf+XyFsNEdCMtV0Ja705tLX9QOVR47cu/OWG+IbhJ4M22dUTmz/nA1cu
M11zVTETgDdHf86I9AKjS+eYB0NYagYZu//nQf7MvPdy8TlAXCD/l3NGcwelAEg3rARotMe/ddMp
sOMlyK+pPwJ5x5UptDfpRKO/i7hbiGdj7qQ8S0v3kY7R9OmXnY6pV+MyPl51kq8gTI5Wo08UDkRD
sVVaGMMnEemJE7k2n2b6/eXnhL4oe4K0pH2sFJJjV/qdVnCL8VDfgDGv9hMr1qvdzRlB9NEPhWSy
JqK0ovJQGiKY2lrlxbl3gEx1hGb/0cLSaVAy1w/7ON1Himo77QKU9RqtVhqBHDxUuR3CmBUhDvUA
mXmqYSXHKFvZf7sdo3LApwRNl314hVMJpXhC67sCi8YZIo8n+I2paUb6fbvgt7zg/iwAEe6foPBh
30Zn4h5ucT3c4NcfVdd711J0/WSbDE8ggaCXrl6ezIjUcGa/FkLRmtJZsEstuFF8FRfG19a9wfpz
qBUUUvYq4078Ut3UToko7lBfiwnYTYBNCU/xKGO9hznjDSQE90k1vLbZ6xauwQMcdF5buMUH+cRP
yUvqdSsjirE55j9NYhUPqPDnPvepJCVmIOkkuUqQujNAzGxwPdcu0i0wNEUUCoMx8sXiXojpE6YS
BWwM6EAm7fu6pf06R09NVq7S4ZA5NQVCfMth4rZcAWiwYICrhgOaKOgnQwGby56o7r/wyovaZm7f
LhpyWiCMpZiH3xl6d5z43WHB8Uu0wEpVsVMUNj2cXVOM5/EVt/Uh3f/I8qlUMj9ktTcloouVA8aT
ErFzl4mcvhWdgvjjTXYgqs0BpbrIw9T21Czago8NFMQ+1W4BhGxXGYOsyn5NKpAaMEbZzvHWZXaK
E6R58qcbL2vyywfNiJzVzaraJ86EYfPlwhhYjhMNe15dF/tzwHokACaUD0y6vReGT257ytghO6Hf
ti97NOGuTrDt0XBhY4DIehg9uThp5/63xul/t1Lw3Bon8nEH+HfmPW+la4u4svUXlK74Wo8Vr7bM
cPHxG7T9Zlxta6VsHrLJzUPXfXzhtzQe/ckPEZ5sgu27YlOwpOlSAGwuSAcRDPkeh9s+6XGUm+sP
qbQ7duyAMg2uWc2uKj0Vsl9h/xBFX06wz8k4OjLN+DTgrTEcTqwkKSaRrE4yu12xhOMJ72/MHp+s
qXt7cRJF5I0a17h5ZOsMdLTy+kCvRrwl/zeMHVTMotIkkgVWpfzFuxv95y0U7TaonqCkeMNk7feA
ZsUs7nM1jtdkzC+rNHUBF/5bkrhyRjhrssoU2sh1ng5g0/T8sHDmkRkHYNhyhtOWNjjthmbACIQT
tzknLNWpZKApsu7l/GRaR4BozRslvmOsQctWmjmhWpweLEUWQ8jdYasT75JkOUFnrD5WQoCmLulM
6xJ5+k6wkeikom8lD0k0yzhkkd+iihdDzdzNM3ToakjCyg1r6YLm3sVpG6j8Fo+XBbpiKVlmw9ft
H+XShyRcfbjgP92JucW68GrhZcLFb5AJaEpyZYFsCjSrdeUWmUKsLMeT4u9qMYB0NwadXs9A7bhq
Z/XsY2kjkATzyg4TzSQaWG7U4JNGmQNTruWCpU1Z+ocizT/drolBB2xWRz4RILhm5LCtkS2JrOZD
kOze7hM6xyVRqQ5eEZPs2ewSrXxYNiypQ84eIfRS0lRWSYj1Xu4oKKp/1Vc3VbJqJnyRIIcxZlro
+EoBevx1I8VVbb+eZaRd+WM3qgoKhxzAFBaoAZdQ7+6rjjU4lvhB4FZS6juNvUOY/UIU5JJpM5wN
h8iagcnKzCy0QmLzx0kzDNN6BfghhNjhRcYpIz2Zw313pDo4BoxNd+ZNytOjSzryEvP1SwOwF+dX
QxFyjEteae6EMjTQukrksHFtGNFosBv9QeZLCYCaUtZrL4Z1r9EFxHN4wWNUE1p0V39DJa0CG571
X8VwgvGMR8Nf2qdpXW/QkfoyquiM5NucoJNG4lVWcFVRmKS7MPr8fxqk60BrcvzZWRQD+FKNJj8R
6Hs7DnqnYW9LmqnayxxokSTunHNvpL9hxaV1OrRX5PTXUYico/ckBq6/ikhBLmFHsmMUkKQmXWmo
0S4A78kTnTy/x5jLJ9jtCGmm8Oyuu9LBAvTsKxDDDqY5geBHbjTfffi9PcHu7yIwOWbUsW34yCOc
uT3FM+hqWkpzoE0u7sWjbVJcJxRP1ownD5Qr1icxS47aXKs88Wd8pnzaiSwG/cFgwMqNRn+Tg9lP
428UoAkGRdxCnlgnZnr2VNZ+LyiUNxb1rH/aQIe48CtddPE9VZeLHFJjvvvlOeoX+w3NRmgkdoJg
FnZUi9o1oXd4JiKPrrzXV//p8PlGf5ZizSQSFeRt7RLurhW4wbVm54fHNKfilgDLISxYdWZl4beh
cDRxPgQkQQQoBSwRuRPX6cnwan3/CwI+C/xOMUldKdbClOApop2gA0BHszQFmOI82iFa42lAB0lN
5oAdzuArwmB46b9aYQVD/2WO81tHkUwL0S8YOasdt1i/EZsKz+Ohr9cvIy7AhtG7qfOVTmAxgnL5
6G/Jmp4jxokoL7VwGIyOPgggkuAnpwsOVqtEt8cKQZrXXgDlYXc5yTj9fJtJTEZseFTGxSBSE7Im
LkSL5ENHNUAuKnQqJyLvR3g1/e3HYTdenaL33ykChIUil3CKAv0C8l2X8tQyzSsRN4+my2U1dLBm
dBF5oF3C0ssMqB6pBgesABts0Yy1Um9H2sRmAiqYhBGdWPumXutDAYzcWOupKey+qkfTr48q2rye
Zx8A6W2ClDKPBzVA2na4TD1PoI4UlqqDGSdCLna31KTNc68Rygxl6ePPi6VX6VT06om0D+pa6aBa
a0zDJySBxQ60FbDxcEsSRlTrL0bxCnDTqbhcneV3gCZn/27BXQr7P4hHTHSJ8J+ZQWYO6Peax4NN
O1eheBXjEon7+PXBAdQt8UoGLoNzo89AndPxrD1MaJ34yrhc03WrbuQ03NdodUd1MvkS+Pb03G03
8Ss/fvlZKSpXg3dNw2GeSX7sU1uE1UXYvCbG7pI8qv+iWyv21nmbRXFFss5+gGBVo99YIOHHcbjD
uE3MYdL5iVwDL1Cu1caIQX9Uh6iBki89OM1cCAdwJA9h+88nzoJJgWACrdCCP4sVazadndGx3Lts
oVVF7lyh2GpFgfQTrka06i74f5H6teEuP2Ba6TvnqSLErcOagTzjqFTo4dueOzpjNAGjeL/K/sro
sNsZRSwA7WKjidiiC9MOp39E+jvNmZBEDxDvRJhXHvHhynqO8VQqSirr0Of+tOl/UMrFSIEalYcZ
jJ2lJ0T+JBo3aTIpp0o6OriQT1WK6x4qWEBZFLEdDupt0kFg04D5TJngucrQ2YyRrrgZX8oUhp1V
3tg/DOd4GoFxjBcUvHrQOYQb2Fo+2U76XKPGoHj5eYFlJBot4X0jKqd6xB0ippCVVLnKnNwrNkXD
mVJI9aTC08nPw8PDlcH61D2jbGEnz+qpweF77Bs9XbXkTwagwpN2ea18Nu7V1LmO9LSNl8596pfe
RvaGqcE4hsXOX5azXXTKbmLNhEfzOZYFLZvAYDy25b67+BtQzejKLqctH636Uaa9yoMTnn/Uo1jj
a+dR5IP1DX3i4w0nJe8Lr73QA9XAS4rZd5Ul5rDK8fEE8s5ZJBi9XxThOsYSRQnRBGqP/0WXf5HR
2JWEYGNqQsPNkM6+Gm2d9C+FMfi7nHfoNiOPj0SwqguhgOaqaHKca443nS0Qzy5LjZkqb+1vjwzD
CvgKqQUYqvDLSwdlQdkX2Uk5Kd8M0LpQU8r9eBjSzyswv7BJI95PSEBtssgAHTveSldoPRz/Jstx
P4b4Xw16bm33JNSqCKsdgwLBkvOrOjUO4VJKy32axhLMj6okzupiM8y8hcNErWQq2Ipf8XVGx/oT
ueLrD93NRuJiidSXdrlga9226VZrjSjYxhkLjVF1Al/+Zggmga/rrP9/B+3iJRPduC9xuAyq35rj
aDiWl3ocn7s+NVW4f2CiaZYx0NbENlF8PcmFMlw0TLga8lLGW9a8jNS+Gqs6uXQ5H4h7zeOOflP8
+dLBxj2jkp1Pc6dk+vX+VQwNqktgKyW8iIBki5SVN7xoKMbqun0wxR6q0roQIQMqm1OU/63Pr5CR
3ioMcAPnELDhYHtxgM5zD2m9+82ntBq9XMTAaYKJijAndOuPJjSogZrSI7vfHLPLHuaaCvIHzm/0
6mwGbUrilPRS2AOJJ+w0StE55WcUrmfx+yfTzGiuDbFTo8hN+Sf4fmvoHodrZqnBELXHbbRyUl5s
RQPOTAIk1NI9TavXRrVxdw89oM7CVdA/bwFOu0MBy3ADuvSg/Czgar49ZMDNPp1HrjaRYHq2OwkJ
5zyvLL+lMwDE1waTfGu9CpvaImGYTsE7j6z26J+ieU8ORf2GWXMWQq+bfSEHsKk98fV0mgi1o8YS
00yJkiI9v00iK0XJ3B/ZGIpNyzzcFJJotHl2driDDDQAnrfx419dg4hzZpxW8/mIPo3x5rw12+un
YO7j9iYkcM1sjDy/O8PloXIB0c2RQSRRsp8LKbK1X/QMe241ybIYW71S79a6Whu4vYKDa0xopALw
3FLO4y6TCdyBbRLY9V2RlhzaQScCrLQIjHqHWr+XGYq5rszZlzCmlv3fcZaE0ZhhTFLWImZWfgdW
BZwOBlgJPkAEC2U5PqZdBuLx/JS2HZ5TaoAnB1WHyFQQmqK1hh92Op4g9gHdVD5ZPTER2+c7EZfX
60bvZhj9UbqA4IAPeokTq7IhxPZuMEdC/wnFJ8Dl9GFk6iQNHtkwynf2Kq9KvQSxHuRXEL7AZ/bn
K3bSMHF36Z6n4unAH6CCekZnyUOmgHvGrjPRHEaGtGraF3k3ssEuobE7EGqhSlr4FMI2nQGxumJ2
mUb7JXfoqfRdd9Fx/Yj81f0Vi39dP3ZNCPCTOaEi4Ev56ZzM0S2WEscqBCzRl4cVZYsv/Q15/l3i
1yWWVnksarHZzPuyWX2bjrzOe5elxMaLWkbzoXE9OCPPpfg4dpNId2EzyozT+k+6ls7EDpM47+Ka
RNJ/puwVZC/ahu8qangbZiQK+T5VgA71sfMhMnBzOHPyvdplnlc33/qaselvq2dDWt5+IuGRbdV7
oX+55aiUGZmANzwj5vyirQuAEelf3pQdXcuON3YnVubrZLESp+9pArUnyfUG5DWY+fq+5rIUkszr
ZlEHEmzPOaUAEqoUw3/AyixAqpazdk4YG/xM16X47ur+MegDRNWzuzJgyrUMVHsXhNAHTwUVazEE
WJDcl2OFC51mENwOjYD5nzelX2YP+UybgBGpmGuWjxLDcCGVdX3eGbwzwCWunK9IuGU4J/tJ2Xrd
iDlBjh1WbdSjME15ketvVrlf/aIAnV+CWX+VChCx25Z5TIlmpP8mBpujM5Xt0FnEmeiMrRdWsJZ3
srnlbhz/GmOKePZjT0uoTVDgBEoIra6ea6v0nnr4nYG5qTYQAsVgza5U/k2XVFXtNT1Se13VgILW
ZMrYija8vp8GUoQRSdmI5fN0ezBwCAU5XtcPyLhVAOhDf70tsspdFZ05xoXjnHQhxGE7QTOSJXeq
xLjDuDNVrAmsQpSIZaYNoT6YSLpsfRf13xWapBkitd7cwpurR5FdCeqfTxSkwPrX+jQcEPNKk6Pd
NZaAR924/+C8w1vcWoFJuiU/SWKuDrWNBc+fp9cvAs9yYoL2kAWJHWNDpmwhPIPhfkUHUxRTm4aD
O67fWDSUBsV8/3fq7S5F+rJA1r7ZCSYK8nVHN2SgfzFOrtrWcFkSqUZKsrkbvukAZ1D8xGHQj12H
7DobGPRyekz9iedL7lKD+/IrivmErk8cApMjgdVUmqttXn2Sexu8TJXgVEv8bZv1DM2Qg4oVTe6J
c0DC5guq2ZrRgeEM0UiQVyJhj3RIEqJMZ5et7IAZLI0Yh0QfZ+Mo4iGKoLlh/QoJNoSVY8LekzVc
Z2KOvSUfgqon2gQonJ/XzhufKR6f3xqzH3uploa8PEKblgCELRW0C7GGO7gdJBLMHcaB6lK4QW6+
B6SXHqYvZcwpZ+EXbN1sU5vW5z946mDmv5ITMaGvwyci/GCR+R0kqiwIQ32Xz5tsOQI+COsSLb/B
OUPRpMDcQfAMB9JM5Pb8rQsb7I1UvM9jIFm9ZiouwuqaNJINJ2NNK2d/VLX+xdmSEfRb6aeM8koz
pGEgX6kABrcMHoKOiDjT2PY+WvfXVlTVc11Yn8Gb24wrJD0QWX2ZTZbc2QYzYrdd2T8XsdNvZc4p
qUXycurrsntLw/L+s/j+oA/oHExH2xqjc2SEAYVSsGIoGvWvWnNZdod9oPQjEY8Kn7ULVcdOtJr/
OKFHoURpsOGOhbk6XeTTtnfQR27/c3yALoK6rj3ogs+uMoPB2TraFpszLGSsL5t68i/Ab6xrWo7P
Dl6+ArPu3eZzGdOpYf8Mu007fyVrgUN13pvKd49WmAI06zqDZ4rZqIVi6tQdmys5qbZbmBL1prcq
/Qh3IlzVveCHMkCJYLJBp+9CleniR1NxSw+WACBsNGe3BUYGALSvm2m/vx8YdnOhiMuv4jwvU4m2
Z1NxczFnanMaeTA8JQwoOPF0dd9RLRKjwz5DGH74qHKVA3CMjo0mvH0fzf5fQ3dLPRrdsGA2vyH/
nNQvV8CqKVVRhH2ihBs/IQ83/QXAnl1cLyjqP6nPXQv+KvulZdzPjLuysAC19jdiOfyu0wYxkO6n
JqrbTVMKYD35Mz0Div1eHwTuYgTxPO306FXMTFPscYKxQwebORfbLlpd82TGYwxKHINBzrp7uqG/
B9dJTOfylaAayKroShwSY1YaGQCom77L+wpke/cJY6FiffzetBKsg9Xm4UiS57Rh5mVZM1s1toHR
rlwg3PedzfJnLqO8N1WVxUD8M+W8vNkAcnDDdY4IWu2j8QGla4svh9SXYXfAl7v3al56MOIndIe3
mFKFDpbhBqLiwxXJTIU+/6iCqH3Ra/RynB2yx6exFqJUNgg1QrpyyQ/f3UrxfJzlAvipmhbhbg/8
ck3XAJtjP9eU9lfaLCcwNHnLKdJec3JQUme0rUiyrZHECmmoHlZtIVm5oIeeghL3qvu7djjK/hwa
yRB2R+uigpWQuO3HsxPvR+oSmPzlXhAek4BwoZLBmlMoOHDhWzF0qLJ91NrMc7mqPbhvlPtMTqOP
AoPan825QPmWpWzx/HaDrzH1SwAgH/mTmAkqeGqHiqDo3KY1gPZncDq0SuI+PqUoOMWmG7M6u7hF
aV1kUnRqxllQ73A7X6VcAU9uE/voOanq60NJlNV2e2DKyogXfe0ypWaokJal0WFyppl8ZwAO8EQK
/wwpLwzY7oE03vJM6QDkdcqxbh8/XEwYWhSocXJH+zIbz1rBsXEX4xjThQZ7PHYlK80tjOvSmBcs
QkGv9aKyPTNmaVoIl+oO5vF1mm0AvMOJg0+kJi0dnn0gSeFES+zXcpnTwnQlw+Q4RVkYFf7WqJQP
hcvdJLhn76nFGRSoRYtnZMcAG1ny5v61sLIQotaw5kN1KfPioFpbalmE4olXo2K1jhTNh2Lt3mOR
KPAtXxSmGTumavSWOg+SobQUwTg+GdgVliQZOe8KFeEKkIzkF2Yow4rNsE0mJ10gbgtN7i4xQisA
F5x6L6vaQNbw/TkyARsxhVM81xijfqk6nXd7Z4/4Zi/jO4R/eRzyUdlK/XVGf4YuljhQAua6rSCC
Wd70lmA9wXJhKpG3E5M0pyVL++WQb84M46eP+pEoZYUPYeKR/Ep5+s/meLomM14X0+/UTRhEmy1/
mOFDZ5Nn6bMeisYZ/+ny1GOJO4KpGKM7eCuro9rX4DxaHauIT2nrJFSwRqY5aPfXsySpQIJwedvC
G+2E++L8lV+kPBXJHjp7/04H3E+kgsUAA4aeQXiM9sa6HWglK+n6ZgejIRaYcdiM6ksqhWJ+Wmqa
LKU0yBnSt1Hx/FSiOi3zLtWBSxWPD7gF5UW4nY8vljCQDxNmLAnyefyAADaVklNeVg+L7q3mPxwK
WNQkj4llVvEoQpKLCcZM+mXMIZXPly3Rd0b2pvdwQbp1TJ0gvnCuZVlnQLKTNEnKp0p59Cd1BVmV
QwHT9HvNkrx+4lNhue6/Wld3t/IJVSAokNJd9iJdJxtvAuAUfY7ClwTw+JeYdDUbZj63opeLssar
bXWcQZJv1xvPA5z5CO26CeXL9IAKNa1VAycP19AQ7cK/9zEXqhcPvm84O5nQy0wzKCJyPTprkSlJ
4bBVXH0N1o39K/HNn7tMUd8kN6e7lqgHev3dE6Xlb6467dZpcaI9m+M3DO9Kigbx4oMF4FlPOcXh
1TAsRn61XJW5DQxhNAQ9LLQUlect/s6UgJUSxA2kPWrt04OKJ4p4i+yK7p4E6MH3rm17ChL1xL1p
J6ggReXdV5RrY1IJKzAVmy1Igox+cwu2F1QiaqU51GCaYYDZWOkShj49OBEFfPPDDkD965sOIIOP
XPiCuCc2x1L9Rrz5uQ05QOGd0VcFj60c7+zdDgibKjrywZaQYzbKuHEFGa+l10uuvvvjUbd1VZNl
KHRVFAh3CRznxWF6e+L7L7Y/SpwpmmVR778kjo9lt0K9iqugxUj87ZyXyi5h2n5GBQO9snu+Vha7
5zKkYcVYyrQmRj6992qT3zhkJFoYErYjSutx3gHBrewcEnhaqoFKHfHp83CNYjrvnvjxD38fvmtW
fCW0kHGc8QynUl3d+7DnsAnTRwAOioqsWRWw+9A+hAr5NiVo2JsvXCs/esTHEz51Ny6EIrt5go2F
aN6RsN804d/5BXy3kANWYEDDptqcRSD5Vns+Z7iIfks9ogM5zl+4JmrGw9KJhos6HeTYG4+7HY57
jumTgsuT9uXrlLIOs8L2own1Oxy8WpviGdpP6DE4db3OgYjjgEo9bNgBoz1VEV/PXQOyWTnysGMB
7XR2XFzYbVKckvDvWp0nEdI0BTUe28IjkigU+6pjrh3OpXfttu88yV9X45w/CY1esX/VJYterx+1
4miJHMV76vY1ZzV4Ek+2M+q5Cbsw/tF4ApBaZY26h5WKI+Th9UYRGozuBsRAgpr79TkIaXYHpyFF
VdwSdrjUY0fYnfFIbNTUsXrGPwmdOmnjLZ8j5/iwjofBx0q5hnXp4KZYhT0p64WOCsZnoQgT9dmW
rJ+bTnGNr8FOKi+ZpGINQLKXJjDawwTBe3ltT821ldqaQmniTePBnfzBj5Ku8mco3OCRMMC++zaU
uYPAZUZs0tluQM/vXOcZn9p5tFz4gkoX7y6Vml/uDPpO43/da2/t/jqSObtPyh1fPO9V73U0TYrk
cu9WBYkQMkGsgH9FWoAsIrbK0M5i4udgDETqC3+JW/gBxF5GhRpAB1yhVYm9U5HtkTyagn11b4w0
Aq2GzTuhVs2YoaDv0HAPdyfXHeBJTkinl0NEg7vi0ZwTgGF6p9kkQuIUoKPvi+fxLsKGWHC70v0r
VEMwuhpkBDxW5R/4nDbt+wFzXTvuYxm95FDbepU/lO8CDX8L5YLEIQbtLj3lPJ/IdYzvpob45hXT
Njz3bjU/I4beIX2IIQ5GiEIbbmwnOWs+kRswt99U53vz3XT0IP92LkAhzguydLazsVXXxUgFhohP
XIcHaxqU+A59TirLkbGlMJ0Wt6pVOg+wYpSSY4/pTHF9AzZiCn/89lpA57kNpStuDTvgdw+BdXJl
nNKygL6jiJWu7ttz0zLkeA0qACtgI0o0qzsagg29yl71ppodMA3j//eqD4POC+1dRDM097Oj8T+a
Mq3Mhs/9XYjUcw3OlEOssX7jjEIc/0tkCM6ndDuf8MbEDuzDqle3FPW64as6lIm7hTQbBMBkuFEo
tiWzaP7H29iw2AbRqAsyoAtTEUwnFYw0OmXDAVrierzDGHwcs9X8Ir+Xto7iz+hiG8R3YZ5Rq5yP
N6GAUrWkNABF502F+IxZgqReFUqmUrVeSsLZAXmJn4wrBxHTcfldt47/Mj3fRTsO76K/Vnn8bkWy
/NoqFlgdBn7FDu6KhSqaV7BFvRC97ZEOTH0IlFGeLAujA+2pv7Igke0s44kfdbK4zJ4ZI8vcDCJM
OfezB1a8L4Jc+HvHJx7EcEbsPEzndS/z9upHMSbv1mtzjShmac8tA7y2KtAgdoDaI09WV2AEIgvZ
lIbEuBa66g5v3JC/MU1zADtackfKsauJ8qO83cYkBA3DB9918jJyryZ/GzK+qL9YxzlZVf7Lol66
NZ5NilreXjWNgrJLKdWy1Rqwg0nCgTA2/jhz6/wdMS1b+r4KGlctQUPsIo2w5BRr09Y3kIk4D85r
GbOyqD0KM86wW1115SyKOiZZop4fUk+DOQEzURDfXd4KGp7FKLR/tZoQT6yFxnAeTH/gVxQ0Xvhm
qprjbq3ZCSw/S2hQDAZ4JiAYWDSbL4JXDbl+Bhg2LcHwlkNdFnU6MXqZVu3w1Al+KdXped+ow1B1
xK7XZnyMxkVWvybOwgIKMrBvKDIAUMkihwTvc2KEuIskmgBqOCMX+/Hna8jJGRqr65CxEIS0n8u1
QflPehe7ZlJrNkd4c12fQXZ+QQY0iovSGKVO3hqyYFtmP/Z5hnaU8AJh5VAqJXaKNWjz+BHW5LSz
958ezYIwitxDqF4thAWYQsfqExcfMFKW6Q8CwzhQG85D67ibCqfYgeWrLx/d0c+S233SIFbd7kSm
JqVrnjFCqNOHBft0Sv1HQ1+RASTtlZ92JMylZazxybtwH45qxKl1/ScvaCd+8VUnwhuPBLusmlap
C2dj4PjgEu70IxvzBjkQrq4XQy54Gmbt2XgFAmtLwoDdB6cUSaOaExQFXJ3+d89lwDivS39iTGp6
ju7DJxpNbXhFY8LiuP9CD08VGKiKRSkc+d3lir0oMFeh+KBiX/IG77rTvkzBmmjnHbWMgb9mDV1f
NPBR/SWh97dAmJWoryyw+I2GycklA7VB5iVJftNLNVDcpp8NB+POE/6MENpHRSZ7EoshVMQ2G5k9
ENxwUzraEa6ocKD/RIRhv1oTtX6m/qMhIR74U+27qMb9sp8EZ2LW1aIchr1uLSFZIqbg+IHM25x8
9Vp4TfGFUHctYG506zhMqyv184xVVW7vIb8pNDOvc+JuCwffwFP7jJZqu1XNWXGxLOi1rGO0SILy
6LM9Uq1TU8/EMhQQlkwvTl+YAFuI2ZXmS+Qi629TtpFn9tEim7egXvzErpEUUPK1IOsvA999852q
O5CP4nZttf263O7W2QMqG6pZIU4XPUBbwVGlXGiGOg2SVSkp+/RD3UVi2CZuGlx9QOsCQhNTDXPs
MUgq7/f7WGIK3PYiEe8rLrTEkUuAOqjeYdqvmFMFT0hWZmyzXLenaTuBWmMm/X4ngRHSowCvWHzG
x8k3uG2I3VZuGE74hGhpih1EU9jgIwK9iEZMOHFYGIwjZxdRdB67mnHL2dR3x89EztS99wHDZ+dU
/kWqgIimSxyO8nUs1EyYK2SdcxNNqa1/8NY0Y3nPn8IFC+aP8l7WYJR1V72YYnjPfBskfv9lqDfi
Ms/9rrHhvKeqTwOH6v4EmoU5rowCocarM2zkYhDsnbGAZ1EPv4GjzWkCH2ynORlwQK01ZWE0Mjc3
uMf0KcQLKDncClK2jP3gRqvIZpuIWYfiEFPDdNlv08Hy09YCKNWP9krqXOR7Os/3SqRj3i839Xal
HC8G6awSk6ep7QosNO0Gfgvo8WEaiEopGU/Hj8Hw9IvYap7gr9plM+daKXg57EhhVaegAIU3taQn
lYEbO2vUppQUB99WU1rA+b2A/v5yuLCPCgAy1Zz84dTZt3P+pn+j0I2FczntLJyGOpUvy96BJeza
07yrhZolBPgQVsm9dCEL7maPjPUdun7G0meEHzA2lj2IbzAtqS75s9QgB3ziXZfv5/PBH26H6Hqs
/0sOAEqsrbdKdyhuUWaRBiayqh/ZySMxYCVemQMiA7hK+ry8t+X9wB4sopOGn85an8BsTXbE5aPF
2lTiVEL+ov157ZWAiQ3WtW//kV+JPw35ehFQbSlVJyfxP8S9HYxp9uAD3kH5sFpX+qZOFG7oc2SJ
PBrvWf/sbRS00Muqc5VV/5lj5rGqTG+rN/g5IyeoOVTUblbMD7znC5Kh84n46EX4LadiDfM4D++c
P+K2UltC6vMc59IitkoR9xK6YYT8C2d9CCt5e5vpKp9xuZJVBtcxXR+pjKQmgMgHvlaG+0XJfkdr
dQbCVob+2o9lm1BcmE6CykgqhD/j1gsAuPTOgjxAUT9K3A/0yRaF6VnC76f/0Atxj54OBSsfrb3+
id2NK0tOq+CwougcehpF3iUeTOBEwTizKPLujyEajqu4ttCCMC/zLXqTMXrMatnbjXSNBx2Go043
/Ylk30+eCqABCYjj+TJ7MZu0+xaKVrEMI6KD4oAm7we7E2JExy3ZygPUZTECqp8tnn3ueDIq8cAJ
JV1fvRIZA0GVEch2qihc4eBIH17RCBK8WgFcO8o8p3H1DKadx/vv9+jX/nTYna+GQDpERHoOA4zg
yN65XsKgXXjVIgXkqiGGiR/gNBYmR4/7xogsPm6ywkTHLH52cVdynz5R/M0KL+dHnTMnOI8pdoGv
wT03qL+2J/qNeeSbflT4knstkNU8XyAi/HP5Sxgs7l35GUw80vxlYhEUyjCj3DG7/fNaycEdyiAF
UHTNhJQzqXX5oohYkNBJU11lIsBPVfWft+wCy+iN9+oLKRHV6ieKSH6croVisJPpgCkjdUt6ZRMZ
hWaSlf4+PcXaJy1pwokSRlujl3Sj0oUg3HT2ien6IpEHGk0NeFZiHgn6oDnnhp3VIkAtiwUhZ1lT
ULnmpfyu/hge7Kr68AxMVyiCriWDzOTt0kDqjfZsFAeQxaCRbKcZHsjor8U1Nx2ISkXfQu6IeHa6
wEi4WVdI8wwIFRtwStZLnAL8QE9LOrDkAw0yj1AcR0AV4jx2hbOxLvtiTJMxzcJ6mei5BD6O8yJ1
FR1UHF1ehjH304irITNQmjuFJn6EcrPJmqeGJydFLV5FK9qJtRHlu9AbfH5lanmXeUeuwA0nVo2G
KaiTnIVeNVnXhS25zbzVpWDcBAgJR1ib5pEValiSzmeSzWtegosB9Kyfuv8oIIijU3Dst6plvgPz
TOjd/mQZ+adhVb8c6jUQhtr3ayO/j582bg2wgIG0ypfuKgGhez7JsmBkxYwdDZlwid1BDpIFZFNj
wiYyouPHok73TjuZaMqSy5FhrZ43fOd0SV5yRe/vVOHhYRCwujXf/JGGtRW4k74SlBQuII8tRdg7
ibI1gaFZNa4siavZQ4iBOuX17eBKtYnpWOHBlwpqEsYQGqWrKhsJIzWl5u7y8y8fMrV3S+0INv9Y
zh90sjFFOv+cCDg1b4jF1z6JyjzS4pLdD1pgoyYTI08l4bTsyIgMX5ngYL0W/aM6O9gVK1WToNDi
OxMsL7lJW6IeVdiSibEqe0pd1QW/k29WlE8TBdnSsavBKFyFA8HXa59Saqtcy3iP+88QYj+pVyPr
Ud1j8uAjSsbjS1p4pAcwgmgDGCvUO7CjyCcG+2HmQ38ju6w9SQdzVNYIctdXouKdImU8rIDvuSzy
I4YGDITWbimtRv72ark+7YUESZ2y/EKlyNha51PUr1EopRXci+PMXWsMyao/QfxbBY/9w7/mpwvY
nGJLbZBY+Q5lZzmazdh/d+bNZz2geYP3cKWQJ2SrS5bStub//hlXbZHgYyQ4Icumx6GCbF2Lnz9z
4oHUtRRM1Yl/cRIQ+0LEebdu5uZn1zx0ByZvV1yLluNNc1rlHRkqxnhYCcdFDMGe5SAU6Nmu/BkN
xs96KDXYl8BCncboz29wxurExx4lTlwGpODbd5TMgRZAvzZ+XQlMmv+8AL1rbuQbqAP2TrqsYtup
pzFYT8NuEdttunkBPQkr/zhhXkIi0RHyDqln66aUB4A+V/7fEAzShhZnMNCKTroHIOM8j+LR16ep
Wm1yFzXrKIFRFVqlQ5+Vx9ly8B/t8KATb0S2tiCxcZUEa6QwqpQv8feE9pcC/GavRcnHKXjj7aW8
xc+W+bKdTEgVvKRcrihDTH26NpvFBx3EsIYITkq9SSX1HdaR70EwDILiDJIvMS8WuXP1r2q57bQD
LEYjfn4oco/DUhUkYvE9V1NLPfmncE/cltGM8RDAFSya1NujAI04Cnl+E9TeYkAzyScKhddtBmKt
Va9fhiV4700gqZV6Les818gYHsgxvlF5OimCVNy8YQWqCOVaU4dx737S2/tW/nGJl53EFL6Oq2CR
u06crRZBArhkfJkU5DKBaoQ1ZGNoPDb5/YLVFqdVHqHJlNkDij3ZxIOHcBZOice1f28Noksz3FTx
Ffdv2M5bYyr56fbxTjPnNr3A8DzV6uPtXJDCROM+DV14jbfzV9JhNvyU+7C3QeCMKXTyXRd4QkL8
9VgrKa++gr3fliLFGCbaZQ/mlfE46lO3vppDOH78fknaurC3LR4bvcq5/oZnt27RzrL1JOIHV4dq
7XDkZJ/myQrfeNroonqH8MFwp1QB31/7I2jcuzU+SNLpK+GTi00KEwf4+QQWGE1B7W4LN92xeehN
iuQlfa7o8LteZEHRzL8dK7rsQopuk9aiRU0WegOoCRfhmdzfY/nZoZQ5abzRq/D1nZOflwYCO4qT
ScRJP3IeetdM4TULCZakAfRX4Xf/+TWE81E7F9rxCsVoIwNdGcPUabZY3+R8vQxLU+cnOoM4btzs
jVhpeFttd/j/BhwLakOM1nNZT37nGQsXfMjfrWa2HEEiTki6OuywIS/Y3FuVr0/7opJcOZK+rPNq
Dny1+T8yE0fl9AhoWcN+rl6dzz0QcnaE4B40Z42eBpq7jNwCvpgAvlJwhVhiO3gXcaErq2xD7ENj
BNY8EFCeWTvf3ESJ+4kPUi/NKpEMT0BXU9a/KB6PDgzs/IpxerJiR1yA1jXnqx98ovqK7H8yHuhz
ti45K8s8A4DvvM++b2DHS2QT8nGDXDkpWaTN8VEAbKZH70n+yEZjHGchjy9P/o9tc/Ensiz92tz1
gYWkURojm43rsAQgMmTJUfK8MwG26UH4+T7VxXhiDfC/pfUi6lC8cNK+92lI2r1Rz1Ge2kGHTDkR
MdZwsv3SANj46nerE4Cj7tH/QY8gV2JhUiMXcMEFwujELH+MPjENzVdgKiy1ONR1tOZyUUUcyRSO
ARa0wak6DAkELEj1fs06+MOpuYTaglIPfxtICSXE5Xp+uZ8ID8ZAkTejtkeoZWgSxoDJX8MbleEi
084hiGXERbiVrZ7NXvKqKv1lrGbvnyZEpUVEdC9H0ZDPiA9gCLGX1xc5nbeFeTSqXNP/Pip6nnh1
7xPN7Mv2bCjSfKZU+R6FAeaeyolNdsE6pqkpPv/CN23wnYHUjaCjhegP0m8K96K/X+Y84tpvEa2s
0paMZlTLkaRms0aeYTncdS5m8QP9ECeb6uxFBkgtsMGTVANxIAgXv3GSLqPzTS2FyniEx4DN7Tso
bunfik3REJrFQdBGqS7yWCC5Wc8=
%%% protect end_protected
