library IEEE,DWARE;
use IEEE.std_logic_1164.all;
use DWARE.DW_Foundation_comp.all;

entity DW_gray_sync_inst is
      generic (
	    inst_width : INTEGER := 8;
	    inst_offset : INTEGER := 0;
	    inst_reg_count_d : INTEGER := 1;
	    inst_f_sync_type : INTEGER := 2;
	    inst_tst_mode : INTEGER := 0;
	    inst_verif_en : INTEGER := 2;
            inst_pipe_delay : NATURAL:= 0;
            inst_reg_count_s : NATURAL := 1;
            inst_reg_offset_count_s : NATURAL := 1 
	    );
      port (
	    inst_clk_s : in std_logic;
	    inst_rst_s_n : in std_logic;
	    inst_init_s_n : in std_logic;
	    inst_en_s : in std_logic;
	    count_s_inst : out std_logic_vector(inst_width-1 downto 0);
	    offset_count_s_inst : out std_logic_vector(inst_width-1 downto 0);

	    inst_clk_d : in std_logic;
	    inst_rst_d_n : in std_logic;
	    inst_init_d_n : in std_logic;
	    count_d_inst : out std_logic_vector(inst_width-1 downto 0);

	    inst_test : in std_logic
	    );
    end DW_gray_sync_inst;


architecture inst of DW_gray_sync_inst is
begin

    -- Instance of DW_gray_sync
    U1 : DW_gray_sync
	generic map ( width => inst_width, offset => inst_offset, 
            reg_count_d => inst_reg_count_d, f_sync_type => inst_f_sync_type, 
            tst_mode => inst_tst_mode, verif_en => inst_verif_en,
            pipe_delay => inst_pipe_delay, reg_count_s => inst_reg_count_s,
            reg_offset_count_s => inst_reg_offset_count_s )
	port map ( clk_s => inst_clk_s, rst_s_n => inst_rst_s_n, 
     init_s_n => inst_init_s_n, en_s => inst_en_s, 
     count_s => count_s_inst, offset_count_s => offset_count_s_inst, 
     clk_d => inst_clk_d, rst_d_n => inst_rst_d_n, init_d_n => inst_init_d_n, 
     count_d => count_d_inst, test => inst_test );


end inst;

-- Configuration for use with a VHDL simulator
-- pragma translate_off
library DW03;
configuration DW_gray_sync_inst_cfg_inst of DW_gray_sync_inst is
  for inst
    -- NOTE: If desiring to model missampling, uncomment the following
    -- line.  Doing so, however, will cause inconsequential errors
    -- when analyzing or reading this configuration before synthesis.
    -- for U1 : DW_gray_sync use configuration DW03.DW_gray_sync_cfg_sim_ms;  end for;
  end for; -- inst
end DW_gray_sync_inst_cfg_inst;
-- pragma translate_on
