%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
vWxe9Gu/7RiQSdpJIk/CeAplTvTE4G5FwkmwtTyoM+JEWUiRUYSdWQ8pI/GyZ1WujVFZhU8aPI93
l1LcOitcnwZmdp+SKclTrlavJ9T0O5wGTytUjAxUSPDMLWozNeiwC5VXHvKy/b6lOEO+mWBJall6
FWjEOgjECY8gi/3dDEQ1iypIlkhp0duwgTohk9NMFoCfquFv4FHG5q7/xycomDGmLDRXkxO2WCn5
5qgiFMK/gfipXgg8eVVQLWVPJLmi4W7Mhv2hPAS+2HJ+rQIsfR5WuIjELPLZXWgHYe58fHLsFwmH
zU9nCyST6XPVrK7QlpALmqzTWPYhcmLkTgTG7w==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
j9UOtOHj/MA9IxyyZvk/TZH4TA/Xo6T8sceuJczxIYU6MfRXEz9WHtA5GOHDI4RM/nx6JDUl2gBL
Kx2a6oTKInjAKtWlW26CkYnRpvtY5EXJePVK7YFId8iYCEVkVthQlr9Rm0VMqjyB9lrKySL2Xujz
1+lpgv7CdKAJ6xxBHH6fZSoYiqb3DzInEyUeOMNvAw2yzQk6uyHYSMkSkEmSTV00vJKTD0WNUkCq
P89Uawss5raIPTBC37VPz9RmeIcyJf3FcmS/KVtw1VEukZrZnG5hvQkk4smqvUlx8P/rP+FYEm9g
mNL1GPlu+aIpvTkm00JfBlTcgCK306UmH4ZCmd9NhYWKZhALvCXnxI3u7W1LuCnlnHwRLCArAp2T
zrqX3NS0OXKOzgCHGmaFKORoXxpkVG9y53IhK+wow33TOinSrwPl2Od/UIPZxXFgUWFX6zLEk0HE
7z+jpIumeK2DBNWMDbwfQk6q+ixC4/2oGzPbud1nQKV87o/i5bERwUCCK8TI1F0F8qIAuC/pX5EH
5TYkMYOzAcXLLOt53cHTQjbu7YGzv5WGw++YblyaDZZpHHs7W1j6gMIGMPw6WlX4Z1E9jUHo2evz
FuaZ/h2JmIcvw86HR3NRZ4Q45AiCJrHdDm9b9sGCvs92Xnjkn8TkCR0HwfjEm56sX343VzJBfSsQ
w6SYq6ZxlwXPaR90/U106gefcEAj9/PR0zXc/6rMlL12j3c+hSrfOmj9CQ2/X/PrWz78YBiXysta
vJARd43XxBLT6vU0kQ9o5xl/HqjjAUnYDPLoXaNJvU9Sh8CGsGEvy0yZsjF+qqqlyad3J0/ag+1y
YxyyUPYdceAIJRYOa1yxnTkmk4+Lo7efl5m0dibnKhiBoOZZLQf3rPMmRsGb9MuxiEOepWhn5L9A
vCxqAZlM0Zn3228V+H4RWRNgYWdWEnZ8C+rmc6hVO1W3ZAoIbTCjslXpXYXmuptuhSphy9aNdkw4
a5fVHUaK0zobeTH0I1DpthKkHS+wajhFymzp8kmYdAkoetJlyzl2qK+RZE95S5qBsuZ43TaMINkB
ffuYfVoMqKkVqni8Uhj3V0511y9xPVOVbBpDgvU2TEvUyBCV7VpGvyDc/sN4OPzmWiDhAsVvyRHP
d7a86ULjVekMyKM6ZykxvFSC6RTImHpUSL2p4veIftWarlY+lIIEBJePLc8oYuQ2U3rtzaQsrEM+
TVCbjexxlvbG6t4sqcY7AJ7onyOStLKtsY3VWN5RBXjStn6Tevdd847ICRnjlHxVJtBmhRqYe6RP
Jk2GXo/uO3jobtI9Mz9VOLhpVTQqCAUdiM2XCW4e8jPaQt2y4ZdTorws4EmDV88TcAyP5dzaKdzj
GEFS55Z84RtdHMuAY55Ft250Imo3tJ5D5oPyTXpctj6bTArzfUuZFa4+UkO3l5dSNvabDqdUJcVX
XOEWkNbwUD3U92P3ht0N89HCriRhbjJ6+CDBSF06KjZ9iHt+LnkHqlCXMl4MeQOXfZbch3aIZedB
8GB8b1yAb9CQdIQv+n+r4oyLNEloEyHWBFsr0H+Zxh2pTV1L7jCFDJiy4Ph58TkjpU7Qa2i0AYIV
iVIPPe984XU2HVKt58ygrJZN0E+swqxx1x6fb1uUudmWpFdWn3E4Q3ROzjBvG6A8pc9+aPUkMpMg
h9FfrCkLRLAxzlQ9lu1/Lk+UKRp/Eu1oLj9DbnE8oeXJrxSW+cHw8k1HVwiP1Ovfw/aPR4kDDgLD
mNyJBfsxFny8nXkhlbfWEM8l8DJCVeqN3OwxKo3WWSMvXZoKWN5yiUMhE57vcbdbOazbfTaGMdON
8ALToDBq+g0wcHBMYHiXDt4vEqlpJkvgKcug87LzD1ExUR6QNVnhxFIh2ZFp0MrR1IH5yJXYg/PV
ZcbFcpr8BofK2ALln5oFZABfO5QK/9AvJ+I604A6h8pZVTnSO+8EN78tdsqIjSQhkF7PpW/CsZNc
4dQwkCg4mPdHUj8K++x3ke1ktc7TLd7yiVMufk7YGeDzwBJxcZRa5c3FbqvuBszZOWJCo15J8TE6
Azk1HNlGN4saLu8b5BoGe2RBA8czwhFOV0aW/SEj9MtckpSFMdClNeBpdZNKk2Ji23mL46esOaR2
3Le5l0Wig4mTfvy5BX5MA/iUoZfTSB0ykjYRgBKnXFngYHadBeP95QVeI6XHx6wffmSF9oiJih4F
SevLxu3EWQLGgHFNUZ6TKU9Xsy5OfTFL22zLQcthzRuK0bIi3pF593aG1Vn8ZTB65vmy70MXZDbg
Rd63pgtMWpc/CS6iJRo4J5g3ssOKLi56gy/A9tC0ouiTnp9OqnZyC3I4y73TN27BstK4svPBNzbX
XzQcutyqXYD5aT6GdPiU1AFRE2Jn13LZf8Llrl488S6Go8QpGObTdiiMiolOBvbodqTyJS5vxcpZ
R5IcnMZeQIErfZOE/E+DmYz3xe8y7n6AUqyP1tg4bslkgmhQtgZ0cP/70yI9KXs66k7GOOKGXG/g
TpTubYat4ag0awYVE/yBXFx5pHxPQHIN4ueJu+ldq4BfP9k5rsyjsn6xfjChDJg/E4cq+xkCKGbM
4AmZsz2ibvmbfix5/3jzWSMVx+32DVVHK9XVCP/Rd++FLNvbFoEuHnuxGgxmoyDvRYIHaQ3FyxYx
tbBKIqJmyxb3lABHb3Ic2qAKm6iy/6SBnSXcqKLs2/9Mx4mCAC9RIjiRzz6USNhawwdlXvgXEA6L
m1J8nck8pLDb0XmgMOZpOcHBY0xlJ2JX+WtpyF0CwTahXa7/9cHYwV3Jk10ovEgL65GgzUnACGgw
d1iFyXEyPBONcdIDydw0Yvrv0K0RyZidDhuV2h6JE2T7oh1wS1J2soniNNvOvDVoo88MmpRsEY+h
xXVxCVSJWcEnEpsFM1Njzxjie4NNLD7EB/azWfzXhnpuUkKaGc+L3cK8s1AwIQG+jfTzjdHL7MxC
3uu8Kal2RvfyiKx9n2oVru/PLtrJiYld3yEiPygrcsl8mi8FJmdSW/sctxpOsO5Zo/hCgJtOeeXw
2UXd7PRhdQ0EAnJ20cm7o620t0eZTUp56TdUB/UO8wCL9338UE6EV1JC1OgJUlq6wCHMhpYzvmeO
X+WEqD7gLLBLHlDO1aeeRbNUOJ+2ow6Tl7flK33nxKGq7qD17D1xcH7CKxw9S6pQJ0tC1jqIA/B3
WuOx05spt9soraSgkPvGj+LqhThmCZVrJFC3jjZ3rfP9TAJZc/JodnMJ7rGtUgNdfXF2pzzjbM8i
/WsnvvwVItWRIbmWSEdgIEMwBC19/ba/xixRlPCz+pnvri+gsCkbkogw8ck/Iq6CK+DBChx/1Eb1
p5p5GqYoGy//h1aFE372l9Q6N+pW4RF4kHwJkqzmyAXiNjx+yaHT6FiePR8zITLuwwNSMAOwFW8g
7XW0tKakdFSmASDuSJxO8RxLKUoHQwM29niSvbWLPVjUxwzeGq1o3msEyHHeh9M8UxCq+yi6FsYb
KkQP6FuHr9bXoDD+ffUT/9nWHcRf6vlG0ZY6krbQEDwm6Ay6Pmqm3IiW7exun6nGhwU/VafxpFs4
ThjpW4827sDuAvs0SHKZd3sKEKyfYbM8agf6UqxHQepzZZ8UCzIC5yJ1nSYB6jPflH/rgBHIapLk
hVQSPhq2/kBQ0t1a+e7sWa/3WD3/jHYrab9E7bwjg+M8EDiaKTm+3GD2u3+RbXEKqKGXatURewps
N6ZxmNpkrEiExccoxni89JuOlj3XzWD1h2enHtgq1duxKF7jnsztT3ZYUAcYxYnZxxgCTFTAX84f
1kQs54NkbmJv8l8n9WlOhxg6O/SPlIZP+HQeHCsh+rqZ5kNFdglDiVlqPUuisTGneMmbdPHjrFgT
ttC60crx376uECB3GoorsqbhN5vIUeGnExtwNYmHv4SrQwkTHQbWLRyUK3FLbLdwpKj1o4d7Y1J/
1KR8GVFUxOq1K58OJYmTkqRVYXm/upCglNVini9ifz9dBTlNorFLKVfkDROrz/cXNJ/KMR3Cf0/i
ZSFswkAFeqXM2eNk4TI7HxsMb6qK73uqm/Pu7L6y1vyGasHQRlDPoJqL/S3fI3DNd/yphcEZ02+n
OLs0oknOyyOqjPft9i1Ka6hslL/eydVM8mgEU8dM782NR90CzfjiK8TjAHYuYpBXL7DBViu+2qvd
F08Vgbk/DAC1dOG+n86NuquHuDMH/mPzw9ef50sWQrwqSoDUBAQo2BoE2o2GbyMPaZCqCZbYA1gP
XhomTtbkbavmg7C5NmMnCZucDyIPBsHGTPuAYowoePifqIsu7nWfakxLCVBLH8htdmPMt7qng0Ee
38x9sxRlLfQEBhJ8uKM78wPUYCpJ/G1poxsV4u1HxNyUAvCQJmD4NgwnAk+YMpNYacAXzLIIzA1g
24CwpztosTCq7zXABeRM6HsS6jhMcROKczqMVEjUO0YgcZR63oUYV+WTieMM1QeKLSEeR+qdd7+9
HcAlUlMed/T+YM9uw3OEzNakpcyLgU7Be5Ksa1q4DN2LetDCln+ODVLDmw7b3hivCKT42eEBFNq5
pZrLr2+43Fx6mHiopYZ/3eYlqWmn/1xfewYJI4tQGUbwecL6YLPsPR5Z5jOC2h/leSoGppbJyZhx
Wesm3LMMp6SyMQ/y+DYJVk6FYczJP8C8Fhf6nmw2VHgUSb8jRavSSeVGBFMfK18Z9ds1w8ls0T0V
duZrSwxCpKlL+xOkQkRWIzsfxEyUsqShjT+3xgMJddj0EabnDdgneGImtzMSevFvfNn3SZ5OAGxw
EDvbEWdwfOEtJId2yGh2TbQJQmnz+9xPVsJNrtXSL9VFgkYSb2L1nzntAHyRvWKwsXgl/zmnMJ6l
l4WUoz9iPMxSBKUgOIEft83yQUPCDrDUzKfLv646OEb9juSc+yCcb1Yaw3eBoNnvlcQVqirj6J6I
OD2/8VWnEIi7i7QGQyRJKr5QK21FA4ys9Iivw3lw35CRf0dhcyrO6QdzbtS0eppMk+NY6/ZvyHdS
8QkSsun3WMbjFJvU9rZkqIsOnZFA04BOWQjsVrlMqhtitmToSECa2Gg1hojUSoqRoo/Gh/lw/8zw
8F2WG4ntZoLLLDzYo6w7NTNUWrSU2v1aiZMOZT/fErang6udkpUy59LaiakZwQAG5y/52SfE42Of
cGl6R/ol2afZjJgk3Jn1Uqbhf1itMRN1nArUtKKACQ9JBtHFat12thoZg9QWOY3CyItKoMWMfNjs
0p7l0C/65KjiSRS6je3VylcktzxWYSJUhEwBKk6UqFSTcbePwKL0JHCbt4xzDIdqRHdw5DXw8+6B
OfIX8R0VakXoT6qKzjHZpSWF3EzYZ3YeCbQVhra7G616qJPZ8SaxmjxYuoVEfU9RD7e8yHMvZbCz
DVTCxe3KEv1qCA+lTwsk58U7+GfG4nGIFRMQlYclW2ityOshj+NKJs1yKhB+j/0YyOyJO7ZIFikT
uqKHaQZrEo6+NpCfCPSoWuDJcvqDqeaqvUNTucwx5cAr4tSXMa5Qtl2nclswdD9AtGoJZX1zEGn/
3wGeosRm/J3Aho7dQmMAc02U7fErGijQKXuPHE6Y1zUlkwz2dbSMMdmauq0++6jlheB1poBVR6Kk
lIr4yUkh48TwWm6tsWFbclC1FYjPdyxiLp7LYK1TnIu4dRMLnG+TNX0/eh6rsP07w4X8MSDU9SPd
hKE5aNT6TLUMASdeB1p5YLJrSyPxqYpaqGpO4ixl5GLd/fWSLknGojXisiduaoqfoN+kDbLtS93e
9y5BSUU5cPZifcUNFSry4doAQ2XUw9ms9p++ZP3ovY0PL5EqDRqOtPbm/s44uEtFsYZ1hbpMRsV/
3HHyEtL7yB3tSp69OGORS6/UqLtiGtwQ3RiCeluTKJ0QXMMnOCLHsSepqt4mg/Q5yBMQ2aM5cnEx
xFyNA6h62S6tA3Ml9yiBLcVDjrm8IGQJRIfFn675zFYw8/dCtpXVQXIBSgkLe1OAaaOoo7lytsOC
O+rFkv/JKbZWi6aLjLmPjDTB4sEbzLH06FvGvh+De+k+uwpKnYOIAYR/Raa1z7vANqRz2PS6FypI
nQjLaW6z3k1Bg+cuMfGADf0Eiv0XCQA+756nkDulvPhHa8C2awh4iCwdqR+6kHTgHsXmho+WFqyi
HHPC+L8ziyGHfByvUsUo3jWXg3u16LBtlNiOMPto7A8W564cae7EsvPfxkYUFrzjzh6VQvCAkQEG
XoNu8zKtDM8X+fPIr7s/WTZQ2cS6VCjU1kbee5wTKaKoUztWr0OL0p9Bc8wIA634VL9uAKHmi4Sl
NdnugSn+EztvPkXwh7614NAcDek8HvDQAflXy++ir7dEKCI8jYgOQtgGazsgGiDu8HY8KTHMoXXW
wh0glsbEecoxwSCtICVGqG9cCdhVFiD6w73SbXKsU8MeGetL8gPFk6Ut6fukVeVF/0dHJtqm24mt
wEA0aLehQQquY5le2vzdhi8SBG3a9sEOPNHT1UnnQ3m5zKKiy6rk31bkE9io6+HhtHAKQHCPcs1p
93gPScpQRFyAmZbjo+jBmkqTXzEpVN8yrfGGjs81P8f/d8DUNkosI/K5e8BfHj9ZpBygALdLkIBs
qb6zEFbSsJIy6qSlbsqOb7y6MViEw/X3CkTX0WwPXum2XmdgY7KrgWCobTV2VF4H3qce9iaEkdxC
SDTeZBnTTWrOY5tybSZxmTAy6tNvcmfTvecc+O+DLmr4KHNktRAg8v31z6G5cz2S6F9+b5MtnpfQ
aMAOimOqstHUOFzOYd+BOEML3cF6gNT2fqa3A9qbJYz1zyH16nPSvTJv1zFqWU6/qilicjSHFQsL
J1UktyLl5qJhp97a7fzaaGzI5E/1yYpGkdJIeMxXLdrfIZzHGwd5NQIlu+jOvOPrtdqTYNR8McTH
7kGu+BxjB1vuufRlmYKUjp8LfTHunaKeXg3kLurWcoh9AZZ1rBQwnwbGU0DgtNM8aa/igUBAl7yG
nssQcHwBjIveHaIWIFPELBURLSCMcwVAOuWu8BGyMHkAhSt8iDgEuy+JaukSVbL6PFRh+tQxStny
zxqH+5PyxIuEu7xKAEubEFxBu6iZ+b9uWXneiTt2JsKW8kvd+q+6HFCdBqi6Q0W2s2qSxZBuLoEb
FVj714c/oSh0FKFsK7hQ5OI2xJHCGrzucB84l4S3NYpJRFQMEluiiXt5H9WbjIxSKFGJ97hqYBbc
UIrZ5h3NgYvf9f8fpVLykPJ8wSatkcMGfqxAlVRac+5MrMyhgNnmjWdWGGQZ76RLVFS3cKKW/3MS
ttsuo1YJFK0UDJsm9dbmvTVgqXLR4CSbWsVClx5FqiDzVXErJJmqdb9mGIleFCDJpXed98wfMfxo
XeG0R9E35DfdRIz0c0VVzWryCNt+Bllf7iUBq9uwXlxw5Fn8Ydl9xgbomIqjz3kB2NxUrqQgdGH4
pGdyPLFauiXJaj2Bn/61ld0WPqsXzBxalLHRkn3NpM1hkCGOaotCbv7PRMjX05v9RZrvMUXMO5bD
RVXAMJGgiwBc/CG4+4lQ4EEjbM8kF/sH5x+4pj/T3Br+KFwAKHOX4ej8MKMDvnu82+FrrMvH50pQ
Cl0G22JdlxqECY4+fcXlyjpjlq/bDySuNV65IEGCC8GkmeF39xArpAN49b0mbYUxwfl0T5xMqrl4
qOGaC7hqNZG8QUq5RoLgwtpW95ISfG13XMComuh9dpzI3pEl3/TYwCQk1Ayjbo+SCQWZ1j0V6iK3
gxj10DcKOUiof39xKGPuYBQulb0gTwaufyqPXRCIiDbw/pqUDDO/8k60KJ1yx4qGmQk68JGod4su
v/lRf4XiUgLIfavEixWKmJ7A8Gv4NR6mVaqMRWVTKIcnlCgaHIsG+Fsz9Pao+7MAVDzEuVLIbv4c
uEqG24ZPnoZPZWpQWSTzsYs1UXz2tAhD0QWOpZHWnaMClnzWMoeFtKAqO9nOvPHr99YKBhgaGgb1
PaG6xHD68edE4ceUOHQOdpwxT5Nn1TKwzxEzhueMWwz8yma0xyt1LtNq37vumzBwKAadw8fEa/4j
0098neGGGIfTBoMyoBypMyAn60ZDGVsmdDe6lD6l+CWZD7ZS+utzPt4qAmfpqWnvAr6ewbX0AZN4
y/AVHcioIrLSTl3X4F5OFjyxFnt+eRqocBQUSjMfUhk1UDEgCKa3ryyxQ2hkdBQL9yu8KaGjTyoO
sLJR63ARzdhlvyVSR8PXBi2KiVWpWwWbnuGk32hAMgKW4Ep+K6Kkx4yQ4SxbEbH/k/An4etITH+V
cAZ/8W/XznirPRCQaQE9O/BTtdp1bDR6DnGAyraD6VQSQLd4lqJRW8G3dQVawyjZTfEME+EXYgl6
tyy7N+UEWMoq1LZgs1ThRH2hMjisnBfSFZbjv2Tu1z1IWJZdVVRxS4rlkTiZJW0LodR3RYwH1K21
s5uKt2ivYlbZCCzmIXkcDZM9UcblP0gr1TJK6nazwnJHX0iacKp4ryhP3Hn4GckZYA1+nYgUT/Ch
eglHXuZcGnTy2r1mITk/py/ddHlJXDNXd5FSXaLeHLh49SJrsWzcu/r8F3aRfUZ8rkJ+1qtsKr+z
DkwTww8mPeJW19zG3ET28LDgyfv/r9MVxk5TEj3YGcrNaGu1pIsW5TFwHC+b3wYWIA66wel6LEtM
6eiHZfKvaxallYhMEbM6RwOaDhLMYXTor1TBdr47741NbD37ppG0GqSScEqMjNrImT/mnDNvfR2w
ex11e9ItNhqpyTo1YkPTOS7QBrpHEn9qQHf5f1pbYdMCtV3DgOmtp1lnKv8zO+sQFP2nDxdWGvGG
hxl4IJpo3P9eole65j78PCHXBIrrHq4OkThyvqfYI0oGk+4Uy1QqguZVl5jBCQtkcae1Me/VV2bG
nCnc2Cc+ynDHnOvnHWG50giSlX+0N2w/EWTCQMhlnLXpfEzugGt2BrnOtoMH4Qg5RYZV74YujMof
xDz/G2HC4wsjyEMzx9OTGDK31yG3qb4t6s6zEsw9hNVChdy1qtLIV/xqSjTAdsnZsAO+dBlOEUtv
dQ8+5vPLXDgwlHoGM/gTZKTTvzHtTDeLkxlDub9N18IFhS4I7mqLhaSZ6wC3rXgHy4kva3OMnQpd
pCz/ZKl+ENBGt+j7ir2sePKs+l+/kEHs/K8zwWOYrOPQc+9M4Ttwfr7lNEiKiHohOpan6ITgglEp
nXfvuRzrzfZhHBSnOzrJyTxxaZO3xoviGnEjMujzumfRnoW0ervdurdpslyx4iraOxxGDbSGcvyl
+aMp10iMQvgjY0iccFIZskikTwTHk/IhnR8tgIf6nYdbTZpnLGEBG6TWL06ApJosdj202Omz+uDF
r66hxv/aIuajiCP6pqdf21oZS/M2KK87hsDfWGrsdfcJz9hvCKjXVYGjUu4UbU4OKVuH16kn4nby
nXvcGArrcldu5oQVHzRZZg0Zrsr5L8wLqU1bwt0Vyi1joM2wq9YunIAOgOJe1dJWpl6xgHaH+dfr
ncdsLVRhUVzBBXAeOfpTDhGcpz3jDiYyymlHErebilyo37z6ao7OibP9YCl2g+xTWzuBCzd/qEVl
pOoybQ94wskTNFcS4vxvxki20mCUYVVdgpA5m3FJYAren/bp8tTYI0HZSiGypfEGNgLU8l/bkms8
SJGZflFpvs+9Ufz7S54iVFcVQ5y72v0ucsF7NILbWH8H0YnBWJrWpJeot6f5tOB1u6V/rueqwTAY
ZSmTDc9Awt3KU3ExZJS51YCyh5EqiWzqUqVyY4o5VS/GdCVUCopXEzvJMHVN31o4TWzN2z2P3+tC
XHGmPEeRCtJTD/aC/qhlqjeNGkVwsRxo3pOBsuQS9mmB4NJNWI2x2imE+/UPgYCe4ldVmNCDceb5
AxAd8iQeY+pl7QwJtajF1eff8AcRxnYJSc17JcgDaM6kztJCvLFclHt4RuE4B8jfiNnFb3N8/b+v
9O+n8b80aGvbG/npImpmU+Hrz7TK2QqhB+UZXooOOi/tEL+ms5Z4IhYEIejvhZAxZBqLXKiOXB37
iUqupEaA6W6Fb193f7dT3Wh3n4MHeMmR2VpfBmL+/BTvMdeqmW7UHz1mdI9FgAT/Tfkm85mvPl2v
DhQQ1c5iwqWj53hCAOgo3min+3zN0+nbbCMIhJqgvbgjyW4INX7dZ5BhZIy0JjdENRYmgcYfGaFw
jE8WKTJCOwwaqkIc+/d2LWYaz3cAd9juhkjYZrqqo4zbzM0HXNB3lRKCcvnoxaCr8Mt6m08NM3NA
9cRKLTILiKDcY2qtk6q1QCcBw3McvOvLqcd+fA5Qk9Damd+wZoVJ0qQuxLn7ICOPd2jCHiviQlVe
E984yh6gPJno+kSmxSr1SxHpFc38B9Hk0CLar05J34XJ5EWNYa4QrySkVzqeEFaW9z0V72xO9pqw
M36Yhp0PfZ9FAO9Mg+w1513IQxHm47Q6GVGbJ4EQgYouro9G9NNXNHxO//ionYjYjJdxpgEK3Sb3
0s0K1V3z4FtlAHJGBM7ObTTtuZZ5LsAYI+ZhikMF/bQoF9WispN/DY6DzRMRfg2nu0jj+kOlyzWb
hxxR4fSHkGItXfLeuurol5/dFitSRsQ1lcmo0DxtyyAXXOxR0/v3mLamPPdOpR7kFHVkvyK1a6OO
meqGcnp4/Jh/ZgRMbnC7mmUJF0BnY29H3qS8w8ktKj7mhSXhQ3lnorc965UnZVa5O+ZIWM1WPhpw
ZaoWtTqevVcaoC+AaZHWmv+6sOMW5yrYBF8BN72v4bMZLLc5d7O/W1ORLFvt6QOVyr7p9fwXSkgK
6IUkgjERJuSkqhJeoKQaFf/74IEoR4MZGNpIu8NlU2iM+k17a7vGyYatEBf4p3OBRPM9u5xkk4YL
FYH2GRulHbCqCrkqHaxAK3Lm/8ZrcBMesg/KBW+0/xAq/G8Gcy22suchQAFdxVOcKlbhOhTe+uCp
JNENqOOZUpvAyaqaClcBguEhvQI292qwPT0v1Amsecc86ydLpmsjpoMzxLrD6XwTLT3tiO7Mf5+R
S1x8k24JbN/qlRnzhmX4QLJ6U24XzzCt8Yhh0dsTQw3SzHIEfzJg41bB4UaZCDJ5uBciBdSmTVq3
Ypn65kGbIc88ttxtUZ98BW7r/bCFH6tbvcKSLPJEpONo29G8z+uZvoQcKogXEIWQJMGHgZURNmAB
exKMeA834f7i1uC/2MTd3AQiWadTTmR1qRj+bVBoa8togt44BRUM6ElR0mksyxulCt5284YPNhIy
TBkcDmh6DfL14CTdagwVHhMdJcXraXJDgVB0QkEV0/Dy2NlOEf0fWG9jVlqn8GsnmR5mshBj26L2
UWs3/2m03dwWTtf5U9Mr8oo78FjQxMzH7R2HBrUtqTqmo3oXPKdx7qw/BFSZfIBOeMHdHCFzk5Bl
zqyocUXcaDwXiiG2rVz/6p3gTZZmktpBbxkAsI07GRfnP3lJ/mdjta2bQSwB3J6eFEwEtQG25M47
NY4XoCdzRXjS7lLNQQVL5Ti37ZFY/FvA3z0+MMzk4UrHCxB3+8KNxVkWGEBIP+5buNj+ZAAV/w0J
1tYuhSfUWzqXn6H3Rl0DxzaxzyIn+Hjko8ddj0q1GckaM0mLj0J3ir+wc8iIlT0Ixb/JJBW7023D
BUaggL65fgaoUlYrIKpGGIOhk3h5ofDF5hi9sIqJO7bS1qvj/jAVOh2rcwM+K9tMHTrGvTpg5ZOl
L1T5Lq0+MPnezO0EyguOpV7COwiHdyyE3KaOHRaEdH5ut97YKxRdMGsf6zflD0DRTPlat5emJ3UG
3pUCHfu9FYMumUq8N4EMh/oemRaAidmLAvL4kIOjHK9HrJfGQbWGC+Qy/lTf98PcL4owp9VOUBs6
bbhCwhK/FFWvlilA++OlY7d0gQZZI/8dJj1D365l3Ug01tcVDZa9r7Jg1ZAlk1Y5BusptIa0Q9BW
iXV6QLPMHehl8+y1+H/TsWV6OAglXKJKYiTky1cjyNEXd2Qrt1wecya4gG9Wm7J4lQUW29aU1sAd
PWqhwqHmHht1rI0MVddgwcopd/wS9TCmJ8jxdwvw03e/CCtY96c/cE8p3L/GP9oDX/ylwVC3vDOY
DAo0vu+QvgBLhVGXOs83Z3DNqMcBNmTRU2HVWxyhxkPh7Y/aw99DcO9+6V7HpWKBOrYaiGjZZmEn
KmfUbV/cJ8eFpMffCCKDTx6y2vZFOg1/MCqL89iP1jmHVV2XwonvpZjjpQc4xYs7tPIrXKOWIhGy
btvgMoCMkwCW+OIfkID9VbsKazdvIXgtpQhyj0kzi1LVuJRYi5ShjHt6hbIdzSi3cK2Ky6fkuFn7
Q8WQBTmw7tVkBtzFe9D8zvmoImu2AzbtvnqSgE2/Em1JwYkgj5cReDo6JidpiJ1UtRn3U/rc/4gX
Zc8aHFUEMB4MmHFroPozz8Md2GV33ycCrRfwahHEUovy07Z0RrsdHUAFmb3aJNHGyjEc73pRH5KV
l/hg8T+V0QQocH42rMYJf+emtAA4QZ2O4QT8BGrdAxi5GMMw5jZMy0E0xwOa5WgNjvjqXJFfsdAv
mvzaVVsuzeBu2zirhl7lsQ6N0AZh3pwJ3+T50VK9ufePKujkGg54KKhWBUUPYoW1/Ft8bsLBFVsU
ou0i19retClMODsbLJ4vaejvRqMmwB+r91OB+E7VYYo14JmjY/n4Tj7OJO/FlNs7cQiZ2oOuYc9k
PMfqn31bJKGnn/oIrAfMekKb3e/bp7wA8yF1NwVouKW/iemtlmANghgiMQJXsssk+z9ha3N37fVU
nAdfFwQUBxprtCTC/h4b3fEcF6miTIxqenRqpnI31RvSEJU+av3ZhWGGuZ7C8LbIHIJ3YBSTjq7Z
Lw8Vh0LHmbJqGmWr1UVu5jtn0nkYJy+QJ17y5MBdTz3T9k2TBGShUY4McVKYgQCfMfbwZytsr9sx
SKHpiZQNPbY0PmVJYOY27EHuMAX/1kvmgbaBIF8gPY6tQzV19CKlnDKLFc0wOeX7YtXOPfhV3QRP
3i5wA01uYBQ2oPJ+CxY/qdG6Kqj2HCNCHz48LlU525x+8WzQxZhfcEgYuW527Fh/AvuPKcTQUCwV
Mc2LHJkuQUT/lhovTovOU96RdPo3RhCwQTa4PWre7aH1qm7b2L7jLMbA3KFpI/PAQFFszNgnGB5x
J97U3fpNtYsNWzYtigU6++E/MxZXVJs06+RfZ9Gfqh82dhkseoWhFxzoCpug3zQDRqWajVaZYitM
hAaIiB0oA03aVeiDezHkv0NvLxYEI+Mrw9xtdsxY3MwV5ap9YLCZao4gRBYjmq+W7dpWPHhos8hp
VHLyTQygyZ+mwJPeWwYiiDMOukvkL/2LvDFCcnJreWbX6CdJd39LFj/fYdbCssiNgVj3ScVz5vo+
w9IZKg1ifFdDnqJfMV8jWa6R5PKIPlWWajcyU3+kdimK59Qf7k0h1ilUpyaGJ8HZBdwyhUjcWiMJ
1Auv2vnkqRpUsSpbt7h9tW1ZqQYlAZ9s5/+hYxPLPHrmdXFmE5LUQ5cam+2erQoFLt1WhSfzPrB5
0QyOJlJHDUhzfUSX9ht2jRqOJ10pxN5TkhptV6DPp/D5Kr5D3riIB++tp67NgyzcFsgQR2209/Z4
WBZQQCkHJU+xpsLGRON7yG8G099RN2EMxp5EaeMCmjejDQPpyzb2Q8oGpu61dhmBDlQzmtq7ImC7
FC2Z5SAuGRT44e5sl2YQPqJJi8pR1cC6uHhalEI0Z1jZZQqHdVTWb6eIFqkj9j11lZNLOqoai2PZ
eLm1VXlXNdpoTWLfT2M4Ihx3hm0wnWlDYDlSXjAa5AO+mUcfO0TaIrvR63hfXDRfG5e1Mn2cWO9A
HBbxvAZewg+VYagbduwK6BleYWLNpz0c7YyKU8n8MfECBvIKP42Tjmp+yA97/bUP+B+XVRzHhcQY
zp4UdhZ5hW+lcLg4SrMSxB8tkyo9fzW0LpdReSZIRbRp/tpdQhAB2v/2MKAJUbRApCjaoagye8vS
uo4dyHKzaX06zdpAUOV7F/6lvuSSLe7asBXHT5iIvx+ukdP4Ual5wwcKyEUDsPbb17Lhrg5kFfoB
8V+wliEpvD5isj7njqgSjXSTcyWUGPREzv/n42WPl6ssHUgARs6uOUblOPaWNHlP0TL024oTqE4V
w5Q2Wy5Gp+shzp7oCvqDDDOuOZAMJ19fha6v3mTYEIr3u2hmK2dKxYyYKiTvf5h4D7rBgqhARkv+
6mmdC5CuH9p51wj7u7dMaH97OJuTQ5TaGcTJ2ez1f20xSkPiMci8cT7/VYS3B+TpFTkIU0txRkDn
71FU4++eQ9/FjUEEGEx7hRlNu4jiaXV5GjWzt5/492MaTp6IFguwd+V58zi/6tUGJFChtyUVrnQB
jVzuN7sw0MOCKZICA++YAVZCSmAJFRhXfC5BM4uRSYjI0y0DE0tF0/VRvOep2hBk/81dqLVEc3LP
2GbvuGUfDOUHfRh229mp2pV+OtdYg9b1waGkvoY0TpQDVcXvp4trX2X55LM0cz9qPZGIcpat5eE0
B0rRq9b0K4f3XmNSz3Mi36CL5thsXmVli+iA27qPL8KZABRnsrX7WzR2u6fLtEmm6X3ngb6v07Pg
BtITmfuMqrQf3tC8wtU4EZkdQsPy8gyhSDJ6FOcVa39T/yQUUivohbOVqY2KI7NhSlcO+gttG9ly
V88oxSqbJnZGYeCM4zs0jDO/D/kbEEHqImYnq7iQiblC2t3aC55E1HZZae5D+0FhWHEvfHW+ot9h
EOi+KAgPbzzXSocPUn4msi6jC8U9Plc3BJOkIEuXr1Umy+8/HY4qTtZvdFEXSw1/TV9sYy5ZTjOV
VzIlmBMMavhf+haH3zCusm9diZ9Yg4NXKA5usGODkUbIkhGtysnGJARrpTnFBMah+C2GsW3EWD3T
/TULanDUIe2SM14Mh4koOgJL1cllnrj9bBh/CwPidejn96pJMnsML/X2e9RZdEgG+yVjdEUnb9iL
VV393iwGwhItF+Vi9zOeNOG90QG2/c2+asvLp0VKrJTXmwNeCexH/B8KyDNEzueqJBrR+dUeuTja
FezXaBIQMvtucynUZ+4VagAcXKmwarXa69pa4mptTyNrug/bMZwMEVldz8tDHxcIRKHyWLDSr+ND
ua1fCqeTLM+MkvKO/JGL3LAYqkGxWsljzz3f9G2AuWpy++di+nCSu8TX/N21v6pyd5UeJk6jdG7G
592EsRsb+AfIZHo/pJFlIaOzF9cMqmSZDr2WTmGS87Wkgu58HV16Nxh85AljnC9Z4xjWZ9wvXhUr
eKGt4hCWRJdSARC/BhetgiIt8IJ6VO/MalLVMhS97QeNvYjRTOkc0nxKekWjNz7vRr8M5/ay8YzV
XDMMQI68BU59EgSkHE9liaN0RAMwPt4cCTJOaLJy6T5xA0ecNh+o5Q6HLM4SYnFA78nO2ouDQq8A
QRCJLhIiWFhxig3+rUAS6wVDXWyO26zVTl5bN5QFJbLIp9HN5sAGovpwtCxAo6UoTl34XcSj3FYA
dP9lEbexrsQlxx06EteyxssefgTHh8cZ5RJwGhqpjKbaP5UX7vR/Ckfje0xT6+zZbM06+Mvzjbv9
cGdPtO2shptou9EAa81BE+YzXn7yjvaExBOIcfthGS8OdsR508+ojIkwISt+h+VdB/wpHuOVPfnG
JAprK2Su6ckvQiZEBiunvzo1s00tNL9hyE4wGeMUZHUoKMjO1kNe2WALjMW/VGoY7QesuzpXSe2g
zDgYZnlNzfCnkgEl+vmzU8uxxkSpMjCc1SZgs6pd/I/S2lUU7jrbRPLUmAYs4IYtqOJKmWQcq9uE
V6dEAFwulK/PFngEpSCMOHRXGldPivdoxSauQEzOP5or4jNC1ErJwBtF0AIYAl18Y8yHE9BWMaPW
aFczZzMi/yIXxksB4cFaowXvpxRqvuTF56NG6752Eo+6sgGX3g4V5SYcrBEXSCCvm/+R1vsue2zK
yeMBHL+pAOfl9PSu/KyH5PeNAc/bdxV16G3S1H1x0BsIbCkdkvvdkYSS7TKaeNuwHP5Y7u0dCyEE
oAJgtVR0El+ajZEVCN0EBIHFPa2lnziAQMwr0o8jWVt6PZq336vBIPq0MJtRq5PQUoX5fOVnW15/
0C7wxfji5gNC5oDhh2D88VkMom6WwCgVapUgPrAkZU7yAvcl+Zyam1m5dgUCYrzoTsyCTPLWWJjR
iy+dtfKz2Th40vmAyVshYoQcL28Hw6KciFORkcY2+gy9C1O4l6+LLlMft0gO4GuNPZAIwzHcFwyX
4IoDNrZyJhFfM4ezb/1sPs07mQr4rtY1JcjX8cst6pwj+CvvXIzLY8Etqik5LRuMjPWVFCGQVPfp
SCAYw1x/c0a46QKBde3d1W6tG0+UjYypQs0Ev3h+aPifuU7lluEi7SO+Va9zrQt2PDtZ1WHQPks+
BoapqavgKqG7081JrNrX4YMQgv5Hyq2cDm37R7R3Aeof/xHhNsuu8JaTovf8cqQt3mZHML3K7Ww/
gmVIYQio3XwFHo4fzQJfh5eVNVshBrcfG0TH/DJJkWoV+uTkWVi4uRkmCARDP6yfb041saegina/
+11GVBjRW/bBJsrL+PkaMaz5raM9EAvKtSCqW4Wj2DrLcPn9tmpWFfMEJBU4QQSDMeZxE83KffMg
m+sAndBQXV307Tth+qeOWovdVMqKwC0Bw19ve7qbQg7bA68eV90gZ3kJf17JWt7cWDtte4UYqW8a
OSAMgqvmC+YZlRp9GmHNf1jZupS9zELrmKYWQNYZMnkOH9R6YCsq297V/o0+oyvUPdBcy8wAGD7h
OqDi9uFi76KX+5CCjqqfuww38Jt/vwT+2+A3fQ1/qwpWywQAXk8/oRVIsxKo8aATs8Ki+khA8mpS
aazpc1S0lIRGlJHYCKeRubh9rBgMTatrLJyRjYbViLpYQy99DLDa/UVLEdZiC9KUVUKMsF79K54G
tv8bBtt+rXSx2Y9wIUuvqWgXx3P65wE6XByFon+jlNktmKJre45f1Qs8c2KHAxGHXPQubxTHLP0n
rFbq344p/ttaZLMdNfv9bNPq84L9k7DiB0mICDHtA4TGJKLNkl182UtTSVybQByJBBVY3uDpcT7y
1ZCkoKOp6N0z1cb2/X0dwaQ9kCzhf++nis6F9PS1FfdY2C+bAS6jHw2au8nksnMwYTJ3aeNgW7wW
BcDN4eD5mKMblkHpb11MGHHQsRn1y2ISDkJDjETQ7Zg33CNme70EvFu7umqkMx3Zi3hU/2NCLtF8
6vTacommWZ1D+TR9cq5wQFhQf+BNSfqqN7S+7VzFhami0RI73lWR59TlotEgqWG6NgFeiJ1xwHDi
6xiY6t1ANJjA8QtlVKOit/1aDBYKsn7/DQ2jPibjw9dWEzK0Xz9R4vV4EHs6tlOwOFl6jGZGUtYc
kn7AVq7zirY7HoDZiw8TjvesdQccxqQF+JiR2Gx3HrXBGRw5x/J0zm5T/S4vRWygAR8P2KHhUFhd
TEFFC51cwMbPeAqaSZwKQUr93XRuTLF3jydllIwjxmBfpDtutRSmETUmbmgjAF/d5jXZbGwrNmL6
TQ+nfyG29mFOq5nlHDXtuFtRAa7cjGDQI4Ul6zjJsp7MWn6jt855vT2p3dL+OzPALoMMG4ZCWo/5
JprqubED/39SFveup0dBGXh3LkjGIk2+5mB/odoRW3RlrqHJS33X+8lRIzwhDsaec5oosbtOJ9wj
KcHuurxhMFWzUcr+gsgMJ/LkV42/k61ihGc4z2gSH21TSKhd2VZF6QZKOmPn5ftKk/yxs0j7JX5H
WJY06fl4LSP5G+xMbmPJuL3QJOmtIXTko0/kvmuXLZ3c3xooFr2wxvawFRR+wje2iBPtqIIZLtBK
7uk2HJu8SofVGCsgu+QDhww1nSnS3lIAd0nT7X6wwqdmyWgKJrIeBjzxk+hw+viXuYacqBPweaIT
Iwy3WLAUQRU40WvbjcbNRUymRCVsTGjkcXWnL1CtwOPMK8jPd3PqaDkW73GMK+lGu9g4Uc8QB/cp
X/2cuUJN05gRHHiLqCtGZPg8Ol7O0ZMg/bHjNH1fkOrR3eAtscqfa8pWqCPle8LXtee64ZSWZY+C
ravnzzaSGXKZOlQ2Vrj2a/19UCmUHg8SNiWposXIWTwMwB98/vwQ1t2xafz+gR2rJeoiTnBmL+WM
KpIQ/xKkHbCsBQ1x7/lgNW8ygmvb8udQfEODrNqsExICIrN1KzkdPGLbzj65MXiD3aTZC8nzPy3O
IG9+xuKqArfyoVWfjapSZhDFPa/7PYm/DtLuezHCJuixS/+11kqoAJkQE8R6zbpKkyA4O8GmJKJb
OIxEpFFHCCncc10hVgKi0jOhinIDqqWzuUgSzrBIKFkJFYyN4G6BWI8KPfNCe/tMptkvOB4efgV5
/jr6uTiqO06k+JHSNsioy1274QMcBA78qro0GWaDLmA0zh7Pw2qGDTtyzGJ0jYtwxpDNGMmEbR3t
iWHIuigqsdACDHf0c+w/aFIdGqsTSpUAFCbd7Fj5/2snZWUTHzUmUcJvE7KI65GdqTRkXZKzlmKT
wvHfyUh/VFXUWhew+K6TsxQuthJgWnZHAYcCeZQlfdcQz7vqNGt/69j4od42gDqNnV1GORzOf1O9
Saa/Nta5+h/xROERzEIm5rMFoXfL2z3CVZu/OgXxTCVBuZCbd9nTenAVLON2b3NeeSxUEhbLaI2R
VlbTSRZarbcDv54OJ8YlQUqEztzeE6l44ir76c4iMGdvAW92/efFagcRCh5vROTSb6WMPuxskbSa
0w0IMNUxGHkr1T36E/Iy+KqizXYHXgiTxwHO5zMUO8lvIvARMQm5EamIEqmVk+jGHoppoInhowxB
xIMxQqWi8zt6eZVgnARbylm7Xg9LTj82SVknBx8Zz7jjflhfXeKzez8X9nTUZ3ZwO5ufIXQb8DhE
BAhW7Kq2hg18WWmgxGAk6pIyxbwN7yH7Ruy8mh3b0vOCMuGWrnI+Xuz+8XrgIWnHi79YzZmTGOGB
2km8r3nVDfv42SI7Hk7fHO088fmwxJYGnpRhFUZc7ZcQ39KXxErIS3RJ3O5JE9BuaMD4Dp/Dm1ge
3TyW+dfqZbNvexFIdhJnaJMM1mJVqAeZRv8lZW2PP3cgSY1N0K3DWmRSF2ykKq18JQ5FFfVZ/l8M
PgvdAGvMrK5irgkf2ju0Kx9pfAwf4ckDI5DBJyvkmBgEcrWqa7eWTn2K9N2vAi8HgzftPn+Ut1h0
GhJfELtskov4wANaKURCzi9JiyFsszuERVKAIqZ71HaSfpk7J0KmxVp4aA6EuqgcHIZZHVjJ2GLk
7Cf0yoGskheHqH18K6RB92CyXue36AzWmLxNw7sbcZ+fF+wmKtOR8AIKMofT3c8PYHvCdrAubRqv
9SL0iev0+O9oLioWUa/Xa6aEvu4Z/ln+Vga4Hp3lL7Qm3ZgSgdo59PI+3OMVId+A+vXgMazvWiZN
IE1t4STm7hJ3kwdO1ObotrG8h+wK3oE8nvdsVxqVetW9rN2cwv+YBYqLh8sZSW7BxM2F2wHQc5Uv
XqMu4ZISDB0a6tt42/8I33wGwvOHboJPxGgxWLzdx41L2RIDei6S0da8zljNmFl3UuwExBP6dPNJ
i7lCtLiOQtEE4iN7Q8SAo2K3RbAAPNLkyP8j3wQTmIBocbscltHNGCRQ1RYXzumgSoBDlyOGpGBb
GReBDUwucd2K1gzz5IlphUmacCi/4JSaf18sgsjE05WhLAnoGY0f2PTp5O11TppRgHZDKvc98y5X
Fc3kZvTbtvBeSqqkEjtG68uBraUCzqcC2JgxIOsSG3AKqGZTUpLH0uIZbFRelY/1ah+uazwUiXsn
T1EDBY7EP8WIhU4LJlzPL89AIP1Xth8c65vw/oW0xrL2d58n6H4mC1dvlXtRNc2dPy2SGkcSHd4E
OZsMPbeIBrbcx0pKMW1mIPol8ckPgdvXSZ3hcLRZ+d8li18m5lZnyw0PcTsq0PNMTdpAbtahInnv
c33dSX0Yz5x7UoXbKEHJVwDuE4QiJ/UMZf+Fj4JSGGKV+kBnwRbtVAKd4QA9Xnnb2YL84i6pSovJ
aOSOldleHQJOovfwZdYgHjHmXjH8qOnC9xkE34gyJYxHPoRmC0GgD6wWDAtABlAur1HkZ7hMN5Gg
XWt+bI0YoAJiQT7R1Pw7NGyTcrt1zKlJvbZvfmD0/DNvizjxKH9Etu7B14ia/LcUdvMsHxvjGN+Q
/ItKNgM3cj8h06lgG/hMJSfU+T+T9MDsO38cqIzs+dUWPZ1Ykw1+LVDo2KagAmHD2FlF+Aszsa/n
3gTmabX9Uk4or+YqwhcEeU4Hlzrw1qImzsCDLd6hSO3kg00CcNwY8DmtVNqI4wP8x6e7+xWae/Mk
EmIpV1X8Nx3+mlHOxRdoLpJVmomlTBbm6D8t/2sk/AS7uYytbyCbMILY3WtZBIZ/EfBU029uXHYO
2clXSp8LVMyHhELF1ICtq+cbTIjTGiKVgklldQTAcCs3OWbyEurh9MIP/oQLHqllTISy7LQdHAne
Umf9aoq56yUr3igGMfzZtPHxVYLzST2agLo+tf+ytXM1zY8ZEFxf/y02uagJ+mq7+fOsEMSZoXJk
OzGaW2pCsMAwSRQC0k68HPjP6LlnbnbIHVS1ke/keaPAyL9gMrDsurHZ7uycS8pDhJt4NElb8RAX
B8zko2203pwSXr2J6OWDxKPG3K4tsf4TlYquTlhY7q44NmSr4QERbkPeMwpCurzg5IN7+G/q4TN5
e44nF8G6ykj+84wNN2Zat8sYgUy5dC2+VUTkfMihlPSWtF4+m0wNrS2Z/Jn1nwsbmL5ZmOn3fBcy
60aGIik1sg4NRR0fQ22zHKF4poSXTv58twPhuaExDmLCF9W+5SB9vvbZ8lDL8KQiuxpycpUBJatk
DB7528OLH5yaY1FrHLbgbw2Gamrm9xsmU/2j+KnkIqD1kOozEhY9+vEd2Kn/sUhnr8blwYay878X
gQrYFkdwmjj/X6jgqsik69md0iH8vWZHXiCcl0J4McJuDeQb63KldHENoLgrQ+HWNp4JIqGgNSx5
0LMKuZE9r+YU6Bsu40MtCL3WJXCYEfGbEen/Xb6SpSw+Dtb3dEyJuwMCG4vQFauBpdktbLGDTj/u
0ALM3pKsNINT9M3PcHjroH0EVYWWAe93IsuS7f6250ZxwlZr38p+aRYTNxxkf/GYzZ1RChLoWzsm
ZO1RlwBqpsMMSuR0qlE9YEe/Kw+x/R79fmid8ydVC4D+4yfwQBi6riErCZB186zEqMbL5TXjlVlu
tkfsnwI4hzs6nl+ihj1oGgfqBQn+elrrWnsxXyNnF1Kgs/xL7XQ0BHOt6GoVx1DB99iA0mgYwjzH
EkWPmV5Fe7+CpPnZJARjy1RKtUNQpo6jHvUOq1wZa3sB7WbnbSys08CsR/Q+fidGHs0vf8NeNodG
7ykVC5biaIFH7ODIg0kcBylL7+VTrhYoP/fXicJ10YGcxeozGLeyOfCs7Fm4+Gnchq1hL//aWjpH
6JE0rphn0HeA1+2N1T6sgHcoOmQC8/DL6PF9q/yeHgMBkqxKl+kk9c1CHFJeqAxsUsCGtAsSjWuX
qVr6X2bWlGh7b3ycgi/Ss+0INeDbjUCmrnbNiJPbm3pJCP5WOnppJCIu1+vkejSmAImq4FuXlWeb
ZAVQxTDCrASEQpwNFisnUDP+JA0B7F9t+WkRpB0RqvK1i3vR7DBYg4UMMelMugtNHKMNsj0o+hlE
1Xj47+rXhrcjljawVpvw4QnXq/xcC11T7GK6yb0CxEKwalt2cDSj0kF3yyHULm/TWVbM/fEgXsi2
m1PHiDxg1DjnfswcppZVJZc8ahJ5y8TYSt1vHAef0kB1r2paClYt0geBC7J/SYSAr3W4sb4QLrqO
sybkRey/ROkDUf2qjIG0JDPUe012a0yLk2NGf6ZRMg5ZfeEMS25L7sdAZH0A59HWwlcJhH4PwHnF
ZPpC7U8wprUv3rsA1CfjyBjzahmdBUpNYlqljlanihQ9JJAC3I9+tmSPuzJJ2v9Vcg4qOXeMMNVE
fuPlmhYxvgtKX/3pCNlNdOwXQqsRbuUQFLB39T7n0P8ghCgD38UYaifidBmVpWsEf29l3N4wiBVH
GdxMMtRYRww+lrB3gfwmlPYaOlUXjrFWVVed28Qj7Q1XHOriK3TRwylpl/0z70ixQAZdQri/6LAQ
OPU1GIMqXZkT7MVuOQYkp20SMc36euD1GtkbK8Lsz2CHpE1whKuKEoUWqkdwcGczHo3cqvimiSvt
pCfMFim7aWGb7vfMjmJ9b9ABV8aR/NstJ4shWFTiqhBOsKaj0LVnvlqJDQInMV/Yl81lbLIOEjMd
PVMmPv6lFzsh3P/VpZVirC7NzwK4w8Qt0fWnN0PN8YaqQPvkB9lCoEd1ITXHzqiO2rU5U7AoAKQV
NIHDFnNeqOtIqZmTCmEy+ZIYAxfjvJi6hsVETHoylvw1PhpAGeE2osq+HlX/XagyIaykL7hQEufb
3wc22zfD9jJs/Bbwlb6OxVtKoZ1qdfyNUG0U7/kwtlu02rVtNfYtxc6AZmpuaArB325WJ8Ay6pfT
01rkH6fwXR0VocnuVw7ydE+JgOt35GVj+eNru/XcX3EwLBa/Rap5f2//3P4lMNXXuR0QUQ3eGj66
zfGOUKrMtxAZyQieag8D1X90fOvhozMv8x7BneTv14M9S1UHmCJq3bwl7apMzwnqynadjij8tmUC
eK74ACNKtJaZLxQOlBG7oiROHMoBU//WMrmVF/ziZTaNvGqtUsRw01cUhx024SxQ8wkeIfTQqESI
/RXm/FLwiQGsUZhNaqzG4Q/xpXYRIMj0VfDUcNX3aOwJrT11oNtWt+Nku72zoMP9Gpjg5mzguRXW
nTekoiSeRwcFEkCbp/xXtzKP8+c5Uyf6MAbgX3fGzXoHUoa92YVNQ4w0/UHMc8cNauHuUq0NpceJ
XiluVhNBX4FhoLwvOrKe0SiWucjdruPgBQXvLNRqC+GDr8rdDk9gIGpcZ/BsMHidQWZ7cPLKkbeR
5FwoM/VLa74oulsguxB5fL+Y2wHLg0UdZfNtw5B8LeFv73WlmrWCIvW5UG0OW71rxGDQVVQ4szXb
DGVOnfx7a1jQar8BSkW+04St4A7SfqG7rWYDW/azMGGZ4pIUAHkUzxVu7omDtw3engvHUeFArJQM
SbuhqPAgavCdTV8XUx6ZoGI+Yese0fypW8w8HQoQVpdfZEaBCW3bsEXmcWG+FhhEPqA2QOlkdT77
ht6qMER1noLZLLfx9nd1CTvTSzdZIqU9wtYIhjh1CalVdlAsxmYgt4vJnPyyzA3fO0UxsKVRoKpg
Jz+3NB/V8Pprr8BskK4b89HGjLv/ctBGSKctsl0Qnv26LQhuLM6rt++As6FGwjIixEuNw62UvX8D
l9KrYko/cfRbHSUd81V9G5xYajduOXtTnqQZEzcBUmZNKS/6rCbK3419id4leseWa66DewriEzGL
cKxPsrcASeZJVCvDflV4YiaxtE3pJ72wlIRxYwL4IwY68Hp3L2wnBDUBpd7i0hy81P6dBxVKR1o9
ZUifGdVA8OPJ0D5Nj9vBpBEX7nWomFAS6fkKmyjx0np3pokMNwMdTfvkJCN/2jkBStB46fQgWZjC
YVJAQUcXiDTNv6WvGgCrpC51EN0xxZ0nj0fZLQHv47/0QEpGWVhRHlHAYWkFxbwTqjt1H1VAkAtP
DrTQMKcc+Lne+qm3Rf0V533VZFkhop5Sdw0e/zn3opqZJ2Gb4217KPBYiUEUfpzagBxp5P/q856C
tIZmqG1BQkBGzMOrGNDgWpVB4KstNwdv6wWo5DI1RBWo3q9AoVUclXzhEdm3Ijh7WclrUgfqwmsT
Z6GjQ36uYCc1lNyA6MQ0eR81LeJFkmzSx++6VhoVPL24SSPVZKqWDDjrLWKKtUAGd27FDv06NjM1
obrnbd+nYW56LvqoAPBKHCRK/2kdwWzARMrLKU1duB+JF1mxpTiGtsBu2MUD0V6qzbvu1YiuJlZU
xnN+xheN2O/VfKALmOl9Lcrr8tNOQPISQRjqflLzpJpdRtthhWRfsak6xJ9XUUF+G3mBNnlsUyGa
VbrBixK9Q8BjNCSYUQrav4qnbG2KXzpPZqKulCWHioL+9XGuWkO6USKVk8lkLBzbMU7zVrGW85Nu
UWqSI0mBdw7w4txcuC+oaoAD0EMKHfJT/GZZknhxzJC4KkX53/AJH+/P1KXxJYD6mooIcs0NANoG
WgrYr0X0oDCzot0wvrxry5dlSeNj5dEQT4kd9TcmIFgjqU60B8WlGJtFP0K7dQl5tkMQ81zoRLXT
SYV6sDi1Byzf/jbJTL6f7PoBGTDciIozc9J7t0shW97AmtMLTqDxHtnh8PWSPXRJX3uiwc1JPuwT
7mL72F9SWGUnJ8fi2vs99M135Ht6vjU/oGaYuEH/aTIuIpetQAoDXfFerm50hzWx2Otbt2iW2bm+
VmqrPdwg8Cu/bef50Rp8iXfyngVbZ2K+rLZgPdZli+ndtHyEsz0EA2QC8WCpM+E4eq4Wb3SJFTGc
UCcwlBr9w4pAtYEvO+GeTtE/84uUCY0toizzFXkQTbl4CfVoyol0WkS1qN21PLgYyFel/6qWg+M5
FjpCS4jh2qRGLrWv9OiKoaEH1b2kBt6AKPYfjhoeSyH7bOdTIxjNhxIgd6iygNO3rMkA33SGxfw6
D9Z3j0CdH1KjVI3ViOdO2P5cSB4k2Av6IsZAwCm5ArGRWi7P5mwHIoljweGur6qBZ/gjxCbIE4tD
w4zsQcHzlQkloxjY//eWGEkpdXiZaMv0bUDk9N1+rzDgYiY4/EI/mT6Hqx9TNOOtu3lUlLsoo/Ni
UELZWhktc8Ba6Clv2CNdsRXG10rqFsjuWUC4XHz8DtyJcEQp/rHgzN57GMQkv8IgeSuyST2X9WDR
PR34VvqIbSWbLiDFUTYBoGeaS2p/BFWCCtTJXLC5G6dKjm5tyHbwxMNsMXfyDVWssMC7VmeozMa/
1/zaPY64nRlwtk7yOIJECZcCs1a8FHtGXzwVyiAEBlXUfMfC/SEP1DsbakwYcECNlZYGFoSrL0Cq
xCn7drmLPCG8nKQl6ZpxuD73CAg/n6GKUmWT3BEL9xOBxcb57Ubc8j6DFaC6TLFiPknT+s/bFz0J
vP+Hs4WF72dMGQ8zl0EeWhGHmR+YPsDcOMHSTZpSGS1t7b+foNbkwHjMM0TexsxMoyuhQ7uY0m3m
eIfQLzX/sSHQk6QQyY88Yh30RvfHL8AQCO4olWYXaae4/AR3M/5CyBFiEMywlSs9XcKgdOuVx/ly
Iq59annIGLoQ3yNOVMhkH357QXD8uq1glJ97WrKwMq7GCzylGL/1Y1/mOgeZEPWurZRc6+KyLdjQ
ABLjH70/tEG15AEi8YwHXDi+jBneuc3Xj3M099ZnVYLSSTCoS6OtntD5JY3SzZSPu+yi3y2/mUK+
81csIO+2myZl0r/f1Jqq7jyEV/+Zmrk5CtHoNK6nAMGQHgUX9lf+MTQbdWBlM2yf799ov7RIn2k0
PIR8KEUMEbasf4Kvpnca831XELvpTv6mOyALlxKfJER4Y3gMSlv3KBuaH5capMs9rVPn/tToYkb7
+MI1N4n8UFuMRL5S6/PO+cJofZMweXFCy3JY3QrladP0B7g0bhEsBIpck56NOieWwppWxxUdb/5K
NrjIeuNraFkrE8NcTC2fFn0kNi0ExuIS9WUw3o106JxhtCyagxAwEJBnIBuccrh7tkR0BU/PigAw
10/ClITZVAq5WK7s6nX/Gi8IKqioLmEsH1RdIuu4ROfarYdgQwD2JNjYVecb4Bf5VXKJYsSIrj/Z
hhiflE9/SWzLOh4jjFYIRP4/GIpFFjebaM9ZeS6yKeFtkuoAQd70lsJ7gMAd3cNq6bdPUwtdCgl8
X7aw2kpiHvyx6Hy4qgN+Kr9EAN5KkJ8kySzXhBtlfo4Yw/jZN0XNs4XDZ8mPkNT8Nc0aJD5XPyZY
zmwEXazWV++tZnrXpL2/tlKuD7r/xbfGpEXvHK1qmWY+R/Ew3WjXwW4EcduMvQYQ7LbOPHb8KnvG
NqTGSzWVOz9/Xi7p7XlPPof3bPuSoYPCYaauH7TmGzqfBT/lG+7rnrwhDErDqTR9/PxvoQOJ29PX
OciCDFGCvKa3d2PBPbo+z2py5kQCi5cpU2Am8+4mlabXXT27cptc3ikB3ZrMs9SZkoaxClaHSgnM
0le0cBdkiBA7a7mJ71cXd/IdSohV5T99vFY9QOFyau8L05YP1PFrg/hwmvPAtee5CdDXZl7a1EFK
XcljTMZuaQghYx/Ouf9A70vSklLDaXkqN/YV8YKuuJTfkl+uZK+eSbIkGm19s5fDapy1PXhrxLcT
rCK2T3CweHK3+CgHfyDsjQFM3HK/+h0pkD80q3ALwVRL+dEyi9ZhVAcFG5wmVIFHw/lidrDojJxg
Wt5wybe9XDjdJrZWmjVW8RyHJ5+4BxOZQZ7H+Sm+KlHCjOJq2zEdFPF1vEJLXBUXeQv9WfmxHQEC
WS6HRbNcwydqC7jqB8hbfCk8ymT8OavXP9Ges2hLsWPlZCa0imQkImTeX1bfOxX4j1xpQNZcymZ3
zIkaXRcgkOc2iPVuPn+0XVwzUQ5OmYuXUQRgU2/VNYeXVOLMp874wMBqIpvnMfVukKQEq6JskzMq
NJHVUlbBI5pnVzkJZZrCnEYidPgqYtWP0pLZTqLYOZw3h+y04WJEvGaeNz59bk2UJCI5P3xxkFYh
p/5Wfduq04p7ORASjZVTs1v0ghDaRPaNue6tVd7b1vp3bsq86+CcCSSqLuxSNnuH6ikJRH0MxbAq
fVt6MwrbBBsz6ECCVFlfPw7m9KCXltQTLxwSpnP+1bFQvfp2TvtrQpiu9NMoBip3pd/kxBwhumg6
mFr2Jm7OGGTwCNWwMdNvBEBG2ExJQVbPT4QMidrsPeErj31/aIa/FndBrM15hac3sKMWKthX8IqC
Zuf+Ku+BRwRjEksKHULpRFTXNcsUEnW67UbMkY2gBg4xoR3MCtYRdvGy6/l4tsSQs2Hj7biVq/75
GPARvephz6MDU/PcR8q8dDmKz9di1LZ3rcihonCtS+wpVSskEy2Q6t20N3jKrpbgTkJFoksHXL+E
TutI+SCjw9ySKtj6pItF5dTbjklbz/er6TF8fCPhS2vKsn/Zm/RAwvbFw+OkcQTAAdIbEtuYP0Mg
dJZEXySkV1AbWIb/pxSDhf32I5wa1ehKcj6szFWcvFj4QnUW21gU7ZOFc41YqjjqdSdwp57R8YeI
HkfR3QhksUB7Wpv0r4Dlit4FDx9F8z4gyM5YHhICMyD8dHRAd6GJNnSwWoMFCq1N/xcqLYz+LtJJ
JKPNwdp1yUfHK+hANmMyg9ylxBtfLsCcyQZ4fnICQkEE44fpd0VEmhm5+BsnJR9C5s0p/GiLhz7H
lok3AeM0hdRrwhvn/j7P2bSUdBu/rBxpLh2RRE0rrvPvXjgHYc2WKFzTnOAdCtvrlrE4VRlr2MWy
W9eoyLs56+XoRfIdFOQeCwuJXRhYmxP3QtYlGacsp6ohsGOyuPKSku9HXOJOMN4N2OUvj1tFpbys
xLrX/LkNsl5hV9cRlPRUUKH7FDRp+FsIq2KqyfWoezRP0CjvrMQ0s8wf+shpXF//jb96m+8fQBPu
mP5B2GOx6V1aFGR0NrNAZ0wcg/PK9rhr9oiwgGUSPD/fPvuInFBMEse101FSBnki5RaBvoCsJ2eF
QyfwPlyGIgztKftoBLndaV+tgdl3uFpgAwIuoSh+pPfLPt1QOZ7BVzI0x1pMPCQ1mTWR5ip/eDyG
DVKgvCm9C7KXVjKA/x8fqaVruQnL4ssCgY6jnLY8H2w5X0VZDJdldLoVfplerw51JjEkvGXvqUvf
8V+8l5rOTCEZ/FbsdBHRXynssdaIW2sMK+BA+OzHCIhWfgeI+uGfGaEDLxGXuniIDWNLi2V6Nq2h
nkZnkHjjTHnG5Dhml2TRgG+MxlTl2IsplIFLiV5ojNmbc5RbnvbWG/gMtXvOzpzeHmsDSU93Y+um
r5vfkKSYi/PhQyuTsAfqynPRle+8WnuEF4B02UPyyKaTzBlXfrBpSUBpxN760aWl4jRyqKdH+xXp
mB64mKb0Ku7kQoEW0ShyiG2BH22GC0paEpMUX0i2yay6pdRaHBEBoX8De+iAlKRRpKdCEeiMxME/
LQRIe3s0W/THL63qFMxVl0So3fk+9IM1N8fVK/mHhg8qZ+58nFjAIXmqov0B2HrACORsLiz5Q7f9
R4QuMM9eANOgH28vmgirNdARMCaQLEfzuRDZ51vmgr7K1+93k2xVffzK2DhFbCYbjl57ReiTMtC0
4JoN3vwtvksTn9Hrw3ZOsguNQjOBTvT2zPFsgZwYisColUPZr7Jv6Xn35aQZk4qfk7xXEGM0/WiY
TAn50I/ciFurSir7MmjK7LVqnZOU9gR/0QDyE9sIj46O34P392bNcMOGMACYyFswHPvyG3C4JyCo
ukKhPxprN5cuAgGKvURkmrmur7xXJ34uIuyRxDvWOKjLzrZnZwa5JRxLfRmWX/LuY2BrmtxlEWDG
1rcMX+GauNnPgXZ0fSzuIJ/DrjUAxY6pVaqck46lD+eahhVYKPAwZCuUUz6YKz/5pfo0C+5xYV5j
B4IHzywbkGifOJla4NHmyChTasHWOay1e9lO9g+jjS9UDlBaol3+Xm3Md/8sqRFVjFwe/3Eu1Hu6
cSbrL5MaK5hAeGMuhavKTpa0PdE8EZeyQTJAHyZnXwk1hacBFcLGFL8rMv21KEg+MUwhGOLnx7vP
EpG0Ine0PNr/Hui0UJ4aicSJj220jNHdpGTtfMUCfigRy0apdy6OU5nU7vtnk6GuSMhdxK3X7M/B
27QAYrq5sgmHtI3Cexfgzke0Jbz4WLX+QCvlBmmADSwYqoLh4aRX1InZCiDNGf33kUsu6whis3lV
21nXu2e8O0FvVISTGyBtCZmjdpADuDsXReQS6SbdoJAyxud/yJk/2aQLf2D3YopO9m2OKRgkHVjG
pWse5G0Oan28ciArI8JR9aq1TPmU9eumtXhElhe1cec5tM/q4yckNxhwvHxJS5XpgJWibQ935YOh
ZDT6d89dtI1S1VtLVmH7QvABn46fBc290lUgT57AXMsqvNOP0kZmAP9NZaZZSkIY8klSdSfg9XnD
+bGZJAGBRHNy/Ji9kv4YDZjQr/43aZYlNkQ2Ti2p/aWsgCDZIYgqQ0D//O/f9DfxHX/7Ak3JqRBC
1+A30SXI58Acl4K8omWQ+Zoga+l/zBzLmVwviHayna3K2YFX+lHncp88wsbGGvLZKCzLySCPYghg
zK5RxiOpxETPMnnZ8OgNe60GF1533nHUtnWCx5yd2zWgU++rgIYw4XtCksadYn7TECNienYte1lU
bS1r0aiBI18E1QT3A33ZNm3YljEyuKjw8B8tK82Db1WZq1zbilS8dxrDLiewHWueknTUY5ewIJS+
TOZvGC5lKNjqsnIRo2QkSEMrQZREI6/EN9kZ/LLf8Xo0Ufvw9xYaiAEyeYgwrpjd02Y1Se2fkmeI
7EUjTzleYCCRMxh4C/VeABeFNL7C6peQ7dvo4zRCf2TpWqmODreVP/uLZXKyrglbkv5oVEdRa9Ul
azRkytC2a3eBW9yL5kQRpTTsAqezIz6xQBUokAUQVgmHFwic/e6Huu+MuFE+IupUnUhvib+odXfB
ZN5XvctKuASYcCI2aKlhMKT4ABzIz5u6k6UNkJ87HAGTKozMm1AdxPGAwq0jeYek9m/eUzDUK/b8
/OMqxljqB1UQ/341f3RqjFmTvGS2k2s60JJq5LyBfiinw8Z54irpgiXkTy6MYrkNcjFHlL6wkk61
WUzgpy7UfxQacprt5gBl/2SpnRPNyDVuWYpIc8Kvg7m3bjsreO6HJ/79jdKDXv3kS2nT3B/OfbKo
tYIXcpWN0FVdvc4cbjblRQM54jVCX1sBWyViFd3H/VAqGIC9YkAWYDzQ1f/BWHIE0H3EM9vIjxQj
nVb41vgYSfD+nTvaXiTn51A070uDWnEf0RlgCeAiUlg4FTA/vP2PxHKXXQzoPj4DcyR4uEBkVFcg
U/In8BDhGs3GKLVHoDDH+RCE1GcAQSa24oePuypsn6ME+GWo3kAxeaOm1drS06GMafv8hik4yKi/
qxzhFdPliIPbhgURooANZtmFDoHFjwRysGd+2aqjn03oQYZl+9dYZrYjNzXNN4ZFGYIxxUL0kPx1
YgHuo9F45mdH2YiXPEQ0C5/rppw6v1S7/sIxnjqtzL3qF36nl2SALk0CYzQNZETZ1pBcxNGy5kau
uFDW4DJzMpEGdbaR24WLAjdXD2rVZxux3IdGchF31MQ/xe1ErKqGBKSjvRYy0LWJwTKWMu6qx5p5
20rp+pYRG3O7mAXnPa17fMCUztXeRqPmP9+uIK/YJPUZdJPPkMN+Zrmq3tGYObzOlbENc0T0a7xp
kmXtP8GSmFykwcj/pNbuiOlbbry/QIRQcfUmZw0jzBSa0iYjyBkIb0KBXfEOwfBJRVt7Qq7+uylC
q2O663kGm+0k1WTVd8w3+yAXi79pURdwTuIs4dPMArM00eZCaQeH9ccNSrNtb4IBdi/U8U4fJGaN
bHu1Rj7AKITUaLsFXuR5dBJRcx8XtZr7yPtc7B9G6arLi/WF+tTMei56Qb2Wmmzu1boIqVPI0x1j
DaAJiXQsP/TipXAndIWqW9jNxF4G5AvW2knVkqU0lN0ov+/joFiv77TEeLA+EDzXHYf3ZWXE/mBJ
JtnYygZCDKt60IzT6QLHZYViePtF1uIvuwXHpS78Q0jkN/vmC49+9LeZ1haZgxZ4wDh8wEIu+Zv9
FuqKrZj6Z+1UazYjQc4J52WCpz7NrSgKYjkN61SD75ohcm18ucf/GAJ8mZf7rV+Nuk/WX9dhyrVE
bECtWlPVQ4pkT+5zY0vudsIoLHVZwlLE3S1o6JzH9CndeEQ4ywi4j76+5/R1HZpVp+o2XUUty80h
4Rt9JaRDAqX9haGEwZwg71Y5z19qrgowgSheen6OJY8IRTBQMqF76Wizi3n9VJXgbYPM3rNcfyCE
T/g3zccJPMn3ulIAdCC12nEwQbkOu+RJSqHZyZd6Q79TBm13P1Sp1wYkKTtp/6MZ/RafC3vLGe7a
tkfSbVGzpmTGcWK4+q2/PWn3Bpv4yhIAgyQK18sN28SCtxntnKWZii84Qh6jDI0mAa5pFXaJ5U8o
7t7u8QK5fvZr2AOfUrX5t4zRfZGJln29Nbx0zCq9EhMyZ/eP9hEexJkjS3qc2Sg4/ZSjB4n60DvX
LRqobQLhAX7yXVgUlmpxlUwBtMbJcGvXpKnS32ql1ejk264cUZJiz4+LZfoy3q0+24h0/uSxBzT/
a1Z4y+tUPdSOEL5gfxNSfE8ZNqIFB7fu+Q4x9NvYTdkuMdR9Ht7s2wqur6zrXxkAdSn4RYlINBuS
4YTlZRhPjLpn7KN+WRuJKlj41qwmLo9aFqaNGQGrGCpv0IeBVbjZBNp8dMMaROXwliF2+I891UUc
j/lTRDNgTRLTL7sP0WE8xYvDGrxfb54/SSQAo7TgCxX7Mu4l4S4KAaDAdmABY6g0BzkQ/VTThsuL
8ozibmQiAclMAYTGFYVKGRliE3mENZBfPrhD9QhhYWHx/+z3vPBVwwQ/dfz7L9xgKF3bJAK2Kwsx
9iu/wa5T6eF/Vg98rWCvCBbqKsDKqMnzW1nLs/QrhtzzChl0CXRotIKsFsTMMPgvtK4Ucgn5DVV0
2niwBqic/Tj2FQISXMv5YM4f7MYZb9FwAkl96Ip3/fvYDpU7Sd4Zn6qKe+Z286IT0k/xvuyumzdo
vzbC/DxCYViM9pGnX9y7z2WzW2J9RrimYRSJLsA8pgiUNcNbHlMkvMuUpHQ9kXYm5LTxLLPfLv1y
I7qonDuF5F+88tZVICt/unDpusZtyk/NIjz2PARg0VxdeJItQweiqu9IrXtjAPAc6z5ibINa+SN0
ISCgp3YfQ+terG4+kKiIOIqVGn3RuhDQjD4fkzQ+WIW6ux/NV8n7XkHvxsWOdA84N8BBFZv32axF
NbF7mLGqB28o1w9dVL0+IEKPnMLPm5D/aXyk/P4dm6UoqeMgfKOd5vX/M/iUc/HAm1dVMzjDxiFg
w8KhzJw23WUAvAdWqOK8V/WjqStFLnXXNyG6mg6u9+Vd6iVf/VudsMOb14MD4pm0RRtMNRsDM9Ho
PL1UY4F1X/L4k1PYy6Z0eWFoSKMsRI96YQz5QsRkzOWnctdiP86E21tEuu+/tqsCcG0pQFhhOvs/
fWbWJF1JNWLAMAPT0oJEPL8I/NGzI3I17jxEXIHs3txavdstOlO6BZdO4TmimgyTDvOdz+E5c2xL
pcn23VaOqoMHMHWZkFVCpfOJbgdm68+HZxpXbhR0E/TGkCh0h2tyIxfQ/rSzyckG2hJp4r71Zxw3
dIPV/2fVq1suXVh4UCzW++UMVb/vL5rxPj0gJvJdExTBzgWVRaq7SgX8F5igGGfoWf7/7Mk4G1od
2YLB65I2jCGR+WSO0ziMlzKTTGv2Qtqm/Cn1eQ7e5exYuDwzfx0S1OApkZLj0cvehsqIrOjcsuRk
AL6lOt3YzR9QXbZZEc2eNAwCX0UMturYl1bFLb0gpfmYSLOBkKmZ9JZSUO93/mSe585hnEml93TD
acsM0wu4JRKeBLHCNbJ/0kzKcDcdI7nocW7epS+cQviIN+IAbhtrgSWC+qzuzEjE8PqqF+Z+jCIR
bP0kJTKp2ASg/5+6thQXk7XKvSeG+kEAumXOUWGw/pjelI2OyzB3tl7kmY+ULOqQxS7gi1XEkGmh
mNh85nb0BirH/bqgDWyvUd8A272PTNnTV+JJQ1vM+NhuJgXk55ZpIT2L5cK8FIjt2TgiJ982aaL5
CeiG+gTpJLs1Dhf1BuNs7CHI4KWovotK4quaflXUTvUzo0wQCeLSSwN3CNpmkJt/KXwclYdCHKUd
JYPGdPM9T8ydVnpzDiwmXO14V9HxEB8jYpRG8Je445Icg7XX6QaUapk2SBlCvBYfX1c6kPGh3f6s
P8V5V/r2kVl1jWjyCgfsHMgdJauXFjy63FjIcZV67Gkz4w8V1bYbYL/e5ZAFGDwUdhd3GjKlULe6
3GslQmBuNMT4hN8bPsaRcFvntZ3ngovr5kw4PqXfYN4yZnqCT1mk20Mm9HI+wWxJit9VFc+yK5Df
YA3zt5HZdjVmIpVUzsLqswbM54mSSEypyM7NO5VU1rQEAzx4ob+o7MkoAhKnO3EgthudPeRmgfq/
ycEW9iyC0/X8bctbzvAf2j6IiS3h7gAluIdmm4VGIOPf1D9fa36dQpUnbcvCJziGiEGBqroFYkFH
p80sZ0T88mT+YK0hTAwr2tvjTI/EtVrL6YDZBZhJ2PkpJIM/fS6nqekZ8JQolLACHQ9xz2D9ru/l
KfYgysrLqKUADiVvSe4pUFUb6fcI4UgVGn9gBxwEkEdL19qZKftIO86AC2/PoVorkxfA3OTTW9Os
rdBcggEiRuY31gmTGXXb+bOEFkEZYFJ2HPAfaiep8xFDTZrN7tdpNRv19zuxXsVBe8YEBn/J31rP
pRGX/oeUatx8DTi207ohNdhPJs7EOneY7LmmWNVLSHgDI3WYrvSaVSjAJEG6iKjU3iEf68lo+7PS
O64n8aTMEoa3UA3wu3JrRxe6iXJhjRjp47iJVibedI2yWV9IfPHRmWh2+dlxV+UZljMXscGTQ24k
ev4LvGzhinzF0l/3ceouAmX2wsjrvchNg+8sG5O2zZLgZRGKoItd2Gb4x0pLYTIPBRla9nDv2Q4f
0SENKGdPMPaAHxww7ApBDW5T7SZVVWPhSEj0Bai9nXwfR11UtF860vFXGih0JOkg920i+KMtmKiu
4eGlxax2DbwORmM0AQAGTAYuexBlFv06ZjVyCYXt+UriQjwwZtE+ymKawBey/cDMusETRVm8JsJV
iWCxmaOQUV18cc14Je6P0RmUGSCqOVHkKX/G53S8I9gVXvbbnwXlJ0uIoSH0W5b5pkWeVNGsN0JV
Y9wwkvKHUqgVpUtKye6UDHRUj9SnofbPzQb6oG356PapLD8gNDtMAHPd9HrPNo+z6x6g0h0QinSC
teuj1GFbnV0xaK334XmzZeCU7GKjftk80GBfGB5XJAf/aFrfKMh/QZJMXD5tFCw29uxVPnmR5dux
OqWNKr+dn9x545G7kErzoAYuDnk/O3OzZTz8ABPbRfdCc21QLHfoW+OgsZkQqbmqRcDHPjC8psv1
19hMVEwbXKFxydtzxmLRdimeITsFEiVg/nN6k+vYSg0WwU3q5BOCSmfPj3k/qNpXXNuVUa0BzWOz
uXe3dD1qPd+tPFF7xtSrpQrRMChLEs/NBjIKG6rLtWxSLkN3aQeiM23R39MyTXY9OjAu/ORdvy1F
Z6fl78EraAJv4n12GEhsaTSZwWvdJkB4/D7nUzDh7wfrXLnD9h4vUMa5pdk/bGlHotz9PUI/zLzq
18dF505wSBpa+0ipPBKF/FuZMgW4HoyegRepW468I4/CKDGblz6ctyldbvVvgmvyZ4j6EtDKTc0k
9eMOT4+XxpcsMzMORySe6fmlIeIDj+VJU93rw+Y+X/AIes1qGXs0n/Y5sjblJdwc+JIF9U9pDnRB
sR0tH7KQKSN7Cqpa7g2fm1BCUywuF3bMY50LcEaOIHCd7UrOug0G6yTI4QRF3B561/w1CRwVFTlJ
pL73T7TYZt/cKk+qQuvDpv1RVjk9u2dor0JyMiMQLWmzv0YX8WfEJP3sD4rqewy2sH9+lCK/CWEV
qz9E5IIiJtJbAwOW/PGAdVxIB/lgalfbzBKfC4maY+xrlAzQVmvErnbRvP7R5BP5HTte71VyFxt9
+107Ddeq0ruFC74nzFJblTKx3IQ/CrErDXZKRNBqjQdWiOH0W3yr0H8lLLThaTg57WvAEm/pTCEH
lyzkJTliUYDNHLp+ooNvNvtkMOzVsRoJd4jLE2D0OFP7hufc46salu74Nb9vC46tTJ8qVm4hmeGB
P/DZBWDGJI35+BsAxzdMlDsr0zT1UBwDHxxbVGbGxNaIaT6cBJSS1Y+ZsF6nR9P3sjwqQF+pczG6
PQmQSs4wojr/UJjxwhRtDzYZKYKwHrkUoNGXjZEDtKj5rVmhGaENIDc5hYSfuOJ9TYlOi4FauyBj
u458Jtkgq3HJ9KiksSLMg7UC8MR3wsSJ9TBV++z9AW6m6ZPQiGsI8zjl5MRvwxXrW77utCKiqp2M
79kKOFJGYIdcr3IcLsVTZ+v2Yf8VC752rHmqYHyHTCdxu6TszKYRJS8Z138XvaWkMmKNNtesonjx
dZ4VI8Lm4Sblemc5atP9Lg0wJYa6BgqURKvDWKdl0G4Gh7fNbMAFSaQiJaLQ01KtKYRUpKjYcD+a
/hvKp2fqUdym0crIuUvi6pubAMIfh1h/QmKZfnrI/NNFAmMD6Y9CbrHIhLdOU6nwLxBJqUKqzKDg
lEsN7ZoI5M37/SKBejnMFyn1lL5I94qtekfewM0hU5epiXzVnH8u7/7aod62QULlmObHg0BdmTh9
a023q/eyy6pcs9RdhT+6ExJj7whSVcmo6FPnhksNvvzfmvhodyWTFrLtoLfw4cQq7oFurU7NNcrD
NDMYqyy+EP+MMEyjt4DtWSGkabtyLpqIIqnf8Ce/PyfUjf1rK4+EpilyqrwBV5vcLvNpU7HEklAF
5b1HxoOImwOWBg+3sBdVC1yHg2GC8o4TToagF7787LPCJJeATFrmExMy4XyY7s7+WwK/uNOJCeqh
GtevqND3f8hiOL5lRNRIgvmwS8bLaN5Xe8jIknSw8K5OS2Ut8+Y8hg0NuqYASZN+LwVCZwUZmXq3
VlBXxHVVmhufW0voDtOduaLPgD4oK6OebrsvW9SxbHvgClTA3VOCkfDNiYWGYLg8SrrSE6sVw4X3
eKnJYJBPtuCHxAgGgpPgmsVQOa685PFZ+0b3YEfZA/6zfYZnxGzW7+ri2LfpqkN/8X4s4CyE/Q4C
DLexakJv6Pk4UmM4mBKHnz0snpq7wA5kSGkzndwwvTqDhsyV3o1ZrUjk41BcviS0otl8fKVTkv0J
i78P4IAB1zOr46Jgl+3IxPY+a8kyUoTp6m9Kt3yNDyidSBvZ/z9uyvtcYW2BvjBRQwVYhwsNbAqb
flqQ5qGQwiIWQl5w3ONtgru0zWQQbTAvU1pAjfOSEepDNiHGlIxz6a5A1rpQJwbsmnpyoEjXqSJj
TASw+eZ+NuUXdN1RT1UEPzXANiqy8c9qcO4WROKlC7iRzaoXBaaL5e+4G3zQYGTszWnVVoYOVaCb
BjAtY2f4094xTRReBqvAKYsspgGh4aTwbVZEtBiIen8Cx9XUJfTRiDq5lEf6E43C0VDqKQdzSWWo
zwHPm3q7huoVBOqgpW7KdEQGQipToDgI8rfyOrzZTyS8jUsn95RBSWWcZrX2k4SWakhbDsoTTj4G
5u5RrR+V0Fo3MaHxhofV0IfT1EXiaJ3zml3FjGol+krGbxhIN/ivNyTU4w55EApCTVSqqSdrZ0lb
M0d5EZ3k6NanOyG+QOSNe2MfHipOsCyhTej6J10Hke+XyxZXxA0Z5RuolOCv1RwOv6ZjNIh8Z8Uh
lwx1xQ8Mbk/PR1ORXJnuLrEgVUrAcsPolUkjVLZBusRhbDj3ADL2PRTa83SfuD4eNdULn7OdPcld
jGnp+OKRM7XUIgch1/iSQhKN3nYGb28sbKX0sYhgMyslM18GGDXJm9j57TuLLaWeynxRsPvTitgu
gKm0LmyQXdoCBEFKh6tupL7q9SDG+FI4b4mHkH4AXSbvd66S1fx6J9eAIiUBfuioW5mNQtFU18z2
SsvlCAQ4uXC/zz2Y5QQxeckGRk35BzBcOOsJC3K/ICBdtIj6T7DMJsWvmZAX2+8iQQvq0mbjPlpT
pwZqAzGXGpFNvkMFgdty55dD0Z2ThP27EZVo3Dxz8x2BRJys5Qv9bcQr7yfLqxJ5vBM6MfxTMXOh
3iXcUfseSUbkUleiM3AJFk5Q0BSAiyXVUtBDWrsXzZj4XbJArJVcrmX034QOWzIOdUjNigsJuaE2
S+C4RSivE/lSn/Ze2dJjtGOF5qj/YFbPInldhbOmBQu5ZdW/GrOMWw54hiNIUBDOhtIxD8asjI9V
D/4VueIz9oTLBTRXkWFm5Gh29suTvL8dp39iEkTGA/FHWV/Hft+3ahDRXS9XKmSFDWS7ooUlFMbc
dN8L4/IE4G1laYkFZ4T48AZopMeVN2cb8TooOsu1Wwjei64id66lXVhaHs496+YERi3NdZofI2Cg
hXIlzpt0qLgAm5afIQ2/AjL8sPGj4cv7HjXRM/m1j/x1KG8IJSBkdUAWR4Cd8txqPZHk9O4TUJQb
kQMi1s0MGjHWE9uNGLQfEeKolaKYqGMtLoTDm/ZlOw01dKmt5P/0awjf1tEIgWv2a7HobnNbvYdD
xxctM/ABoYH6EXEc10Hvd+bjuvnK7lRCa5j4t8Ryz4GWP5OTmlNPpD26lYeea+CIt62GKKZrhOk+
4mEan5l+xtuXekBq1o8LCN3A5BlZyjqBfBkxpCYtIR6l85vBZyUuYyyKKuqOUlNSE/cd7a8leYBx
2l8eILv3htg2ioubYr5I/yABrONeYYhrx1oRUhWht0b6z1w/Nv0yAoKqflO3+EMjxb1Qyzn/9IL4
GfIPjP+jIS/g307BUwv4Cc+uonxQ4RCgFKHpykJOOL4nSn6j02uDvXrenLzoZHX+kYdX5IkMllJ1
7xvk9v6LYQlfjSJAe3a8lrxk4WB1GQYA+xdFLB3r3VAhfGt/J7KwvmOhoK1WRbsCbnzZHaNuWTaa
Fsh87YZoG1qggBlFthzPBUFmQGlnMvR/Vl363A9/wjfE+Z1eE1g42nG8PGCwguQ8OjZz4sYgSfYB
vca8L1baOkIstHiMBoug6lPFMJBVOWXOJWenmw9uruXfAamhvllJrjdnpBdweI7O9fxky8AltZVi
1UkGPBqDoAGqvGw63TvxP8yinIbDxhUQxYFT0v1m35ovsM+zA7v7mCJ1GCcARRtaGNOwKyvf5oap
uGMLZ2WgE1nc0kg0pcY0hH+yfoMGG3nfmViKQJSpmGZMKfJD4njAMEZ9WqkOLI1a/ME5LWErHjos
HU8BjqJlSJujJpMhq459YBbzkaKWXl9kIsJBIiudTOrIgbPyECOA7RaquO6/WJfW55rIJFNDc7ah
jei+quTFjVLm1yxq7SVx+dFxKS0mGCYQjc7I98pZpNLSxdTIt4xRsJErz53nj51aC7ZQlV1188RV
x2+eYZqqE209DpntD6rOpHtA2lYuAtwIcPvzEQVoV725Mc/tCVDC7b2vpjq+60GeWI2M/YmSCVtW
3DGqwLRZbPxHI3ttBb66XLpgQvMnC53Q5rB/I2i6ZGrUXH6e5cnzm6KsOuiwOScBt3JG5QucS9U/
L3Tg76NKo244oMDyMPJJ7SFkH3XGXgj/Zju71nceXi65x+LHctryDDHjYG3C8qaoj+m5uaLBpKkv
3q0QZ4m6y9jUELA4yjX9ckH9YZGgIvbUo6XP8GXU+R3src8ap5/TcdQbluJiTYpy0H9EUaqAC+zM
YblOO37R9LsvcQydR1va+AZmojvoj1pw9++i6kpDZZ60R4E4hPIG3iyaA5qe/A0i3drCxwhAi8IG
VojYTqKgWOmurpvK6gzGiuo1keoKm9Xy8MTYul7SP1g5Y2exbRLFdPAJiS2dI5rsIPSKhti4Pic0
7sCpVyvs3e3cPmEMhJoo7nxILZ1GBWXQvZ7+/vGb7uq6BtcJm0kUpzIzquq5PdOO4pHHKBLQNRak
N6zjDptjU+yMWfv6mFFFKPcOauNEbz3Pat2RS3jrxKS/g8pLaANVbMjXVwVincuwSkyU4w+C/BGV
gV2qAdYLrgyjnvbipS+2PJrCvPmlsvQjcbVASJ558b9eHfhdarijK8iYP0f1eps+XJ2/MJRyuLVC
8pk767IpmAnMw3VSqswgoVMrG76o1hxLdtav9S53DZSlCzsT5CojKC4Sk7asb5bMCHoe9iE/oVb4
7v8lnNkH+/v2Ge9O9VlRvW3+/NTwPogwBBxPN7ZwK+04tJb5nZJi9JHJkOKAcIblw0x3ZdjwbWMP
AtaqqI527YdlniW1/sD3ZVsu/9JrJVztFm/7SWCbJpT1Tr88FVci1G5GVNN/X77GFx24rqb/q0Bp
0GdCZ2qj295fivHpv+a1sAgDafTCc7lDY6SMO4Zt0v5E/Q9pYCeM6+honVFxYmS5t/rJRkDt5V9G
glHbm6Pon30DUB4pYJsKKyigiqTVqeohmp27eexVYP2WB5Ca2I8lTs10sVYkgaWOyLzlodhxKptA
AHhocpNnc6nKZyQ20GPoCkKOwCxs9ITRhxcDuKNp7nhjYkOnoD9+uI+NmGrYZOisK0PuKoPnKlWS
1wKGCKPS19GFjDtpD6j40HUHBk64V3SeJf0X8eqoeORsAY+iTChURqi58lhAeQI3PxsWlebFnEBt
oEQpJ0KvbCmvq7+IxLyExgBCtmPk23ipx8y7d7XbPiCgRTNpUXDLZhezxCjG8b/qdSYdDf7sF53D
QHh1RcaD+q4ag8i1bGhgexbN9+48PGZlfMdhxtI1fHE9i8vZ9Y1cmzAP4stcPrek7NtcgZn/5v4F
RsRH6E+Gdw6mqWJexrzx0APORhAqwQ75vUmpV1TEY/bPiDqNcksysYs7hHn4lllwZ1PqkzTzzJdc
fRV1p2lQr7kzadP7RTRjPRZtHL5DJmyxntMli6y0ri4Edeil5UEClk/GKYMSHjPWhXcZsEIRaMyJ
MnaLfNRkuDQiXAoeElQC4QeLUzUWiTl/qiTPqQDu+VqfCigk4qBHcJeBoZ2gW6zziqtUwKb7eAjV
vn9B/YmVxpb5hzrbECTOAh/Hb22CrDHtWegJdIVS+q8ArpAeI+d35DtJkfLGAJ2SLxQPZF3EiLEl
vFkSo23eGubLnFwux8mHsAe/2T3ZFGlslmzdBEbFFIy/3XWiKVLWqq3URYh/Y+6IX103TCqWIonK
uNos8whK7/TC2YSDNQaA/hbyV4JYdM7Q0GkcJrIKno/pdNGl2oaWn7Wk3bW3VILV0xFyheUhU0o5
f/PpiIg4o8qDDjSs9lDzrgeIicZkyYI1cHkDTtYSZ/m4l1V2IdonWZ4+dBGNN0PY+met+c264nkp
rIMVt6gMfkj6IgsLEublK0DVrrIRNUM2++9CCcFGYYJ5ON+BiWcb17Q9i1UKcctVfk/CYgmtAmSA
6Q0l9TeQ/OB1CPwMApH/8aHfCePvHd4ZkXq1fjeCU73i6eHGSSuL5mqBucxN6wFx3BSLSE3V47q7
30vlY6eSRlRN1hmyg9LSVpvS2l8n9f83OD9/vZWYJIall1ePqYTJOQrm/wop+Ccton9J7fP7tJRm
rkhka/x31LmTIZM8J0/WifdNHyCqrApfSLYeCSjnTJhQjX43Nl7rPhdFE4MGlOLYkJUFfzlv6zJR
NsFyF5ZoSZ9PjC5l56lPjeTXxPgim0eH7uqjaoYGfcGtLM8p9apTp4jThojwM9R723G4Mt8lFdgf
hI8RGyNR7QkYPwSQe/DwdwwDMqwGGmU/fa6YCzYNouOHpwK0XFEJXk5PcdsncfWKJVQX5mc8+z90
WUNYT9a5HGnBPW3urlq86a8Ph/SYnlRKZMyVvb9faTqrNK5okUAMlgE5TcpwfdlJYH5x09zh61w3
MgGL6GrUzB+lriAIunJ2JoOlA+5R1ElTRPDglFCaW7vy7G58oKZonI8EIRBehtCOIqQY6Swc/4Hz
sjnn4hbXgVMkW6O+xERYMBMbQysvQDhj28/+7sfA1YkM0TpwYQAkJlxhT2O5sUTZMgMdLkiQhAws
GNxR3HAkYbEdlLF7DtZFD8d2xzr+HexZSftxjwAafoXq/L8jhCcH/fBHHmLsxPQzL67JND80+Del
YZ4xww0EzoqoMIceHZ2bBNipM3lZJGW6v5C8IJ/Cf/yjaQ0QnHM7udFPFkRSaB0UNBKVshhAh1d5
tKUDtKoxbHBS5Ea6Ba9dpbfBRbbRmmNTG3CTGQUASYcRnZfxScR/z5EZH7+3VkO+EZa58v7uzssP
6K9L5NCfP7MnLfxhG6Ab+Vdho/Jop1EidrxxGhumgzY9IzH+tkjuam02HU4Xfm76B16qLP2x8URg
YmD86XBp4zaQW3h9/Ydr90+9/mIxVPC7TLXmCbQ3U4e40268sWY9EdCh4ednfOqQcZJStxbCMkAW
jD9vGS5qj1Fe0Q8wgMniMNqDFahxLcqbKhriuZzKeOj9MY4DFbobKj/vehcGxwmR+MA8EszA83nF
7LnmMrhmfIVH8/q99WIJ2X/kpAuXGCwltNh7bu0se2rcx7bbXDvDqusTIISARvBXeDjTOAE2f1T4
GIlN/9F1NCK1KQMLFyfyDEffg//rRasORO59CQkstwtELu4VfunvPBfmj685ShwwYfemnN8iEgfx
BmEwGJhc1kExL8jWYvAyj0KXVXP+tC8MFUrr9IxvfPFAiMcNO+BjypH4oheqLEtIcgVgeq0g2xOA
XyTJy6pYg5U86ULcPph/T40tFbfJlGZu3Rhmm7RrI3pUYPjDe723gvA4rSbmiYx7Z4Vb7gBNiPGN
+nFAZtjO+qe8F2sAaHONQlRbZp7EwrNuuGcdrOC9K5HPO9aZ5/9v2Gtm1gIml4RIeCihlgohCEp2
1d5zZp+rNys9r7BYpSoRE3+Qufa6Y+NJQ/N5lfRlwdmhmVL9/kl6oNzmZeJyj9QfIesD8osHGNTM
1dRQcjQz6a363i0hDI9rndo6P+iXIOF24FS6/wrciMBU6+CQKbYMSUNyVGQTcJFwvyA30ruA3iBx
Se9gogCFc2p1ZXB6M+K5HhRwERCc/L1olgisxD9N27PAeWO3yzbtwkzSoyeEdEmGJnbbDJHPc8+X
2Plm2BfzKdEhVeOsmPGBWL7vIvh/vsugVMu8e78XwPq2rxlyPY7gMvO3Hoy8nvYmfrdK6VGZKO2Z
HqHOIhbxceUGJqr9ERFzH7iD79CdyRykGxZzzuNabqwYe4zD1TcCRQOgLluo2dy4h9FbnBlejipT
yh3nkzaIBN0x6D+w6W3BE8CwsvQ3k/lMTVYrWCCqQLd7K0YWpbCiD1H6VbBfK5scD+UsXiSgYcTk
n2owjcfspzobFHYacoWO8A0imF3Pj2DumN2x3XZrhKjD3DSnDBBAeUP885KVuDWyukUoDWvsHgPF
UHFjOSXLteyTOCXGh4wIlxSkiKmypThwzpBrwadCz5ALMQL4oTO5KeMsNNWb8ojzGMMgfzIuAExO
qgsck9qBjORhYfLWCZogBjyijP0LL2NKHYRtmAEHP8NTBy9PimLJl8Sph9fYcyDO6BsqiEGPV7Qh
kGcJeKMf4alXH3/SJJcwVr781qeFzeGGqu1xdhTzNxrfviOxTmCT35ZSjdhHM6Rc3cMpJxj2sNel
QXgcwvmYjOQKRUsU0sTOwJ0qux8y0bWE3xRAS6TtzrwpAouYnA3XTlmjlveuSj9HUF/wvgq5sC6T
RSZ7ukrJrOglI72gcOXX2T7t2PNUqkjXW9EPF667PGALsZn+C9yvwyg0wo/Rzk6qRr9/jj0iQEet
SNjks/MvGWMwky6d68GMrlWaRnyinl1VMISswl2mnzcALofsunXNUCUy0+pVRyPpI65s3lMXYaAb
Ybxd6Cpc2LE9Eb7fM2cIKN9j/Hq+N/plCzVdaTSxZcrUJXOE/8VUZXkuQ2CwufsKK9kMJ3abAa+t
RP3kI8TkttgaYl27gbzyX9VlqvX7DNllZMTnpU63TDeVPDb0C6ijvIctr+TBYV1oo3IzjUPV7hcH
HiGdUQCaDhK+ggaCvEMe/avV5ZthjMu+KMY1vo/60Wo5sGTqg9uMatt8Ds5yxxjRTtszofhbqeKT
L+j9kCmFMEv2UzDwD+dFgegSil8CAoJ5aioB5y4+8thBE5NYgLo7C9MKUEEnvvxsdTmxC9s0ipm5
JmT3KHKpCfmphQNozUFpDUsLU3aaBeFj7gCV9ofkw/RyqtdbUrtmJKMzFfHTREH1Hkgzv0USna63
vlFnRVbEp/boleQbTP4EpNOxU4LimfB48dwdsNU/NhzjaOUMsxo5uceh8BRVXbpn48vJmXiif0NF
khZwaukz1uewfD8oJbBrNi8hT3GZWac1U6/ShqSLvGdXNBo9wVa+oQq//7lI2/DSlKeRjlS03XJE
YSUdmoKrwU9psuMKhX8/YgvswjFt3iRAMw/nZC6msT9Ip+tv7vnSA+c6e+dRT1KrcpFvtq1Rnq29
HNF6Uf4DF/ZDvp/Pake3/MhAYpKI0ABSu7WJg37A8Wh9U/fLj1yyGR0PEGpbcodm1lAZf7UQHVvM
lIvC2LIh56i+XpUhif0L4umJ4bCptCacAc/HrNDHhvJQ2OzTsQrH6qM0+Rdt3TKpnmtU7AMzdtge
QmV33CCAxBVoYRJtTpb9tIuKWYepFAGGyDGJ+4L46W86n7f+X2Dk3Rq4fwWu+IVKGGJ0VhgzDILc
TxT8hyRGVRHLkMoul0SnUq1WNPeyb1P9VqKftHOmRPgp6j2WdP2wajpytfN60HyrKhksOdPmuqVN
Dt4m+Fdc3PA0pRHx4j34dDlGOj4/9mwufgtBQ2wY3zI6g1jRotnQQFUEyO8HSb+6uw1bcvs5NW+S
8KOFJZVMOO38JO0BE5UkfMAY6HR7gZYywh9HyvMWOH2NyvExDzjELu4Y0OoRTMB340Ne2Ob27ghK
TSgT2IhUCaD73Fiqg/0O/PUrQO+dADb6ufSt6a87NhNDhUmWT229FMz+ucAU6fV2yjpqRTTE2DdV
J536YHDDV8WOUuYZPnVLaCryNqlVHRyAqyqhPquu/UvHeMXO6P9oLza6GiKg9ollPwjv05fY8CXL
nzWMHJuVI1/fOd6VaJgQrCITHT0tUiC4mvQdho8WOEcsOIMaBsbZ8epJpY5xWCZm2r3fcejps6Q+
MJ1rdnEtxgEB+DabxlPYhb7T9W9mBeGMLMH0alY5R6uqYRabOA75B1TECuUrajVmVudWeXwm9RDo
mu+ZbP6yaFa9ZaFVhMcaRQgnZPgiV6qRJO9lE1klgQhJs9HjGbSSOEpM5lfJ5sskvEXYOyfDQrAk
gBv7IyD0kys6Vca4pX8m9ozMDNuLuoWQAIetNE6JJnHJO/Bo7Hl7vJGh2fDdDfE8ojp7uL/diE2Y
E0lzub013kuNNfafDZQEyRp2I4t7qQIWNbqJ8xzpBi18zDs7qKDV4WQqVY9e17rcGjhNrz5e40yf
xhgxnHKyDo6Yi5Y59cQal6jpI/iex/COdrTIeFUJro8436CW9FTifKlj48vdZopbBCqep269yYcA
RqZyYd5BQj18NShXr2ISvzEt8kYDEZl6dywmT8qoNw+url9eWf3UfFEqqLeWY5x/2u+9UYBqy+Qy
g01/Is5klQusS5RtkwhgenJK6NCh45nVz45j9ObvC5boy/0io/eYO3nHBqCbNm3NMmo4NB3QdbQ5
ivBh89OHO4BjVcLb6EpATibHK0msqCY3S9yGzCdQg3JEEgddleZ3UHkfTdVJrUdG1KY/QcHMc0nw
JUInMEHq1VXYqTyrYSCtYCLtvJXK0262Dl/Z120yCLvohi1y4rqeuO8+w7LNjXAE3UdY6FaRbtEb
yhZEdr1Inc2YVwowGjHcmYFPwPdn/xXxxNS+OzA8wuiFP5C4qYyOuSoXFcCj3276eJXTlkZt+ihO
GxKzE78JhwOvMWbi2R5sFojC9SCx9vws1THwSXWpyxNLzggA0r5nHeyOCI7uj2NrsP5b9tkJJ08N
QrBUaqHKuRspgWcmxsQqSsWHu7GhNcrruKtZComUGmaHJHcZfK6yV6uSEM6VYW0sn1UJRBwWVfmH
QM9nifr47HzA3V2uoPPFrAC/ASaTTvfx7FTAq+PFB7jzTGLw3MA/av7hNENrI0L+t57olilCGr2o
VaeQ0GTKVUzY1iQxnZK2Oqbic1g4lcpC/US5yY8TwNKRWZ7sGKlLjfdcnQ46dAd9q80+7M7TTHu3
TNsjVm62/z2r2vEGT/1MnFFtkuwCQzTMxducG83zObzSGifV35CN6wh3WllWrZHPdD4cy2sZxsuW
hR4LQurxmc61RB8k2zCnYlB6Wi5L+85HoGmBkRaG2yOb6JUKn12xaY8/9rwHpgQPvs6/cDGM+3WN
yh0yE7PG0eY17J/a0/ke7ybYd7cEaLuGslQCt7/WLx2jq8yOBuTx+eBK+xDwtF/1bRZHkLh7CsEE
oIuwJ7JLYb/CIlUH7CISfmseDyoy1BhC12IsVdIPNZrCgn9yiWkkmh7eAQSrmLQ41Hs13/xGcMnK
AiK/hhFOnfzhTj1SD+T6Zcoh4UGWFbisGVgUzewGtG9grQ12xIrtesJglOwGEseEmmHaSEo22Jg0
48CYrkKz0HKrmjorawqgQhLHzlqcxpcuvvi4YBQ+OtOyeKGD+TuKBmdXuNZ2ZKITaVQDA9Y/mzkN
WXU1ud8QOFyUFGrTpLAZx4nWpT/3JBrI0OxuOiVP4V74bE8AC+WmbbZUu90cYB89REDQB8bCX9ok
PNpXEqGIte5TeqyCRNlcXA1JBBjJ9eFeG1HzUXP7MTrDVMtYy66Bi5ootvlRMo2w70+SAsNvaVgd
xf8+G7R2nQ/5kpYIsh0pklUFSGKy5O6Yyh4BQQ6fjCDoC0Y24TccFoEPSZpScB2Mg8NOoNWoe9kd
kD0O9jlEtZbnxZ44i5pPwFzp+/Y5Cw/vnj4zOcP9HqyEL++YWZJDvP+DX4FqySTQ2GVr+rqyAM2e
VRu+iGHjIfb7rhxn2woXHMlcmOkQkCnx8QR85IKGzrIgG8WPDT+Q5DI0oYREtp7auGVYZUt+Dene
DIYpaE+3QWXO9IzlLeY2Ljg7ojblYZIwgn5k1kkVwM97qRxXecIGrIRC768+0Ll9QyzGDeNxxHlY
+JGf7YCRuP9XxybGdsBmPOqbdmEONkZzKEiA0xLd12d/zuTIXjPTKMIGy3Et9r/6Y+rw6CJs+hJH
yl8rxgXug/dnvdyvuDug2FgI9VfRVgFe6S0uFxbqL+4ob6ShBgD3eP6Oicg+unJFzYcbS23RKCL4
RjDRetrd1LcR/ven54+2XM6I4FRrHy4kF0agECpAYjc/g9aOzCDnN8ZkHDUOWM+YYrag0VlZu/lQ
w1+pt1vagJ2oVRRbbvCEOT8HVu1gHM4nc69VzSBWU5Hdcz4YQXt35tSf7nxXeaTqmjLDRCtnCO8v
PnUCW9g+lD8Op0XYnavkE2n9VTljzwT920CedU24PA9S9ANC5DZ81yskyReQRKXaL3PF11GcDNqw
5Wn0chSBX4xiSFDLGtfnCdzquSyqdmP0XOvEb/rAOh/GPnyFylNCUWWxRYY+smefFHx7WfDL+Fk6
hgyKlVaSmdW+9of9qXuCMYr/Hqrv9+vbWArr/n6BK6ezaEY4aN6otP1Ih/79PbBDT7vVK6aTVPec
FZpscyZKwG8cb/zT1wRjuCgchX0MbvWoSdeOFdKxPZ9mSfYZJmgsho1oySH6vIxesl4rrMXNwZgB
U8A4U37xzm43Op8xVI0guRQ0va/2r/VFw/YBvtQDw4RuAyLw4lvjlz7qev+mRA8EcB7j8eRk7kje
32LDxispgrzXT632pNP4BN1elHb+5uNK/bXCeGqfy6wafWiPDMrbkFsiAYBEA9z+CDcj/7NFMXp3
NfXn4Q6blb3JgpREo7EmHQ9jPTvMUSzkBBjd1eeoCD6uqFT/G+3b+X9lZQRTLbb5+6ssjHVGBFna
MUWbYP/oXAk8ZRsyBejhB5YjXpPM7XPSNikuszomc/13pNyp4Ifyak/L9apxcOAtf4p+ujAbJbTy
+hnwEHbHLuUwjeDmZNl6gB0HVv5+SUb2XJ4HzuQRUkv8CNsMyKP5kBFwKdpAMkd6LFha1QuVTbBz
Plf28MzqKkr5OqnD5BreNg6VvEyy7De6ErQSBKY9CSwPE6Gf+QbLqLGDBB9ecjxfB/0dEimEcIIG
qzQiE+ITeiCOobZHcqHHUJVngYs+hwgXuBU+EDPvcHkBlp0Et2Q86ffFuNHXB+m/UWE4E64tIFgY
64iSp+OT0DmxLs8B9gdUKM3qY9+n/KpGVLSxbk73vk6fnI6wC54D/RUbeyPZ18Ep/ZvyG3uSTl98
Z0Np/N9LL8uv5NLur4gKmuEnZUWi3nXuOoKahREXP37CysoQgniMSRdjxyaSor3eVvgL3UyQxh2j
IfLUyyMq5uv7H9qviLqJqg5ZOSJsywigaIWU8Y964xNz9MXOvfqoHf6EnpD4FVkSJ/7s9vqe4BUz
6UgHVjq36Ib+O//qh/ZxL/Ks6ZapIsTmMjCN0HC67OGRd5rTOu9c1GGbmLqeLWSi0/rDv++pQi/Q
sXUOcoPlyJ5C3R5ZVLgdq+YMLjLJmnDcBB+wPVaVSkuzOq/nSp7cHZy25OlBfJS1ipONlFqQpxPQ
c7dZAUpUXPnUGd2IO+Wi5Qdl/+u+uwqcO0m8zT1N43JCFx1Ag0Z1kJKL5SleKpAsHe+wxN9Idi8Z
Hrzf6GYjUQQoQcETx3plAL3fkUtvi4Wp4MmSAbc1aN6rB8kdHp1TMCB3VSukOPzhlta33YBLVTiI
v0rAdWJhZ8tpLZfcm2hWZ0zAcdUojWwsxJ9mH5J3JmRnbikUYE3T33I4GCTLem5qgJCFiMMg9pTX
1LNk4TMrw8GWWXSlJcFguQ+6e3SRFd3MfVTiK80mVf7uAoPzyuDQ9zdLJR72X8iAGKpA4NbZLr4F
145KpKl+8Pfndz2PMpIVIKGQIZReWSbw4ZIEO6xQKA1KU7ZmI8eCsbh80cUZYJ8fWUU15g2VMrvh
3GeqKgk4UloUFv2ZUE665HE89UjO0WoTTArvvrgWR9D01LcOpnyBrY8bMEQzJxZ+q1M9/6TMUMLu
golXDTMxnIbeh2GC9RYrfqgffYELrKb+BYNiKQCYKUJK5L7QprkM8YK3CkDsFDPlaGX0Edgi5qCO
mkaQrajoBwEVzS6VAPIsBCE62f2su9MYM/1xH9IDTTxUD/t/Du8AX1fJDiiwa3hSqgdRj4k1yH3+
jO3TDdERMuImFSE/6VIWwNu5/WqFB4yjHXAu4/c+eAH7bmygu1RpGtgFEOro2OZ4/xAyoYQ/D6rN
6zrnt1MqjZa+FzUL4ccoGDDXeehvsIPrh1bsI9sOxVymoWcFfXek0cX9ixgh5rwHu0F0my2iehj0
qKNwQ1FIcZxwHeiVEupVTihtZfimT2fap5aE6kZbiW12aRM/fY2F0mkTxNL8ixpRWSN8oXfav0CI
KCTwNSM/tr5smnCZP75oSqlzTYiiKb7Pf4/FpNmbrwRCU7EEXjc97atZ4x3h0WGezBQm4Kkf5nf/
fYJHlWsXonWQdj3Q6aXDXTdkUnautsV7HJ/zwfF6PQEMgFebV8QFXwFp6cHrP1J8oN0/hRqE/f/z
wDJiAPAme1/XvOymIad6yH2XX7TiWoGIDune6v94xy/0pYTTALq2A+0Unykc7YhjdDXpuYkc7KU5
4JMw7uvr8EHJc4xYhAKOp0wRWhBoVpyp5qzZtRLrTK4ah42AAkeG6V4z8GqJTn8997VMDcJgDwM5
qgS/pE49SLwiv/StYwZm7f5FfWdE+CKxAOJ37N8FxKk2vEFAoJN50C0ybQnqjqPnF3g8rnIV3yyv
2qIRH/qd4uN2vqUloi+roDp1isT5i1SSg6EJoxqTun/QHx7hb/zm+H2wmoJZ+eSwiCXIRYIVW+kB
hJJdQaBBkUynEeJ6CpSluR5DHS13H50M1qAVd1WJROMX9HGhKagFcyyaBU3OQK0AWQyGnjcFpLqu
+eDraQbBaaygzQRI8MPTIYaJXa50pJnqz3QeSvvgaauoFiIyhsj7u6wOkBFGWDw0sDs+aX7bOAR3
Vss5PePY9Nn6OixWLBrH1lka91MGB7MR4/5S9Wsu8Mx3L2K8cgzwG1lxCn6ANPaC0riQGHou4aQs
bm6WFFUJanjp4KxkBmZ8bx3jL6RASz+LBMMjHwtXWPpjuAZog+fkqXhfLlpGEXC0VW9+UFKPdQ8e
JHMnMVfBlZ3GMHvQWIiwNWyX3wW9DmBpkF+N9wgvhTjmnxLNt7QazLkxTaPrtPwcZt8dk0QF7vx5
9fGgnPKEzgBCq/4omLK52YUgWa+Sw9Y4wTbHPASWZGq9/luimcH3ntNy/seHfRsxrPLmUHBGyUW1
qIJHyGn3gK4PsgoaVkVTanB2LRFpbO2994p3NFaivgz+5jWUSZpwqZ7oQ4zOLC8QZRl6TfKiJSgv
XXr6ibkP3rptLitsmkruR4rw9hY7mdB8JmWnqOjmkPoe/EkIGXxLlf3auL2LQp9mtm3GsC2Pgsp3
/OWbJeRL0Br7JBFkYrGClomoPH8wJYQlqrBZczbsSN1jCWU2spBsSL8DDtydHfvbDe9a91Vib6VK
VA/KBGvB/p2Gm/8cwpmMw+HFUd/cpRS0953BnjHJJPOa/9y8ISt7eBeaAGNkk8VT521J54POA6wG
OvJtKgPGLbUUuqVHyx/GXcxy0SKOilkZnslq+W7mdNTWI6SAYTk298MdNvuInbq/Kz0adRL/xNlT
KFKBKNujK5C3H/Pk4CR3OWxWGBh85YUPAXpVJGb+2iExA82IsQYNDgjWD14pEG5MyQ89FNcAuxk5
34/7AiaRr61P0lvgegGclx9oRim0GOrbGCTcYhzhx/DpNq3b992i5esJyXBXj3qAAJyec2JR2Uyc
zLUG70HGWwEYiS413ifguShrYISbV+Gu1sapQtr9vCe/aBejeC8o3BR2TxMEYPdcE2JX6QBEX0C/
A3ehJBelaFvoivdyGK0eEY7BwIdmX1tHjTufzNJW2L8TCge3vnSTfvuDC6Eb7lyvEzKEFu6dM7T0
OwZVd2jdSHJiOyoNks/UQoOd8JQQ0zYgMnkDjUTQDEWV09/zQVgIJNXwrbHClE3WwfpX8qN4YORL
8CSi9JY+Vad8IX0Bqgc7CN0ZnHAE5MEqdAwTgqiZqaJC0zD3qncvgK3y1BObnuQfM4xvmCNJExGD
mczbMFSdQLX0ZAjc2w6kPHFouFYEgEPWu0/oHID8f0lJsm2g93fNb1hJvCS9HWq4rCw6iAvuB+bU
wb0DxyngBYfOwMMXV8KBUxdv6nzpoYTMObwnimkJEdrNr1B20Ki+yuTtMQNimLmuDgjjWwUxEhh7
kx7WI9v7K+p0LCvuRrVpXU2IpDJmOtyCMDOc050kjKua13H718xc5eXJdSavmbheHutjJuGRXXv0
9OC6kcqP1uQavtDxJ7hNSN1M2oD/CgagqUW5FwoS0dw6i8J5pAZXoXFUbkfvr+98UNEkXsStSg7c
QLqXVq6P2eVQPS3KEacHCWCnvrf9fyMMRmVsNxaRZflnDZ5Vj+4+Z0oPTbBwoL7zYs7FAo+cYMvV
YQgcErGTeAOFtvdBrgn/Bhe8smAd8nJCpURk58FEzQvImw/yVoeaa4SWsNkKBt9qnDvMTiBYK207
DLAYk8yjPC2SmQd0wHflzsMK/ORJ9L7fcYKr2YMIWSNiMWG6VkugAB+tGm//XEwm+6DnFCtAtqas
mZ5YwkeTMgiOsf+4O3Q+CTWY0l+vJDMCWhZZIY/HWhS2fBjY/0xUv4PaPycVabvs3FJ6paWj2Jpc
mT4fkcp1q223hHwg05xWVZl84+jEvYwQ2DijYp71BL27PozyLnpVxCrfqoVezq1o+J+0xX/CEOrG
McE9iX6bJa+02a7lv+ily87PPVNxKbc6WLBY4wWOBDXjFjUppXX81DWAak4EybDqnbY42NdECBBZ
KTClYdrB4BayZqdMAxamVVPKCdJGXE1PeVPnhcTno2T7hiYg9qtxllo44fUetkpBOctgbHU6A0cD
wtpkM1KGBKSY+UxbqZ/pMotIDCYVz9mt2xhXyLw/Wbr9tKnRML1+hdEqK06gtncI04rFNQ4CkyCe
rCSAKlfgYvCCvGMPPsardooX1P75BPWAg5k8vfTAvEw/wjFvsi2+Tar6E74iEZv56fcwgp4K5vKM
wUbLu0txJTryflS/HvfhZRUFb3pD5evS3Zo2+NyggyGELV4dg5j1pD7VToO86fEPIfRIJXP58QJf
z/JdZXBSy0eqK5zmwUJ6XbwrcF7fHmPidCQDjRWnrk4SS/qwEXCXcVxv7455l/1UA2YKKYjgnXb9
y9W4hhGWJtPSiHo6OYfd2ACPosLf+3NM9rnFyzJT3NDqZR7ik3IeX3nW2lVIEjajpWeFLx4xPmOF
DK48cDXi0nYD+6ZSbTQZalm52Yrv13+kcnLmtORfJs95siUiqqBAvmJtf/X5hUyFnldC3ywUW+qp
RdfbXq6W9t9NIbnBZFgLxxQlg2KMCeSoMK9bCs+uVDZUCptjCTWOVHk16F/Wcovh82agJAgAduSa
+zCnpHoztiUVHbcwiE+dpCsfrPBQNCaHlRbFENmZPPDneIUE2CHQ2iMz1lvrxgEKutUTu+0G0xuJ
QfVcq2stIZNXfZFv+SimhMP4ZZrptLXtp3INEuU/VIkOHRoiYwNMTaI9KmY+SwNntkpPm1sYAnFL
Za97a+auW2TDxrvI72m0jLJfXGckn+z522VTL9gjr58QoQuSD2BYZdz7qJhaWSAvOvmb/mfkUpaf
dIgHn8QhD93S2WbIWsFRhPw3/IWAKrsVx2Wv6tPDVy8vVXoKr/prFfUGAB9To6coBOYra2KdQebI
r/HJZABp5+PTI6I8rXamH4iFuyi3EWyHDHD1VpPxRQeBYTGGeqyL9s0z5XbzNbiZklbBcV2E4clw
Jv8qdiXpynvnGoYkwlhkEOB13gO/yKQASYIUArPQ+bPtr+T8c2cFBWfasHuUN0/xitpCcMmN1l1X
nsMdGn+rkk3bh8fj20H+bpx4GyND92rRAjqqUdW9M0//oUfgTsB/03zjPAIuiSt3XzlNgf9KtO0z
fpVX/wfXHx2U11JuOs0XQmFtzuKza/5KbU8g+E9YpfCyInKFPi9+IyakQJRcWkTcCihOz7qPT9pl
HUq0+ybsE2JOEF8U6aWAigY73K7SmT+9/si7yW4B3wPF9MFHESqH6PTUZY7ZkgHBmRpnu6JKrOmO
wYaEpS+C1owmlW0UiyN4/pnrZ8Wm3Uk3ylOmTHlpEz44SLBGFflT4P317RFa/8yjBIUWnUb0pWxC
jOULKp18OAo6mqY213r9DfOJigtu84Ja5OalV+l0OJzBspyejjdfARTBpN/evOxWda6jpqCdfE35
qfA8a8LwqWU2ZStKzTPf8tGtM0zhv81OQZXZDCMLKvt9g+a3eePY7SFJG93O1jpXFWnFqwN8Qq8S
WUYNxqy+3lVz4nJWuw7qbQheRhqBGxc8RE65/yR/ciEf7Ic/tM2Uc2xVtgwsQ2LK5/2YVU35cHuu
z8EPjKfW46mFe2MTnR6OMLTaUJEZV5/NSv7m24V72L+JtSrFSYqwbhaES0ToCIGPuu7S4qxo2hHu
lacS361WcfjZGskOcSUL3xsTRNZAIXR21vhxpwAR/u4rUF2aEnFXILHDVq802ciZs6Lc9YYLYfvB
mJw3aKzLfhAupOrsl0iLSupqnVlyV0sRL/9SAVjB/hxc0wzz4CXXR+61oGlRd7tV3tSyZNPXG/1i
OLmqZyq2iDjkHEOmA00mV6ljp2Ifgp6701QoaonzoaFRXokgzHm03v1ufK9wrBgbKuMgxbnywK4I
NHo3Q0F2VDFD76klsNH1pDNqyKOxGvxV8TKJRkkHvwCJFz9mMVYqmgBP69MHstr1mcuOHakpQSxj
laNCcclqPEiOEHA7TMuChkZbNNsg/Gkjw2JvkHVap0bSv0webB96ZTVXQX7McLWtoHSW7UczbrS/
k5PUDgkWot9BWExOVrT4guuHa/SCvvpDNcYuU9KIFswba7vbNN8tb+rvVCVWOysl4lGIk9lEzbOU
avDrAhKfavkrGXF2YQI/H8I6AHx2JaUdTZVADOJvCBceLt45r4T6mqjW8L6Q8V14WcvojUyUbzdW
W6FvXZk2gpaLXfCj4tdB8REFY/NzoIMt/triRxNut1ruSYNlYTcK/bQbQPxAgIaF0qoQmq2QsPOD
+Gqguf3L6X57XMvxXoTVtx9AhPHehERybDLpLrvbdZ7EaMSwP4sbSLZ3kdpIiNldjmNenRmPsfiN
B6ppJtJauM3uauz/bZRoJJ1Dnae7hfisxJXZm2BlGXqu0R889nwakw/vaXtq03yGKJ88+BfzKBxv
cHQA/eGAsggbl722tvcncziso3U0qWe4bdih2apd9abOvzKNoK3ViWoxEZqiWKStWGAD9Jl4LFzr
lH8GvQ0vZGMT8wqYFBCiw49AlEw+dc5xXR3R9lWJ5JYhmZ/5Uscf/f/rW7dIUBRzXYD7y6Q/I35S
IwLWGR/WVjdqniUbxrpEY8OtyFFLAWwggP855iJSYbqTgXJ0JK5vpfROBQdAlh2L2MtwbKy/g3ad
kVvC2zrAXLsHkN1qvW8hzGyU50lnQ9qZy6djUXV30yyJHlP5+4XN0rrqPTnXESaQ+/Hb/KGS6HzJ
8JusE0QS7UmZYZzTL8qUm/MH+BTu/8JrrJ7vnpnEFwJqeZWaKSfdRnboEvG6kZxibtLkUX+iNsu7
jiyUpED8omyKWNLDqCGeEuWSjnXz8uuHuPvq0cDV1U6AP6hJ9NMc3hp/WlpGbTkUXjapLQSqj2Rz
tyFefWqOYjrJC/IZE2mTpV7ob5LePSHlCyaL11v3uUXJAn/x+5HIizHuoZhH3PVl6PG8rtjR0aD8
AVSMnquzu9tIkYwXEtsPkz/5hOC1KHmzbNw7InSQTV+iymVJiuAUThqxzAO+q2NyBqcA5nBjEukF
h5ZViCkxdpMMe1X420V4LFduoZ6uC0hDocm4+ZrCuI5g+AafD4/1Dp04jz3bcUhKw1u1GnBSqGwx
/yERzzkV188CgS9Nl8TPlbyKEBctiRX2fWzvS1xnwaXTiCdXHbC7iwI69MDXcgpaobVc4Ev0HoVw
ZG2upXeK3BMlFcKL2wqR26jw+/Xnm1zx7RtqtRuOQ1ENRm7dovsZhtfaD935KIyWuFyx5cleJ1PW
Fhns1Kqh+dJn+nP8ykkajJLgCvprsn+8FOl9rwc1Cx/zF49ptFt3KW8BeGHg7rLr4dT0/1NQM+tz
qzXyTY6vs1MHVL0R14kikYWm0rYS6UP2RXq2F3M2q7s+69mFQWcW7qdYmyeEoO01EH1yUwX7FwFc
KnwqKY0QH1GwnQKewG1dY+IXY3DZPt2EiK7D33OF9MTln4mTBSo9WeNBpYNrcrwtUK+r++EwNCZF
F7YGOs02H6dyH2hUq4cSMjSJpt3ccmCaPNy20nwH45eOdhXoAE5Wf50iafgkbrO9/SIoDgI2pqyM
tOczVg5n4M2REkkhDsP1h+VfqgZ7zIruQ2EH5wAK3oBlGZwKQTouwhYzEzMV925k6KUidEyF4lRc
AOtVVQ6h5rhi3X5irOPvHvhdgT36Qt9iURkNmeCOYUlSLsrHOjJpXvprRg7sGfsSBttjmwR8eyzF
66gDw/i2uuBJ72+jUfPNe/vAJtORY79P1kxpNBvrvJU/JnwGOJQYn3pCDKZ+CBSZfk0CgHAIRwOi
gk07Vwq0R6xM4kgnHh63562wGNgbWdHHbn9aeevrVOrVGJmy1IXRhfykvbPjGwc2NV7vcRSo2HhS
V1XJptHpQayI7Wz5aULCShTARejCGGyKmLdwk2BomfUYxS8BfN6eWPPUdq5atpGWbt4Tr9K2OX51
Q/52QIJyd4/S4E6GyrrzKa8J9Fd3W7ivlcuO2c7Oeqpd2Vy5etK+G+tn+v5r91m8QhpVSLpmPXEu
UkgyXrIzEf2syv07Cgsc9FR0wshf/BR5AZbeYeDFEWIChwz75X5nRVP8I2xibvlK8Q+xXQMuxOpp
1FvrzLNN//DoyGzH44QcsIQZsV8HTXog2lh8+J3IxTa6//jiMkeUbr+jDrUj+t8OlRidBjK8BUqq
5l0He4uGIYpr+RIeX1fWe7kJiL1NL4utRdV5ab55ZmFzE1R2Cck22UZUxDL+JlgpbkjJRh4vkz0v
cyobpO9HoU3QGvDhWl9cK93MZjYWmDc3MaPfOa44UOZclnURyXG1stbQ+6SEGWupVCuvzy3hmS5b
2eFI6koZiXF9Qg0VssknuP6QUWi9sjZCkDyBgMQzvn1E4Q7g9LwpvC7TzapOmCcEBhtLQ3fJhzJw
ixaqtQGCQaI+H9BrmjUub8k0aih196aE3Iqq11SwOEO9UOTUpdirIcXO14NprExQjMNo7TQ7s36y
fyf7FeUy3cupSuJDoUhqQdTsCYgY4OVUycZRGNX2R1KMI8yz78PdXGTffCG4t3V8ZpBlEXjBTSKt
jzaVFp5wW4bbvw49phBTMbtjErtqwYzcEBJOrtasB6BwDiJDseczc9/PFFLKYIxnoIChklw46EO1
5Q0WR6t6DpVw3H0lbgwlX8y3803iA/EGH7/NxE2hfT86WKMOAssajBdHUNESTKaIrI0riFalKePO
uMa3Dn/WHpq8wb4VGLxyThw8T3JsxJ4sDG+kduy9mIo5GGFkrEY857EcvgiXJM+9q/4jKNTp+jQX
4HGQhga8B9jPexo9ESn/fWfz+CalPD8YqZefe28ZZuqwXrhHefv8BDZUEjnZBpzMPrHY3DWTx6nz
2tU6V3MyvtKUhTnsJRF/afttfMUltI/XbvzkSyOrk9LB1DTGmmGAHihjGj3BsQ1LUD6SGshzFViD
uRFcSsFyAS2EDSQ/dT+uZNsD+3TNZWApxk5I8/Wxos5UoyfNG81z/WhR4VSugZYFjpqh7KCtA2Pg
yxLF4BqWRyaLVv+/Tl0UH+zgvsyN20MOIxa0D5hz3wAjwZ1Zwol0JkQj+fcgH/dYlqKSC5oX46ys
2flHm0V6D1nBcxR8bI6XuYK339DcoVllXjL8Ko/N+hcZgSuKLc1vtOCvn6wcq8LChYp/ZqIgBAfw
J0tH6ggdo1i43PrQ9kJUgaj31v1Pdjq/YbLwUviOzpbdC3j/3kFMd4kkqJ2G/Vgn6hM8xI+niYGF
Bspvu8bufy/06lASPXVUZ+hHFwkkjG0AphWpD5DQE3wsrjIWoF95PJnAQ3Q70l/jia+kpKguperY
ivtlYR+cxTVAXDriRrNKCb9xxLjkrEybI6vd14miTQBJA4H7ZpyeMpflATv0pZm46IFTliOVHg7V
a/95LnRyt61KPq7Bw2PBXtssfcwDuA6Kq+fepp+b6M9GjA19rim/OPwwsV+RTNjk7YRO9QyMG/Ue
SunL+a8fRaLEg9RoG/FTJ1Zj2UDlg/Fj5nS2r5mNEfr0P4n5FrRZi6yN/jKC4otvc3WnY6R1kTbO
H8sgB8eu7oWfbpN6P7RUIRCFJqL/x4vhkcbPT8mnKinDGbiB7+3X+P3qy2F97vI6xFILeWYbjYYe
+gWNxFDEn0M6qkDVggIuIZ/h+LctiUfDA4AiFAnJBStbIbXm282t9ZG6QiVrqwT3fnE08e9yqNDs
E2ksPyQtauFJhsw0bY8BkdY0lIhMblxO1lsG43XDbjOJUzoIKNSM9Vxn070CDA2h+VUvb1ynmn5L
Cwx9NnDqu+Pphml8hp25sy7tyY3Y0+r5D0LGGVnNLZ1L9yMcn55hPMTbN10yOxEqGC/Z1CN3ChGT
4ujqaWmjhURHixpTTgAMud9n3OIXmjLuZvTcyQjcsfxRgXUD1CjdBDpF1Wj2PQbr0TEFMsGMYlXr
VYR9hb6Ib3njbfKGRmnpWfSWsbrjHjwpL+AeXm41QgQ/MlPep+xrlJd7V49vn3yEoNIhAL1T3CK1
2LmJRqSlNsIOkICQr+LohrGE1eBibfb8iCWrqXM93cgSdgUnHWNYTlRefLZICk7tYJvrkE0tQX/O
Vj7kjlmsgwZl3S6hjx2kl8d5ge+wJ8+Wba6d8KO4uNKuzLPkzrwu0O62zH7L4rttTG7/fj1UPzM+
rRoWKPKFr6zRVEkUCgt33hXmHjcID9zr10DZ6VofLGOgKsRCUjkc2LF09/oIMPnsR6cJc4pxWBvO
DO9fQl7zymhyiLsdS7Cx9vOcr9+6/4i+ITsTYlEoYTs9UqKKUyEAhHENEYbbXyAH3v/2Y22lhEo1
XJGIf7mH1rooH10U4O5tGCmAqsoASoCsaSGuB0uk7s8M+n8s9omTjT1i7zlLcY/fyT54oR8jDxNR
T2jLZ8GqOHV6s5iqHo9afoVIv2RmaQWvMZJLGbUWelwkJSreP2ODure8DBN8NStgf5dyNKEaXhal
YkLjHW7Sylshw1NRRau0TRTlrCIDV+QNES3UVVINq/PLuyto3IZuWstycCWi+FdyjhN7fQZwR22W
Ky45krQG0ko1tjaGmA7zmfFKGp9gW0XPfKKtSlE39kW3ffU7VsQykCn0krio753jyvNzMciihroj
NRFQ8AihvHo983VETjPySqsXB4M1hCvFvwwU3u36Yl/mrdT6GUwqGGxrXAf6aiX8Nr0SD0LYyqpm
n+h/S0YNFBfGBJlZpYS4R8uBnsSUHEUSK1H/PTqvRu/h4i1lly6F2O9mPgVrARFYkoH6VSqdCKj0
xeDrUCgSWzWQEwLnqJP4gmQbO1uLmeOdr0Jg8FV2ppes9ddtOg8qR3/njAJXLh0CnS/f3Cu8u5Y7
TvPPHzdX58fb0B9Vnu76iy9LzTuSRyFiuezazSuU9VsCngZ4LYDt/Zi8ruuHamZBGLPd0mvelOhQ
h8EcSLUVCF4lNCh284StMFKaNS0TBS7sTVEXyMpoIZozrJaCuE9A2bWtfNSJT1cg9BG33j/nwsE7
yP7P5rUN63ELzZ7rZnY5pNQKLIi4wFFHSaV3px7zp40unDIulsMA5u3AiOoWWe0uQcLvXXU1lfBf
9dFuWvK8PDkx3m02ADM3PI3n7tGc41ayxQX3h1aaKWKO2DlG1QE4X7pmSNdYQua7Lws2VaMBKj7K
ajpCOlvJqAHqtw6VaJUAaFmPkv/tP/Q5Fa+Wpz2OiaYLUNLn2GgHmt7CTYIgjnftLp5TNZLqww2m
V9tLeNnfh/r3kyZekxF8LhYwrDNFUJBz67mivvZyGoFSIPCccY4ZHgJ6zyVPzG4wmNPFryKdPfmW
7E3OgGZGhuXkhZIYgEJBRrFzkWk8ABTSOHNDmJgnnkt28VZ0Pln+So/4jzeIzX73xCH/js5ZYKj0
ZBSqKrQ1+7poNBOtCG9mvfFaUQrBUhf7sk8Xp3Tp0awLy8HUt8owVSWu0P0YuMV1UhVROzQh435K
ARvMN3pnpvKaFUL8Bu0gEl0NGcbN/m7RJJeRcDHyEfSXU6bXTIPKyX0JqyU7mTyVhfzF3yYLY0g0
WAjO0/NnmxMMEYIfh4X6NipcddUXwgs8LCvjy8jArrZLI+BiyiTWFmyHqY+yaw94lE+fcwxTAuMc
Ybg8Jmc88aVWqSnaOmQam9pFn3XQ5GE4wX2wWTHRVtKkR/buZKNrVmBvm7Rhuh73Tw8Ph7ITUPgF
jiFW/OhSpvHrDrGPM6/4sBJ0XOtaOeqVoVPEXfzIsWFJVomM/VXcC67Dhv1i8fFnTZBc99VKT5MQ
8uqrVzNzAmk52fKsHKnvVT5oskUKoLvSc6ICcpI1kngPnqVCxw52881mL/XZpfRyOB/QVtKqEDkx
7WiJJ2zgpMoukmAAnEiT1p00yTBzIBOb1wQiGM9KnhN2Sy0WVzcfEgocfqXs5Pf/7NP3EMWLGXxz
kGoLE4dPkCb7srzACKOa6Xy2yqrgec3UXQa3EUvXh3ufT1g0VjcsJo+HUfpP2rCiqBbBgxhiohv/
wBe7PeOVFVuFeZBpknK1o8M3Ud5EcGVucT7xWscR3LMs6KIbGwMCvCAobYaZeXIZTFa8HCXh1kb/
EUKHHSbn9zcgJL5UAON1yIV3gpDvBlbp7byF4jpQnThWpIH/rBhC/L6sMg7FSBI5xu/O3HmD4pVg
0yJDHv0qHgSYQioALI0+QTfXRsU6yZJMV8YJpInb7D7Xd/z/ROYBx5agrEe1g2ZCB4dIP1NNxGVc
2mD2YF8NeSidt9L3EK2FD5LcBPUdit9yCI/eRYFAWmoHmnUyYYarfFVHUFr5VqxCG0gOyOEMujiM
2LS6Sc0R4oT6z52ocKQfRd8rcrPS6aFcXH7x5Qn8BuAudnzrurbOBqxg+UiWXm9Txpul7ZBK1S+z
xh/g2PC0BnUxjM9D6nLM5jQSAg/f0G6zaXd78/QI6PuX3st7pxn1PPGuQXkc1IlhyO40oHusdqT1
J5Lp+/W+nSPJxeYgSAhu0ThaAf+R+98/ov5+vagtphduil2qu4x159cP+oGsxpnZrwekK+BHSyg2
sWUL2P8KYzAHTmqwilmGEwNP9tB7Ar1lfAuPRp1wLfXscKX4oP0XtJlsnUGPKNoQ1os7LJ2hOAvc
4F52aM3cAboGiy/K/csshj3XqYonUCg1pkUlgzzBrCfeWjC7itjuCdN+fOy5KpErX5+inCRwyWRZ
419cQJjVyVQhM/NGQ3Dm6OlgL+WIxAGaAdYfvtSXcq3lK69cx6MnbzXB6U0WjCLFXqGlT/7k65sd
ieJpWimxcfFPKqZlGIK9bfKbB7fBlUUZD5c40djr3itN6ltti918d5JaCrZoBhTot/m+V0Fs2L8W
RF50HV5Y/ZBr3VyDbVWxCeTC5wCw2YvNhtX7iCobfALpxjSBf6PEt2aZpii6AJYCritNBizjwW++
pKriNzGDen9EoTg+qMtfZqiSBO1E5X3xIUE/E+1kyoikcF2c+/XAgKplmucExe3Kk9hnuk7XoMkp
JLXwe9jTa2F3L7DKjFWbORmV6F/tZQgUrPbuL925MOqftodpyC90aO+z1+TF9Nptcc4BVufKiGBz
ht5g5lfsSYUbgiqtGjJ5yE6uojZnLOQvtckcqiO4W5IGpXjDfwxkejuVjVjMClyNOUCbgNPMslKw
W6vjp5oToKZwyM0QwKlcylF3N0h5Z83s0g+SASXGId59taZf6/wsel6FrLF6aZLWS6iLF32qaZCF
rjQIZ8SOQzuC+zaM89/5njOx0U4671L8qFlC5xGanScu8pITyaxfj+3Bhpdgk0+bQGZFdj4I6czM
qOXyq6zFBiQGtkenSUuXdHmMHfDvo53LVYRWmsoBPm00yvs+yQyeqNpX1wu44HwdeWVveNi2DL+p
5nBxKm5Uf6L9r3PRA1T3SKAHPSC1X35kqYS/my4Y4iSQvkl3PJeAEzE9OEQOB2AU4yG6IMurjLgp
p+721F6uakm+fNF4RJ/k7V8tZZOHJhSQxpLpKHk8NNWCYB3cUZAd14S862jJJWhPbMu2ySekF9Vu
YN/2CSksJflUmKlbuL8MFhs2VjjpgNNAJkhtqV9W1IuByHlDfRhqecy6SSZYKrx87qTT7U42hsG/
uZbXn7seFBKIMINnOiMYm0O7E/ccIdrU7ee8S2kgV7FR6SRciO41DhIck6o3Px7c2xi9rSwKRpOk
1fWUhqwx+nqYrvDE+au8tAJeG4hKDd662YDvKJszZv4LDb90LI5if+/sWzWEQ1DXkh1N4FfxDyc8
tqPuamq/4EdM5kVZDbV3cjDdoA+AlvN3ia9IP9cjfIcaz7tHytGSqp7QyVAjP6n7/wkh6rJgSiNC
YyLiF720Kq8S/+PiSu8CE8wQDKA8kC6cZOTzc5FYqBqSDwTbrylWucAWvQbeunFZllUivon+AtXQ
CTlXnKwe7Mor3h9HtPlXDSUlTfqrhwfiQuSBLwq6r7fILhf98EoB1NgHMFgNJ/prg93/M2fwOn/Q
dyfJPJTnpmVL+78sbkMvf6syxGkM7s2LtbOMmig4qTY45TYW5gKrpuX9CG0dGom5cDnJFxB2RmLB
+37+IuIdNAY2+Cf83vpGYXinlBRvUxDa3Oup6PiijP4ikDlsqca29ziy9la01fP8p+1yn2E0wXCe
7dok57ZiTBzd6apEXgXdPA52qopBomPVekxG4TfI5BIzOevgElHNGjXShae3k/FmspySzrwZLJaI
X1HIWiqSHEh95AOuPAhZtVkHvilwYbL3diSlisql1D21jWl80FzMf5uhTQuiYLcqwoPOTVQbEJUy
cWc7dOpGYVjywmBP3ZoS5DR+Zg1SFmf7KfU4YSHba/en7bpeNou0yhdNRuM63EuHGbn5H8MecAmO
c+++q69NvtJR9qawR0q+cZVe9gngK2tM8onx4arylJIurnDlmdBUOtWbY0kCnRtWKWdXYRdXGWld
Y00VmHjcxODhM2Y8HJHBkC5Omepr4+QWQOR2a16HmXt/iqtOWHip6uWGdrjLMWXsVT6uUvV/7JDP
gJj9EsL9Kr4poJYKTQnnknv1Tyd0WflcGuAY+iK8fVJeyA1m3EeRtc67UQr4gcONFt65XwR0vlvT
+wkRFhghuIX6/7UI9uOoPnGPcFICsWgga529VBRynE7dY8B0oULlIDwFLzoGa2GBVWY6stJU8A5W
zo+RoxkJG8ffv9PINYJzkmMrlx+Cb+MgpymbwlFM/vaNh4W90lIbqKH1UV83sMK+B4JvJbim8Z+a
y8v44PrBMsNi+ckyEjIrpPdR1IcqGsFJNxCIzGqRjprcxkBjT140jpS8oE6nt60EQKu5GaTsOpvO
Yg97rKeG+WO74njVY+XX5mnOZFhkSBWmbsxV6SlGaO1GZA2Q3qRJxIMvF+oRWKO24YFkHeV65/Ka
SvzZHL4JRiRRc81Pyv3m5JGLzZw6Ig0aulOuOqg8yMnnF8mvFcoZhnkLUkCfpsD2ZSGET7NHFuqc
FTTdj1AxVPxRzptUObaBZJJq9V2/2Z9kuWaiv0UyLFbEUCzlX1UMGN4CI0qFBBsT+BEnGBUYthrK
MPTh0IDQ2eCDsVbqHysoZRxKEM3M4pJnijo0cXu8odUkvhpB+oBPgDjdzmj2lfToNjCmbffVH6rJ
0d8c8Cs2MqZ09tDTLn9DzUZJyKMwMwga47433Z/Qm5pOuGkQPb4Y9TrwWx4JtFVmViLYRr/gD8VJ
GewMYmENSkFCvi+DHCB2TgQMC3ZZdTEggRvVZsrmB5KKiXgWUbEF+8BzaT9pw/CId97Sj6CryOLd
mn/fL7SCQ7x/87CRH343IlEXWFSw4eyOlVBC+XU5qlwjGNqgLa71OZs9jUBTkCiXNzU6pECFBlXo
XuqAxAZ6paYubae88B6SmwiAEk4hpWMWZKWy5/dsUDihbW0IuRodaBaUEiPYwTUrc3VpJ73Z7XQP
FRTJIS500rKnP6skfXrWE0bgtqXfZYGD5wxuQ3BgFMDk9ylVNtJsqLBikVIHqtiOKgnfzaApYelF
S4ls2tTmqKowcI7K++OlaG/MThMojwaWkshbfqJtBzQbAFQkFJ6GMMjtMWU3u2sTyX4xBU7rRjxL
XL59+EjDZUozcCnplbDewdhoI1iHTgqa39289JMg0JchWipIVHk5PrGippMpswpiHdurfh4HWclM
M6qtzgnF/oS34xnem1NaEPM9QdkTWt3ezmSWdmdou7YBsHmJxNxFB7M05/lqTtfzexg+ouX+YdfC
6dHfVoX92PMoc8bqzJFb/MPr+i8qDdg6r0yQPNkffUEdl2yxP0tICFEOwgrStcoUWf7d5zgwYAWr
cQPS+5rTN+rkyNCn/UqNwhbQKV4lGuWCOcutelk3fRMItsijidbuKObYMVzU3R+qvZks8lb0kKsl
mfxMwqKjkxLEsUyOuIrYiUdagmBUBMMnfFslkrCw6+EvMEKMaR5a7cngV1NjKs6us6fSyDhwhWgi
0WcmCy5aR7o4dwZXc3WcQb3VZthSDpQzz6cabBY3AnerCUYp0rxxlUpiz5dXkM9FwsUs76elTjOS
5/h5hxsOMxtYiWP2I7Qr7PLrgMjluOeb+aW0cxOGqzuwTl/Iv+kjYR9uEasMhu9W94RdYYoR8cza
SgAcmw8Oz5aA1qU64e7GDLelps3+DKC+TG3NGr18eSwQ01dBUMXrtFZgsfxLDYP8gOXiCsvTtegD
n4JDOhNXokgj4hDLR2pqTvSXb1iOQe27BNhzCzn2kbzpuPKVcViB/hg9ZKrZ5eX7uxv+K4x7e5KQ
filYNt6H1Y16ZEcSrAi3mIxEdzWndAjaJxc0eEKHCOxiZZoAq8JcVkURLbY17FnW2i8mpXaTsJUN
DnzAXPmE6v+97OuGQBMEd/yjRfinxPmfpsvpeYUPjSakpQrUYrRWizKieJfA6KoA+0SGVk2ACeGQ
BA9DHix2LtRp8iAqEXa+VLBLiF0DbfbCoxWRYns9Md6sFOQ4BhIs0iUG9YcRGvOUH5XVPkNGT8dg
HsJ0fds/kvlqZWGRA0Jt45Lse2rOPZcs+/5WCLYhDrHUFgXYuHN5BgvBQkF3SyGtBZaKxSd6K1ma
PDNK1OjBB3YyZBoVJuLaJrU1HMyostPdUXSw8JDd8JYpzsbxQVeyjrMBGhbem9B9bwoEdoqtjpWC
RafXh9gUC3dVnIQ8bUiyjPd/qXBrlATLAMg0JtvXr4B+ZX00TH1tjPFJZLoVMWpud0AUs8pCZbEG
3ZTFiUvNIcoFYZtncy6/gHC5FZ56xjwyEAKErT2xC2KmbijTzULfdRu1cSo8h8u13FS7FSrPJwhH
hNS5vuMPqSu1S6SESa/qw7UIhUYyGOJ/sQH1e3gdfXxv6kklPIBvet9O/757WFphCNzmCiRzP3Jo
QvXiBzJRB9MowxlKi/XpYfIHmvST5vNow/rjpj1bK9xl5WBd8IAxntBhQoyrjBuKMp6RcLSSdDtE
KECCOrZSMCE5oTS0uPcdAQoxq5W1Q1hDW2s0PN937lkztCe2DyUiQ1dyzVsJjeHzxR/9dw9XF+56
gvSPLenfvVbaONRf686AtzaIvyzb/i0upIr0ElU+5S1E0i2axeIMYJyxVu0VvsNHK/gyH5XT9x82
JlljTOlNNxEXA2bVnYTde0dKXwdtQKkY2E/790nWNeTHmvYtCDP8YES4cCBrezUBXc4sUWwrx7VJ
r5ReDcENZfxmmCMyu4zuKv9QAACbCA+RIr68woXwzHdgRGUhOECL7SOUEWW2u0VWLHVaW9OX8ePB
qDYBraY5IfliJeSBpYcvGZcF7ONXXeUsHW/OQUAvLbcNHc0x69JyuAi1g69RrGhbGnqqTF/o7YGF
7MnwMg5eqhRk7nrEC4ag5eu392ZC1s3xMvk/BjDUk+KAStkliaoudGGmM4G9PK1NdXZOqf1+LNQm
QlOPPKEpN/VBbMATGKcVnR2veZOTxsCFp0IexrICu16hnxmYMhA93vf8C5M7v/Z6ThZJ5NGyQaes
yQS6U0hIFxQlNhhs4cHHIeju0D1nQR7Zg9d2xLoAO+0EXxr6H8zlrONKcV7aQJN9NcYfsWywOdSj
zgqEbFh0v6PlAIQ0YdHitt+9VQoy0qDZ8XtiNYSg9E2nK2CZaxjdZViyoHBBvx5S273PKBiyweQD
EuAk3CHltFZSQom6sx2qEN2H4RjdpjSV4gsQ8E3JBtGFlnAUOEpaL33/qc5n4A9jFhK7eNS49Axq
xHI6x3F82zFySbTHbsq4IhqTQmwhf8kOOzMBVIMfRyP/ALHzRxGkmlLimVsyin8eBGg3VVhoG4IG
jBAmjVuFE5nRpWLumSwwqVs/OrGeqeJnwpev7nkfCkGWlOT4JkeRWiI+iW7S1HRhIcotFrSc4o+3
HvBEdrHQlWK/mCJt/utJM1LiI8CT65QXGJPJlpGR6ML1xhYPhz1lJ83sSjyZgrX4NurUKGc/vd3U
uv3DROX3JAkEbgpcxaxk/PWg/Tcnfze7RLTf33Dzb/e/0hwdAOLIdlv51bYa+beDUxgI6llnXmX0
X0v7+WCz/gH/K5zvzOB6FcPsdB9QR9Yuf7Ha5ksPWy2EHNAaO0wc1ccNNu8Dl/u2tsU9hwyJMp2Y
bzkT0HGurqst+o4A6u+LyQL1oeswnvcgiF+HZ64M5z452sAOJzEEGHJ2HRqGmErwQ14o8FJQAixn
EbAkf1w+zb1AXqPQkFwN/AHKET+YE3Ffi3tn8Axq6lO7gGYZzQQkNTLb6Ic2NM4P/Jmw2AtWDBQo
mcu4lamkI4pobvCdKS/tK/UWUoKFX54mTpxvF6rGfb5SwY+uDKxwnm5aqPUh59JWIrUpRkzUmJK4
3Zqst+R55/3uS2gbbFVq329lfkqy01SdC0Uxh1S2tvSiMPZ3ngnnFmtCOVMmKT0CpxaIZQTHL2gE
BRJpXk74qvzs6T2iO8kpDV6OctqlrAhcguLReE+cnt2HVV6cF8nJvO/fTosD/IbFfHd5N9XZY89T
rOinKdmDbzM95uBSbNWw254My4WnztHPxfap4SO8uKw+I9pFdU5QhwGgSCXPkJfcxiWIXNSPECwy
GLLiCb6bK1+jaCtSozyZ92nz3K0HZA6z/0X77cGqHIk3BotYCz3khdTgX7JIIxSn+5O16oRNNgyn
4/dgX9De3eEUVrMvt88bkh70UwypenwJSW/PNv6YkabFjfFIKgLtCaC839sRWng4dzRVS9P4tlDz
H8B7wHl1tfHogIXfqE2H/GX0U2lUy654TOUYifbMI5OwVL+GcnguWe6PLFpcNsEzgzf3XFeCHZhK
rO1OnDW/zmXkGClXg/oDKk8Ow3IIvIEh1kwEtBB3bP31+N9+MZul2mX/f9P7fCy+ua5/fZ7X4AQN
KW6kNyKXmhPkAMveYkxnlm3L7Y8DD0i/CADwUDturJNYPIh/qSAqAQX8FZjR3y57xT8lTU2Ipc1s
nZy9kcZ/oHQlQKwIQqnEYiesb+NDK47RzAD5giNPWWxt52bho8SNQnGuba0dpj2/sZSFHE/dPwtR
sv5/vMnPb1XnPSiXPysq7M//3IoaBTfBajtqmarxnlGVLtiytmaOzq2jO0XkiauIX0ZkM7AwiknN
QjvCDUsreAZemh58aDeWjkwnWc3U9gpnDmZdCK/RCZEgFBAZA3KCcy72pCgFlnw8fOypOh2Ycokk
WtITUwNL/Zf1PoMM1EV+OE59FtTy/hkR45J6Qfl7ClpYrkolWqRjpjxXKE8TX+BLIiq9220TcPY9
dMPx2tM70viB5i91Up3lfMpRQxZNzDqId+6qJmWDmb5n2Ko4+g5fTZMtjF6CErp/nwBVt4NJHRkD
R8KdSYVb/33pFA379joEQ0P8paGhhULmVZcvGO9v1fPeDCdt+xGxKePCboi8jPO5OQBqq1jOkqgY
PVnt0AaSwL05McLmGavSY9AXbQI9R8Se2Jzn/RrX4xjGtIJ8WPq1pgSY+2GgZCc9tiLq5rgcz58y
lmmsQZo9IMiN8Q88yg3dF9ME92OfQcuAgWqn8zunZzoHEdqcuD3g+xeb4KeWG2wy9e8Z7F3H4ZVU
3feG3Hmio/+1YPkd2/leraVXKbCPzhLmUBSLR2oydXoA9lef8SXP3b3Axw6jG+UOWag+KfbxlL3+
Cx/PTQ9yZsxlh9U52DSk4MiDBxQh87fabnqtTJrAzmIOinc49VbTdm4yB78MWXHQG1FbJXhfdn2f
MdcL2xLmJoqhA0Fzu4Mv+Mbie8jhtwoC56lFYhYanoX4+8RQobwm43UmoXW8W/Mcx9UcFHTgg4Bm
L6ahFIjBoEFM3ktn4RGW6a4vQXZSuSQUdA4IrPVb/0hVlUCKnNw8Mc4u3//0iPC032JmSGPFNq8I
PUeyE4FtH2LnTsCAHH+k9Y8lYVPgFqoiWB6QdC4sAxI7VBC+kIQjPjXAB+3vFrF8DF0PDOWk6BU0
qG/77+wrKVJDaTt/Kvm2OMVLil6fAKyiAsz27i6rHzjRlrYT7TNop6ExZg1aiIuHQyr2SmuIdBza
IqJdlo8mM04HfYQ3agX+JEx0L1wqiaBqHPw2054B7brGdJNQMLqtp6VO0QFHYOXQo6sd0rnVBHsx
mDKS3kQn4GYiCFObYfZMyn6M1ArcrNFZsXmVA3oN0ZW49yHCZpSkA7TFyjkK4hQMl8UsnQsBnMXv
LcXLyhzmKm/lgRF/UgCo7IoHlFUWs20x4BBITJMBCO9bXdqvgZfvJ/AtxywfShO2fX738/UuyOXJ
JwjBj1fwcLmBzt3f2GfW/PTIOHCo558u6fwo3IypUeupOESODFmXtXaq4sm/00jk8u7T4Xw1X6pJ
UHebCqTg+GT+MDAEnJcpFsBnVK1zj6MrQdCCLcJ/eqSB2dPDrVUO3JvFOBEU1FxCBfFdCJtZk1ko
D3FEBIG5qgT1RcugzTOXJbqoQLXatjZ2lnzVkZuXZDmEMWE9eZ7TMOOimOrt+q1AStfeM035yB5u
CMDxB+o0Uo+HLcyLszYgWwndQcschZyzc7nl96ReRkdmVxwM0PpUaOe40f3ktQf3WPK6aI7bRuUC
WrUL1+RPLJoUbQJ/RjLIrM/2cNapHo6qlHf31y4v74QDvIIzbabA8sQLrHInYPOttC2yvkmn13bN
B44taspMq7Bk6xpUHtMtrrkkhk3N/EPoTZw9ZCvzd60P+vmXtmHoiZkoHz9aKrwM5h1GHZIdkc80
N1S+v7X1KVIWe3N+IhivqYWAOUj9vWwkgcpsW23tFIHCSbaJz/l5/pFczDuEi0h7+oA6p8Ekkakf
0PIrZqpkyWNoXGrJ51hfJfUOCxoG24lNwqbfhP/RGry5ez7dTo6wzY/BzEmZbeXbFHn+0dIV7Y26
XvwP4HhF9CfcZ6n54S+MkJ/sbVbYLup8rKFlRnmZY32YgPNB78jnAxKF3SXbhwjZhsQfI0W5d03F
VAVvqvM17cYJzyieptWMbL7KRhYS/J9RkzBcsGX/KT2BoVbfY0oL0ixL/FOS+kngZcj+0BjhU9IM
BV8+T6Y7sTe3wES3JDpg3o8qomxZeSu1MxbdFKwnn4I2926FAmfDgfugIJ1p+y2yfZPlUtZz83jy
IeoFYugW/DgHbzEEFcCL/zZj7rnYnPfKg7gJaO9MU6VY9tEss9wZ1SKu54XuWIKfF3LRtx74aLSK
TrbUrgts4fxC+CqWBVnt1KxLwMDdBy/8KV3uZ2tZTiAiP0X1NZUtDRTlweEJbKvRPf1LdQeHB+8c
DhEON7pqoDyRRfN2YlJ9cpCcYwbnXvVmBIPfjTYYlilg1fIQoklS5zwlJ8RkwOQcwBWWKSi4BpKV
XVHxMBK/mwZgM8Lz+UN3cbEzw3blixu9Gqc7Vq0Yd9nzVNe3khDD/Zun1ogbzOWuFaPVXzah9VpU
aSYN0s4UqpN6YCxR5FxWBrfXAcKUy2Mlvsn2IQwdF+eylBKsvxIyXap6TqUnBraAWPv5IFyuE9xO
fDMoZvUfazwQXLLztscfjPOJWXnxDBAIJLnx95QYSmgKvspqVYZ4SoNr9V68mw7mfbgk/3Y7/ic+
PcVVl3b6ovPBV1L/+L4I/YCjjF0+H14pPFeQrnG1Y6qpSnN9nv6Sj9HMrOTWJQDNz4POQIa6OqPC
jdlElK8WVRnriIXcQYfNwea+BhmInxI5yxwnwAn2cUW0E5stmib6qFMZV+38493qqRqZKsFnvR20
CLiDffmFc9RMxGuCQQlYfKPOxsvf7fR141yOop4Tl99mH0kN0jcmxgfQn43OttPXIWnKpv1Tbc1e
pgTGw+ICDHv60gA+3Yz3wrEPaadvyvyZPkLP/lWu8aCjVr2iZpTcOol7/QhILFdtsdvPZeP/ZuRt
YB+XGj0BBPeFPCBOvqJoLS2gvUtvwpLlnSd2JV8vgNq+utHZ82q+G5YJxDVqI7A1f5cBWIPLvuNa
TMbzM8p/tMkSaLEtmtg7Q/P08W5ee0ODVTBXiBKfgdWUyVJKLrbknyNpiKgQE8puiWY3e/BJL8I5
Z5/fE5mXHnSSmcPNI2L4TclASz9rIa7cwbd7CKj9b1bPeUC2l9+RkyhAALyvAxFWp182VGkluS+i
++Rmj1UBWmY7uGcTMn037JKgfoiNMhSWgUNPH9uvqw6Lib9mfKWsHd19akQQk3fa2Aw0jMOcMDbJ
l4B8qkRACHwrjelWF/+gRbl1Z4LdfN4zmB/3iiodkaybqfje0EeJMhK78DX0XOOSFzrFwiKJ6yXe
Bqu8V2Qre3iDtoYhT4CmM10xrHlcInInOaf47EeWi3egljihsqb+MerSFxVwDBWhC3C62FgNlfNC
kjlA9QAnNFDuKeaxwEkX7oQZMF4qNjKJ0sfFRgRU+a44+1r2PXO81kMnF50YYxuWDiJeI83JWOqf
Rb1aug8dKwlqGXwRUObrDoe2ZWrQtgliyWNhmNd0i9FE6VcyiBDObwsgEgVb36GeRpp+Ui7ahpR5
N4kz7anuHdPvKi40xH6DBXFA7Nx9TRoj3O1+wlrZg5eYglLUFJqTXos3JKcIgYc5mdv0jYz+fmyx
ezapZuBoGUSGebAZ3/Rs8PUvIVOaVN3eqglClmDucj15yG/5fbAaqf1LBTFTA3HZZk9TVuz9AEzK
O+0eEQPJVZeSZk/Y1StCukc+lm5Mie6oyZAA6H6gIJMY5uygRtV68P+gez5e1KYSKwwvblcELoqO
W15gd8pJrgHTJwnX3wRw5EMUz764k7zuq/rA4pXlOcSgqj31jfCZTzC8FXkgN9wb2KgdV7cmEj66
qa7CdIRl1FZXV9Ew2Zy5efwoguBRgu1PVtxvf/m1l94XEDcF7225ZoeIGtvcogLzLRoQ8ktS8puq
vYuLY2jhtn0eGSefC62euT08zU3FmS5hZYo/p5zRRHLqfn8xpwxDZzk0MP7pCqNZUBPxsh6/r0nk
r0wQis7AcZc6Q75yAx65dUcW+x37vZNvW9USfYvQNvZhLGOnAyptGzZbcPuM82tyeYR8zW0BRcaP
KlV814nIGPHWIomMxUoLxMHMkOupdqP1jc4DDZbkRa1k5dWIgQrPKDKrCvDzmyHzVDoMz8CaFVy+
mEQEqS3h+ntqFGqt8lLVGOUKNfwcQzrMbz1jN4++4ubNgZAxrodXCVHlihMwmNglLVsnGg5e5v10
E0Vyp1J497zrFU9c2WINtPPbezs8Z1Cn2ZrnybmS6A7D+HE0TQmx2rWQg5Th7ZLmzZxSCbuBNvAh
12PipsiZ4to9mEMDNb4IlaglqJfU5OxRn+ZP8iClWvQPPmld5ZWC8e6qByKqZpSFl/Z6uT3fTo7+
0w5dbMbF6X5p4lZj3ZtjCPifFkyjqDZLsH8wQ3NV16tLz1/n1LY1aSupsSxS8DOSVnSy/NYQoirF
DS0ew1cHRq0AZ4KaEaUpvwbfrnBSLrzysI+X0VFO+PZozyqHrCeR3OOFkTwD/D7Dy1aU/o+Ko3Wj
bK9uR2W3KdKMKxf6G2DqL30gPN4iHU6m3Khw3OocSVwgiAuXRJpjeVIstHlD/C7Fne5dyRHDX40w
r9ATStVBu8SFx3E/9zjV1ULTVjnCwtVC7fNaM4DGfqs5ZYKRhHE4Yna+1wlBCFrLEaDQifp9WoKU
fZqyppF44pwVGyD2quPcD8xMXvwlsUtZdbwuaLwAMZndLKhD+/LDYcUsG5xnpiqfcUmclahiu848
puBCimxrRCfRlhXuv1XlwctdUKj7KxbcSAWqq7Cf7z5Z+roOS7DkKTZcc2oIi7Uj9sTy3i38ReHS
TPoV+9gDpakAJngLMOHns4IIXkdeTq2YsMPV7SWKYZe9aptXe5mkPwJPQyK1ewsYTrBzj1HKw6Hm
XGS3JFMXWp8z8Zp/Kb+UllIl47cAuP30y7Vkzl9tSNaD+DG3JcL1LuNaUGPja8yALpmkYsTLpAOw
2Ra+QlKRNcR5bQ6aZzU+NVLuN5qJNQA4+vR77q+VnWJb0KRBNpQUj2cTOUryBZkYKdvhwpiNpIpe
4m0jsWWjnAYfUFyshWTj4euLwIEClRD1T9UOmkTSIb0jtzuSApZh/95vyvTKj+mJvrMq9nGyWzNW
gQRwWIucVsVO59xEqRPfpz3Rwb/9q6yOOAEW9f9gXqQ2lys0nF8WyK99uTg2wakP8pKP7vUIU4U5
bs4ax+qtfyCqmdZa7BPuWb9rpft7UlgLEdvhheaHoP5G9vCpd4RbIAN/yQds3FCKMr8fR7WHzo9u
DCOgR39/OvepN2eSCfzVomuVQf/nH4tcYk6APYOWvftsOXN/Zk1EG7K2DSpFGIJgoUOV5OMVz4Ri
fms1SxFeHFPrjL1m5mchNcsw7+KvZH9cpBJ5eyqCvVin82zm3/GDdAVl0hAoPS+QQohBGPuLl1uG
+AJ5X3zTZa53FOlv4grpDU+QffcErlrO/y7EHmK4LkUIUGjEXFSTPqqApnziMTqXf6vEqWxr0jVt
JoLsX3Eus+l5gBnjtDJ8x31T5CVNTgj8Ky1F7X7Mca8c1wgjvlIyuRuDm5lslk1Qs/xn5W0zCArf
As5wBggKPSyB9/9qXtHm20rv5pmM+V6JqAyM7YXJNSwd/O17BR4D29DaNIgiwAJnPaU1SBL30Gme
+1eAzPzaD6BwyWKTjXfG8jUHxjF2XoY04DkF5cf11wOHP8rbqb9EENTl1Tt/oMFSFru5EsGYZycH
eAa4kj2Wi084RQdQC/AAqLhF+UMrjpMbveFELOaQpRDLO8X3boJzExM7Ajeg1cUPoxxzpbRSo/ho
u8OfzwLXVZ4vskvBxsR2x1nx4N/+BI9W+0KK1nXMmcD+jNkQbqBb4buHPDhBb/NW82gDzMUH8mwI
nJh8/pXhylRFZqsJ7FILlw3z1LDJg01yHeFjJShGxoWbJshjFWrALxfPH89oM9rcYlCNwDM0hC2+
XA8bS02bwtojEVwpnS4UgnvVOtZcUEMO66WDGRg7HtAEa3M0iLsQUOjzl7GDrP9aTMIpPx/W2FeZ
NEoL2AcR7tWiXi5PC3/A1nZnUfUE25iVtW6iZ1GUsM7pO+7SlzFKiE2l87GcWCUJeKo6nb+zMvdJ
uM5eXX/TkYFSpsZJi+QW8pfLc2j3j8T68U4vKdFkhI4I5GdpNsdiCMwN5S6Xgbg4wa5pNAF5IH6e
gB+a1u086Tl/bmRnc2WlNQrKnKpyT7pU/ZGg1qiCuzGe0xW94o769Q5Vig+r37qKP/L2VxvyHXEk
BNNHFe3uTrfBfK7Ca6gOrDx8BSBkOXw0hhPPOetDWua16kWd1dI7AjRpyhf6+ZGtVqjn1htYeLrS
tFS0wX3LIOTZv+5vfFCkADZQCoV6bZ/6cjc8wHJqN2jMq+krewbc06R6DkhJ1WzDwvEviVsw3VSM
vAmX2ZRWihOkJFOITPnKIS0HWsu5AV/llEPApYXt4vkf0rdo8ZOub08rAhP3BzPi48ZxtRT8VMIG
hLJ2HnWKLD/ul37V0DkS7YKqMjyjDVmXI2//WGvvM5R83/+V2NkU23vNkVcV6lR5QGVxASApwOsa
V/iO08MKXpJtdOfru0AIZiU0EEhaSnoHmPChl7FUACMXwoM2WFVo/gNRF3IH9DjOn0X2L7a+lfNV
zVR6V5aSm9uZvjHdJaWMu3jSVpX0YkzPy5YYl3jVstjI4YPr67iaAy0QI+by/1fqem9hav+i1lOl
McAFpvg94aEeVCxNaAdJrlGovz7C43fJHdsfFQSfgO+MgpodXYYsobRwwvvDUI0FsFu5KUeNAEUv
Q+GDMeiblDw7FMm1O6y8gWjKPfbryGcqdL4vPvTrDdlYTzNND5p9h3GmxO5ZkFmbrEnvPW9mmYqD
nNxiU8pMSSn9nPW0/DA65twYaM5u6Ra32VBMyObCfpXI4BxcwKe/FZs2meEEYbc0zsKErgpWmRUL
ANgCZ0oqv5938qzcRG+N2W3OKqvN7ZEQfUZcDuJH6h8IWr62Me1+7dgNrGjoyQAUTvVvT4PgVZ29
Rz9rqMZWaRGm0mFzBmgDcX0IJfkPAP6q9LOXZBtQGUW+MU/TK1zMj1Evej352Bb+MYf9i1Y3LhA2
JbrCmf+LHyWs3CasTfjHU1LSGyrjdrWZ46sVRttL1EW8VKiXW3ly3ehjxO0dXj44LA77KP+qvwku
H9ywnTBJpsfU1sAON2lCCV/5FjP7lB0mBimIdhJDEvJCpJPbXY9mGNMUWrj6yXK3ERxLu3mJKTto
x/j3w7MoPZFtLs56sLLlqm3T+k9WLeoKaO7UnwSlsieSSWQFAZ8LQH3BRtcKGSnlc+/NYp5Y+PZt
N4OnbYL8LhnL9fzDwtGy3eg9OHFd0pcBSVWzgIRe5cXimpyZf+hSZiFu9diXf0R2GmwwZW+F0pWI
fr5B+fkNoIBkuPcoS8nDp2wDf3/oVaFFEUkMdSQl5ApuoGEPAek9Aimw5YRLu9wxZ7aK9G30UMRX
baWxzbT8enpdp/Dk42/pwZdw+lXXdM3uBhpIFRmDY8Wg69te6fFLIKCN30GqOeVS3g13Iiz7GiR+
3YELMag3kv9QZy6y7HPRWNX/rBTGsnhdK3xyBlFerFGaIWBB5j1FedamDENL5kyUo4Y4BTKoYxPt
H7LALYHfCSsVZOtw7jtRhZazlfsQr1/+Bo/xjuIg4cTulnAm8ZshoN//wN1XWqHeQ9ti2CGirmBx
f/Exjf1IfIbXR5RPQk3yTdNbYiwkrF8ccKDeFVhnULT9zARwrozO2Ax1l9OxKW8Q87wcggKGCdVg
5GnarQV31wJf3tW2+BtHf0hOjNT4iavi93z7iOuGohID7JH3eNw+KvbQJZGGPLWVhtyu2LBr1OTt
5b9SDUsAH+Hw8m1pBhNFoSD7p+b3TRDcgATO7Lxnno+FGrFL7PDWi1YU29Q467DadJKreOR5nVAf
+7Rqk0bdp/7TTVK3a2BHJ4+QPRgC9KD+VuY2pCgip6arj7fCIVrjT3l8wb5mLc+2cl/37lL1bMO9
A7rlGVO7M4ypdY2Ljklti/YX4v6i/B2HnFyaJTgO8JVYpDfvuYxBYwKWT8ZHkQMYQ+/Ar8E4vkjc
KhMYYwzTA7AvBhWNLTEyZEXsk+vIjm7qIteXPjzHWMySsXk/vyvLieJgcXduQCnmyV6EnDqFgCcw
TByAuTCIutaTc9zRxQWZY8LuFPrmT1/QwSBByaC6/iu8ioWYlm83uhdoO6XqxNM/tyVli17Sib2q
silKODhkJo1XKgkcSMPYgwlyr3IeiPCGBNGAHFr5nodCvTE2eXG8ah4Onkgq7OolrlxrYOBv3VLk
bOD2SSwhNSW4rwuawydeAufLf9k/vuc8WNwWK/7ijapsae5nWrwxbrC96MZos2p9FtcJ0WAiMjmt
D8FMtl598H7tLJ5OGzyWTHynxdMIHXCPQjcVlHxma3xHQIf3/KFGAWml+NyOv/Y6pRJGIdIssZYF
urbRTVML9JVZxjnNztXRjwcqt7rtgOrnSpcJkAgYqeZ6VjS/EFyvapldd1ka2zwCbGDnkeYi2O6q
kUhnO8EJuNkR9VqhrgiYXXth2Bv6Rdq1L9cTHbZOBAAxbBKvtBwtlwz9YRroN3W4TwltSJZHEPcq
q57nNNy4dHM1CQ1OHMHLnzOW9yWo+3v18PKoUHtrrh68z/dyvkGaMejWaaKcPOMIyeqskU2+EQmW
fZD3poCcYC39xHAp5Z+aS1Zd7tX6/zthkJ8aC2BPiz8KMrSBon5DKdc4j6YrmvQsaMmGluYrKqy2
e8T3F8DjVeU+b2JAIGhaMoHcbpWWxpSUPw/cx34vjnYRD8BKADjglUDWGn3PdZwFortVSjltHh7a
XeQjZJAVms4CBqe8HxWSVxGrtAC2jWlOR1MhGhfOCrppn3KyPBp94HFllAYkJE8vN1ksCIvSnJ8c
8aMFEkOEHCkP1QcLIpXTfm4yk035bH/347KfZ1tTltUZZ2rhaCPOLAlOO43OImZQbxfye2gsv8x5
nc/59A+PuKRr09EMFM+Lak66E9eOLeJod/nZQaa/dZ4fPfIpuJ0/6TrokABsslOSDilmpYDpYfqg
HYtgBzzykJyohRDRQd9/EbeaU/Gg8lr7lOL5ccaL+c24COracJHjdzeFzM0NM3YJd5/75Jz2TqiX
ALVcjfhuWLF5mkqCSijF8sI25cMRL/oYw+C+rcBeZOwG8U3Spht8kkbvPoE/Lkt84YPqJKM3C5R5
X+fhbg0S9MEqZ5jGdWtIa3Pa1Zja+Oh78codPdmoE4YIE6zpkeiK8TdqCmfcMEdAfOPI6xKMhr6A
h/ec5pTG7aSefH1yKC7vUr6+UbEMMIKzfo95tSnd1dWQR17hrjiEVsRqLK+vyxUsk6BRRM3l3FEV
kXJk9T5PnKKk4RJ9EdaFUSresNuz+O4O2J282GlD1iuoCzd9jhxLnXB1DOVjUjlvLQQuSiIUrzq+
lMD6zbVgXMp8VOitS+opWZ0Y0enhTbf63b7SI2CPdXlmolsOqxaxiZm6qsupcmGndCY0Z0vDDR8q
cKtWHkwBoJXGs8v+9blWb18Sq5wiFqbsWH4ManTGzN47+HnBzg1XSKItJFRLtn+nzN+i7pUMDJLW
kMGupQvDkgwF4ySCcpY0/depmXN5Q07Y6H9zqDKn+EjJBr9Z2H/DrsLa7YNdGS/w2pfYmOIGjsOM
DK08t2CGCrcQp7B61EEqLEASIXIFcCJjD5R+yPYrMqbSFEWlNyojzlAOtkF2p9fGBuqBTJZyr2kb
UtBCFH4qHWghAe1V6LI2Wd/fLtpAQKtEs62e5c0hDh7u/j8A7MZJgG1cEuGPR4sivDYQhX/SElDs
n0Nzt1ljyP4CBA+FUGIsymG4JglrgNWh7JWEutpZtHzD/J4BluIMnahVOF56Kinp8jCYKugYHIrM
ME+EqN7hJh4LeBSK9atd4iVNswfTzYqLPwm8t2cazy37a7fp3kxs5Wp4C66baK9/iWkxoNceSUhs
Jodv3OFQydDgkF0jl07UTm5DRH2wsrSSzNZo6tonUO9CnAATMAIFwylVdFRuWV/3ZKQBvOkn3nEG
aUAkzH4rR8/NM/HCGDLayhUWr+49Yh5GJBvtFXoKcUOyGlIG81SAkP6rfFqhVILijm51OIFTyGlN
63D7Z0KyKa/LN5CjA58fWdfceUy4CatcfbMnFtqBtgc8AURysAGwkwzjjKgvlp+ZrCiC984u21jB
OfYEHpwrKaxA5M3hgKFyLmZz7oih1mS5yMsE6pDhWFX9Vyf6PCWE2bLK44iaMXsv6zso+ZKM6f8i
6Yyz3E0x17lIamFnaOiJzD1Ok7Grm7a0/d8bLQJH8idREMffw8/bXvt+HDG2HD2rHH6jZ8yryI5t
LanVCCHb3/HAF3yHgzSkDM9Jg8JXTLyZxZ8CTI6p+Afln7Ri4vNpWru4j480mXLU8IYUTKIaAfNm
GTlrpuyUMh2D9CWwqAVZ64l5JzJz0rCnJ8ISkVo76xgH0YvQJ5sS7id49XAwaMiAcZZU/PL8ceUl
MBkr2x4HEttdUjwSulqr1qEjMiHjEx4Tn14aNIJxLUZefRTtMZJeGR5sx9UVeoSqQqO0UZozlD2B
CQUZlzITx31O35CmpBPdDGWaRBfCchfvSN06a1I/NAXfJzdaNb8E7FoQ/uOWWHegDhKsVRtHwoo/
N4kYpQFR/C0eLUkPKEnBk6/KxbFM98JJWv8ZTKtRRs3VGECfbLxUzqisb8mv0x+pgc/jZPZiBvts
Lk7z4mPsFmvL4ATnD7idno6W+a6YWg1NraL9FW42PMkQ0mPAFuVYqGLd+RFTiXr9utJP6icChMn5
eOcVXvz1U2CfqaQiMsvwkssiVKUNE58REh6WNYcBapwZKeWfk+I8sj9Ibl1spkntGKoZWaiPvcQA
qLVruBx0F7GwLCCsrfxspaYehOMQAlXYP6JtL432+S7Vudciu3XMW4Qb92Q3WfjrEcV5lInFd99T
8HerM72OW8GmFMG1sDD/GHBzWl1UqwIG/6Lm2w9aPheFy5VWoSsD3YPjWRli56pfZ8Dbtse1Km47
cn5uwNQ7jDgw23foAD4MlH12AZHG09kULZo1MRMQOpRI8OJladtCPQhCzPEEnCAgk8q95XCT7VoC
je87XQg4G7+2VqELwapSajihG5so7Yu3u+dQfRrGyKv8QlFnGxHiaxU5hou98Dd1Et9IRoRDijnd
1TGpZ8cRJr2S8VgQWtzraYsfJzxnzb3XZUui3ON8l8DSZPpgPA29f16WQSKM4KoNMiBXCggCvVdj
VWnNxxXOAhV1rl8yXU04ij+k257aoQj1p4/MBC0rGyCkBY3j2vy51kt6dTX8UHEln9F40WSpjf77
ZpFaPh66y/KhJB8sVZMVNuhv1YqL0Gl4pVBWhcQCvnKduh74cIevJbl6J7YEDxzUTmufYGD1NuqE
dKQS4dJCfxA1AvXp/58zz6e8SNd1wl58kHaKW+nmX05LN1e3XK4dX8om0es0Gy59oyQ3Tj9fq/Wg
2f3dEe/Znfuew59/sBgEusUk3NwYLoV66zROUYg4SmYOIG2Xcj8753E8sRnCCFf5xjQcYTImEV4D
ybhCuZMjtz9Rd7rB1ms/AQpf05qXRk50ShVh4yXStLmxCYaTlbNWInpZcS++qTAtvyFh08XNs4GK
UfTeJOsqsdNbVd053mLfn0+yXk39X6G6ApJFIo360uU/YVJ0ZhGsjF8VgaNuY5abitn6Tz0z25Jn
7RlQgVb1vGM2WT21yfXQYkOwGRdh+DYV1LS6Ggl6c4KPttG0IGZc5j0cthoaIvMonbjJotNyxDg8
kumtqfDPXfHj0w6M8y8apJdXzpiSFseoLmhcNmCmJ2rqu3HFDsTmlwQNh7uy0+BBdgMkmkaWproy
wz7Kl2rJiVQOrJQBnaUo355Vs60n8bRYXKfggkUAaxzHKFfyqMvVgObZi8w1IdZ/uzLvWqyKHgBw
tsocnF1xQXesqI6nYEceHxVWmVT9yCeqI9XdWgWIBuBTkr25pVBn3ffmXMgVlAD5MVnt5jnSC6dc
fVqCapQYjHWSgRdTeTHe3uv7zRvanzE1gEcLlTj+vnfc9LaVZzvRSVU2PoXm2PqqvjKdVko2vJ8B
1yLieZwHcCCwKEC+1b5b3ibrprWlxLCiYA4i1R0BI1/XNqi4gFL7xuVowf5SaU/LQZtR15p5Fo4y
M1yyQOezAU+hQdHTZrNvGm3ffPXPfy3+g5kAWjU5Xn125KdHlO2uBgypU7KzpeJ7ieLdo0Vjnyw0
yQNhokABR2TK5ZKiBgPLiF7SoxF/rouBZVkVP6BoWJ+eMiKwR64lhqEh4lYvE4cQTpL9oYARVpKS
8zNknYaYSZ8iZRTGnIAfmuHeQQoxRAJf9xWX5JnEDegv60l+Pjq0mW7ZYYpQiO4SyA7v0cQJgc+h
WtqRrj+eHYTf9XrRlOvy+AfrILfVZ0m8mlfoe4MiCL9KIMvBX+akW55VmEI8pXBrY6kS+9YdLqRn
rGexaYvuDa+5OocmLTfnGz5cOv55wKFARA/0Ns+/JvYuUjQUJ/nXeX0v5QlLrOb01AdSBqvYPBv+
kU72tS4ML41OTPeB45ToMiUnRaq85l/9lW3iMC7nL1DG2B9aIE1lZZaPAI9iYqqQqnu2LC3Um5rg
u+sNiAsKPi+ZsfV0wcSJrGUIk8WwQxnDSWF9vTrPCtVwYG2QTbp5QOQbJvtG38bvlMdlOnIC93zS
GqEDd+Nvd2egdvnL3g43fIMdwTsP3yAN5uCflQ1pSitDMolejAFEPd/Pt10UlVv1mwSzy165S9K9
zGIASE2wpXScBZ2LEO7WpRa39D5f11SD1nvv4ABVazJ98PsNC0bv5wCsTdyV6t++XUJWLxVrYpIG
OHrwqlvgYssxO2728D+tF7kiIdNuQ6n/MiXrFKYhKdYlxPfiJpULV8H7RBl3Ir3siUdsxPI+sPPA
zBYctRcgrxt6hlnb+ZKWy9sK0YECl7b/vhG86zlmwyxzMecfYYJkDQrgkr2P9Dci6tA4PAK4j5gX
Dg8n2dPcL7WWrsNZ7pFycw0IL0SBwd5NxcWuxR8HeuJ+K5pUAxyrErj08SHVGdKgTl1umrLlrfLp
pd35BdVdCDG107d8R/JYcCdoGkNnwTeCzbljsS8T3fMvK4A7Zk8fkdIrMeXffoQN6U8dKEoLsLly
eT7g0nxmvd4pMF4pz5NRrWEEMamcE8qgXvS+OF5KqgCe4F0K5j+a77WCKnjuVolki4E7YvrJbgsX
qTxB8JiyqOU/gUb49l2lzjwhtVh8o/PROZWhFv70M0VMglgP37ywuAeWw807kodFERN7mwdGbYBP
4Tvih1lw7WfcEYAZpyZzy5JVJkSFn8CPpa9uql2xEs2eUWgJUnMdLvE5tN/B2z1gcKAP5UG65f55
edXlU+b+5hTfmNPsocbPMhqYewFZlwNO240IkPmSC7Hs8c5LTCWlV29WmnU6SHceDb5zkLESEkm9
Qge+jrW6eDTR/JFew0c8it96TkWLqkv/McyLWB9LRsZKRV98qtpAu2yFT5pc8CtE6SYSFrOClf3i
9SWOcalaWYQtm3lOQmw7rx2QhqKRM1w5fKRps3KAmbdNKB6LIPWYg8Wbb9exWgumzVqof1JuRYGS
yum4kKL60Fe8OX86xyVRjpjrF8qrw2P6opcprBC6p4GAw4fny++tzBQGGo9U4h9qxUnSYeyRk86q
EbRiC+BgrpiLzQTg8QJ5SeRDko1wpnf/7Smgv718F/lTLByUMXQM0G8i15BVWbCoO6HPTNiRXwM1
uWj/9QlDOG6J23l5qWXIpeXD9ZaLwixA+HFNGlxY6W2aIwV0wVoHPTDFOCSQBpaiyQucVM6Gp1M7
y4xCN67u9pizx3QOeDaUL20ZbmkgPYoR6UAIu/aQfiAX+sRUxBYkV3+fkj2Piq/+Sb5sClcPo1Vn
Z2GXhc6CvyFEAgnjZvJoK6syyIqPa16u+MUdi5D0aaKOTKc/d+fDyf9e7R/IwuvD2UK7oGVBgBZx
yqszV33Auvp9M3i8DIbrK9gpwMjz7Lqf8hune7SbwLsqcBzXQDkIrt6xLpDZsjqAzomyxlH/wGF3
CVdcUpuN6VDqsoFAsiN+7k6hY1EUSyB0qd4MqQtLlBmCCpGDgnSRA3GJtTbZTipG70S7xUMA+/F5
qL3eY0TcWXM+M2PqCwPvbUPx+8yk85fETzetrckIh385p+DAK6HlJZBOTs6YtTh6hM9DJX9uTSEE
sOC0UgpOyxnmq/Mkmf/lzeXx8/RU9KFEm8jliVVLqEN94Tg6tm6mswsiPcO896Bc1m6/sY79CwEn
3I00KchAg+9AdFLE2DNw8PEVRxguhYzeC0WaszIPfRy55XaGLkDH9K4uNVOMY7KzHvmX/QkADdQe
OLQi8CNfSR5yExPJpZsjo3w8rC2YwMWkv0UziiG1nkvOobq/NBw3QI4z+cW+v/yP0Uc1NEX3DHOL
V+XoIvhI3QdGFR7P7Xc05AbaQ0QukolVCDmU8pxQaL/BBr0ulEHbg7ml7b7PsUYqaB7FEncRlmix
97cH1KQCWRf3aNrF1j2sve0hOVF7vdOED8ZGeIH35SBNgMyNYNucmjrovhl+Fe0HTbbGGeYIJfHV
6LWumKYudtz22FZlBuYGqPJUBQaixpt3m3CItuKNs7bmj+R9Qp81XQZXQRP5biefmbKMLxa6XrOQ
3sjVhXQBCs0qQsHJKyNPFg8W14uHO0cULJlMU5eU/EKXPiuucbFcgudyKEpIcwH/jvPwXHIlNwOR
0wK6gQhIGmixkE9U+Vtd4m0XCCtjNlpqgSiQ1DU0Yi+nQVmu5EPze4AzlGt41PWKWYFvyKqPWMVX
uGdY7MkwpzA11ThqaSgzVRdCRYxmi+/VJmcIdjpaJuyO7GyCVZ4YudAND3/bqdJw/7QP1wfTrSQc
TvQUsyUjsBKdVxAEQiejKjjEIRHhuCYmOQK8bxnWGILY3o+tni3H0g0tIJOK9IFtaGPuFaNLcB5Y
jfelmDaelNenJyC6O0sZQvURlVNslUGXOx8E3dgf6Em/SL7zBZx9wMwTBzucnFO841uJ3deq6PHK
fgZ1GgBbUlSfZdfwb99uxJcOE2xaX76yLJbodI1Cyw+anJyaAt5EuB+1t0v75vUNLYzVy135rjmV
yZwfkp56GThR7mnPJkTqNIIumDjxr2OpxK8ktQNKZ5XZdxG4T/jFZDmgGyKddRIeTCrifGWIa9bk
7fDEy14e664/FnS+5imDxIAHOYWCG9CRCNF4BF16VzS5J8JeTzxv1HrHUy4KD1A8uE12HwcUiH4L
LoRsVEgoxWlGNVjoDy1KcsYkJCTR2OVesij9C4JSMMWsIZAg34bjIRc6l+0nwHVUrWyP6m204bIE
9AzGRjlqawL3+gd1Kf3C7LMOThe/xOvmjsSydpW9GoxPCUpQhitOU10aqHrypQzG33W9qZ4Z+KU6
/wnw9gohZQMfUWV38pmC6jvDnwhiehbTryM751i0r8R92/Meyag+xii6RTnzI74ypbjzxhNvZY/T
YsFhf8WEP5IfIZYuxyQVNbSaT/H73Q92HRfTf7H1713piY2tFLv2CS0TedxeDDhsnYbhDTZ2Y8+z
/PDCBr+5bA+0s+XY4ZTtx5ZMLcs6ckiFfJebeCkwr76oA2JtzHoHXHvkLK/N8C4lhDYQQQkbaXof
5heO96deftd7Id51+3aA0uZtIpKbWu139hA1c2Hn3H/vz4wXSLq2/pjVOhYABJKFpp0pGtfHEOzP
qeZRLmQ2CqkOm5qgbrvZil0x1jD84x8RyNar0k1ddV4ZmSDQJy2HCfTs5ouseAAFZ5tl2VRh6DZM
9FDcqRV+swbCw856ENnaNGpvZGxkjK4ULeXm+iZf8343JJPJr+3ngPWDQfjKYpz9LNKePRp9xXrk
Vwt0BOLpFhWC8pukBb1UwWEmT+t14aaiRxgAw7pCMJeSqm+IEl7N1C+EJxSO/10aiAN4SzHmR3KG
ZVNJOIetExmINc+8g/T/lMyBFp5Le0E61MWFJ2OYfYbszVF9SEAS6ZxiayQReiZlLCrxdnN2v8/S
QS2MUdhSKF34ActbpRLc4ynH9ElHLcz39Jhn25nW+OHl3jJKOOj+bpjsBX6/gW0iF1fHoFg+SGPr
Y3FDS0I51xvfA2MVtQoadH5urkrPOojhk8JnzuZFZq6dcAGZsNmkRNvlVqny3yAU6iFEKqUaoGpG
eKkvgX6o6f6qAUUXxNHM99nLbA8WpAgDkEP8jGVQs1bsYvhG/0af9+x6at+jLP5xouaaGbdiCl7E
Eefd0/8TXMymyJJKTOex7An4giknt/rEMbqz7yID7HX/qphU2CwOsJlVgl4exmgfqiA6oScbJaZ3
y5q4ktHcuKHfDzpAqb3Di1vGGHJyA8eJ/rr7x7n5Ia6+mZ1ARb1dDuSwdCI4hQK4mUL68LxE1vOe
+NGEcG4HEN6hKnsVD5EvAdjy6PslldFMtTNX6mQ3zh4PsEcmjRNpetFa0VEJZtiKxHKn6XMSP/zN
tJcEGuCjw0lx/Z4zn0iTwDoGNCoJOI3tQ84yOaBXQaYvWsl4h463O1lMlOm/UcJSejdrAM1MvsKa
BunDe3+L+1h2Rp+bzPB1CVcfupj888r7EVi4frtAc39JN35ZEQhWopuYzWJ5tvk1iqSMH3MwPWGA
s1W3MYLXuohXGdTg2zH7ReWX1WydruM4ZRoLryxhRrK9OhsGETXvy+BxNAJd7ilV0TzCaUDtABLk
WaOoinjk7XP5RvTHUCmBRHK+TGQ9kkki9LytB4VuNRQID/c5F0hxo6L2YImLtu8cK8HjUgboRiSm
/8SgzYtMCEqDcYquPvZpmtG3rTh7HW1WWyfHzifZJ7hIHvm3bfq1Q5IE2VfyxRx9ScvmWaodASMK
XMcqlRpibCCEC2xN38UPSv7vAN34YxPE2UV0Ce4t9rch52XixqnyKxWovi+lZ82MQQyNk91gpkgt
nGImr+M08feBOur5osqm+66rpLVmrYhXHcGkW+bGEfzXcThN1aaV6mjCx/XsWuOb0iRsKYlQi611
5ug+sxZIQ0kGATjgSrnukWt0Y3dOgUZLrixbSyn0ZK5cWl33Wii7sT/HTIP/mcrffRGfY1pZrJF2
ASyZXR+oKDX+uyfgBAQNz4wI8j0TMb2gv/Qn/Yo81NnV/dH7/pEKb+ayUne1OOYVfDL8Oxtk9vSh
Gzs31NH6ylMYu7soYE9+HKQz7dLx7HxAOmKm0CIbfiU4Pg8cqTGQJazvcBXOgOvVQ2+a5iaG5Iw/
E3XOvZL9s7LJSjAFoKXsv+WmmNiWVjig1k708E7bOVi2dMyhENeffzTooROqIy8a4X/fyVtGKolP
XdIauCcOa+LGIL+kYpIFEe9klh1Y/e0DTmzsz1oSfMsCSejBGlDQiSgxIM8LYZl8rc/Sfdvk1Dzw
RntxJXJ9iZXUaux3f/jf04bg7pwaC+2VTrd6Me5GSc8ZU4FhvswYhbm1LwEs/KPXTAdZBijTzpjK
4/ME/lpDV89Ku2onqHZZoWYmgdLYe48D4gKR8/PKTR2ZfHnL0/iJPFkH7UxvtSNVJdnTrEbzu7QD
atCMwqvpiX7dx2mwGUAb7rSDpqDtWClpaIAMnLgkeDIcQuQhh78ZVkQWurKD9QqE65ndNAY+VAy0
2b47zEpMRB/rZqsvJqFb1mGzdULWvUNumJcbETTt+gUH2XgppgYwdduzIYz2aVn/ZwA7rm/yb4hg
/cN2zOQ1vOen++wh41KD2L9jiEZRWPxbKuqhfBBN5QOIf6iE4Dmp9UN6utPmjqPXWTsvfEapVxt0
cv0WweWUaZGbQ2r7eiKaD2vxZyb3Tm1Q0RkL8gB3bDs5A9BPGXWHjBY8KKP/sWS4yFPAyLuLdsru
1B7nqUhHX5l+r2z5X2jXGJN2BorwuKazGBUL10QUCDVwG52THSI5O7wlfU+KdG/bEfuLXTH+cFgs
tGdHbN/WTZpic31sQmdAeSU3DjJvKKhVb0G6xs1blCfAsRY/++PlKYg8Hy2iE7CGiRczJk8LirW4
3RloeW5QFs4VNX/U8hJzguN6Y6h4Oo1/MQi3CZ3QT6bdZRRXT10Dbp7wtk+W2jjTNk3CSaT0hS6k
L4LmMtVl4XF8gCAssvZRnsNGkl5Enm6Edu0t06WO9jCiICk7GOomkNu38YKSrDCKcakcV7tJrtz5
Dru2my128Gzv/9SN9gt+dkCKtopKlG0WHvduwRrexkOvFvAPEe+s7yA9TiPs7f/8HoeWuUzhflIy
xddpffFfnvF5T6fFMlfof3Ug6tt4u83v0Y4xac6MP36fVdCUHKhAfwcQytWQdiAPmb2XyRALV43W
T/yyMiPexyDDsiPBscCloMIPr/yqXGw4j2rQ6cGLt+K2EvAkNtzBj4vJ0MeT1ixgBfIShcDrdcTN
OQ8OXAg0D/9mmwMImOlykEGkTBOIIvtUXbRIuuLQ/idf7ivr6OYIpxpB5xpVT4x5VjS5jQ63aMr4
sTJDjQfLVCPXzoQEHjnnW3y3vImA79dWsm81U8wzxnX+z5QLFRz3TtmurFNjI+LqTuZnKjijQcQd
6X8wkNvb3fJUe/BN4V1zD7yEaV4dCjWq+9C8856BIvnGEBTusaKNiN+dDzVVP1kFomTUM7P2Ee81
Ibdt3t6gh2k7YaIBh2oobrO9bQvqforQn0xKPk5Q0q+gc+pvnilyQKYeLdshGsp5Bww36osdCD+X
ZS8Ef6SoyYLhhbyU2YHXqizqPgT/OKm2ijoK4MDMn+TTYhkVtUtuixhr0ixVikqN3gCBDhxpTfdK
/ZwLF0IQwGPtPoHfZTouUuB8bpgRz3C/fecSaVRrnS0EXyCfgHF3dvXaGwAVaEvPVWMDAuR56oYY
MdkWRpC18M95a9/3WSXKKPLGLtDvqQVwYzdOWTsSqWhtwGQqoE7ZEtylgqS/wBaDBlJMBL1WP8fH
GhGvcK0cTi/z4g5r7vAJPBqZcJam0QDC9i9tQMsyi4AnTj+ecCList0TN98bXmRbdqMkUVrgKe6f
rLmbjrJV3RzXP1OAw17e2HTbk/QAwHEANZ+MKMCngHvitIRCdAjK3NfDiw/VYXthWwPZy58I4U3r
6QqikE85hysWkTSA46lSQJtrmwRodoZgb3kWorsHjryNNQ12ezAEB1Csribm7M9g+wR/i9lSM3A4
y2dj/Ot1vfYVCAwxO3ZL5aPGUJUn1gmfUWiT1w09jm9MTf2Lb5WZaHEGRWFeKV+1VKGMZlYaCeLq
eyufTYqOLG/APYEqtmyfkJ6X7jvF5AiY3cevHnmUR+206ynxKrS26Xcjo9Al9XKHkCRnxlIKGcYH
zgBUVGffPq1zt/7/B8uXdEAN6qDPQjbyU29UONfYxgdAcseUiGcSQcrKgU+TnYgKsD3NRx6/57YJ
NgYU5T9j3qfsal3JSbG8MGL/gBB7fH4ZIP+pUNatL/QqNB7wiLIz4Z0jisdtLYNitZ+HE0d9qdYJ
L9sirSffGZS2c7L61XNQAD9v2unUMAaqrdwP3UtArl7gYVP96QUoS0X3wxhQCZzInXLHW55di+py
xxtWJfoWDYx7f7Aw/eyxzdGmvm8wB+nX+hzK302+U8+RTik4kaNoFwoK+SynXTXzV/OYo9yveXzg
NxtAgSBJwAaDOzquKkax6XOL3CErzv6NGwNevMzACmtvQkvAZRh2V+9rkvvpVlk0EzTkEbipgMKy
7+ITqiuVig1K5LiK5mvZiE5jgblHuWvcWUdUkWeLpSUb4u08NQkHKT3fsmK7Rz/x0E6sgYv19Uji
VmnH97/p9JUwf0Tbz9RGNOkp3bQPAVw30NibE21uJkAHmC+UpY8tiMA6z2t1WbBVaa01rQxqZl3M
HIo5yRlSpylBN0gegi+2H8Ni7Cy5aIEB/0hylyaUVHTqggdPYaakwc95Pp1x9t/8Zmkug+p5mN0a
/ufBP5JSOFzHtSKb/nS8oOoZnoBoMhiYyU0g823PRqK63q2oIiHuC5IeIbqJeNJjtHviGELbzPT5
UoiRHaguihiyTnNZDihNUjI/OAMSCp1G1F6NsiQTYlntzollTmFES4KrcOXnN44mImf+zwEzBRIO
SwgTqV+ang15GaSAwsFRGGzl4ef/VDPR9qL0sFJguCvH6KiNMjliXbpyzEj99qLPnOM5rZedZkHA
A9quucM4WUjJ0CvTmIJTin6pq8FYeg9UpeLZFQW/ArvCwEedw+5HUI+UHzKHIh+PmMqk7I2m2CWK
ZXkg6syiZv6uu1gqd0BY0BDE7fMMMrJkWmkQg/nm3UaZQyYgLO9YapG39O0m0ekmpfAYThCQkTzX
TYFuiP44GlvKcycIzNRqGGD3p0hny7YmR45fcc12mLLDdqB7OSUrZeqeut2MqLE7PYWq/zEZdDBw
T67KKlfPmVePTWRCQjnHbZNLlPA8SPwwZtzHk3lveDRLj5+bJH4O/7NXYC+7jtk2ZmP+ODavtOL8
qd/YuCu73JTRoRsMTjU7cqc04bs1CoNG6zO1QpywLgVl8AEUk7KUBJITTIoG2AERTiJNRVxJgF54
oOu/+RTp7qiJXP4WAImGnmSWhl7qmmweTxoM8LkoIPtI+FnNwERBBbrxo2TgElhyesbMw+T6JCvh
/RnVK7Alob6+Bfnw4N4r8/GjE9lfC0Qbl5gXS5tGZ8/qtLXEDWEmKNjajRHR75wZUcClTQFi65bA
yFdmSjuweXznaWYGit7QSgkxxY+6VL/6fg+StefT/RbUbx4RJReG4iLkejcDzRGKO3ZDkQPovgCy
n5OxqZCQ+MJFHTt/TmOL9I9lydfdomlstR9filf12lUBW112speCGeuAEr6uKrj8XiW+UOj3huy4
XKCfR8HjnC4a3/aIoub6qwUSCdqF/M0KnlXTRqGU7vuOgHousUpo1pMjFc2S129BlMUKD1S9DBsq
nD8e0I3TLYEFvVog9ZoHUr8hkta/owBzwBLM+3tscgkgogbE22VQBjM8Q7GmImf7HYgF37BsH8zn
88HTlEU3ctK2AgXOCVVzZ9SwRl5KBYTGEUVGesxC580O4IqSmP9JZVmW0AAtxkQcTNPvD2D6z2NL
1oygJuQO5rvyDRuNRVR8S7XyNk1cO7DAhuu15Ycv0uLyWq8VNUPq4tFTKfc2cTl2crjPdL+nyrLM
DBRFXHOwTboTfO8EpzHDOwPSteYVtYDGdE1857nUfcRfFtLFPXmTY+n1Qhc4CIRSDtpVCDY8BGEz
2Qc1/ASEkXgJpDABuiUT36Wlo7475BdEtb8gcVvGVvfghxU69bComjeUPgvLw49rFP16eAh6lPp4
zyZv9RthmN0P/rIY0ZVntbJYKIwzLr4/913rr8SkXOX4n33+tZNIyIDI4LSoUjNhgv4SyveMiXj6
BmZjow8bYvp5Ht/dCEIso9IEY+pNOxD74KSCXVYy7NcP1uALXi+rZiaDxU2ogeyZv6QrwBTFVytd
IgahHZsLJyxtrPekQrck+Yq5zXDRYP2yFUkMzrsLHLiGlHgF6Aythe7m1goZDDCYwWfJd7IzF1Xb
pnvWkPIe4oR14+q4YyW+lqiGY7W/cpRQ37SLSNsEvgV2V05bRSPu7dYS4GA3wTp2IKvFCoOAUInp
lNDOwU+XRS/PuPsdz8OIL+gefRFpyGuHQbOjDJ2/9p/H9VwqkuwsY5YW2FbAVjLBy3X3S6NIM913
N0b6itNBUvfCnhM3aGiuXihadHrPbdnyeZQrmdA/zH4AOTa31/dxKxI2B8bkkC6nCMbz94JoTdIn
fCsvR0LN8A3joBr+sK77/is2CZM+PH3v61MruRnc8XgFxAy0QOjbl2eQ4hXWZE1wizBxO5INrxHD
Pl1HSOtda1rG7wxIZBGkfa0lz5JcSy+p1Cn0YMPhIWWr1LSW0Lq0FVrbWy2NmqGu3ms5L6tD2n47
FRvA3Yytq/wiH6c/zHIiRXxxF6HdVOkbjYYJiudE+4LZEiRQRHzx75lF/R6Xc3T1e8GsPDMI9iU6
ArbL/E5zjAjDwt6rMAQ5ufHC3lrWN4XHGhLm2TlaiSoai/zauWlXcfqdiWr2W3L+elpP9OZh1rLD
LPXieHp1T/h7yDS5B/K/6rsRjqwIu9745tEB9diTdzR5rU66wKxADH3q3mdF59Q0OZmqYsEWwATE
RXZFHdIobzQp/CSSPQKivJ3DBFwVOQLsUtpgvtPaKs1gByAvczsoL/WBLDLL+qgN7fY23xFCKJzR
8I47L43m81wtrYtLePOmzJWwFkSwLxdLSH1VmjMOHIWmUOepV+Gm8m3JAfv3c0jkhnTXkmKg4HGL
wkp3Szz4KjzrOcwPgvfC8hVl9j4XWtgkjwT02BqfkgpKP7CJt5DpjyF4COp3uqUkpbHSQIWHpyEZ
WFL1teldBcYjvHPw5fkg7N3RITrH/sgd2sPT9k69Gz8+7Zs8CR3SEvaXq6oGGEIDyf9vtYGrvqf/
iHorEFtDd70Edu/+TTtVuYRn18zUBioeM2SKdtULnzQ8sxfz+74B7FiAms8UBMCP5/TKP7po38yk
DQATAkoQirsF5w9rPmaqu3qZ+0GCpyBdrLmQOYgZ9eTeyZRKRn4SfopQ0iOULMhsANSg2O7YNrOa
fh1tur5oaS1IPIkVhuMcFY8Rgsqn9DIncVBlhtysJHeoupxB/Zcogq7DaMFtXc8M7sgPOh3/ts8X
e/r5TFbVS30DYd0e6N5dFdCOZNGoNVjAIP7iKeTgenwm2/+C6dreLlfOi4vBvB5NGgsEezZzB+iN
qfesxIwRnYfBPh1RnnX78ozgxq9yBSJz1FHrBLMD7bzWN+2PDY4OA8WJVamUvKE+UyUw0VYW/L6d
JNSX7nC5NrwTiUaVGGro2JwkJtRvOdGI+a1timmVDWT6nQBg5wGdcArc108DnbDR36Oi1fO4M2Do
017GH+R5JD+DlR2x36EPD0ENg/Ji3oFbaSE8FBUc0HKNNloewJj6zQjJLsmPpu4dnkX0YrvESRb3
Y1BYJPsHuYgjCTANEIJzV/Pz9VO9rB+/cnroXePqZKczozLuAYaRt9CIENO6GtgbbxaJLuHDs7Ih
9EDFUrWyXsIdQmqDHJxD3CKQRlxAd2C6XXigWMmv4U+Q/eUGxb/NsJWsZyOV798UYPFuSmcD6XL4
PTWs/ViaEec4Ra8SmhDf5IKymhp6bY/G7/COjnOQuci3UuIeDOG6j2paxMpPSwYeCccdZnz1EZHw
b8zlT0RB4pr3bT4NdIQzHLF6SbLcMyXA4rP4XFuWs7XJQ4I3wYpWL0a2WE7DexbhIGgQ9zo8aGKB
uADM0xqJ5Akd4rYSXyFMpeO8XUoOzLN5Mj/udI0yLhw21jbsEBuCi00uFjmAwpudD44gDuBRUL68
VvLzI4vSYVGmco3qFiCS9sosud+0gin5p5U5fLHmy1Cw4vIJOjAdFbT/bUmL/ICjub5+ulQ196cm
3sNRJTvmFrOCAW4E42BgyabbujskmbZsDhVuod03eBcS77bP1LDdXEgQqGp5U1Kl7MXGKLSgLddA
TH83zB+fJcH3L5gkwkNtNguGLrOHaDqiHe1vOztXXUHItjQR4w4GOg3toDCVn91+9KxHU5Bb3QGi
ZZJt3Dmw0c+upgRLsMkpd0IaU1W3Q9kxyuJ/amXPIlUPJepqCzGG5STLuZvKb5IgpqXdQzxtvdHu
CPPSxGk60mxS+nBOIOzukfowkRwTF5k6UN6S7v8C5/EN5Px3Q2Oa+kTlhFBguB+I16ol4RR11GlW
1NaZqGKzaoaF2YvWbokTrpB5Ge/yiaNSAdC7vz1ULhZcQhczq2TpdxVKG8URTdzQRC+ItpnxKOKi
4tewcNcaKiEU2kqehzou7YAgcIDHQQrvgxOV0+QaztDl7aehFvcmGWur/pMKNLqfbDPCvVPWFEvS
9PMFqoQ5+Uk/VLAv1z1UNxbvoZnnpyzJvuSX/wqzLHe2ww7+rncX4fdYdQBwAHk2ZSuz54QQAZRk
4bNPBXxkqWKQBFMMsQ0sKVNhVL2sImpennYp8XmOshQfpFaoEqSoRsZhaDpSPDXrP0NJddNxwh7N
eTLYQFWWXnVI9t6Et0sLZlwpiGvCJIgIP45y/paO37QLssqNE1x8ajOdPwcY0jd8vYJKOAqnOnHI
fTTH/wPThRSUW6+xswmXu1tJuLSGTi4AVXJeQKb2ahla4YcgWg7EJA7DB8BFzDVkcmF1SeLfF6XA
oClPLN0zB0NG9aWrmmRhC4RKPImz3RXtMLm5DYFmAHDD9uBrROIxv3aiY8Ov8m9huGzi1KHQJKDe
Qd+7wiu9j67wjQtNdMMA6j8I/J1fD4bwHJ+kmex6rP7y21zZL0hKEPoYmUUsI/zeUW9yUsMetRXv
O74Xc0n5FCPkcRRXR/Q5veEflKntdNNteyAJBbZfve4oDHIwQTYiSqHoWujXHrlwiS4KIdmMj7KV
9Av+A9LZelpV2ZH/xwciJz3gbTCLZnU+ToSmrT4j8fT5jVdMlT3REiRsPC5wHoJW6uTasYMJC1yj
w/pXR7LbUsT4P6UikMZYWlP8Jh7Jy1apSdkAXVWfm/5VyHiq8SbaB4Jtnh6PBnBMMnYaJvWKE9Nf
1u9WtIAgZ6/LdGsGBEi4wRaw0DrrPH46YuG6Lh31cN7Y6Qx1AENBz7vF703oV7kFNEPve6H1OpOd
Xa5X57YLbRlin95B9XmtGxg31IsRtgGoXUlFeIcq4QTzofaY5okEYNzWlPST6WrVwskRvSiNM4Nx
gIHv7w5sgpGoTquAHVZzqP/cigtVPgUXCq7vUMSWJpXCfn6x1FBf6aTmUFg3NU01MMKGd8chjSt4
7xhE1hRtbpU0AiEzJ7ivaCkY8qpO48D0bUmgFZHvkn5sxJl2HGpvVqP66pvpCHfG+jN0gdKlTZCw
l7DWgD/pwKjXc/9PJK4aGFU6TrroH2MAII9IIh5cqYrvyxJOs1CUFn6ltSAf9FSOHLfgqXBoo/Aw
HR2NWkftGlBboM1zT/t4dzDaHwRFlN8BR5HzBcfSzX81X93LPZjoVboG4Erfsx9DDn7Lik/s9znU
k6EeHbDbFTfWSa96L981kky6s7139KiqrX+ELyG3WiJhkrCD1xrv21q7nTUyVNNlikt537CHlte7
hnuZc+xRFbcZR/iHjb7Qt6uReI179T1Ozwk80ZJWP1/bpDpY6uIKgavOm0yeNi/9ST/rXmf0Kq53
zTMkBK0JYPyjZZYUx2/kY9I+AkUkZnuZiCix//WxRJJrOBE73bi3nB027SnkoB/+fXFjKae6XKJB
BsTHIiCE7xMezFeWcT8w0Aot17QiiqAXIMaTbARmi425ZgHdFAFwhkpQAvpMT/HnTGDVCOHrawQD
eZsr4SWiGqKt2taIRhZPHZNc2PubnWw4oUPISy+UNeZeTZTLqhRhNoOaZZoQu6y+yg6OVW3BdIXx
y5JUX9zn8ZezAYl2NMsIBPMQRY5Mno7M89gpMSDIdtXtZN16Yl3Orm2e1tS486rugMmbCY+kFEEA
w+ft4yeUtrLoFKRfoV7aFzGREaY62P1dRI4YVleb7Y4NtKeD+whw2c2p0Npg7xhDOlj8qwHaJ8o6
g3U2H7+CL67QMDS7UMOxjO/1YskGfe5b1qpRTKBg3VbXzlM4Qzsf+fqA/ZPFQJqzty/i0KQUCAo6
0mppkbWBW9NHN6Wj9q5xHhSyb36cAD3nRhkqDa7uTXq8gtOTPuEl29t0HATVqAIT9UeIcHowZNpv
puaFawJBdOS75sFZWr2Jt0ezu9Qb9CRsRnSPFYo7RMQ4j0crjUqVYyhpM0eSpotHl5nJpfMC4kt/
BXUjGzugP5RprCJXVJ28dJvv7INpFtu3JjhvfdrZS9lITm4MhseAWlS4EfYHtBf2jaNSdnTO73ER
NNQmhBZkoBZ+PGyLsYqvcqvmabo7LcYEMqseKWYC7g1SboYUfLedxLih9KYgs+Jv7gmTAVAGXZBR
D8NPLg0tV28ZwKtx7jSkh+Gwfy5D5u5IBcsMO1qYchk2h7E5lvg61wjC48WeQV6HWkEjqpQ1sD9/
9bZa8wt3UFgfBKk06OCZUAwdDv4nhQVHA3le/3DmG1L+OTf78QssoEuZZVKyoepuDzV+5imqQkO7
A8Szg5gCVmVi5gGVzRW9l3wvvHgX4sur3SSrxSUopMw8Fc9VRoJCfQBE1jbt4DmbPW8pOiDBs+5k
FemwS23XLmSwFOxpH2gNhkoP7D9FS4ka7mX6xpWkaMuu8cZKVHzhqabT6tydUhTbVTTpypLVYI7a
nkm1hZvwgH64naScgcYUrH8YHa4NALAodO8p0iXAXekpEBL66t615prXI+LYCF1doTEBk417WAKh
P4/wa97F0m+irrZNgCPF1f338R0Bs/HSsCp4aVEtta1x67/Etf1z0LdgDFmO80T2Ky4VyI+2Lqyq
tMWSuw6Hgzo54aIzdBBcal9IB8jtPMx5KL3NgbE6+FuqOuRvct4fFzxwkA24XohxcWtry6YuuvW1
KMA32KZg0/zw6C90oVbdsJNKWKlz9rdhBSRaAmUqOIq+xiXPy15N0RkVuykpRqJlvSJDuBM+uYOc
HIKl7CGpjop1FiObPrt449cut9RWSoS5eYEI6MwAvRqCTYXlFJ/eblKKvFvyg4L1J/dYcSyAN3bo
/5EXV4Swb16mmALvlhKfwyaybLLHVAR2DGuGv7Mg/9ZNEjSQ7jHCMZXbbCvfBiLgNoXzzO7OrLDw
MSNabIBbB2Ji1YA7w/o8lJznT4V7XXUmhM2yXVvUloFx08KrTLtjg1HBVFUMbqTE8grOPCg1iARG
OWNje2o5aVyvNUCJRaTfngooybCcU4jTOKdJMVn2D5OurLsIDiOOeI69k+KT0G06asCHD9puFxPP
ZANyvofgoYj0bS/ZO36wBKuE0r3f9FpHuu4KaHAxni1y+iq4nsrYj/ZGoipCiLJlgQSfzQ4UfDen
/t6/2+/KMbLqZ67f8I7jFW36Gj8cV3M8Pkm3juhLKaUl3JQnLTdHRo5B3dps9XD+inHfeQO1QndR
xZ52IUFmjpRdGs9S64HzL4c+s30mKnN6ZEuPmCuMDfGQNoSxF3yvutqCVfLfu6C5spWOBIkgNcLf
D9gVcS0ekTGUmJqKu6R03iS2S8vFQv2RYDs93Fw9b7+tFP5TUhPBF2tOtUqSup74sFfqbzOYmPGH
gjL0p8u8gTPUMbrb3pYPeBPQKGKpl6HxbNfSEspaFKjNLoDa+6YT5L1wynPMItZVECETZR+LkG56
qxq1omKiCXraFJqpaeATrHTeWijcuoq4cbHWOGjgOG3/mjh3zJmBAC+rDBhaBjRgHoLEZPNywtw/
yHM+HwKyI6zTFA0CfFj+Qad7uNsn43pnAotLnzBUHfDEXHYPla2IJkAUG6zr8rzZ+B38Lap/8IXY
fNS+MLuMUaA1qg23GrZoOQ+9EuTRMRNgfNoAWyo1J+lf+N97T1gDqZE/hCp3XRgs159rbEYp7D0w
ecBMlYrflunXaLfXd2j+QPwqDVqfAaEyC18HGYPvNlvUU+DxN3X0Pgc4dr57+NKvEPbLMEPd6MBX
k7XrpohZ48klWmSpD+k6RfciOwokd8ySFWmq/6E0MldWcM2Tt/PcTCZog25dvP3Xs7Q8aMzOMtVn
AiE/WK0Osi/D86DcpyzPvdo4Zpre7UB466+VYaDVPKYKIA5pt9eom9DjEUHqBGY4kc/J5TD3R1a1
wmWoWRPubPOEPPkQTEIgANs2bMjETtok7iUz4fs3QO4bCEp1F/255Muk6RXtoP8Dp/aVhYQKaHQu
lzYii38a1WpWu7zDFb9wZLHvnD4XbTa07TUBCJoOfxpgDC4n0VgG4nMLaZrHntX/7mBL/IhTy22j
fwsgzSnMJnjFKdwLvPRKLW8sCQgmVinalEnZyApwRx1IzBvZXAWKyz3Bm7EP4XILqX1nxV5hRWjj
2IcEJToztWq4txZPpEMsP4GCflFn30jk4bsXcZ46QhqBmqRypuC16VLS2BUD+WBsoqeLv9+Ci44R
YxAz/+R4qxyTKlrYppowzGJO9H9pW6JuHO638Ph6tkb58rj/rRY0Rg+TyzZhzS1tZxg9hKoDErg3
XlWHc8a30Ok3PdS8SucA7c0nZlJeqYEfU+47NhvFBOSHwZKO+Ve+ktKIfqsJEsoLKLzQNW6JqE6C
N+w15kVM3Uph9QDHW2z39eJCt07DJBbTvdqXZFj6NVtHR6cStBZ4YTPdul3ehuZR5BgbXB2Q8fU9
FTGutHFFlvs7LYjM8SKyhvj4aWyylDNJ6SpKwT3js//ibqWV4kkdOjZG8QeRqiACbqKcbZb04wWC
1cuthdmG0l11UOsy8/ewpt2AeawlWC9OnQT+nkP1Y6RA/EVi20LMA2V58GbiVfcqt23n0gHpgeV8
mjynnMrvQrC8OXi4XxLgRuGc9c5EyeEIuaxoay90RJgmTpbmk+ehObpmSGmay1+EAor3iCPFuiXi
4GZqUZaKsgKsnshTlndYwfzkAdkoxv9npE/tg+2vTBtjIFImlPER2KCG3gTvvYOvRc9fu6bIh2mr
YlvYz4+DWDfgDD35CHJAYfoHCtwFBFAIbtfNfs+Z+Lo+Q4W5Gmckmbmh50PWNVGxaBKWYo/nSPyQ
E7RoV7FcrKuandvOkskkw+8a93gEVSH+nPut0AatGdd+BrReSQjcAgv6wzEu3Q2O+MRO9wD16FgK
XCAM/3hJ1XscyTUANc1bGs+g26C73zMqHuD0pp9sPfSW5BWjsu9woYkqroUYNSBZt+GVpS0T3a+m
ezaQ7tqClw/ZpOTMmBPMtbOU3hyAKSa5+YyJqJrAtxWY45W7jJs0sQGhkP8+z2gANnlAyDd64LIY
VQKNTsZl8y/vGLNVfcaoEt/Agdb8j9tL4c6QOU6RrxGwBwjlKTqNAyBX7U0G1+nJcUW8dabCoY4v
ao8D4EdDMIBz0OnDn1+5/C2HgulvAUDe664X9WQFOIcugHorsFIivhqKsSvHzRtwEHggNsdE5iBC
HyU5wqcLWnkXOuLWaxAZdeQL4ivjynvoqBRXqRpEZ9HifEEj4IjT/h9792HvYaV02UFTvOBpHkYq
PZRGzPqt2ktRhh7P72L2yqXHErdpKgogvuLYpbi1axxsXaQhOrrdXF/N58B0vEtDLlnJmoZkhngZ
Iub90VP9LX5CtFpkGHnX4UImSNLacy+XtkTSTbCBHSaoACxohBrIwJOyivxot0aJDzzohjrvn5jt
aUkdxjuVVJMqiLWIL1/h3FqGthtz7fUmFZEli6Ia9LX1NsAOOmco+KCtZMUwFAXTqT9t2gOKUNFO
LFxraywTC/H0NWnzap41CxZsASzNZYQ8uZfxxK+1hEf8U266NKlMZxhwTjeSQvLLskxWoYCk/Lgt
bBc42nZRa+k+KlH+TOSisD01DEHscnalxrdziCbONhua+pl4SH1ruSl8N4AkSTAEhI8Bdj7DmuhF
l99oCgD0z9UokQJqPI7rkd4qJR7WSEwtu9w02+QJRGYI8PGJFZy0qRrAQRjpjBzYv1CsZqdG1rOl
qyvcs+KoKjdN07uqKX9AOxdRXr3KsCTgXFtBX9ie2OwB/W64Q9ZuYB+P2gE98aIPNo4DmAGhaJhY
YZn8EI0r3NmYW7CmsadYuRCbvhJnNG/3M2QPxRTt2yladtuZPA/5IJaAwCyhuxHKa+jgzFNr5jd/
2ANKqc5coskBTuooRB/C7CblbOd1xLxitfM3VAG2MjnSDuRddXngcjl4fKiN7wvejl6hb9UEX7qi
CeOxTEZfcTwTQbUx44CG7TnHhm/zWRrDOqM8Pa0eQRv0bXGR8UqUjU3wjNe4WrmlfiWTcb/hJcvT
Y140NwO4Vi9ZUZplUWJExHohMnbIa3XgXMRe77aZWlRipCXG8gRAu//pFDhculE8L2xZYNU8Kq63
1mw5sAm8hcbfeDB+Hs5RgItT8vUijToUszch4Xd5Cufln83StjsbOD035mofN44g3ySEzAGj29k7
kUKaIaxiM6m4z1qkx6oDYZlX6qZI8oC3Yp2TrgEQjC4PMV+qMKR48sZPQ8CAsMR7iuc9OtKAG1XP
x78GD7if5BgiIdiexDfdyux/0xjZSZpY/mQ982MeWn8Ovxj9JsjslA5TH8ncHGANXJUZrrh4oki+
zD9OCENtsoHogdIULsowf9m7M4yWYzDgdLSTUNJu2cYVMY0vFAdH2QAFPUh+Qe0ybPyX4Xx5lbA1
s/S4SRa2oZZEDynnTLbHwtnfrdiX2r8IwQXJrxLMIKVuQ4aUg+x+7zOnx4IAbzEQyFDdgB2NR2P5
6EhxHg3clU0gxlvWfDTq7MPIaSVdFL0qn06r+4QR3IxPEbJTj9pimkKdlzqSWXJlCB6IGy23N+YJ
5DY5I2eNm1lkH4sivmriT63aEY6z85Hq8dnjwos7SVGshLiXKrbNX5clqFUX4CawjDZ42fJWXn5F
e37ErDKOPvRNdLfb1drfxonVIqZ/2pSZtQmEVfkrCNgpv2f6woo3AmrtxS90kzWqUyP0IfzFXtbw
tQEqFCBYUfM3jSWmMu5DzXcyxP06zgr/+R+G3hzxqoA1LU65q93ff9J2ECuLe1VvVjkCCP5ewC+V
SVDDRCo6631AhWlt/50JHKJIyN3R7wKEwwcN+U/KIYUK03oyHLalXcHraBZJ+Bhe33yL6yBUUVtE
5zGlhVe5AR663Xo7qsXCOtMk/x0qUJo8qvU3PuTrWZ6KBQkmMXT7EvK9tCLLMpMZALv/S9qmUPKT
5Dhm+p8FntA8xqu7UKtKOSh3RcoRE7gp+htR7LiQNj7KX9LxKbPOwmNVAsJ8DPkU5tZJf0e1VCTS
TEpkxmWKt2fml6Aq83/zhjH7FgvQGUZN7IphFt/2A3QoK3eVgIDNwk0TFI6vIXBoz7K4KL+j+IGg
t+JsavWUUFAj8jdTMznJpDvskW3sQubS7/po8oTCdsAPZvcGN3GRhzscVcokLRuGlCqL9t2UGrNl
O/sOi0wGtoEuFpOSYdmJPVqcvBZdLsGBPPtBnPf6J/r4ksaGjdBLUjsVZWvgy3fWWend5K5lqE6m
Mr81rCF9t0ipbpGEBFEmnnfawsyl5CkuVeE1GTNxl21q2AujjCgk8EOYxY92EMuu9zbOjICF6ce6
zm/jQeGtrliWqViiR1xcevQ8UOeu6WrEWv+mxdYotZiMCzxT2xr/myKsCFGAYuaeeVzvykH5G1vb
6h/VyRX8axMCb4vlODYcDVaqPLBG65tEvv2XhEAV+ysot5v1+3BcJpSS/vmarD24V+1r6B+/uFQl
bKiCkoMNgir1Q9V5CS8G+qG/dZx4pD/mBpKU5Yd1KRJcwSwWAujaeIFQwaF5S4kzBbkmT/HW5gLk
i7xpWVWkXXNI2+2db+IQJmvzYpITgS/V362A03BHx7aD8RpZc5EcUUewT9wz/UqFD8jmeecjF7pD
3p2i7oaDDBSsEBMGpfCK+5/e2qqZLsitCVzq+Q4a+kUkff7bYFbwgWkMCAY7hF6kilfpmPyBPW/S
pYPpZ4Mfb1G6WUYRRCSSGBiiF7/NtdQEB7j2mKtAE0ddknPgc4Qj95uZHmj8ppPNo6myitULSElQ
S6p2QI5LdZj8Gx5UvodeRFjA+Nhj/HdnSFf9jurdq3oyrz0ZXrZD7v/jXm0vIFkOR9XiPF5I5auL
0aNuEpbjm7ay9t3jnRud9JgkT+BdKfvltVxVj7kKNQNB+rpiwmfaYI5mbQ/VNjMEpytgXYnySG2s
hCLCp8hpqNvI+/agtut2Io5+QgqpqJ6p1g2wBTTRmiXdfiYmJLlVuytfXMl87sboLQbQpo48vqMp
WtkEzr6srHggxz4Gk05V8GIHTejKGRSRzzsU+M2R8CVkcArevVmcao24EclagoYcQKOg8gTzdAEK
Ay9iUsjUjITYHz8Hz0D1EnW4lPa5EH1/tOZgi7M0/RNH4KHFlnUTL5e5dCp4m0t/JVs6N4ao/KGn
YKNlHIOQ08o5ZJBP9eZwVoxpYjSeWkFNOH3wSUECcfxG39rUdEXKfEuH1wxcXtAVWx8gTfPDsje+
O3HnTlgUUL0DcQkpSXRual0IeC4XmG0egs3+BBeh1hZRpQ0vyD0jugfpgivCWBr/qn8Fsbf9u6qP
rZ8KioaTZRXn4x9xG4wJpOhq+Kx7Nl5N/2KzK7cTDmK59PKNOGnPeCF9P9Rn3zBag5LRw02CV4c8
jKQxJJCACDly+gNi0beFU1bUupc7A9hBZ4aWlC+uUKiBj/xV+uTEFd6+a3MKlo8xPTyZozusI0fV
8B4T0tH7Fl7P1BGcW4U+ICDrD7HqXRGB5kzev2mSd4wu3wZMYi+3TdAqhNbMvg0UbQbARn0S58gx
XyzpJpaX0NBpTx7G7gf1z/Ud2o1+y2Sn9zEqlNiTrOeHZNka7FiDJif7iuOBt7WjjfeQcN1V7/pO
DBumvHbUy/a0c3gT1u8eVyyS80d8dKozwC5Qizs8xfdX6/uIrGK0e2ewG7QkdG7Js8f+Ng2gXuDZ
QMfwjnJlJYdSEUGsX/hxhmGeCUF1hfDZ06sVlbAM3H9XE88dLH0lanbnAMgIBTRmZ1o7AhPM/QGc
xqI//i8CqfpTgWrTqq/ehzlCyikpxi7lHFXrogmJFu+Z/+Ac0LUPZcmZ7zg20z/jtbKBn4oT4K48
CI41wkkp4K5LoTlqIneydWXrpivbWD+kEeeB4tP3o8Cz/b7Yjdc7SdaSzxkKKN8pFd3Nc3XJSljQ
MJ5rCW99GAb7mTkUXBw5gaKXQvhb0/2mkGKTtFRM4gBo1CWKbK2TG4HlAe0LwCTZJa3x+H6fY/Yz
rddWht2fsxu1uua8DQ3BayjaKJtH0hQcmSK6HV2RB1XH9TwCriCourfEnd3Cd6s7eEW0ByEq93jE
fxaKgI8bGQJuXBBM/inwzgxCrYad6NmpnLTK2pxJXlkmmoQ3HgFxfAmsqXpVygJgH5LwyH79q5fH
GYiHGBCNQbnz2IOcVUhmPwSR85y+jEekLBiHonZCu9wx111wTxCKjKa2hW8t09Er0jPuOm+OO3hM
pbcvFiRdsAysU5TezP00r/qNmuOhVmpW7DpqIVdK/uQxWkGQjcLLw7v0v5QXiRVlKg3paXVnzXZh
7Gtrix3ArL+6kVC/gJwK2DieaECTfT5IvR1LC0+0OgjnePle9EcJoquSobD5qqIeL+ErhRs/d6dW
Ph3O04M930dX7J8x+tDrLR2QizCBsvfOT1+0nrjj1raYTLJggCnHh9kcMF/7HChnARrj/d51AFVC
w8MdWobEfoOwr+IH+UeilpanIfzY+X7uBe77ewT2irX6f8s2d8AsC/zmnlBM25sRrYQwP/uYItSW
NXk8ejNVR7ymqlAv6DCrwbuLVcdlfSSD3ktZIgc/1GSog3EHN6+HYTC65olbLoNXP1ssG3DnUwW8
N+VMBWV+/7tdJIlJ98oEz8L3/tUrT0YW3PQgNAyHsJ0vLurcv5CwbcpBaVsYiFuAo8AbL5KCOhlP
Jjl9uJBDHdz31s+UKc+Sbg68J5B0WAZ9nBXwWvRBBRuemntYkzEotGreX0kYBtb66dQmR7ZEs36W
Ql7S45ST+k3Y+2j2GyUkqmM1vSHGZlbpBsxn8uBmUl7MFZeRKCBdc/e9yWaqzZJOjxQjjqR3Mo0t
R3w+ncSYY8sI27++fWyGMFCxaIIZLDkSIv0Olxsa4rgSYSvajJHn1UXMKnl51p0PwumNJ8bdJS9/
FP69BfdDXCcylKJycR8IF5+zP6aFe4uJURkYcHv2NZd6PUtKULvS57tTeON2FVjse/M1PlGPp3Kc
P61yF78qE1KOknApr39Vhbw8rb5KDdg0pSSZAuXmRuqcO2zK6+Md0g994cP+bHNO67QTdm7YPwpN
aIIBRlfJpR2l0xnk4marqx97KOZw1+BTFHVpPZTIN+6mtBLb0TjGbMYajaUFRTsrJTiv6JMmT4Qn
WNbKLloZREhQC6O+Su3l+Q0977iuGZAfCaDrPypqB+56K72sUk/LpMXJ0kNURFVnK2dQQNlgQbUr
ykDO/xSrchSignCftcL4GcCzQvDcyDJly6vw4FMtIDfgo14zswU86FH06LeCWyeZ0TQThvMnKy8o
A6e6NK3mEgq4O2hq/+YQZug+9HMyv0AQJzl1kYcyncLVbpzjDIgPJ7mMpyfPWqxjT7AiTS7JOqpY
NO421mnjFBGwxrsW/Rm79msq27di5vLPGVYXERfdpMWlrhzZvxPX66wV8yaqxA0PNCgKKH3q2WDE
JYro+6lFANKQxZaHTujPhaxQZ1mTZYoye13q26zcYucx8p9FU3sQn91FxJVV6XR2K6OSk+2YgwVM
pg4bKBiPZ0l4CZCfZupkhtQJZJQc7fX1woYWBJmz2gxhGg9sbN4yzbBsiy1wG/9779WWGumLANG8
OG8BTU3FN49FmKWnn1obEQFx6szQ3fJNU+Iwib1Y8LH3ijtRpOSFiS6lRu3oV6W0vtnc3Hg8lXfc
6LeF5FzqxaK+ryW3E47my6cBqDeusJCQSZcZ+c7EE76cgza2vJaVm2C19nKp5Bs193jfjQ4ehECK
fI+p9tSTD2gfPhEWNqTA38wvShKuTdU1sHtFe6r8NJd0KkK8o/fsjme6PxVe5rw84eZsAEVeW9RI
rH+WuIA2kb/RDLk3glY/jf/9dyT5Dl8uFPtipH1FPsEbZAk8KV/x2lOcUGshjn1bM2YHRMKfA6e+
OHcBoLrILH2W8bY0DTOsv9MzFyFI8y5dIr/kBnVIZBlcwtb4KL6rMoX2onTPPiowU66K5J25D5nD
CWwbfHo4RxGweWExkrHQuG9HDOH3xhDdnD9rpIuPVzqx5nv9fyVJ6UgX4+mL7RhZol0r5/37cVQg
DAvbob3txm8o/HglGJmvmTjquNJOBGoWfyZfMGeUtBig/5b511lxorZQjzMCgjvCGyj33Lm6FW7s
GmmJtHv/W0SKA5p0mMO8Krn6h7xaeFpgVTrZ3bMBK6+gt+Z2i/gDT6IFmTL5ACSkFTjXdJyIctzv
hyKaK33P1ZVGGdh8bkBB+xbKdMuUrrp6rXv+8VOEtVOCndrwUD8GddpHrqGD8ufnNS/lBTfkZSj6
LcEMv2erGRySLOHCLFEEz3LOAgjugufrQMhtKwpiPDQJZZAFc3m8WvlDFN0GHSfiTUW+HzRketpb
+/pI5y+8Vwbv1ii4wW1UZ6N8D9SayM3BFfWb4Pd24cA6M0Sr1t06/Xdwysy4NfTT7u9KYy9mIZZZ
cmw9Gq5I8yatT6ztg7ea/bIY1ogFi22E4sk3othx68E2BCz2P4ethlzdbvhCXEuiqOeFrXEOYiV2
j9bbdqBXPAlyO7qDqwwpQX3gmzan/UF7GH0fhnkfvodwQQ1C+UEEfS3I+PbXDbV/rmG4z3p9KTxw
CL4U1yrfq5CLsi+eZwz6IK9ClDveAKLiKWvmO7rCroMc0zlUYntaLO7yRgK6Ubdk9BpvBnffo6Dz
R1OIvhMUB06d3FlwbnkboT5IM4L1QI4ey2DIUdIA8rJAjIeIZpjzbGw/yIHbf8vA6IraEHhHa7mu
HRwv+q+cy639WEwkSJvFwjEtq4RaRXHa0715TRRYfM+vi0ZrIpgL7zzCsR3ArGYdaTkiuBzrkyvG
sv8uRNw4E4Mqu2Gv1/228N2QGtEgajSbx8AY0n+JApzSJ3RRRn5T5b9lltFlAmBPP8uOWjmgyDRi
ateXE39KGoSwcAvBVhQxW8nHRpVYhzlV1LqfIZZr06IZ+tbQ+GAvkDnxAABhtLZxfLIvwsXBzM4m
xMNDrjrpkED4fiCbAWHcT47kR9ROn3bQqfQcX6KWQZaKsEqv/wqZadL8A63YuQEoFHBcJlYZ80tj
QcqnJPqvbKsC4Y50EJ8rreX/Hx46qNhI6PJcQ9VdAigk7Armc1VojDG7c2X6XNyj0a/yAV0v5XZz
dxIX+JiZ3zW2odMp0sCy/hVonjGoWBY9df9xlLROkmuDQERYBu63kMZjpO+GkRNN6ensrYxJs362
dyqW9hwF34myYKXJDWs47mOlG3kUZb8jBkvwJaMTNOSc9DvY7f1IGgwDwd0Fsj+iJjWsiY7Yh3bE
OvVqceHAdXqdCRVA7pyWX1xC1gFlZknPadP1iRkvUfQSOYBS4n2RLwn7hSUPbo+q+IAj7euE+DLL
PWoxpJUEenS0AVwDR61G+D9l0V9XmLES/ocJSNzC8kBEgJM4KbhN8yJVCh7AjfAVnCn3YSfJ6VOj
gH31u7lcqrNqQAt0mbQm6poeyf3+QUoXTlyakN9KuQlC1H6DQvl98dPLlWJ8Jl0o5SVyinn53LxP
kphemUrowOE2DlNJSBqCwC6q96Ysis0y+fk3ZOOc6PGZP8k8PjZfNq+gEVc7SrzUTltnrxSGvC7P
V+Mkujk3DsdCNVi9EpbzOxX6xIlFiGW97pLnN9VDrLVGR9yEAvtmLH9TzOjD2eP/TJW3ZZDkIktE
WPZ7QqCci09XVdT5hj7IAK7hUuc0+MgoKB/s3vrYE50lBsn9GOuqYQ0Au2E6tj1MK65U2nm9//dv
jBdtXQOQHAZT1N2/9nW8CKfvDJuqbJLcOW5Tpp8PIROirgSADMN+ddwr369S4xWVnmOLWhfhlFvx
HknfrM7uXDEshdneZtDPHpeafzk/XS0RsWpMznIjzGEl7zGxVpG0YVX9JWyZY86CIzLHU4Fhxuao
pWZy/ZxmzFKhX4gZHSqGjp/6Ft9QKW83Y0zOvcI/Os1etFnjghUTjFtHbfj4cGoCm1Yg0Pe/SGG7
nbSvomIIIWN+OT0dhLMt8CSTYkOJ2uNjjP4Jcdkshoth5xG2vt20lxxPEsTbz1m2adZrz1+0CK/W
9TnEQJWrPPohhJH7hRvVrFtp1+9MfR/9MuqY3CvfyveP6eyBFig5dmaGLeNwuD1VI8zqOKGeKTxQ
1mB577dYjJ1RGhXVd3jMzfh/r8tgz5hL40BzKEyoT6JZwtMHF55ENiT/XnMHf8bsicj1cEwbJd32
QXssbLFSqyxRF6cA41GhX8ePWNqF+4PJHNCt1wjd6z64ulJWO8guT2q+wOUdFfoMnM1f2SwRsAs5
KQ2rqplHNgzBkJ/nJIE9cSMMYDtnPtSbIuFpP/b1dl7otGXSJJ06mP7aTSpYpR3avCqt4d9af1Zb
nvN2ZkmVt3MnWuuWs9RoLCQsIHfUzfC9IaWsQqTgvUPj1EX+lY9m5x1TfqZVoK4GhREITQrSlF+2
uO0oB2r1I6SlZLaa9HIzdfU8gdYcxmLH23MkxZvAN2QtaqQG2Gf9X7q6nUQE+yFKOSOjQwc0fuVm
pmfT0zvVY9k5xRKQxcPzg13HFgyxU/kTU3EnVzEJPpQYXQ6VILJcufvNydKgQ9HPUmQcwQCPWYZx
vOCR0eFvJNOkzYanXYbfOsmkgt9CYcAJZSluZ4wLPbdb5VJpPw3kwR6EJMX9mIqBZci9/dcPDyP2
becmNdWxHt9xlhXs+PRqq4iNMawcq6GMjgwkR0B6D3bJfasFzS+StS6sfGYN1ld0Dwo0u/TVhNM7
gqDHOpUK2L1Tbjqm+nK444Fx87TTrbY0N70sBZ1LkjtI06c0PhP0ckE6rTIhBuIHSfThljM7BPxX
Sjn1XMfkNNYHtRs7mvB+yQF0Gw6Qq8PyHQYWr/IxB1Ac7GcEaEqoXGz28zv3ZouvDmOz0uzMuNZd
9dRpukNQE2OelnxEBGuRwz5n52xzblZpV4znpWNO3Q72ySfd9jZFmlAXQ5QVDA4qcA8gtzjr78CX
g2LaZxPE//lZ9tBGYR/7GT4glOIIVoKAjKBBdHxWxYem+1vhTpcKr0o6fXtqfwCRri0GOaqy4gj9
c8FJVVmV2NfF/ahRJV14G+Pye+Ljg1iXqbI0mq1iRWsAg2AzZR169wzEHx1DgH1xtvyV4wN8nD61
IpceB8MXeSglRtO5YnR+4mB6WXA00M6MWFaoyJKLQAo4yk6dRSlnF8ifMvAw1VtM3S0fWAE2xOPV
W0N9HppXGr6P446c+Dc305lbzruNNZutKyLyA0Ih7LwjQihwyNqIGMk/JUvkD/K5Tdg6o4MtfhJn
y6uq00JzpX/0NIwvFq7Zf05pclFI3ulWpord+rvMkkaIIAzL9bihcjcCi7UovOHUWmfA+mI00RcC
O7JjoTIXL2Vld39OK43ILU6B6CtfLjf89dvKwIfzGRnJMWlSMaMw9sp4l9hZ5f7WuYxanZfT8cp2
Hcwy85mLyBpyiwqMPFy0ThykBRhZfrRyBOFg+V5Qiw/suXOzs0qJrc7BtY7LDIhs8pUDxMGZgAWu
kUQObz62FLQef4J0kX7N6U7/7oAN32PBqi6HGPnRFIy1us9N9YI/H7uui1QHMReXiBWveh5s0KJp
AAf82EjwX0XUtcXMFIsTrGirZIxDkNcVTyENjc3HOpXdEtn9DbkVn2mjCMMMirXEVYQpdICkp0nt
pkNbMBQ1F6pn4sO/8kJAmzRpnEq2wNZvrnBvkFoCuyGReDrYADYchIigK3TIh8E7IHyleE9m0u0k
/uOlBpCdgGa4pVyTaKwroZCqNVdKfxckmc97DfsxJ1ipLe/aj5q9+AYkrJ9NYdCSi0tlLUFkumiE
IqLiiT5sjBOjaIVmh9taduksDMBIv29ISR6SKLTTdM2SMuAC3bqqWATdb85o+RtVxkWzyAstrJTe
s75xUGIRs/1LdeeMFTLnf7KFUGwHaUCzE+MZikUU6NdFfDR72iqBM8Zd1PZksxudzYrY33m+d1o7
rWjJUnJuuR0Lw0hosayZ6ZFUCLBchZHUEIwRcNKt5GCXgwU3NsKAyKlOV5adH/BOMe+bTL0CQR6E
IUN7Li3YlbV+UeIhQwn6fYFJhR2KHMTFxQh1I52YX6QyAGcd11Kr8ivow7jasdIrgYymbGnZSTqr
ki7XCjuhI0ZgSbcKebgMl7KswDpUgPgIvsTAyKOF6LbHYDXtFE2187aATg/bwxgksCR2N1ChkkSG
E/DjjSgkxqTST/aBmB49LOOIao+PT0iSxNgeaMIUkaPqw5cU4AmQ/NKUJ84ZWLcyIJoKbB2MSNMb
xLm8c3RGfXWYPD1L+0zzlEzcYSL2WcFZAhr+ONUHwd2jeZnRjseExlT+N/U9EMZLeM2Gj85lZL4t
vvgx+Dm9G3nMDY97+a3zqbVias8Y4ut+AA5C1+M6uktSasv0VhmWtfm01d3wmWgm7HeGVSwZOEKk
4ao1woVOVnnHYVe8VqN1VCKx+67Ye2mAdTpbbvFQL5awMTK1A/r2b8gAWXmdyPWl/51UQYND7vMi
XAxFN010l22wUupB9rLu9X4o+u/Yab0N4gygsXWYOV3Kkrt72DdSfj25RHGP4aHi6o8SW70KjAzM
2K8/lsWunrNldh8GVnBD9QFW1ZFSsmgW/Nc7afzGSelrwEhvyEaD7OKfnYKSZfBzvCFvOJT172+d
3AWm+qsq//TkdXa83sIYKAjvrAgXIlk+OLMux8OHj0Dvvv6tykvAuV3gitKNLj7qf9TQtsA6L8ri
XYtdtVAxuPtEyRfxfUUv4xSWCwdU4/3eZoBNDz7IWCSVpbePmQ7b7ZPyLb8No41lxe3kDlZ4mgnm
V6c4J+0221oCl2sTIpB5Agr4d6q42mbhTwtsuqG6/9MJH7ZwfAadKHo6KhMpziLoV7J41Vk6A5jT
4QcyenJdEPqu0oBhF3JrWQnx+n3kWTO3fMWycTGhnQJXhcR3ZsovyHkSPf0OAPoawX30852vPuKe
ErTbj/mR8vSnt8oTPNnLejaR4Rbipy4DfymLSwfP6HV4xF2bm/IYXhEooz7uIshJcPc2NlCUbe2O
RehNMrDbhHiGBmbt/vnHU/Gp9/ZD3ZOVD+O/090f9qR8gnAARAET0BZuvNs5Q89XSpuKvlQC+q56
M7Il3OLwGIPg3dsNYFNrkvA2UVqBzqSUk77wJcWvK99MmJ3eZFrnGESkObWKqjd5h70kC6OIZYDt
Yn+yFSiIyu1SLnGa4AQp/x/rFC+Fdru2H8IwkvDA2NSVe5pIyzjoQd5oOGITfMNTqTPfcFNRu/IQ
92hQIMhHn+wi9IRbAFgj2KXm55nPxxnBj5eX9ZmHTA1XwyTs8dAxydKAUOka22nyHEDw9jNWhdiZ
tDE6937EwRVQn0VeKadeja29Y1Nxd0djE4gD911IvtD1LaRXnHXhoupY3vjoUThVor6VzGV0Ua1m
geUThQATEksXWu97xpXnvlMIcgaXWjB5xvBOBe/KBapD+XP/jm4n0DLQVnrFJk6SVK5IiH0cvdAJ
Hh8jXe463+qUGOtZEmMJIzu9x4DM6U9HaLkQtijUPU1nA5W95Njp5zaBCnzm9epf6fi9nCX8EwER
J2l70Cby7l4I7c/heie+CM7IE9JHHB1wb97k940A+TCIUJGK05oxfN2yhXbrYdcBBemwi+UOVq60
Hkqm44bah5SlQPvf2UuD0cB4B1JsHX5IZqA+noJCKF6WIcly8VPOsD0Fm7k14OET/az7x08jSndr
JJWEcyrD4pfar+SFl7HDO0BWZ1+9bhhQMWpyiosahH+JexVVs+w4dea/YS1gaPka9f8F7dJdT+Dw
gZV6wNKs7qJsT3ypW8S4+iDSo1Q+pO3Bdv58yT1ZqBCPos58WXzoVSJr0HuGvAWrG1Wa9PRtbme3
nB9Qh4GexLQJ7h6rPVcOajPSrl3Z0IZvgngJy5dNxlfSSHVJ+hBhzmyB8C4FGd6ityGVfRfj7Ghc
SqRicDOvtj3ccop11o8x1Ukd6UeGq/dDQZ1bf+HzZkQOCmkkGCornv9IONp1D/IN2hM/WWOs5w33
GBjzBy7o1QMHPa7LSS/jDbxRLXNfLV9rY4oKHHooBSWddO7DLoYqgHacSVjCQNaZ9aA7x4OFvvKI
F4fx+pVPiZti43iq+1jNFpKW1wj8L2G0aus4bqOyK4MPdNN/aYgHiOi45ygQQQuBjcVrC8sJNV9w
nAvMMr1LF1m4l6h5BwG+8fxxHVoydVRBRgg5PtYmlZ5rxBBErfs7gV4U6C4baXdFhao1FqVyFuU+
ovISKI7oOHnImLJ2Zh7CGflPz6cfcJIcBazF9XnVM2PfjvXeUxSphEDKJalBjq1lM1EB00gR1gQl
Pmz2yRvYdSQuovCBVv+4EgknmxBvpzDD7EdMAScuE4UtgkKEg+ZSwSbJ7G7WlcybCcI4NglInxUO
PrVeAm6XCb8PqxLydA0KS8wSlLlB2FxJC3clCYFCml9pcurTf5MH4rgifkvSghh/uqKrvdEbD8Si
J7wSqRslePBt5OCk01Pvf9KZw8RRHBWxXSMuA9wA2F2ba81zk5i/+khiDCCDTCbQCqcBwtSIjy4V
SAYElYgPkbRAAqzwM86XSCVH67EGWCLPhM9H+oz9zMNRX5AADEgOandTU1h5RAXTCJqqquDiPqUI
wNnPsettfkCMuDtImcXDbywqL1lsAHVy+wYRYwfgEx8rgjWPKBauZU4qSwW/WF4GZhBeGam3JROE
A2FhUBEbyGaR1uw6LCGRLgzdJOTqU54kefybhrZT6LN4SyzX4FFE6cJ3DpHGn9rdtUVjMthISQ8W
gx6AtQu04uTbibzOJxCiNPDV/+6TRbKwkymd9/WEN758G+fk2LUgFLsL6Xpc09unK7PRcYePr9B4
NMqR/1o9UvUWKWB5Red3ItEJxsdPvEyHHCsZHyUgQr3UedKF54N17bs+GOfq5Xkb/m/j/kyQpxR9
Ozh4N8AUUDeHVE2bzTcvt3qcux6tcJ9n91q8igBfy72xxjybqrJopzdkYjBRl1bmJHZ+rJkrKWA0
kCY7/pY2DbrAIbKOZPS8FXaEf8pn/jzjSWBb5XbjSSabtEK8nyP36Itm5MURyEaBa5/ocin0odTY
ABLQVJq8fIZlEpgHhjTgr8+owPg5HERkMop57j7k5XjaSp3Wr4hYf3mwnvr+231dwXS3vH4oKtgN
vf10hfnxz/rZHxBv7orFauLCeV5OU4jU5Bx4V61xdr2o9R2RDjWts7SBxa9UFqh2jvgY/V8IVHLa
hhKrWCAK/HX2vZVYG4p0sfDLukq5u2iEz7iZhthf/1M7K2+9DaTsWwpdofao51Ux57l3zo2UXfYy
oNqIxHWiNXxRNgpS+kYjq1XdQ3a+lT+7ys72zGHS2w71Wip6YAv1Ys+WvA98cZxhwQ+ChBx6tPWy
Rkw8pcQEaN2JI3OtEQPKpiuBeAoqSw6/qzpyUFzRsuA2wEfnpJuciAZyMIcSOjdQ4AHzkAvr0nkc
TDk26mn3V66QRF85tLGOhq8OulO1b33fp1KAgVC1b2ZVjeUhz/uCRVwgTba5puH49FT3OSdF3L5D
LiniJww5RThHugZmAPSHW43GTdyajkGSrZ9FGw9G9q1RguL2qXiKkGBONXlsP6xAwhBFIlPrbrWc
VbqkpL9OzwrhwNN5v843kaULUhcYP6hbmWSK7U+5F1SzI93b8ncK1rLvBMTtQi8SaPgcSwsKqPlm
9Xda+skJhQ7IqGXQMnwkwIBwtSIOXnTrFng8fF00dISZ2xKX7Y8ZBa31olTa8PZCnvMrZ2lKzUTW
6dxv9ttTAJgWj8ZmFi7QNwH82NiltqY0Jd4YMDe97sHE6BAP5etgMISPLW7pgDwTLqeGrGwImEm6
ilg9qSaM7zp406W4DP4v/CrL8zrNQlDzEhpIdJP2Qd2bn1XUSZMSVH1/v3ZmAjtgl6NkX5CITVkQ
sZ0ED9vD12aC8olaq+NxbSWyaKPlLKcRpNIjyLsJE4XVPnlv7cMprCD+kojQDH2LiqDm3Vq+dC5H
/pJjO0acanfCRtQMMag8363YPwQWNpjdwh6Ce++p67ojwfN0FZOvOgdQB0ZffuTbTolYpMtFvStL
bnmTcoJmJJyK2gwyZFfanXrjjchHlOlLTMtLcw3Rt8vS68PmIOWPJmlrVRBaITHoGW5bNC4n8tM0
ISG+y7erIQUDDIAF5Azot6ULeJrJhN1xYeLFX+fY391VPK6FepzXv6Xv+kI/pcySgrHcRWglViR8
pZD7LHjSnh83PPRCR119/n+sptaGBymglTXDi6ndpHPt8fmt4L9zRzrN1oHA4aVLvraEMcQRuUYA
GLHZiHKfLHzrccHcRBQC2TS1dPdxZPOHYt5r+PoQoPNGYnnmdChJ8KJ4gs73agJyN9BocVP4A3lJ
anjBIhwDhfrgoZrejGGnS1IXzWGDP4/hy0AXqyjwFyqyg+hkGaGs4XgdBSfAWUMh66gUoMHMpzOO
90TautDnHn23x1iF9yBMJpMLz/gkv0uEoeow2V6pwy8yl1KTQ/w/rEthBqXK0aD/oz2RpRe6LHli
q/IsNLEhJgXPgZhQ5BTk1zTQogwytQFou+i2YgjwQ9jdljODC/YaOKSyrqMMi46/P0XIM+NSxEme
f4oWhVPnFFiWpORTqT2y8Rb+cCtEZT5SgnYXvBZ+KkPVWal2Hpg17bC/IgtHl6o6TWnfa1eQQeVN
kFkLLEKrcH7+KrDm7YMh4AcJbW7qLpqG2Zt7Guk9p3FXJF3SAjrvc4GiNUPEjs7VDA14gd5eeqW7
JTe/aeS9/9i+ez9culA1sXbuNZsOL9YJGttVMvoF1oGJbuu++TS5wMaEfS1vVUq8BQi5RXR7zwwH
JJrI2mr3pfdov0gLj/2f+fzjm6OXpPo2Qk4TuzsmpKAlILhayPQmbHFziemVDiMXeBc6gaQr2IV0
05mdT8zp92CV+OfRL4lYKSyoOAt2CDS6/IRjlDTgdOZQusgbi4hHobeXcmsN3T+0BBJf29q6UXrs
ZJyPXE3fn2QzcRlLCIDKyRogZWW1FzojUA+5tR/ffSvFSe6vDEaw2Ixk54BnoldptKgMnIoQRd0m
WBw8KgJv6Jp7ClCm7jPflVF9MoaMETLgVUdHBcyzqfNyuSY3mcEUIL1U7++rFVagaa7v1mGz1ydU
5TYcNvthbUd/Xc6s6bLaU4tjgnxGpSnUpW+NRf+vfMuTV4EFjnQrKcn1zK15UTLf83c92TtBrrVr
cB1qfzfNRh27ugRKch+JfRtXGEzF44Q6mTq2nGmWaI3fcVFSW8rfekDtJwO6tgcnfIQlXV6jzgUF
DF6+G3JSRF47A4bOvu4p8152KEyiZioH/zrC/eyirDaGEHFoOvcOsvVWctU0HJ8ecL44htgX7Nr8
Wor5M4t1+P+sjpU5LvpiJo8R2cE/1SR6V5eYCJnEefKt+ZssLqjtQBvPQ9YucIplHub0LTMsy3Oz
28wMlqUdrISkJLQpY4HHTnicQovB8TpchkFwsoMrcEsYP/GLQWXRWqT7IvYkKYd1WOsoBKns/tUs
5iII4KRMFBw2wRtXFGzoOkuodHRp+1YgSqRsfJHl2RFSn+cDuSLVb42Of4Z+NDffawdwUW5UK7Q8
TU6mef/mV8LpO0jv2ncIgIlbWyLHjl+tV6K9KA4p9ELx2t9PNwfZGCSvM0zYpoL4N6uUmSty8Ab7
9WpN9lzvLQdl/jPKy2/cLb/qQYwxG6BYT9K/HOc5VH+bZx4dMgSZnFlZ+zwAuhF8yQ3pFXkfqlqO
/AkCHxBWZnCeT8g3EDpPEPU4/w+dLXr964XrM5RDK7gzyBEjijSHvVP8ap8qW9pGyaET1YBNu40O
r2wy8PhIffGW1MGwPOXSNrAQ8dDdUAPYIh/GiMzBKMXPKgHFAh91wQgoZslONFnTb2yJh1Mf4Hwv
4aJpXgLW0YsAUma00mwKeAhAwLQ3YdywwoZow4SG3P1qXe7EoobjLPsoxHpIpHr/ynTH+dPdHb7f
ExRxYbrOLzT9jj1Z9vF5Ug/cNqrPjQnmFBR78EWepfkzZIy2y1ZeABuAVDj/ejhlF28V1cF8cFuH
FzINW1GaDlk4VKoZ5iwk4zdXya31giHGw3qMjHg1XOAckPZXSm7P0SF0Yf37/tdRBl9r/gEFIePe
TX9GRSxEJaooLYthcaMGpiSeV2obOxL7l5t1MYXcXeRIFoU+yhZfmttrngxKsrHWvUPRe8Kxh+xJ
NK2FYc29ZsDK7SqJDJyIfEWgqH7PZ8YJs8sYHR0UH3SeujVA3mpY0IIaNV1IK8WqJTNpVUMLakFn
VPT6koos8ooWk85oLCpajkE6aSKdZbhr9UEJLYsNmcHG/KmJKXdTDB8MSUvCaBYZhbAJDUdVmkYK
cUIBIOSt+z1KZXdg8oqp/3zU5EhhQAG0Pnk9/YnmOWEKDhJfYlFpvDT4jXGtX5+1qh0Mv+IuQtRm
E3dVrvfO3DqPktaDarMW1b1OcW7yX1D7XB2CDJXrotQVPV5HLbBI5D0xxhIdLJ//LI/cNbmystu3
edZ3A8MaW4LZp8DSX0UdSf3B+BTEBxq/JpdCLOSIR91BRxqeIXG+w4XqdzeOBBXiqwiRjJVW6tE6
X3vDdMpMA34NjhKdOt5RW7yaRFSGvF3rQ3yM4NX353/KKWkHqnowFq/KYcVZ8/6BeXE1MvgvOv8s
SXrlmrx1bDkZtxkDyDj/hxr3fHMnDDtNSL6oYTFiyg0vdNGtsZ0/q4YHgJMcibmY/wHHafAriK/a
uW+OFOuy0ogRG2tqzxnlOnb8LELbtJSaU14/yDOs0Qr8lR0UJY7WEE7dM+V7GeLE69q4ESlHzuQJ
r9ox3Eq/buGJ1JScdDdggAVEVepLXruqi49SbLelLiA2419cS91vKtn/MWjAGhICqaiyqXl+lNTy
Kus/l6BRm2TPIiu85IqhuEEKvIgOhs3F4TRrIK2t6wjjNz0ERLcxsAJ+kuq4uhYZmfTBNhVmlkSF
UFVumW4lsylrNbuq9v25A+qbO942InguNu/IZJLzvEnFi+wWHQIRtd4qfCIF5Czh4XafbYcBl0Zl
0EwByOQ+NbUi9Sx9sSATVcdw+LUwRpZYHVS44c0pWyJI9o4u8Tf14uuVn/bAJQJimtImsy/Em5Bo
fF//7iVf2nE+6HrEOqGBJYfJi89dyT/XjAsHVgz7lF7YATjoEnbLe64RnfrzHOhbCPQNgUWAPDG9
uzmIRW8i+CIZSHlvEpbNwcW8DvraurBfQ85w5a0zI+80xeJO2m14Om5TaEmeQ+lHWYPO2NuhEYQy
TqUO8ivxRcVqYPlVaiJOS/EevaI4yBqtmtFZCcImjUkivnVho/5wwoNE6myRpqeN1vUVBQkJanVR
6TMjSM4c0KTzv0OV7vkja34knmDFbQmA313kEzvrjhhDSn1l3u5y7taVMIMg+xJOf3OcZLp872iA
xxyGD8g11jS0vzBgl6+7k7+WZuReedx0DE/GGHMo7noK4/g3dFfQlX1HiArMvWgUky/oEebS4NZ6
IUJj3px7sievmAkTOyeECQfHW8OJ1lwWha3mWA+c9kM0ZFB3cuSxruLXyVXMDUh9/c4jybrkYOeJ
5D4TDAVsE+2j3nhO4ZF10nGlHQuaZkz6ioIAQKaHKX7iZ6EFQ6bRnbe1unaqsVhQ3WjVpQ4zkARp
ouCY4pXPEHs53B5lZydepbENMkJ6ZndwIqaAGr5tR9bvl943WKX2rYPHrLZg/m8h3OMBjqfwDdIS
iNkf2NzxPzyOBBlqhTP6hclFnbIXsWy9B+hVib235MWAenlVhNBU2gIMidNvuHaRS8Ms7eY4UbXN
sLEcyjEuKaZTc8JFDF368jeBRWrfggcJP0PPY0ok74f1anEm6P45/9984zBiP609EXpcQiKwr33v
DLqob8k2nuxuJQXk9FGFiwlSBHxRzxq7lOKx/4WWQa0UwE0ZD70EHDIa2ODQz5NuN3eBYPEtZ6F/
cjinaslRUaMJc2fAn2q3AuS7sW+DRJz9XzhuDmAH1Peqb2o/G5x+pVJM3SHrwBIwWVb6Uk2hXf0i
Z91BHztXQfRv/uptpjvVFZAFAmfbaTHPE6W3sWMyY5nSEYh5ZmddO6FpfCMYNfdUKV7bMKFuFmbf
KFpHelYrVGN8HocGjDGDa2ZquRvKKq5ve2NNLKQo8h9wr0Q2maWOGIkVwz0OI0CxYHaqWAifmGsh
yfhCMyFx3tzb24XVF+fWatSDzzpYx11TFs911lt1Iczf/dTjlSS3ao1GEkoXMgllQ6b/bGCeqK1D
XXAwdiET3feVNmUhFW7N18DGSneH6R67p74+FFXDXLojLbCZQ43I2KJcY56aMi3LWG8B/jAhFcEz
dMcvK6AvXmKdbfJchLMKcmm0mMPNdLxJwkICDRbOjwwGOtAXWr6wJLfcCG5XgOpy18dMjJBJj8+i
3ff6TqSwizjENBV/vxtIrYHOdtVyz3Z4kjBL5oSTmYY0v3fFKBDLp1KzgTkqWBtT/googkxeimi6
iJDZLI9nkplEsbGd+49ib2lTqDQSWzAu7JiQIi3DlHuy0P+l83oo1pS5bwa0tTvZw33hyD9NcSB4
ip6YaOTlynZh2PZRQvn/iIZiw0mzWiWvAg9+y44oMMRF7527UK7LVUHD3pRi4S9Y1kO4JxpvAYGu
ghLNuV1z08frOZWe+ngQ2MoQyrO+7JsLcCd9FMSC0whXgl5ysHZg5FA4or+igN9YFzETEGagzMo4
aCOb8Mq9JKZrCaBajE5j5raBJ2/819q6u2r/vYEtq7Er8S0G9Td9FWlba4nRsoVkIlPCdUTQm09h
wOy1GH+HPmTs2J5F0hNb4DBSsMYNrXnERBRNVYC7AZKo8IKzZS9WG4Unp0zsLcczx/q+CE3JGJwN
oc071MkA/B34iPLTaCFjjy8M3O/lOOX6L8Vmd07P/7wXgHJJMP+abM6CRHBKUdhEM1IHlqBQluu2
UORGPzxdyBMOcFImPbf6AqDJlXNCYTLx0Kpmj+TZ+ylDxS3Ml8/LmB7GoJOIQvWSKQiFjCSjB0gn
cdPdsEgIJqs1p0gnmJTdlu6PVVr0gOTamfNB/bi311CN37Zdt6HbsIyDXlmkNf1DUb6g3FsOfjw/
WU6vx/Nd7xDZhIfxzeXE6VeIzel1XZmSYsgdx9A9toMNtglD0/cfZM0MzuuvUNHJMQpMDFAJgAIo
6dOHLha+AXXjiAu1m84RTp8ujM+l6dAJ9dtvsbW+73aj1Ek16jJZun3kKu8aqLKyYAM7ApDnatVg
ed172HALPqa5cJ0UrjF3OSlhxnzbwLkZ2dmjnsZTLP07sqXR4EQSuSL7t8l1NlhH0sTlN/8QBylx
6MRHJ37/b3ChrfGefw8KnOTTgAekFK/7NUKHA6K5eZOck2nWR4DLXEs02OgDGFT1zP0wvTgwbShy
6Zj+RKmt1uzWXpHqVee4sizZ6wXN8SgkxCNI+63RDSCGSV4SaQZUkaq4IUgd05uFMd5Ci3lZyygJ
OhpH2Fji8AlAip5RzFFhIQZpCCxnWYWLew4z3GeMOXQ1s8K4NRoaYvoR5prCnKsPkpjzMorZ+XDB
wqacLn/OREvuUajDJQC/DHsMWP2GLs/bxY3Ulni6JPHP45JsuHgzR4IjtCvWbglw+VJ2ngfgEfXK
gsaE16xZBz0EYrUTt5OLIdN9qORCZV7VIejmXdqzhgi9D40iTvFJv48xiyQDV/iI0W2oODMfPx3T
T8dunIV3rem5G/j34nDAadPOAKu81C0Jhcigt8B27rYaueqCrGPZdjstrTWEZZ7WA5zdV29WRmLX
QfkI4td+VdnlKOzvLkctppjy5hCdDEaQ9G34GocxmmMGd40DeTR3NUla8Rfa9mea80UtfA81CPn0
wfYYzgrPFIlRkvVuUJBPhvcNnl6dIPdcrDTx5QT7IgUklpq4cyNBIdGoXzx+ROYgbMzCwDhNYmrm
rczWDHlCq7U+9GbhqWOFKrd4uyq+cr9neoGq8pDvfQ9G+4hMozXtdyaKnGjAYNks2juX5/qZEglm
wGkr3rBAMDp60Z3UhZdn+oRrTGwps3q8dK5uC4fhVzX/WeoGAPfKD6wGhndqWpUdzvkeDV33Rn2k
rp5j+iD7Y7N/beWyuW0tIlrnm987vi1Y4CXCAsBi0dQIM0bM9b1R74frYLD2s6W7nHEPY1eDflax
3R3bhl6srV9oHFCqx4K0+0mU+fCU3ELSZRz5IsY8PBsgcjkFA78thPUucQpfAXbieUgYH/dBe9dx
P5MH20qHjoXaWjhhdnPC3cwWakIJbojFYumfI/PoXQlDoFcbRfjnVLR3O5r2yVb5v86Nngc8HI9F
gO169ef/a+O0qofj2J5f5QF4XmWcvMENSWEtfSM0VVOGHTgCmFwzLeGdSoWvUIt2ZwsuPGrB6wdb
GkB9Ejmm2bHzXaR+stzj+fkndVB/P0vghqzgZ+uOm9WODxGU5sIyiMG+ZvnU+u53iWJZ20J7O2oT
7KbKAjDWyVvqNhH6QTtD2QHeYX19YLCxmACSI0O+LpDx5yVTKny8vYZ1Sp7Pylsowccjr13vn4uY
jAxg1ofqBsgtdfZTwILkpj7ssZUg+AyYS8BYznM98Wr0ykRJwPetuNrpjHw21LBwFAzSdrMgGE6c
Rj1mqT/alQ2eT4QGM/Aw1S5s8NS0ouOmktGoN3WhD5raQezWtLmLy2d1R1LxqENzsXdi536/jAIw
5wbGf6VCd9fwDntOoYMteOH/PC0VHeEnIaqHh8WhDyT3OolPhD1wwLzpGf6HN5Az6GM/M5wWutal
NuojvVKPkT7Lo5iS+vAUTbwZDm3WLKcqEYzlhRPyhqh6z57+jkP5bzKWAlpCY2noms3uQOeFK3RC
OJNTZAZBW4PV3oeRzSClwUdBFPNMp6eGKHT8NdoJcUeU+bjid2k6+0MTnbI5kfGab2cFptjHxHOn
2p54zRxBA/0TdGuiMD83N4iC5jp7zvoVsVWi+/NmkNiuX2CarTDXKQL2tDl8n1tUrEUbl/jRnVTB
F3LEaXUY43DPdFduVXdXLLU81jh0J1zSWiq9OxSU5/2Aknkxunv7DCMYBjmOOqTYOXaOehGt+gxd
PqoOSlY9GrBZZMLef4xJXRcYjo1LhpZPhpGtyP15W/2N1rIzSU3vQuYlIptho5EjeEIGLI0S0MAl
QQ/b6xeG2vOhAuGg29tEKHUELrbhHRGgRG6IzN75kcaZDsaAXsRcZXCOX3dCGvOkVl3/s7D31MwX
GuJzTGIK3NwXKhgi5qlYqaL/Jrt3wOAxUKPZ6ZEKbFAx/b7i7DIHrqQ7Sq+pC5DBEb+jE8gwHgx7
58hJYAiEDpCddvsLP8bXDOLnCw6k35hVwuUZAlxCKbRsDgvVEP+3uYDxHz5BzkiePNZc58IDRvGa
KfN/nnogwyHeA0JeCD5x3ii4mjcUl8HW/426ImhrxLM/5Qqa1AWZ9W4rzovxVQIygzO2z67V0hat
9TgxrBpsr+R4Vm5mokb/ohXdLxVTfuZDqoczmC7kIelPrxyL7Mhfa76PC5buPctPygbmREe3lVMH
0CAEOmH5uB68RndVpEx2QOBWY9xwnUop1a2BkFoPR8XxvaruhvDgIvpmIMyfdIB4ovgGLOAT7HU3
rjT1Luxk+KDi4xS+GrKu8BEnqz2nWxYx1AmAP5nDGmSRAm6oJTSJrYEzQjd5rip55+/iNZfBk2kE
eIcHPcmTBX7HBsp1wgJ2fXt0Vd/w4AkxkJjJtXw00H3gIz7cTsaLYtQkwO9fQMZSwvbRyTxRhUQ3
A7xST861LIvrNvXPT418VtucMgNpERdsXcluqQVS+dOY5pnX7+J3fzB77JNdVO46fy1iEZAgY9Vi
Z+2kHSNMQUSG9F1Bz6S/ZU089DPowDxtSUE6LDIFZn5RWBzotrwuEsaqLlsykD+XrjBkt62kfu3v
HK6IzqtFWhBsRcucu2P8sgZenAHhQHcQC8cMFXWpkQEokJEGXmp8HK7Nq1oY07hSyL9z+IH7qPgm
Lmv5un6N7hHJ68FWkhqT74MDv01wcHXRYAqDs6fI/q4pOOygfBULD1fzhgYQQkQKEphV/G85TVCq
mQZZV3jO87bm+3lJ/K/zh3uU4hU8+mkg1WYsy9e/KQmUfBl7sE3X9N8LqiSYpD0WpM23ViMTzbQ7
PnFIaHxdeP4ikCTLcP14wYAUyRf/m0pF+TKLsF7tj30zuERKl5LnviFG7QC8DYhx9PEgpViKlB3g
lhsLfopbI267VALuksxqY7hMCCY3ArsA57cU4hD/EInMgPnM4vO9Oe3yiZYYTWSQoC93ezIO9e9M
1NrVmM9gi8v8SgrdOdMbJpgLxcxkOehuBDVgVJXeDpElSSrLK4BAqFDEEM5Rspp2cHpry7l9BR4S
RslgisV+6+A/GLaXrih8bZODzz/MABqE75yn7kbxwDNo3ZSIvqpHJV+M+z0PIjM2+FG6/9lr+Hxh
f0/g4ZjgsbuP3yMaHo1yKmsKweTfffaRR7eN176GspvrZFJIqFzko5mI9ZxhH3rPnKAlzsgovL5X
fHv4BupBgdot1axL8suTKBuTYHd4syJRc3QO8BtCMcj65jYfrPPVxGeB2MHW/JuqngRBgH0/SU/f
6okesCwDZdOck4ZE2QdjsIVK3ajbrivpYQaoyDVOt4ereOJE4gBJw/8m9MQ13Ur1sU4l7S+cve55
JnbAgyAwp6VKHEKq25H3oYwFd/nEtqIItLiJ2USsog3BJrIkePczWGfAC3U2VZvyj/a2WHCmIj1M
IBI8pQbMCOn1EER7s5O5V1h5ue7bCoTZSevLJG190cWycMftIXLdF3tdQmRJKLPLjxTA9hAjoKHr
81OqcxrJQxRkhnfyLG+vG9HnulCN5Kdeo/+DNqv447urFqFKt9BQLqrQbQMMKnv/sXxV8GqnlvsR
vs8wXjFVdAEGkXzpAFhlPjR4ZrCcff6IE23AoA1eyuKIChbQ3mcL0XW0or4AFNbbGFw46dERV2S6
9DeIVj0GeYB5Vzamn31RbLpXVTPHckMD7fkbWBHrv6Sa6JAbosBOxRHdX/1x7T1rToXTXPRUpM1d
A+EkawNoLoHoj3T5k13h6mcwjTOds0CNXZJnGa7mDLbeTQwS0GoGMMsCfSQUZP4xC4LEn4JxEF6k
1xPvxUeM/1pnfEtWNNjmYWNffQq8zA7U6MvdquFjMxQn99sMenz+PYDsdpt8vue/b5GXJVZMz8yE
Y3CYw3LpgjNO2sAeaUm6xlLdhfGFIgCNdbwiF/AGcF4dzj7QkIwVzNdPrA9VablAUCaK30ZkNHnE
E6HlJhIFrlesaWK3yRb0KsN3u+GiyTNe9AKG8rKvFtVzhmkKCMoU3wyOgtiMgWMpX4Ygss3teWa6
N1fMZVEfQo0mmaFFyKEm2JwOH9cOO+L9B4Ie+FLw2umBxF0YbpaBV36qNP7RyT0ddjfjZiSoPvGS
TQdWVlEe2A93aCjXGa/IJTu7nt1b2UD1+BOO8ndH5Kn+iDZViDxMd4AurPpw3rKjzzrkqDy040Xm
GhIyJ/5+/t2AGxTmTHB39QHGA6GH+3+zaY4XBv49zNTcWlNYcWuhWr3C6/t1poH3K/1lnrcwW+6a
GADxE4TIL23RsbZMnmDqYycltQtnd/QQjwV218v9h6JNZ8tE9AhnYbxXfHf1rLYSkOwbtzI2wVf7
CHn6NV1kDIJC8HT/5YRa9ZD5Apkk2tE2RdeQu+FkCIKfCphEdiKf154UaAnnH84rHRD040bk0kQX
F01uwlBFGvM8JLHqhUXAsMkGSodbmHiypNrm0XEkP9BeqjifYQ/6IRmR+cei9mlZEdDlPxLjhEZ8
pg5UfnjWpNCNsyunKnYvJgMdrNnLW4iZLn8G5hyOAW0ZEx07JrdwhImi9Kkp0Mjq5Q5zu4ptzhuA
6zDNc8P5plSpXErur45+lv8ZAqRYr9ahiDiX/x6X/Kkt7v54yZRoRQWKzZqfenhJ++kAoOed1iU8
536QUXOxPb54BDJEFETVzEoAm8TCCc3ZFWvgmMgN1gJKvUW5Yt2N5xLbDMoaUlgb9/f6OCOTNbaa
xlgSrq/5L48PNnyXj2VzZKP0C8WDXa8WlMPRaF3VrwQfZS9xZ8lbBJvCWSgqCrw4HSJy5KDMI4wO
Nctqz5T1321E5wKTDQng3j71t+VS9401r4mBVYrgZ2kVqglpthbo0uAoe9estDxcQC3Ospo8Fndv
6Q3ULbmTuXjtFxx1k29erbxT3NPKFUJllVCGfddmL9fVFi5Qsz8AZmAvaScV4fDCg8nhT8W7RR0h
2Z9DIABVp3Lr2zJgs7qTNNaf/uIs7CnIjL6vf6zhbginUWvdJdlnAESYVr2wgZSrW/+wqo1yxND/
HlILdGxG81vk2j2HKalCFyfSg7OsnRP0dWceIMABwDghIvxcBmWbE1kghJb1074CtDA1bOjSXWms
bzz4AGTtIcaRnSpVK/26/6l6Uo9SB4MgtgXFceeNXvvB31JdTfboYoDhModFfSofVheT1sJmjQKc
Vo5ToTzI8bL7wX3Up3C5o7B1cVyCCdhWI97GnCvgyFIBIR6CEqfjhYQI/21IqVBV48uBgoG3jkOj
wf2QslkzrW9p1TkppXLZ6oV1W9oYCT//thcI9q7odK1dOUzy4DfW+UFcpSl4t5tssvQkVmQF6abp
VkphIhR7FzZmcXCwInePwhXO5/2ZwUUqkUX3O1p0t6hiMhVhfwBoGULno77sTE4P5+V8lPkHjZk/
39C91UOstB1IvAaHkxrrMY6deaduovPuP51++50jCS0S6wEjDfEQN5Q5q7x0sYqYavyw/uCiL3Bd
t12D8rhvXbwe1JUszR2IyBFvt7/K0ylk/yLMS+VN5idUAle45eCHMA2a/Qu+tlP9g6ePM1NX1VV9
n+cmDU7e+1KUzRFjF/9e/moEgrzMIhVPU32MiSSVNRA4F/jQziDV3or8kPvJddtllfPcEu1Aho98
WkqeX24GalFYnTaV2sRktKsHRQiLNzSC0pBx1zCNXlb0qUgbeycv2053MpfxtYbzo+4nXcOt8Br+
sddZ2X3fOvYRcItgzTsKQResMgLGUi30ahYFUQxriDwoI0QyU8YpGT9mEQIlMAejjzjj4Ku8bf0u
n4ihwChdcG7yk7VXTxcikM6bsBhaRT6m/z7m8UwT77odxC0mHzp+bErGrPWu+TMghOVsbnwh742u
XBkFVkVY80dOePjmB56iZaSXepyxHmm4chiSL+08INjiS/ursU+tNf/tz9P3zKR6GAuRZfRfC3L3
WcQhMhb3ATPV2puG+mGXOET2U/+POsnx3UjyRX5Zpq0wK1qjOivyBURq7UcVdyLhY8vK8u+r/HDG
qFKR4tvqjlkDC/Ym7Q6TZYoDF8tGDgJMnWeFhB65aAYwQ0/JrtXgeG2CYyoykf0COteNZWdrAVnn
igU4nE+sGUggxYHEHLjpFfSZik0e3XowzohsYiJmCnrznlY1awvQ3h0RMm99KGPd2lN+LJ+RcSDZ
WVOgP7BYB5IeyM9KkilZWmLFxdcWi3rkZm2oSxNQC7RnhnzVH43TDdez6OKz5Rm+c4oMcpGIdchi
nsk+p/vrUt/CQSjawjPv8WRENdJvSmmrBARLpHeFH7eJLt1n/j0knZ9sLqV1exkC4EzmDrnLg1ef
USKj/bQ3m1q4SnJk6OF+ZZAHYsqHwSLo2vAFClx0aclqOROousdHtOOvf7ujTrVhbkHJCuzkdkw3
PwSwsD8GqJ07G78Og8zgoEcSc9JoTvfkHiKDoDgdOGNS8lkkgzFv/pCNDOPyQ7ki9zwP3t1sL5rZ
PES1NRTwOK//F3thXu+zXOmNVzFjHMMubipTjNqsBz6tdP1K+yCENKSVjWokZZb1+v4/VPa89xyc
ske5EtsH9LZ4pKT99BXXVCEFc4Si4n2eUFQhUF1i3udSQlMBQDfNUL9RKy9PGmsIAl3QK5UquVZI
Uv3b91xQkde4JsMAECFbSPeQ/sBNmSOFJxNNzPxfKoAbP+yTTKyB/LxmdpQFR+ML+LUS22ExL+Qc
Du8rAUYZ8aMLGlTmLGGnYkbiZFgTKTmooK8RnA8dMHWdODZU7cctt1Hs2n6G+XOwO/85e5jPPqW9
O83F6l+y+rJvIA9f+a0PQzx6jzN4j6uy1byWCPS1SKS06tQJLRkbFEwnTCWBjjUC7dTqiWh2TUuU
9idP6ICp7jyk1eqNcTSGNT0/7SNMharPVyan9UTi1Qg1eoAcc0Kh3gBzA+QXGwnhVSE9/XVB2pls
iABp/V9WsPafMnH4vcs/ohxdgFNHcwm5seIYjeq5H4BIzXEqcHiZw/TUzTvf/OXwhpWungGUmv88
R/Pjz68jFNAEh5gMprQXco69x+FB3V15WJEGK2w+Js7L7+y+r2szOOKlh0ouizKJn6MXo3h4jFpS
8ysZEMv4ga6g4cLKfprqVc/pcoWz7JeaOrOrsnKKkvavnVCRC3fZ4CC1QskOYM3kyLRCaQedNh/1
hxG5Qkg++8azzH4eREeysXfHhNsuG32WvFvTKi3XmY7I396A+ijcU46rv6xMo//WtsBfBWf7+Rgs
WAyZKY032c9fNS/MyWV44y9HcUihG9QmwP+g5zFOuGeGXlcZ75bd5yo4LlCqE0XhKddAsoW3YRou
uMuoybwoIxMecIneOgHtxuu9hrohWuaIJ90NMkcFt9sSOSXO/XWYXkdoUZxTxJgkdup+KOZcjeoj
KC5f+Sq+s8bXXUZzd13+1pEXn1gxTavcbH9DZZ8hsyetSfMLFo7dtZc0j606FFBjwVDGA+o3Lwww
fse8kxBxEBuicK8emLiPDFwsDrgQkUF9qJ3lTXvjjt/dXdMQX7WjZTD/dvm6w55WGUBxerzAkQlW
0bHRElBBD9/Ppp44DMW11Sy7/B9/3Hb+4UNfpHCeX0RU7R5T4+VFPfkDXkcE/v6JNYzNFrz9WKXw
GWKMrdBkP4VWB95iLoEPavgSAROhpZ4OTu/5yr5EjKhrQDEUUi3HCjYPg+RPfiGxSnPhd0kLgNf5
zBB0SDh0ZbyoeeYdzhZmPfi9cBhpQ8B3SpFoiL+i6VYwW9qOozPXQvY3yghxw/oR5peXK3hb9EkH
kekUDFVNDZV2GJV8V5Q8i1Iq98jwOaojLF7ehtz9QplFCKxMDGKU4FH3he0pqqxvd33/eaa8aG8/
NJbClBklPaJ71eWU1nJlGJ9ETBIt2z5l3rcUIyjDqZCgFso9bbWQk+x0LWW64Oc7KFAujraA9ZZ8
+Y65DkXQpzWW45QfrBWnOGRvcNgnODEdwolSEjqPl7yw+8BX7oyhcosXJlOr9jhbhiFPz6E1RCDp
u3fSEMgSxOwAujk9UBnoLFmSQajJyhGTeO6SyoR6SF1PzUXWV+z9iyRAtOzQ+yLqAL+4dZN3JHF/
tMbpkV3cQ/5a+MidOLdtyBtAqdRrRDOpr/bNAH9bE8eleemqnCh9U/uG/5Abnbes07Ow/V1zxGs5
sNGv2W/Q94zEuMBP5/Jn0/ArRqivUfYd46uovEcCC4cMzKnuHsYj+tTYcE+99hgQcgNjb8xHzZTS
Hm8ywXJqVFBxYnpjbVdSgqzTodCLiJTAjmL+YOv/7ycaamxXFVNolXww+7dxCAbGCJzsozvdhAXa
DhoqlvXJZ9qwibJfDq0i8rCAbTW0Cc2ggqpLLrOxffxqZBiZlDff7MX4MkBD+NMHi87+9eCHqwaE
tBjksG0+iIT9m+V8hZOXGhRGCAaQma5t77gyK465P+bfAnKAKJPn08Eqqetjr9whGlwt+9xuXnXj
/WIukx6mB9A79idQKC3750R3v70WNVxDm9IqKCEQt5Wy63laEq4OA4Yhs11T/1/hA9RA4qgEJxM3
IlYtg2gFEeKVvIb6AEd8c3SPes/GCRVd2AoOsrkByiSesNJK6ko+dEjmlGwJYq9/HahwQWuivNOE
OWbAiiy0B+13/KputJJwSKYg5Ue0+P2PKEALsdS/cQLYaXGhwLUPJfz931iHh6erczXNk+DCQt2g
WNscp23OzFQRVyF9TJ3DBF5H582etHaq8SmvGf7A1/A6xY8PVsm799/xMtbxXZLUU5WXPVgic6rk
tnT9UB8gYnxQJm6CjZn7aIGLKd/F1VmDULtKq/Gtbeiyd+0tWH54SSuH7bF7+/sfb4mkokmRfw3J
2YTZm3YYwxs0FYrJMP02pDD88jPQZHNsPvjmX2K5LMeYkSENoFq92y9JXdKP53j8WmER5v8jPsRz
DldXuQHVdmoTJfZe2/PXnDlyW57H6z+LCGEGwX/QUEbT4kkjV+AFSAM0cRHIWnYn4Iuv0A+NY89/
pW8HRTeElqJwXFYhr6R4tmyu8B1csDUg3VnTvdZs2HhsXfoOMEXXS7tpUZTKZIv+RiJJ6FR9LUX9
vDzVlD91Gh1B+XUZrtNXWqWBO+wy97hypuMo0cvhytCdJupkkNZY8fkpTRzeiGxFmO+60KvpL/RC
nNUz6tZGs6uNCnqxcRlWZB3N/pCcox7sQyhERbty6ndb7ie2ghZeTrDKj6pu6gArLx3aY0TBqCOi
HkoPGbQuvTSjOB5adqN96UegMzBrb6jcY2DL01olBw+Pw7oVtxOvhvadiA0+2wL7OOjrGgJNfonI
3LlSmuHQnrIHSDn0oIk6Cuni0HrNtyhREUiX2BN8KPV5+cJAC+uW0wUtlcmDykACej6sZXar/rqv
CPcO+W178Hu+zlbRjw4vUL7llHmufSVcj1imUt9hTDAI19uBRoyvfpFs7Fx2GeHCSBCnjzxm0Ad+
CNBErJcOw67scMaTU2Z/wBRrL6Qhis3G0iHWgn115WTpv+SuiAmbDwRL/uBKPTLSl7gL8fej0ZTZ
ctynYHTlxN1fYz9psoMHNqjtEwLMmpG39vLBlsC1uAggtvEttaId5+x8871L4wIzzWfPqpelfM/U
0YhCdKl9yZA4e1lSQ3zxKMDAGS9H9MDmCxD6WovwxJ83p9DUpogs1J8UDW6oPNGRPpms5fprWEim
LHWaloWYTkTHCtqFqjY2FZE5GdmOBN73Bv9tIpHX9ikKLynxOuMjndoi1p9Q5BP6f95to8Aap+7a
BphGxXGQan1tLdpCMQQE7Q3FFKUYgaPAJqouRDkPFh4SAfEmsN5gXWXJvehCXHulLo9FTRi5kPE8
hevtgr8VH0MWnO4bbpSso2EpkNGsh3saUTKegk+h/h4WcDiHRTVzE5GQ/gh68Z6u0IEjR6OuZv1D
1nfbtH7bKPFwgu1k45TMFHq8i2wETYfuJtmTz52q2XctU9NB68WQaOAJng++TagrarFr/oMK5wEA
+KFqI/gcXgPZxUZs9xtqH89MTdFBeLaZSPcHdx2j2flD9ouridtf0k7/ICk/RqYHXxjy0O7SiMdu
O6MeTqQFTDu3q4IYHlAQnMmo0ADQPGOgW7SK9iAdqqUDR0buW4XlHh/ygMdkG87bWqQij9lTWouA
58wsp0ehzQhCvwDjxudbLjnsbIVfD0HEBIOkXGjox2MTbjtIo4+6AOdIOicH4k9rDMpGcv5RSrVe
o9MuZGzDOdnTo0eOXcZ9KgbQ+jNq0y9RhxGWrdrPWtsHUsZY1YcCmtn0KvxpWNOw0zC8S1PM20D2
8HCLaU82ktIf9C2UP0yFW/U7tzDm/bDXLzX1+xPIiuUSfCfqbm86z+yuBK1Tw2MVaRjgF1ikanwr
MMo1JjNVaLufAkGISu5W0uO87HTUwlaY+ivhbCTHh/7dySzX/g6xZttPfdMJg2ekJ2/ovNTAB+Zw
RRGlVZm4glubY+pPn6Fu3YVPMaKtF14ZkYN3NZM0FH94kfhE8dkAw3MFGdTq2y1lN+qIXmPYKYWq
z1IsT/uHLLS7zesR5ep/7yN4NrBrS5HwDyFF2w+cwDTaP/BeZnslvK8tE53q6jiF9tVVgMG5bYgq
9xb8cateR1Zr5EpT2wEoGqLe1FycSh1CnbqFPVQd0Y/YH8bpCK4xqLxW1F4glTVEMH9EV4FNxl15
txHrrdljG9J+TMCMz6pXjtbWgtaGOfu+ODQBBTUWFUNQO2N604OqJJS+2v7D715u+TjHEYXPrjxr
C3REJv+Vlx7k3QNbL6l3kjCAM47gCEghec7l0cF5hiQ+65ufKHUtp9hXbeS1LXye58LKWvQHYiGg
ojQp+49GVm3TNsmzpo1PU6IoE1tsNnld4Saq1Fon6+IkAyj6z27xHeU1BawArCLSIT9YGkywOmio
hgW2aD4ZZ2S6UbEgQB+XMM6DqNU0qGxntl9iqrIP3zT59fS5/qtbkU4XweFfHEfpk5Pzh75kyndk
fbEZxKzvxIQ/7TnnnlCivtLJTrpvyeuyBSPUO/aqTWO+naUU5S782ZXmsIDtnusj5TaAkJRORnYK
+SaftX1XRDFex69VEbr0B9zfMx/4RH+frye7WPfnUjLRjVZZcnWD4pSN+9NKujDPFbIq8ITJfAU1
Y2NWYkm7VUbgPyKqUEXnW2csufxi50yHRRgS14Z5LVyuobmqKv9B2yw3P1QQybpbciehhK9mjd5F
j0zZYl/gDBOi4iIcf71Nwarf85eKBxlAjRZLtrmIicpk3OkXFBwEl+0ijd8X8oA1dqht7xoOSOsY
qMgyS+vSksTzeRFWlb20PjU8jiv8G83bzHGzWqMWyl2+XrRAR2+kHDBtFF3AIcm8soYUILlwPukP
i4tMDSFFiNKfmFyEzJ/wqheRjJXkWSxPk6N24P2rRcI7Gh0SmgEFMKb6ck46QsPTeRs1cbi8R9cd
/7OoREMTDwJ27cBBB+vOKEeAGbqyhfVLQ65RccRby3XsyMG9hwdTvHcujrMeKXpvyA/AcZ2HOKmZ
PSLWRUvC1BEXnjGjjCpjnB15KtqKP+n6yijSpazzC8n7DBAr/SN12r/QvARuEoIphjLggsG8unRY
tCQf1Jp5KuCmdzP8Z+2FxJZj3Gd0mC1PuE2Kuoosn1HgfzfhZlorSCxm1EX5UlQRcApDvQyP7/sm
sVNJwpc79CubH4X+Yn0eqARF52bQk4ztnabiUngmdhQbRTFrF0F/x4SRHG8bLeUq+byDWg0+uya9
8stSaMINb+1R6R7XsJrnq1PsNxyy3foa1vEJtEjaQPc8Q3nFWr3cF3qq1YH4u8H8i/LLcO3UyJEK
aRNuC5kbBD4TAhsO5ZJOpA1TkVAGHvZ83sjfOq+1eUHHKi0lgeAz2jwNQaVECRuV5X1RCI7Go6jd
028fCoYDkEncJ0EyEGwBdQxDflEJga4sMnClZ4y6/sJFZOyU5u9zZTMe8poqYe0VphfIoNmWr3/V
qm2M7UYd6Wv4zLhVo+d7Hij5ICmCD5rHgwTprpMP77jeHYo87KOgzL01UUQohjv5mmYAqgMVUUsN
Y+uAzNEqnmbTjFRp6tsWbK/N/E4np2KvIcyub7NqWBntliG0brk5U6QnX+DAlQ5vehmS4sGh98jl
WHaPrs0qidzl/P/J4yyL1t99ql6NaRPjviMOPV7ODEePcalSylGGqy1Dw7bVK/jCEzOVCRYWufF4
Jfm119/PLRESq3OSPlfidUrt0JubgJ33APkHE6KBSaOKUNNHmtqb1zmUE1mZT3HUs5PgXjJmZTk5
XZu4nduCucYI9K4OAAZXbDGPzzHX4EI/v+SQEBBeDtEVam4wuQ5JLirpVQy8jqWqCsHjPIrwwNIV
rK+iEl3wPqOqyfpVYyzSAZbI9gXXJzjn6zuF3QC1jteTn+a4sWxbduhqsWgqB+Zvo0hr1njGoib+
0cqNCHAlpu5/O9aq/baI8TLC1ak+RLHqJ4M/mlMl0XjVOqsnKFDbQT6v5iuCNpy2UmZqjrrJ0vvC
ZsuZRGcbCl4rKKyGECsZjjYNTJWGzUVjeb6EJBoFYZ3+P//Kg1sy3Dk8xFq/ZsZy4pG0YP//Nh3y
w9GlxmUs+IGVU2IYNLMMtYYe4KYjqrDJnpKX9xidoFPFfRTUzm63kfMoWCH4LY9gHX32PFf+87sh
aXS5/KXJ2an4adeTBIy8IEsaodxnlT+mke+YCK4Zhq2R2FWX6Ukiu4e6C6Li1BTcTsbYtvQTUYUF
j1Mf5Ai7j9IY3UAGooZxalMh/KWhDEuUdP+QK8AuZ5zBj+bs1fHz83Wq+7uDx92l9PSEsHUh1Vjw
ApB9NmsAbMa7YxbDNK10Ez5Y9IDrBy96vaTZqNyP77taFuo9cWqvffMVj6BNmYenHc6XGBXt/fhP
Pkyw07ov93LXLQ1m6Zrdj7VsKWHmF4+BsxJQspyn7M0fXJ8CJPoNoBZBGLRWhGBRJsQWAAHQ78Ls
ZZs/aO1YgXWiS/3biTuuQbI/qEg7Gub9HkZaPCppAERJ8r65hE1Ttqc18IEbDPRzheaRPXc3Mn1w
1N0jmP2i+xa0+aIgzXeagC/wlkx9YIX/7/Ou5Q0wiOOfA7cNH52GED4cOwey/H+QC0BzNRUjZeHF
EbPjdWu2RkGRdFrit4yLzZn/oRlFVwRQgJzoKnwDrGkCRz037k9Lpa5wpaqCb06gnNDVkga9c7gz
21rvSgPzXxMznbTbZfRdtoNMbI6D81qls/KF4a3A6tpXf9/YaQ0C4D2oQ/jGJUO5Z1WyAwLGWgFm
TPQLeJqEfm40OG5bF8a/Sbq6zTmbIx5KgG7Vw6bA+Fnx81cwPshnhaCUPHJv9YS+QVAMJcatTMi7
eCXgjyMx+wSrOKMibjTlVBiBRFTQQTjnk5bqMIxtuWvztYl0s40ALjMSebkHjz7fz9eZ446XHCwF
SLoOv9AghmGQsqWuLeeg3u2pKw2ivejtifnrAMIk5E1QqaWqpx49m7EffhUTBYlhd0S8NHnjwlLe
NyWqIv91apnMmnfWqW0w6ps50++aGF/wJ7A7Wa7cenOllyB5qB2pSlqrLs9371qc8n6GmqQI3N7Y
Xrf3PwnYt/6UPqtAE+Nd9gdsf57rzeX1Opzf6gVQM3Y25Mjv/ocJtvLm8Bo6Jt12n7vevPo+i1G1
eWB8Vy9RKs78rEyEKtOhzAmBcAZO6xm7V9NI/wQ77o9S0ai5yy+dhFrkv9le2p59AcTgyGkXhGny
oZAvZ4CpMJQGv7OhKSEcPeSdcoUW2VCb7IqMvK7u2hKo567KZT/E71T/Ys/XF7QE25s6L6THEzoG
2HNGBLa6kdgLbRs7+3OBnwOxjCvs6pq7HBzxE616sfIh9Qzo1wDYFjwowXH8mZQ9ZYXVuWEekjGh
eHALXt/Vot6Xt4e6P2/Ge4/7kiPrwIRt4pOyUaaTMN5q/zim4Cvocl6VN5YBpQvcGx4UxLitFnjf
UhnDsZYmVI2iDSlTvZnVL1F4EtZ8IxkMKqjgRhlQ5bcdZTzxOm8bKH0QLtuf/6PRo5vaZqTdfl70
cOhqvqp+v3MGixeH83XuGzb5k68Mfav//N5dBwu6qXYTwh4m7I16dbmtV+korE0M8Il8ejnW3o/W
zr+wMoxACoVLCKam/rfJCuJXOuyGmDtTzgsLx7o9rp3slt+eLDB6umTtRjNspmHMFbqDUsTgJioV
7HujU9zD+iczgGsieafvyJ6AMSUv9CHPaNa+mvGXuUxPnjYhttQ1U41tcd2wlio7GOEH0Ce64ZIR
KfYoQpAm6I0tz+znmjIltNAJzufW7lVX3yzbIf5OmCUiCsYN43l4m0mMcRBLxbMxlOM0vAx1Qu1P
GROhJCCsHc9TfgCQoHvIMC2nGXSweIHfjoV95K2ZYECyGwB8JyTF84vdwXADNCbQHE3Eg9E1beon
1AFD6vyCKm0pi1E1PZUfVADYmI8+Y4+Wb6sNduc6Py/SDxLrN3BzJoKLiaLOETxZoDw2xb2in8ZP
PLkUAQakQ/dzpwPUZSq8vEpEzTGxxaYBjvnEUVIeYK952nsjQ/UWuO1tWolcZ6qXp40IeAhip3WV
MfdBiY51m4KpPVnNvoWqx212RvB+fDkzjD6TfHkIJXdXku48lcPEgTpxfcddn6QZDWHfoOjfPJEy
jlxIBUxYYAoocX/0AoaXGuDX0zrDk12ppSaVQ65ZaMk6R/fpOoOMIQkSHX4yFXTwCvbgBS6rGdOT
s8womFunoY88VcX2PwgBBk4lg0fUd1AkZchtp4UcJpJAHWA3yW7ae5NZreqhmvIPsEG76P94xhrx
Cmm4sc6ILSK4dbIMjJRVd59EdREzwK1j8H+k8OyGBLPrvEAQgNYGzPTZI21BbVVTz1n2BYVdqi12
wCErmVlhUWARwPpfX1Fm2TbyUdOzXCV24AnybEQoZAsM2I0fO3SDsLeAJ/KyOwjw0K8zsJ+FrPXI
keu0bE7wuHnc6ItQJTWtIEDeHSZIWFUzqXVd9RS3p5eNGAHn4CHEVuZVQ7UAjU3uRSGwJN2iPEkn
aZCZFrE+PA5rkr2pgFWYGhEx/uva7CYbWniLezvgsdt3Q5zh6znhYNhmovGXujTesIl8Eifaj+BA
et9cZbPHA15TVULoghjkLKIBEvj+d9TQgJzp3eyRij52yYV038D8vrf1vKQozfvZJHkPuFsWP5Sw
JUVSXcq5uPxODqCmVb6GQnRl7qjm64yrJMPe6AAMh4QJJs2lDavPGoy8fG9QZSavDtTf6hT1qPc5
OHQRU1zgCtlbIje8Mm0Zbiw7sfA55JCSSiFFVKCwS8mBCSVHkb9BDscYhls9Y/0habkPmMjR6l0s
i8Df4hobVlaVg1CO0wGz/2vEIRegFeBnuw2Q6O9jKdhGP3nnBRY+aJFZqZJ8ETKbUZZM8v4lV2ow
eONDz/PQNJ/Nh3bZDmtEMH+NIM+0rq5Bs5XqRmpO4UGuLRgZcHxcPTW0FvCl+PYfuvQ5IFaO3O+b
2nUN++02OKLizgTrMKMO+NdF3LjiRJsczVU+LcYXwbka/WoyueRIxSpndZ72s2n4C0dEkm90SqZI
GxBZJBFRcw+1Z+Y2GkDtLoIRU/nMxS4du83tCdBGSbMdnsAvgyHTa1mYJuIjCUNYKk9/BpnPQFlX
SHXD1xj+0UrMY9i9x87CZDF5YZqJXdMZguFIBSsW9xsg7hKED2w5LpVAJKehokMHS/fHkY9O5F4j
pdQa/kSOJFTxc1C3zVVs1Ck8G++KA5qvCzPPmhC6A6alHVgcQIgoGV5mcHwgNyDSyWhPP8VdDEZd
Zc5ILyOxxQvLZkNrxG6wkIV73r2OJMoTAd1vrBSyeZb5MU2YgAYb0OZEKMUlISCdFqgLp/m58Apg
V6RMCuv5U2ucTyQAFGBYj6pOHdDsU5y4OzalC+bSb0iSj8XWkIVnBfdWdZaFBCJ8KttALJyYaJ3W
KR4PObAlN5B7xr8DdpI3TsPVDigVnitR6iw67R5TYibYQG03qx2iPuPaUBhuI4AmkyG/jDE2cypQ
UGtIwa+VFfTuRk9KIaEFZhQL/JIf9EXcNvLsfDGRNlZ86nq+S07ks8zvi3kf32Dx9PPCCDONtxWh
DiLuig87hCIknF5gh/OSyOZw9HMgvQ3uzLgL09rInabgMYwP33AR2krNfKcxhFXqBLsTdljHhZoN
VHqc89oBO6vt7Z3rzbmK3Jub5CjeB5ykCRTCDPHpo61VF6dv9Ih/xQJNbr40wz8gl+cpyHc208iV
WtXGgBzhF4HotKNhnADbwLAtvYgFeETT9mXvBgpEQO8ld2UkCXwMPrsqsbPkGQruqEDmlNq0Q29P
ZfuWA4Xcfb/wYw7IH4nPLaltMCnrmVvKwxeAd8AUEFjYi0Pz52eqDYtu4zsmXeysrWmCqfbDeLPo
dvldiViB9O1P111veo/rdrlucdqml/Ks7Zs6pz4tvSmWfOmXAQcTZsuvlmHXURse0dAW1HT5o91K
DUOH01o0IxYTl/fCG+5lOnuyZBQr8EtaN16L/iTXoFrcqNiiBHb34H6vpSBEVAKtVv1pb6jmI3M7
eed1l+MgCT6FKKibZnw0W+FIACmQLD74y6BqzWvChgMfpVcWPYnY5TScR+ofYPJjnBeYJ7jXvbS6
0EIQJ+4j7OPZvNF46tJsqgRiW2s8L9/Oeqzr9xB+mP9oVAHb4rw/hn0lABVl8Tt4idAM7CEOdtI5
4IwAO42UmPrcbU+R0QR+d7pyf0XlCZJYikjJU762WzsqhNnf24zHX6SxDcIWiyWYwPchKPhUVQki
UtgDMieGnBtT+E9Dd57iwXihMUX1aeZkUAhIENnuptIizko1MkEB04RqHs+iMYzq+lg/zbWFnwMp
WGatp0aQ04qTRhr7b0AzEnmyryuROdPh2VN7EW7PQ4jAZAskBFcAj/P7efDb2+S5B0QHL3C/BONx
lx5XicEFKsfq4pWGoxpYkbS0PamtXjgxeHPq5YerBpnkhL7hwjw7r9iKvapOe5vybPpEeaGuiCgV
TJdDv+rMqh/mLwOVpYGUGh9NxiKZN/zBsgLwp+GY+yyyzlMoKI11qZX3hVG2dctu3ojA5ewCgrnT
hj/SXkKKuscClxcF2SyWNlSGVT3yKHUmvj9iR4Q69tHTgwoEMtsXg2o1WZTx7IURhTGIGk1lhrSo
jnK67yVXDlaAbLyQcYnMv26KtkAs7BQWwNDM9jsAI3H+bdrJ6uMn7CGEwR8anp38K/ypJkx4bSLj
GdqVeeiCoWxjwzwM0vxGoZzWsjxeoUjXj8DksvATJxb+wV7re9SZYhRiepe6VHm3xsto6ziesYKB
GIbBxZGtZl5Aq+BwYfIDvGBpjWlMFrLH7F2jdXs3zFzwL2c+XUslbehnIGZkOAEcOOwIhOJ/Ex0X
kwW96tyXEhjuPd26W4KcdtMYN+/76G0/CTngQp71xrwfpW6B8EiyUU4zNjI5IIf/RC246WJoCEJu
76NxVXOQmJr6ifKxQvEp0/WtLjQkxpjtzZhwlvK0EUi+x6hDvDzPypCRdOwxdkqhS29hTrOskTzW
78sVMlEQ4C+JGy1Ax9hHlnpc12+SL5+d+uQ3CqW6/5HyR9UP2DNzG/98wyEaTh4HAdS5iIJdCJ/r
PKtMinx66B10F1ZUzUnK22aI0XuMiDv381XA1luybx+3SvP0OqoHlKjsPvNxfa8mZsJUyrwtWvfB
TvjiaI9Qi+Yh50m8frMfO12tpCRkUXR53NPra9l06B4rFi+ZavfZaRwc/AHmfODEADLz+mwRjKQU
Qt7Ho9/mT+uCFo6deIbRJ20qdqQpl9azlXX5LQRzVPvxQq0FoLJuYcfc31BhXa8fCaXDn9othwev
QA5szF/HlGgAdHMfciLq3IPXAfQap5Brjq1vVtpvy9rphQBq3KiQ2tLU/k3tIdfFrzQJhxOY5NTq
RukuRNSuHg0leo7c5sMlIvXsnN1fDabzy0H5cLLeqfE+jomNP9NCVUTBzHHIZ3GkLGweQEmcAoI9
jzEXg9tUWJKX1pLaMb+TzhLVYIZaTOqq9+WU+guuWsol/RnwCMfPrcuFEWoHAGcPMDNumys6HAaI
p5AMMFlc05V0YVlCLhluKffsyihB/pk3CEVlXZ7pVriRv4cs21fOUYj8Q136vbVHMLaEz1ewAyXm
VIPXrDNwVQ2VevGFnWUro57EkfLseHmqQSLJSWTap5BlmL3VMweH7dV/B2qaWEBVmMwu9f+EY5al
hfXh9a4rf9jtKb40l/IYtnYV9Oxufdb4tkjNDwkxqoZKuxH1dJRlWnW+1aDFn9+eTjuOrzotfL5d
CBqX17scW9HsT7Uc3boBg6Kb7it7Ad3H3zv+47LMXWu7vx2gL2WY9+2rY40OqP4RemlPw+4prvvD
7gzZZkYDfWE7sgyaXTsIm0vBs+PhRCJCCbbreX0do1jdJzj54+CcLyB6eW+0V2Gp4hDlgS4JoWvZ
EvLF9dQrpjqTDQwpA+kNkWdzPmnsi4nRUieaUNZxkBzDbAovQkKWuY1HtJtDEiV2Nu9aqvJ87Yi4
VgOGmuQDEkkq3Xe0yWgFbnIA7l5qn1MEmfHw7Y6czK+SVqglI8lIT+i1oQwo9tW/v0+zM336uYHc
KYQj/GJ6FVb0IKOS4nPjJklj/iClNiWa/VI99IovMTr4nv0S2Xf7WLtp7bq6zzv/y7wh6k6T8JD4
SXy2rsh3i1XUXThUByKYubdeqQhQMNH7IyVxoBkrYeeCf32WfXZFaeYIIznYSRAjhmM5NdwQlDim
TY4BCBOz5jC5eqIrItqCBu6Bz1Qn2UY3B3R28b96jWTt8fB9dONHDhFh6A/FmD0f1R9Lile/TFI2
+shqwb0BbAdljZWpGnrWf58/rpIEiaU3pDyBByceYG+wrvPwuq4Jno6hueg6ZXhhZAfGGCMSbsjy
zEps5B/S4qWXaMjpcH7CJ8Ae0IEhhA5ybWkCXBXhhq6V1wmmv5hx6Me92XS0qCQzM+aeJ6AtTAfy
9ZZsRaCVOGR0XRYYfzJbsb7a1V5ATdbKPIygS4qi+pWmZd+5UzFfGg3o2CC9s7tEATC2V8aPotRF
Gp/ZykentDStLW15WOa27SNU7zx+L7LuwofiMaErn7vodmyeVPnLjDMG+KTfEQfjCG7XIvCuseTP
LFC7Ige+3IC7+PZJQXnp+vAC4Hioi3LzT6kB/fXwmuqn3hGg2qD6ie+HChCmfNG/ue2Hl1rriY+g
nB4rTbcIhiQa0tuz7s2voNTc7kfXrnzFuCHe2oeIHqXVTJK87idJJOY4eRVPGd+879RLLc9k03+f
AVE0oWZ996VYt4W9eNuVvwvBVFfUr+f7Ovqo6PalyndN4Vot2D+/QL3Qw8S1j+1Jc3gCBB/SSSBc
NRfCQrFa8RRUDaZ2zEzmpqBJHIVBgwxy5PxZfRP8c3DvFcpk8i3nHdlvnYAPfEWiUOjFLONSgPHW
EWfS9LnfTayuZGuJ3JChRphVbmdwVVNe7cz3IZINAyHx28tUWXkaLIt5wGkNL/cmBFzPBunXVRf+
gznQnpmhUp8kPuLPQsX17HNxYZOiNStJE/WvbysLRV5Of14nlQF65T7cnz5xpQOLBTTbOcsTr3bM
85+PiWYolQMSbVvgun54QR+OHleR8bjDRIbUm8qR+jKD+9h3lD0OVsdzB404seaG8pWhmtERpI/V
ZqNYHn0xn2J3XEeztAGEp+hfdznack4gI8TUX5fxxPznkmO5gjyy5IWdGcwuaqVkBXy4h2qTD9e2
OpZ6VnBTvajxxvbSgoBjANLaZ76oNBrqxPzVYo4Qswpu6gNmkB7ZKsLK98WKcb0AheUGuGd58oAa
If8ZXlezq/yxe6jqf2F38yev/OPgIsFRsjU1HZSDNdztd0wN7TYrmX6NCPBIQvRSq4SbaG3CJehV
tq9hIPZzHIUSdw36xt+knNzFuwPYVXezfjgCVAXvo8t8mXCw87KneGPz+nZk4SdIQwIE5Qm9dbYY
ftwjDEALcg0LTjEv0fbo8uPVEHHGeTcF+fW2AKhLtNX6iPPX4pORdH0d6XyDLYI7o94bx8DdVpMQ
1ObxLM7IE5BGwHfcuF3YYwhDR5HCt6hQCnDF4pWRRbEeuCjcMxH9I8g9sZpbXTt0A9Pe0A+Yh8jx
f8aG2Dmew/3kaDEiXbeZVCi3YSk2C3YzW+YL4hzkprDX/wGTBHrDsFXq4Q5LrWbujO1zqqYGRTXw
KXRJreJYcn1kCw9+KSdWwvOEZP7PVwbQXZCNxlRHirZw4GPYR2HHjbDOVoS0GIvdNU2Ti6V8Rl2D
HrAgGCJ5P2LD10BzyAKnxFsEEQVeQ8OkWXJ9DgBgOuw9I8hoTGe33z/3dgEliD5VKW5zxmDHvyXT
z1oqYigPmpWeR+kJ2BsEORuaeJQZqaZt0gWS9VoCu9xeODtF9pnzfJnDkxiAKYBmtIdFDG0lhcPV
UnzDfpufNiSEG9YMm8d9gsG0HfYS34n2MdpZD6VbpS7dQ+aQkPgYEh3nIgZYCSv888LuOtd2q9fK
GNGst8UF1tLpZxzvgSu5vP+/bZbtx0JvdS2aicGzbK8KigQrIhU7QycJQZr5+Sv5Cnw+1W4hnLh6
KDxzFG8URFnW38TjRzXOVEIhtRHM+5lUQ9uE7dla6AIlUJRtGWokb8+dRdGrGSm7CPB7R91tyQf8
VKUhcVgBs+o6AYHCJ+VqLoNJ5D+Vq5/rqr/e2mnlnr5AOLhSK/jA6TdtIGr0Tr084bQk6FfETQll
YdQWR8KtJEY0z4ryfoCPT//JaCUak/HQx/bljgtdlXgxHjdiqo3T5WlWRpl60hOioiznuaSIvw2Q
42+AR+qSSZ7110bltxt359b2YheQUegiXvJ1My0HK9t3tsBuav3REKyV8mrYjSHlP5srGzIiEhL7
wTFaYI96JiF4Nn4dI9xzD5QUPUYLXawT7Q4vD1tcYrq4MRKqFxlbkmXk+u4qvot7fxzYIHCG4Tvu
yhKURtNPVtxh0BboG2T/fWHlpPuHSEY/hSWnPXrgITz97/J72xh3/4GyvH1/KyR9z5Smti5PGDmp
ReDOyjUhtozqFxmzVWpRtsNFw6uSXbOcxCaBnAFE+4f/GbOmLVy5x8g3pkpCJ7pH2tNf421ph+9V
K8AYOHvWVRl2l3+D/EoItYzt0pNPzv+kH4efQSyy/0Wl1m3FePrHinKNDv8yUanu3GfULF+URsda
A7YAMRq8ZkycobQqYgRoBijGvvyTFVNwr2TufeP7D0ZukfnMGlSe74/Tybfn8w54kduhh/AiNJcK
SCTKE8BSK2gTy0QBS3oQV5nBNsMKlQEQ9/HaDWEoURJTg7mUk6T1pLBiT8aMAzESSueXfBS6bVk5
Oek9Uieeywj0Wcntz5RJ6olwrMCh6g2cataVxUEMnTfjAbWz36kiZhFU7Zza24UMKdohHv88lrqq
x2Y5bW8DXuC3t/YA6V1uy057LBlm2qPamkkybM7xYnhgzxMTMTNWzjIEaIcMlOm9PSH/uUaEMSHa
MRkqJx6mmU+A8xJdvYqYcSJ4WRm2G03tWFNE/zrwOWA/VCyIkJQbqb0Cs0fwHm+xzO9mCJIDtnm7
aVlZ4FDouyPG5KGt3ODf7r7VXQ483mXjIQPAr+5BRjm8iNNsCWBCLxXEm3lLnBQTfSsCQwnb19BQ
12JZh6q62FJmnpmAgF4tp3cc39lAudwDdVeIwnvew89og6u8jGuh0Vp57UWa7uyUWFgN/NN0GoCF
XsLcfAlzlCU6lRZbCCUXhnp6RSJVUmgoZUuOBJ9NQBglXFipX+J+975wQJMEhClx2ZVCdzA3zii0
5FJjKWRqXpFwbXSidfQbLXDxOWJ5ry1MmNt8qAC2KRx6tOVdYsEHB9JRtVLH0Gu/e7cO9VxHK8z2
7s5RbZ8uVCHzwWDdMnKh6KMLiUaJIeBlFDO26gSlUZz8FJkbVeMp8Dd9gJ3oPlL20Y5yr5UudHHY
tF6yk4jyC6G2NRKP+cFkHRdfJD2/cLgd5/0YmF79auN4vbUTWWGVvwfwFOPXZ/oMju0lO3wX2ZHU
uOKRs1PNrjZfJe3zC66pZnw0mNC/DoxHRvts5OsqFSYlH3pXypFnNCf444At9tAMb2vbwA+fWxhj
2r0qhYK8VfPxNhupX/bkoPnNxvFAc0qoWzmendHA0BjOzMXSUG4K7x/zyvk8umHp0QOWNgOlIKfC
KDaQMPSEY5rnLkMtKZjqBhCtWlajtLtYPDw2zNUZS6aRRZWQ9vvY+NMGsoHXOzWfGeu56dOfNWNN
0uSV4aGYPHBLfb7ocHMOJ4QSAHQJGnkB5ec5yPuF/hr7z8iWD3qKidxPapJW8LJoeb33CAD7mUTt
QHjUUv26pPZuRiRqyyaJ0DHsWBj40dgVCoCjsZYpxqIW70jJgUK/2laUD5LGp9DpySXrl6/20sAU
M708fGtRqyROemuwo1e7P5acu1IYtzheGqHdANlMmc6Zf3Y1EG7lo3YI5q/YmkF8yFwSnpdqRBdv
Lc+H38KTIkHKwe2Peke0flsY1t2CHcYsUKBTPMyH8NT2FBtSXfr6VNumav2O/bMroNbXtC9Hin55
JxcTfhy4lqDHFqHW1BgL6pBYVAtXFGn3WcTMsZxNunQ20xowfu3PyQqG75S3964H1cVtsGzQamRM
Cd6o3ubTH9nWM9JBWiP/Z/q0ZwmLH65Xwzcqc9A/Pr2uqTBoU4auzJHK8gEF3GApmwrjz94XWNWB
fqu2G2EA1uQxF/d6q0sWSAJBPJMepFiml224MuCN0TmEiRgEXbmrpBxgkGCKuwc0HIpLM7tu80g7
mqPUjrQbvKrOjJwuN2OhroN7HBg5Vjofq6onvgCn3feTsCzq4YKmqHgZiFUQaUkKslbQWl0KibCb
UOZblW34ruFaRerbBkLHe82d7XNssIJXJnKMq4L5XUsOlV8qlwIdLK+wG3WfuNo9mnvxxPlsIR//
s6/S7sckcN7zRMa0iVZUCA2BwG9EAvJq9e60rYIBJTW0dkKFEI4z+BcPtVMvub1q18pVv2tPAafD
pekcr/PSi5oBXKOg+/IV2Bl34N4uqt1amoNMIKHKRKvPebkO9ReyljhVqF4g2S9sWYxj2VrUhZ7A
sTYhfKP4qLIeXScSbqu/qxUlwjm1ihlUWz9WUChTtzMAZkpp3Hv+fJmKrtDe7zpVXXtd79sZlg47
TgVcE/KEWalyz+z9H8umA9uksXciUxPpt6QsauPi81cumMdHRjHO6owEl/BwGK7+XKS/XeKzYKtA
/R15F+zFBlmiozVbEf3xf/jKWI7E9F7jyq1O/oe+yjMKqEC28HXVYE+cXybuYZtHiXw+CAg2Udgl
GX9lfTfZTB7YnVPu6X9GpMyv0dY01TRIhJ6EaWSffdHdalo5Tcdndf4ML91x66WQWE7Wiygvz+6Z
kvYIXK3/S7+GhV9YLsjhNMQPHeToAGdc9LpAzvnSatVYgz+bIPdEF4Yhpl9Tpd+bjxSyIdmCIjrX
WW791lCDdeQpOXnaBHdUAPIf1TUR/ntPGOuh3VTXRbNKvGi4cbmX04zpqJCUf5N/O6YbvGmYSXr3
FO+vZwdrXBcLlNNtMuWkLulIgN4wrbvyHy0qqJxv3TSDypt8ERqskNd5MAtlOn56NPLnSOYIKlm5
465djYkAoKaHpJI/YoeH6A0MBj+DTktHTNdSkMAFowZgARGg1/QZiS32Zh85/LVLLt9haU7Sp4NB
Z25Hm54Yj2gTJ548okA9XOaSMQcs7MzUZDWnaVKiierD9lX1Ql6mDfxAC/wd+tP1doZxJF2e9eUM
HkOuI1h0JEaNZOdbIPkA0XrBOjcUfearxazptDaCKeUqEdtLCieYLd3E+etGPpqri+Xsg0EtxgLe
3CrCApBwqeBWBDeXfY2xg5E81SJ5SLWH6dV4pLwvCkNpMSboAQhzGn1FngTBRnitOH5k1RmPG1RY
iZValRg9D+biZxr7pJGcK7k0remPGO6VI2uYzb4oxfign+jCtiBslzNbqlbYVNzKPp+Z8c0HEBsq
pOaMxp9EQ6AkuTYJqqwLOq5CYfjAiHvzux4EcNSlav6+tdJCYsgoVI3/Hsk5gaH5HoLwgNdhsBxG
Vk1uGUgkX2QBoKEDCjgYk/UqYd/lUgUsGSb/AaVIpJgVI2Nw/Zmwnj7wofUnSyS/WFlduIytUyjn
1vcXkwyeMz95VDdsCmd/jZ90MZbtvjdr3Rntb+fUTop5u/sK+le/6SiuBy7w4DCffYwR7cN1Uh+8
4bIfw+M6IfCdQLoWjYT6N3HgdhNQ0s5yaCdA/3BtTt0FeZzBnO9FUo2udvAmoIrjvfSaRAadsReU
vBlmR/38aS6JXKswD2kkZ822C+PWHxBEioQ998v/tuqgdERT16ThD09z/2xuWjS4rIi1gRfl2aNc
nySZ39km82+pcApvzE11v0GzYQi7ubmQochpxKEXJRHLcT/xU1IryUxMfM7tWl8X+PHuG8BNnjDf
MCWCRtTozq12k6QuEvz0gUKmzi9Y1ciSogZJJ11uT/6nYXujk7YYRs207GvzeD97kW4+j8cwqsSI
yw38VW+0NMvoh882/uFZ82EdiBs2Ntx6vAQCEWkvbH+xAWyO1VRVJxiytx9C27hQ7mEELuQJM1fB
z4+rQ10V58EDIN55gcxbP59/RGhUh4OUy9HCY3WPa2E7aYgU0/ZIdDhF0XwDvWKeEjJ0Xal/nAQW
FA9F8tHnFSqJyFY/fjFU+Cq1EcUmxELCGPw4wfkcSqcpqaCLtW7NNz0w5HpNnq5wkAezZbkboEt4
uZbl027t0KMP4BZzF357KIzaF9D6T3ZA8QxEW9dTbaCq4SQJM2xUJ1cPRqbTMGyqwh7Xopp02dkL
j6pGRlcWlaDMi9Z1TXb+vvDd9aadkwcb7VWT4oAr+pYE2nhQuPF5Z6O4UM2XOTsEiqQjWItUopk+
0iBfSTg5L9lkcE5Y7EAHbZTu4lKIZ5zSqW1QgLbElJ4GmktyJBarympL9w6nTvhUTzZNVPdwmC1L
FQlxeJ84Ti0zV14pvKIYGM53fpTi9uMwValJHBj9tXRCsga3DeHcuVmmenytj8CVL/rpUdJB/8ad
wsRlYdpKqMZb6tkxOyjEVLXSXgflhFp5PxUKJS24P70+7fVkFXupY8STq3cHnvi6IQzTPrOSS6Ht
BedGKE5v6VC9CIImGGwKZ71Q/XR1B9t2vR49l9MM2LugmKU4nh64Etg6/fViY2YFpG/BkLdvq8OV
Knoz8tyndF97PIVT9eTCKysCHIT1z6VH2xMuql/LvTNBlAAdt9movpRq8u+imVgr4yVfkrJJZUyN
1oueOvQ03LwZqfx1Mf+L1qg8wJHYvEKe9huwDB1hcEOAYY/tmIEFAs8EFvPb4NpI2w0HxSmXavTz
Gngm9q376+gHwGvs/5mEgxKvCTQky/ZY54DyzEDIJ0i5cW6Wru+5hXR9/D1Ii11IJGSFW+Pr4E6c
JhMQP02MpeTog2rEQTlD+Mn3UHNZJy+VmrqoDrKT7cnsBjNbm+ZxMK6f2RiOoS8V8ufLDY+O/FoR
6ANo/t4kaDdnNzY0SekHdC0OfOifjYtfB7NR/2aH7uHwsjRjDpah7iY2HRQj+8Z7lpxpkgohZyHz
KcYET74mT3DPhjkqPhH2wPVxqdXzFmNyQfyJZKjw3Dc8u8jw0hsF3g8cufi6p1Y/h0Wd0nurF1Eg
VDpNHQZS0mD8FTqEijfxq8rFiW0nhBMuOaKdAYwbp26OnTwqZLBkR4SEdHWQ+79SjXQPSTyu0VR6
ETAJb0VLmynfMeWVWALuudCzPdjrDhu4URYKm2mutE5WkOttMxOpHX5MxiwWkX0nCf7eQOtuWbGd
oZBk6j2VHxhzx4Fm4UVP8Cbpsv8zBkythq0p9UC71FCnxOZfrg/OAoUjXH1TRXORf9znL1+uaITW
nlD1eKH6GkaEVPfJYt6DXmGqPbSpTBE/hWg1TwK4Zc4O2Fy7wD9nBRZ8GVnAye2WaLqLCR/ClRFL
S1L9Q1FNnpsKFrSPlD6bnlq0GX9vL42deQu/hsyJ3u8KiiM0TbNPI94o3Vq9K1G8znJNDOTvA5zz
hSh02VX3US96I2RH1qcs4IxkDtASfM4vM3OKgCG6PxqPuWcKMdmgxbYSwIyPLtJw/qBXXuS+ZixM
0vj6CTXdkBGG69wG4IwW8xV7Csav27jBGRt+/N+ShZqIEj29b1ctUZj6qIwclSYPCUWGkdD3qI2A
VVjRrMflL/W5bqX2FHG9B9nCQfMkEyt+c9pGmr6T51eyaeCRDiltQdubX8HCdDV2o98T2WWoSCv8
O8dIG6DSNPynGtA5O3xtwQwaFrSJYVyO75zt9hIEtiramc235ppeivqmbH0KFEDi299vBwMKp2Zw
c9DhbuoA8O2naHcnR8eB73OcGjCAcUBc+JyOy/gS364OlLE/K6eF3J93GQegqtUqEqykPAUw0z6i
ybFRa4D48lKEO4e2u9tbEC3NQYDLTGHOB/8tY1tkGk1/9xSA7CShIug20S2dppNIKi20mCJ7EnLa
/uH/6g6XppVDXpADqfyF9Ltgcq3qCMXE8ZoCcPNo/9Yq3wZ+MaOzeilw1JQmLp98Xm+kYU4iYigU
WJTV0W7xF73W5cWSSzD+bWd5piF/WJjulJgkbjKkeSgNKflxlDrqgbn1aO36+Dgp7wZeQ6WEyvN3
AgNiz5K39o8nrgCwo0CY5lS3ggheougk7+cRROacO5wIAco2PV7g04BMj6mG5hFOBnLuWe2ADN5d
fmAZVwgTmdP8eTqmDBgcdE6AEDeQMs5D/+1O/HMxGR2+70zhDMwwhHMbM+Vml4/mK6pBI2JL+iMO
qDaz3v9zI6SzN29eP7zqqGNymmw9b1l5MxINrzupVcytzforKZkWvlwtrs8q/cUHXEYT5aO+YLYg
VqB3r4X1+TQo434Jy4AH+2Fy5PLfuGnzn/a0R/YcUs8pnkrERsw1cJgKfRt/aSKKD1cyeixNCX2I
Gg6K+vo6eEKZvp+MB/w2WA0VofCQ/2Qst8FxA55zuacTPTEbt4DaC8GevghlodUk9n+bsjbmNLyG
h9JK4TZBKvFR98e4ih7BwReVs8Uy6q8owt6EvRttjeIQxNk+68wysbBQ91VmoQcHWAZKf7JxKnZM
C8I91I/NP0d5WUkMzjexpGW9q9/jTtiU06P07m+gJrUNTqi5N9HE9cU1mq3hNIu/SY4n+RXSRvR4
DqTs0CcxnkV1atNYA9XKToaTX+wqEVnEqeBeDrWzRTj1JNxt5OYaWs5i3HQNsasrXvIfc725k5Jc
ONZSUZ/aOqZunwwel8P7/TmChaFP7sOvyEpXoF2eITWKlSwFUr51PLD+HSdgn3jDuCPmTabfgUWH
t2BfH27INHMtfJPoHSWXnvVxMub48GJ0myHNedUic9fJdT5t3Z6DQ4Dtz64WcF6hItGYKggVlzEY
GqOo93LEa+Wmwh74/CNLaslXHtbeh2oTercBKH2F+fr2PmyAQuWuS4jWhnr8dnHa2BojShv051xH
cn1Jc83m1HhDnidQEBiB3OUnUI6g4M+qQU8GKMavAfqx5jmryMpYNj4SnpH2qdt0DtAb5BOPD+Fb
GSeP2geHqSIs9EaVT7CIi+JnEMkpt6TfX0vXwRPbf8yIklxtaFhB5VwDv+sHDPbvu3mSdMkX4Ah7
FIFCJ6jq5jutoRrzsO+lbVQguplbPKhzv62z/nDQH4M40nEATmBceupeQDQqumX/sZo5TaxWtpq1
2sS6p1Gw+24XKI3wBwfDhf1avmcRAJH7dGWQx4Iczr9Nm8JxmJ09gwvkAovhUkqDP+62Kp5YXegJ
E+h6uV2SOSBLrubpOLzABqgkb5Yd4C0Z95wFD+wu72rxdheo9M5HqkrfrUzjtRvRn3oEjM3h+Jos
SwMsq9xdGPibeJvPgeLydwSZSKjwjrn2aQNxsez0j1vM1YKsM/RwRISNsAPRuk+EnH5R8YgxOzBe
EptUDrAmOgfXKlfgS0TCXldoIESVwppB
%%% protect end_protected
