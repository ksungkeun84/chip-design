%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
DQNv5LJZ9VJxnt96+1nQCehF5vs+olft15NM/O8hHX5CCQH8sQzuZCQqG1HJFJnLs2Eh/I8dtQYj
qJBh7JGPWIdI5JmJ3/27WTB8wHUpZGQfhs0A7g6CLt9mMV3R/OlPie5H73WaQmAV9vDlnQufbW5d
ISAN5ELe2ZEt5yhxM5AFnyiJeVTgZ2T79W4tGLmLQgAsdZccmXFGjx4zvqpyhlGT1L4kRjkpz2E/
eO0lSe257d8slED7/EZs5lACLyCdLD+h3uiaBlnXNZUq5ckpddU5YwcznJURNWb03tTmwlo0JupG
K7bk/1YqrWHwbYHZxqSk/zydOzMehheBH6CrxA==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
Vn9ntUefhJagGHu8qmKflZzgToFxVdVETAOMY+q5RCYcRBixWC4qLCP1N950cLlE2OkfVuT8VuS7
nSq9WVaRjPmXxF7i+JpBTlhxVkA3DLVqj4MiO4zCZGaEhXi2LiRHEqLp0wVQBkx8Z+9iskj/VK2/
aVd1Bx9gIBI3/Q1Iu1lQsiWngBs67XoiM3xSKQ98qd4l6Gzi0zp8JnRjO2kN+PQ/BX30HaPAl7p3
KXcaoYK48KPeZe5HnYRCso7XBZvPZbkS1dQ1xONv4a2ViVWy2aC73up5pIOtJ6YJ2dc2lThAkpLz
C9c0J9vW6AMP6i90zxjYrL3YIWBlH5OxVgiKUoVW6wPjPMoPMq1ViFngt1yNeNl2nSMMBXtt1YGB
XpUgkSk9ib68lr307IjwasA8x5pHEgYHRDuojgTZXT44FuUqyjzVJk3Yfsx0/XpVLuMCMU7QLpPZ
FWGmTtpGezUFbRZxXYQ5bl/otV8UgB3oVKx8vmPucCj9jTbPZ+derUY2DlqGfDf9nNnOpmZghM8o
+jh6btu5sngnDW4sh/gDQEf0ZfsE7ZbOV+CUjmS6xRPyRVzXG1eOGa0qdQPno/FtnfmA0ZUIHxpU
jyJIeMDyQI6qAitOUjihrW8Pxpc1q88DrL2HwzgkTjDm8IhNFPh9njqFOjGeZIcMe9sd7Mgqs9Wu
I3fMdD55GQhCkb/b71+HbwdS3V/UEnjxAsXm2GBD7FF9CMuWQiBPdR/pJgZkPx8+FbNBx+GznVGb
gj6xRTKgp9goW/kqIhNFDqlyqntBT3W/1Iwx90nt+LJakvN6oBaqWBYhNJpT5uKn61KAhUqgXh+d
PJrZqhviuJf1YjIA/AlTpPwcgAzaf0PYj1ELu6wq6I6V5c7UHV4mQl1Fq9YfojFzfBoW7dEeaLz4
FOa79LHHk5yftjNIRqwFuv5qDDbOzxsWpm14RX/BPLaFcSjVmQ/K0DG0bdzO2t/UzfT/YF8opsLG
u9G14fyPbQU6UXBmTJRyIM6zq5sdVRtUiOtHWBU0iCd/Ap/vUfbrz4rHIoLV4VDt5uT8JR1HgZgC
IqMnXiN1hq3zuh/2Oc2xOuncml8pPLymxuMgB52cgwXNnfZ86hM01G+KkdBz/RiElg91zG4LKBZw
JPQdXC8hxAhLj+FLdJlikhRPweFNu/JD+fqmoA5wpAKmyK/GLRWskWueu1OsOdINnHm5X65yxmQv
0ofCvQcv76dMg0B2QglscpCjGBBW1aFK0iXs/iQV6rKzEy7PRV5Cs/QOrIwYozYM7OSMmkSw3yu/
9ZIGgnKPyDkQfsmKSlBewuQ6G3uNzH06k1NWgoNmXlcvNemhPWKwKbfbs5CHJfupL6SWFXrMmUBX
WoydHBf0Y453g/5SeXlxRNkgDUpvqcfA6DYmDj/BcvRnIBtzpcSvobVz+0QFwS4jRmwTAiVb2Pr2
khgUWs7lGmRmLXVNBmnurN5exaniMApjdLt3nAQpPJzjvMjwwZQDmbRJjLO5zu04zA0P5SbLfoYG
8r3WqRNy4D68KVeIEvjXsa8ZLRzILjjKVqlr/zFkJPNwO0t8e76ebfDGhR7GtamBMXPXVf4RZVFu
0FV/Kwq5a1NgpBS8e3+7afkqBVkeUHrhLZUMPhJwsMqX5YiPX2tPEFO5L/sq03XzyDwV6nsXJole
JeOrr2tx5vtxDw8hXBXuHQtTWyWbc3av6Wrwohn6wJp6nBG3UQvKh95pLX+qh7s5xXBvIWI1i0ft
voqxw5vl/8VK4cDixhM7s8qR4ZmyM7Bklkisv12srajkNFF+2IpQidofKvd7hEpLJDGDrgZALeY0
QPLNtN/x2EhZ5fD9J7vGTSZDmGCWGYqQ2MAhifImk8Gbxax5vHgISTocC3XAvgVW+kOfSuNQUsab
T6DkMM6JfFTHD51USRhmyJWUvHlf92oCueLI8A6Fc+2HcT/IC/r/RcYFLwr91/pw23rAZyZNu+oF
JHJ+cPPD2AlleHNadblwSa5nddPyOZgLvqztfFk0h/FRX36B4QZTGCEdXUFIY8rZ5noni7X17QOG
wZAPQdmSaeXA+Ts9ZOlc/HtchkM+GVvqvgQMgWJ6HgI7iUNTz8mHh2HEeARRQJ9S2yndHEvL7Loo
Ny7maRm2Mjz86OhAQ0Zs0itgW6sn9dBDG2Hr9zdSUG/80W3nJG9RzWEjnzxTcAJqHHx4iYept+O3
j7bYMUir7l2or4P4Vr4MjvBWceqXdMP7+Y42S3TZkbxWQ4eEd1MxmqA2cnPyZvt3qKjYijBcBOU/
QH4GNDzmHz8+sw7Z6Gzyd5IVY8+vVZtZtGJ8ryHTjXBABwoeZcuu+VgoTR2VYhAwQXhVBgcllTs7
yTskQ0ReKupJEp9dOFQblG/3u5gsR7xbZEYNa7Z4s0SQBIck/ORN61wgZbylbn5sVaHjEQXHp70D
3ezQVnBvrhLY5zP6P9kt6N6uttY0MWpy1s30RIcnHtlOvluk3Vmy+gu+spLzUNp1pNUDLlENbWXT
KJDme6ZZbYGZGIBZVIRMRmDg6kLlFfT84XEc5xB0H00kn5GU9WTa6GFpHDAcnkuUJZdg3KrKa3vM
odFcwae3pYJO/nu6hA4IcMFbnB78EFI2IV2/WT/VSBTyJMlPOmYftbpNHjI450dZ2pU1DyNTP3Sg
+wKPaj+dt0uALgTWtjPGzxLVlQ4rJKkmSg3Cyew83wccGFCe2OcWQOl+vs8tuCbKhiwIpXIdmkbk
kTMLOlFH9T40PwyMQJh4BZknDDD9KKTt6AO7C7spZyxWk0VQJNUx257PI+lmvQk208lVoOXeWNlS
gxt+UmsSjfDyGYjrAY6GGw+xJQLiGfN3AeqvyyglAfdpy+PvPZ0XP/9xcid8GVcl+eBZ2V4hB9bu
4RSqItgEPZi1VtKc5RJb1PUyK4AngKFE9Pu0haY1SFvPlbysb4cL1EQyvQc7vBwr3Hb+BA0dyrJn
oR92CS/HRNe/JmfJCkdkBNf5Afv5yj/7Uwie4ktWbba9SO2stfkWgVQhIr1fqf0OdvXCcxUTsv6M
UQC4Ghqoao7XUoNw2KriZ5utex716cJ/H1wPkHkZuhaSO1sJ2f2wzpCzbmBAQORjawkQGmKKdNhS
iKrI+dzPROvhhrjloArsVGE6BUa+x3g5fjp0gtyKiOh9D7nKV2c6YSPKd7V6UiO/Q8ALzEGexh8W
tUVo7te9EgvT4CjdzV9jNk33iF2aTbUtUyro6ry28U99P07X1cFMCmYWYVdGuFBz9JO0ecK1MI6s
BqllrC8d2V2tYM7j3vJDo4ixwqMdPpZf6DNGarc+evnYSGpS7HL3sHI17vArrejfya7Nr5kPkMoN
BMjojar9N75nunKkQ5/mz98FCrEGyIKzcXFUPj+um825lMfZGkEp+ngMdmwbOYAKP54yGwTrYCyu
2ea48U3LvM6oFqBv+PAtrLjS35rfqgbIEDXk1expkPq29HDAd1USByileDGHpULibCm5TLmc9M9a
txuYJIesL1EgkOGperJsf7EoyfBCkVseP9nn5UGzXXa+NwwLpybzNa3nAx5yn/xA5ejSt44BfC9B
Tpe4gPdrRiBeRSv0eLkPoAz+KJ8fpQbRt6ByfE4GH5XTuwNnzfpoJ6UyhtFJbp8YhsMJmweLOi7+
SZNkzJ1PKIvcNLhoEuamCzUySlhxkJe4ATR9SyWT0gEbIUwfCb4FGvJEf9m0e588FUesg40n6bEK
vpTBkz+ij6Mzg+EWzmbhQrlk0YAyyDc5K6u1WgQoMOftG/v0owFTt06102iFRem8NfOz+IpUdrKz
MviDX5BOwCUi7AQ0LNX8vk5e0VlibtLEgVcFhi2UKT8eLMKZNtKlODBM3xzKJhjQtQvWYISQmuWB
nV1XFMJDAvPQHSwX5wkaTmSO+a/RTHMe6Rloon0tNXoRsq+tzF6Dof5N53+zWwiuNzDAsFgqXVv/
MO+rX25EgWueJRHgmHjbQlkm9QEcq3zH5TGZt+IRNtQ2O0d4iTvCj5NkoPLvnpGSZFzDg2yvItAZ
LAainBwpTxh/s2n3o3hFLiDc3HBqLZ1Hz/gI93+b0lcxESLoUblJqYDuoc4RukfC6BQrPONsS79P
nLEXfrDHmfQjt3vjga/vPvr3KeXYnd6GZds27C1sWEbO6z0sozZiDOErvzZhCa66cCbxMbgiVYYR
+bUhE2XftKlAo59ninNuNvfbwfDeaniRHJ5tCJ+g9LRmjy5hHcaCVDz+ijSl6pCVkDDxWSlFiZaK
vXog7drKj2iXaWkbd4Eo5Ox+RWYdcB3aUy28UN6/+Bpa8X6oQxSUxX361yZtoMr0hKEuWd3kZPNz
HWP+LrbL/Xq6/LozkiX08H/1UzgvleNHVI0zCA/wdWyNC3dzIYn0zffEBhOCes3JTIG9hcq4R0ny
BfiZKHLu6nkcwQzaEzO6lKyDi7ED+gqmmlUgNUR/okW3xEjIbKNFduyMRjw4NkM/ODUd799mUyMs
FrcRind/skDuVHA7uXiWiWp63CDvpc3tQBaS86iqe/RS1GG3D0/21zZwFpN9SI0ioDsIayk7rv/f
otlV7M3nlDddQepyZlzivpRxOQ6ghIkk8uQMf7U/s4lRPgzxwRFS1WCBDmB0QMv+XxnZuYqzMu+K
9T+taj1zRz/6MovAw3XKTVPwN4JQHTdz+pEXWqh8HDBAJhW0HGyf6GfoVJiG22gCxPWG+8IXISpU
zUe+hLiVXl2bFP/D4j5DTwEnrKRTiac98ycAkEyRdNP9fXFAuLtvOaBFSmYEKmJz775BwhYYE1/l
lgnRIOiDNMtmp0fLd3WuSq8IJ4vOj/rqO69DDdvxwyEWrU7Lnz0TcMGHIL6iCwcw7gJ/sa6jG6/t
ZawB2RUx5sZ6II61e/XxQOgjKQTExR8JuwgLVzKY12Lwr8MkjXZcsJRKW1v+QkgfpP5BopRCUNOm
2N2cLSjPb8oe/JuRwHZ81V/e4a42luRWtwSYihpABoEn0InAYTHE8eGEP8t9jC9jZzM/uEA+GGqx
2mnRqwjKP3RdHt2Uj4I8o4kfN+lO06EuDX2l8fFULnfJiKLvrs/yNIyJo4lkp6skyJaon65P56jl
cNmVyId4iSYsv/3u7BvZYGdqDV40NhV9ge1KD36DcaQ9ZbTfgGOy314sGpd9asYhMmsAj3+jEKfQ
f7+S2VogVXN7uJX6MEoF/hW4RGodHsOS9MyIGsonlUZT7nImEsxzOdeGZCacPjsp+fx5hR9pDLjk
gU2IjKF6q/MwVfLnkzrd7wJpwLETfkRbz+kRS3RsJmtznSQevEKoP6Wq1wRaUjxwO5CTU6F/4+vA
xDGwv2nzLtek6mbxpgbjNlLWV5XeZ5gc6BIZq9ryl7CfvKEs1BcPIh9YmD+HA3H8Z4bdId0WyK6U
yqNEpsebK/aF4gStI2xk8s3XcBwWdvrF6lBdJDlJwd8bFR8G6xwdV7Sc14D39bP/PymqKJ4cIBAs
aaQsBErwTJAp3TZFJXhhIN5tn26VxdjnZwDjtNcfZYyFrvVlEG6AG5xW3JirlTbqxUYN8me8+Q8K
IamVFsl03ECwd8oUH4whLgW6R6KADimmKhNpRSWttwzpIpU1iIH2kQTf4aBQXuOMlSJdQM7uqLmS
jJUFWgHE4GIbXY4fcAVqrjxEGDTy3woglGcRIr7+3zE+9ZpT63JPshL53s4/jtewE8jVMZ49v2Tr
mNTZZCCJiHDhnOOm+awUa8A6za5X4JmsE17Ci0MfwozsFPFCJZojxqUTVQASVKBMfvHBup4lMiHU
qT8irZfc3AcG1DVoJ9urRktpVir0HZovQ9ySNUD6RgD72xtUMdDr6PddtzBumaJEqjGwLhW0KhOX
ZkMXrwSsOsNqsCo1TtHxWS37dw1ink70yy4PCz5DwY+GCZq9682SMHVMdzhFyGsF4E5Kxf4CEV4h
wuwk7KUCBVLH2Th9kqDCTXueM8WB3PyaGoisrTgoPGyfQscoN4K0+0t35eueZXyrCRnh3FnhkuZT
2E2MiaMLycGyj8dKyy9bbXE9Tp8ElELJBju7pti6TRVFBVnYKEpwmnFCpT9e1k0sGsaHB9ST4vmQ
Erkcd6IKLuwBf0tsX6nW7vVJcjYM5BrnydisfpzskmJx/Q+hWzO8NPJaxARza76S9xay3CHLSjec
zGKhA8iEX8vu84m3wiCuQtkoweDHlIhciJ5hD0VQbGWSDxqZjmXFIWVSd18KU2asRA9k7ZjiDasq
TjbT157z+ZH0zEs/BNUYa7YSt8tiOrG/qBEaA2Yy/mjPoFdRGGYI8xFcoFnIiOBUxLjDiOdJfVmj
8yVioAUZEncvMQ6AfR8Fkm7Zkn2YI+nrvQJMKbPLZ050692wn5YeikyaWqn5zq+XSulYHhSkHbkt
hJZ0vGxak0iJ5A0VrUtlK9aOlXLz1CnjvEDwIrTxpOVExChTtQ3Du+oEh2ncRniUrFvf4UuDhsZP
9nGx3TCHTqaIgmVPpNDfqNbvoE7JMJnxNEK613EFWimMwqIb49ZCMascAa3Ok3lR9rUo9tVCWHWi
k5V9quDzBn8s9CDdaQOy8abWzcF0kr+PPAKA0vnoY4inL3ct8IlsA3Bb5Z3cM0tHmkV1S3flgBWF
WtAYs/ZMBmQrpeIQ+HXuuseOlAwBoWXmtyTlcDYY8ISvwQD8wOMh/Fo8YAp8kQctwfyMUb0/4iA4
iROywTBNB/B0XxljmeGybLqMZqz1UuVrYWzQhspLyayE8L81vDYSusut9dNMVxP7pKG1f/OSp2uy
vVHQM46dNU0qLbAcaAKtHEfub142w5TzwqBVU3eH4I40bvoHkoaYxwVAlffFU1Th6rgLbVgDY077
bbpRJE/cgPxPh+np6cVnxFu2q/7lD6ZFdpSpY+0g7rSFKpn7bivz/Nd2ZnMK0f4GcIbE5cAqW6eO
IguBEfDJU2yr4IREDQP7c6t+j9xtgOungBi5nndKDFI/GnZHOCjM8w5FxYscSlpfl4eAVCRL/yiF
eTy/fugxtc+8SLDh83vMj6C0DvOOyaonQ9/RhQ/feKVULYnYu4zhFFPj3seoLAWt/DzsCHvwVxC5
rMvJMxh/6rvcHvOck9nj380fD3KWIiVnkcmpx5o5wSVpmUjMfQVIMcaJtKLOVlLya2B54FPVGJz+
9Gd2eTSGts+Wa/1Ad50PmJ3fCGoqIY99LCPfios/vGb/qlkYFE9HIpmdv57+F8y3hGT+wRnrs5iw
F8i8J6qyimP29k6tFXgwc88+jfIZ7xOSdWsdfJGnxMUW/zclxFg3Jej3QBqyyxoyzsmEWFX5eFOZ
mGfiKoEiRVDqylkui4zS4B5c6RmDlCeDXXSQqEzwIVDZC7hudGtE8RaAx9evgxnSwKokVGrSY0vX
YJqLLfZcQuuq42RiTgVyF7Uo/hY9pGt4Xbcme8QQiiqXEQhJJRE8cQHGRYwWDwWGeMz9/BoDPFxw
FECPSm4VKax0yltFeqdX1uWQ/n8Vjl/RCSbgv9GzSWIP3x0s9I7CCW5Y7JpkOwROT5cDTNLTbIpG
0NHyjPRGMQY/d5F98zItci5ull2+ptZ3pHPZeADTZGvDIRixdbr+tHYyU4lAXXJAeDTX3BNZ+6cd
XaHOzVsmGPyUZMftg3TV7Xq6Y71HaVP0BHlyH7uGgyniK5h+4DT5IPy4j83FGs5Vl0kr7tpUNJhb
CtJuYv3ucMrhsTfV5zBOZuTizQe5ZURYuC7wgBFVH4TVSWkJTLqmqS7Jyva1OlBQAH7KNEg0diw+
90zWMb4HfesYzl0dcJCmxh2BL8bA6xIEszku3yaA1zCY2z441dXbFtT6GLkyx73047KvlUNhq6Sy
Nzhcf63B33Qi1CebCHgIIBT3m6JVWAedHg/WZUJw4iKXs2eHCKt41QWCwjNADz2kSG/DaqYoTbIR
6njdiH1TDes7e02h4Wa12816WTSnMK9ay/RFRffGJXJylN8MQsjxFKvRRfDMEl4yERWi6ZJreBzy
ocuZUW6/w/jGJUYLFVUxKRONpC/gGXYhgZHFK3pX/Y3RVNzypmMPtp8bgGIGgP7SbVUXa8WvPUSZ
6zaW12FILsAI2yjrXcDkD1GB6+JT11dTzXwtJMP74PiKt2o9J+ZPChxGBwOQGp5jzofV6gKSXGdY
EFh2Q1vDhmaCobrIUBxhOlqoOu92IVgUnHm2P1eNW6Ns7sB6gHJZTYaQ93FxMSkZAicgUon+Nzks
XQEC/SRye9WIO6IhcDZzmh0jELpx1S8LLsJfMLwv3cROcAC9HGx8vsJIDKVyk8PoJHDFhSCH7viy
ukMVQ1tUqLxmxxAAD/IV2lnsJWyq2GlTZHeWv8zaILwT+laNkiYAaBtBt4im9SYFpr+c6h+uawjL
NXsj0TVXYvMG5Cc9x6H+/Pue50EfRjzR8j0O+DVYMga9u4PG9kZJfMLJDmjR22d1WjcaOexyauMY
Yps/yBTR1dDmK1qWZetIoC7lq3cS0yr/CdCb7D+9k/dtxExHxiMc9Ia/pQUhgiJfdmJaLUrPdfAv
2/E1ybq0JjW75ABAa3WZtDlAVegEWNeBqvUBIBtQcX/Ti/ip+g/fDeL1zdfEGEkpQYAGUOX9Oo6a
TRHZOKuDT4iOuZw8JbcaLrpHVGvXQOjFK00ZoGgAzwZP6Qxk2ODkMSttSSqrBNjKJU9Xwuf31NZu
zNWYjfOwInfqsVvisqmfGUPCB1nKNSzBGj8tM+rFOwosX1fXOYyiFld8f1qkDUnEFlxJ+xrQa63X
if5re3ahj3zBfkU/Y42p870jOqjWJvVanRXLodVwzISskssRX9WPk51/JaxnDy+JeN0/m5qm1+ue
XPNV0wqp2AQOoO1lOJBy/Nv4NDT06GK5nCYaDShXylgTI7GcZ+BnhZZO6zcoDMHas7+aa4kP7/fz
MLbNFOZkzy3Caz8lNns5cNMIclsKZv2jFqQ+UKsVhv/tuO/dehSk4Rgd+aXpaBSx/64kMJRBFYpy
At/kj7cCYhQg/Rv+eyj62pqUTB364WK1Ywyk5L4P3Uc/64kkvlCOz2UivYu20VNGtFS++frgjuzH
tT8+R9oVXqrv2dufvdxuDR2FlYjljaMUX76iMGbJVYVqn1XXVw3+nlmgAHiLtCv8rSR4tA5WQacB
CJRNTMu7/h++/lT/OQlN44Dtc9FlBhjGT4yu/CKkj3AWC9/IhMLqfv5iJliUj9dxlDwiaBn/I8N5
Zs1zOYt0sgN/gE9H86nLlyWsxFCdV0M4mVBU9EMkO1WxQJwNSvbgUv99K8apBiBawXxLewq4GbfX
2Ua9tEN42OG8FZEzOkRJo+bqPprYPhQOj+tFSXPh4I8VoP42cvxfmGVEHjoUiz7LpjSFU1EUBTbS
P84pO2ttjco2zVeOPvi2zjRERJYiUuLkpnc+/dkfO7q52ZRNC+LTw37tGyN2eNVkJU5N+FCWWA1U
o0wlv0jVl99y/3Cl62rD0cHU7VCwq+9qPnB7+YIm+fmD3dl/bus+TetteCDWYkfwNu3a14hKDHwE
8T1qV5Zr+o/mgyWUXAOBAYIZVJ30NFzu75YH72swBYrMHU6k/QKeXsOMNj1lJWTvEzn/ma4BDlKO
X1EF2+K37vFu9aYNr579VEg6e/cKEa9K+FT1GJfyTcypOTnKqXL8ssPA7Vki5byb8Ki110gP3juM
Cr9eKvV0qvwJvziyrIyqvyP5nhaLVZU5mU971vPTLQld8QfsXLFTDNadZOPtnMaRg3ChQTVUY34I
GMt5yRNixIUl90SxzYxHClDEjMkIuTpCsATCjJtWUKL0MtD9cH/gxlJCaCAvkkyGvHSL/iNGUN72
uCekaMNkuX74gIEkb46xETB3WVHRh9IqaFVdwqNnFeE76/x86vaJZ69Ib3EhcEf4CqZsTMUhw9Zx
pF1UnA5e00LXdQoIGpNj2vIkBck8kkwzr8T5nQAxwDewiGgfGHvhfu39kf2o6sxjSp60tJH9lCp7
9FfG5ap4zD9OPpPt9F/1ipq0sxF7bwf/phebLT+85nkimRX8C94AiB0f2Gsyrx5aNwvZPbddwWRY
sZUIjgrN6uob86o2m/tVfEgbTO7fces+gEIGjiqaKnJDp7zFpOAu7P/tQYwNoAAzkBufeb+vVGMB
PRwsD3Slq4+oKQ34zdXPnWuz1BnxU3+fwhVp0hLTXyz5rx9Q5J6lGscKm/QkmSqO22GWSqs/OOfA
ObsaUpf4u0f6Q0Yqd3y/ULjDRNS+14F+oc90V0Z6SkbkGQsQ5hoqWmGUhFvNknpDjKGaPBPMivv9
/Pb4vUENMwZDhZ6f1X0jb/ctHYZiNBOpRjn/pj6VqKqtfGDrB+w2Rvz/jwI3kWnd/BfwoVIL0Vne
zGoPWtt5mPISnGxUBgx1IPeZusR0ricgPKnAPD7/pKnlsa49/FjA9QKEbMwBLxi5DZOjBqaFnpRH
0Vl3CCvQCHQp/ZBQeQZsqZGg89dQ39doRRfTM271/2/eRAgrW7Nxe3NellXbv6rbhm7MMOYux8sV
JHNy0h/s+7ECSx9Fuczdlh2IhVqKT3ACYuv6wQP4cKblzwg92gdM1NRDnlFRbsua7GvjH1hWLTSf
/FbLdVltXdqX+G96BN2kZ1BpVxj5hJ0d32HejKQKJS8LmF8CM1QuyhfGKHicphx9H8dYmr5U+3K3
YF4e0RmbT9wQB5sM269isAVDey14r6X02mOmXOgM/6/y25G+2ge+4mN/d2MYpEyBUIUvGymzJW0W
T5H3PYaEM0Ca9x7S5FcksZkExB83i4ibw1Fxp9oQ0lsFhrwQmwGTUZpHFfa3udKCUYwoz2yUS8Sn
jipb2W/PbBcEXZ8wM+tNs2ZKIjNS9HDSS9ZR1NHrWHjZrZUJLAGlKOO85DROOLietgQ0axk/dfZu
NV6hNV0KiwxCkFiK3wIvWR/F+kJ3qBJBdVUvukQ+MJ7EECLEQfEpFD/PaDBMNauGcT62ex6PFg88
LKbJQAieVOxb351I0tjD/9pSP2geg1v5vEoiXrAy1g30IZbJsMQGIrWfSM1g3tysjQme5bHXhpSo
ercFIwVO+TewVRyCxnZ2dNoOCN78RSGdRUn0WFidfMEp5FMtcrAJDXnbsyrGDA/zo8JMoJEB3uts
ts4FWv35iWz8INxLYU7zxuck+lB15NdzlXMH4bC99e0k7dRji3xvcLHJ+OEPt7Cr+MUFDtyrAHUY
wm/hCzIVssqfgJnZ63UzHYmc5w/bIAm3NFusyHJBweN0TtiZkjJEl/XPjNp30+sgnPcWWiRJFnu8
ZSJPB1KPNuMMikiG8KKxoahHFOr82sy2bD2QoT6zOHamASRFJHKbersWtoj1Kf461VaxKS/vFe8E
Z/Zt6ldC9yNdcqzNpt029QUd6MAhzlaWy6p/Rcis8kyEfTyiyU8StcFFPiewshEIYhvgmz+r8pBP
R/a4y9Vla6rC7hwi2W9ZFuSXu8/EVvVKh0WX+D9UKxgoV7kfXJrxci4xoWvbrE+licwK7la4RDNv
6NeCcSuBPC+YwbNUfJi9EtdHsCYOEPiXp7oPNV7Sy2glO2UWQdTirFfb7XZ/zRTpEhoYxN57G6FF
fvGMCwAXlV+7sSoFKLUbR9oHFR+1+H5zv3vUDQThA7fDVqHf2QqMjIHUttQq+3OJ4z+/TzZ5fgf4
X2cAoDu/L8BdHuXd+eBINGH8vjFyqNLLRq/qG5HD/jUIw/ujY7RRBXu4j00zSAsy5jgauHs+6fGd
ZC6KTDNOkXLu87yW8rg7sE1sBKzYPPXs4h+GXU6BNjtMtIoz4AB7iscyf6OHnKcssy/AnqIgqJis
m8X9b9Bw0r8mMZIvIr/2lqVeeJQLyn0cMSLd+NMixfTpA7PJ7+cy9651cECVUf9duWlc6KGGaHYx
o3oHGs8zDtKIjKxaepz6KyLWrVOifBqIrfj9S8M6zwFeQITfRvyP5ChdUw2/gJUoG7yQGJs1u6o0
hGPBaWUv774dSv8L9IuBolFHcjORBQLYVpLSHboCqJO7FTa7rDY7GlyjfmJBNsvFJf5Dq7XmqFUS
pNGG2gVf8+S9Eo21ULayzRwBcfhm7i+4ugMq8s+/GRMJWa9aelsqUwmfCb5JUphEprQJpCEvH3ud
dViZrklUJO2oy4Q23HT7kTODFf+RmbQ/iaT/AQrBp8dKCr71G//yUhqrXg0CM6DOSj2Bo+UItdbg
55quIVMJQc9O0pYPl99EWky+vped3DabTLEQR5xG9yWMSF2i0sLfQXgdQWBPmHURgWW3hirRY5F7
Z72MaARQrw2HN4OkdKS18wdcHVJ8de/aHjVfmoX+WjhIsoHnz1RLBG2quW506kUYu4Xh15nt4HON
+tllSeF+RPqJ3IsmH64kBC/flb7f3qjwuhHnq8fPMRhV+RR4aJX0yDW61n7A5B3H0cqB3wt7z/wx
kbGUfVpcqoygqJzpJ2PlK7zLgZZT4/eax+vc1YbKIUpYzjRYvZb29Lic+od73BFfmJKKusr/O5BG
vk8l0dR/KEZXNebRTJixgG50S1KrPDja+efIpQqgVSzT5FH28wfWlVAT6JNkntJXRL0buBDxA5ko
XTnWg+ixkvzhwZkbMrCx4cQ4JlcUcmTTXnBnAvGhXXoDPX/ltRrgJ56WaxzApLwU/HAk1mQotCMc
IaO7bEyGAesTkQEZ3+HcFhynfbUjNKOXSIm/e7F5S7zA853EnN5YoJ9XCfBzd2w0DYnLzmAYalCO
6PwyZjZG0fDHpftrCvDd9JFJ9tYPeN+fJUHXjC+FrSliPJaC0VzShfyr1I/FIBUsxMxnxRyIWfLP
Zs9X6ilcfiOHOMKa8s64AZi6RjO3bTjXjDm94ZaIrDysr6+EsxpgXMrYEjSo832G5ZBb688uHByn
hwyJc1g0jImF+Dk0rV9h+bzXA+pO6WEmNDLMzCx0uTY0Aps2k7k9rxpwIMJtd0A4Sppx8+b/mcQa
YWLKAoEHWwcm6mh7QH5Bmks8p3htJkbdirV9u2zRBl4TQCan58rkKV/6L5ZeinlpYuVAwituT/Bm
RMCfdS8T4SiySWGjKEqHQWOCEMEOZEhQunXBJwcHgpvFL3/9EvJeFrP9hPrEhvQPwjebPv4giEqg
djQtcJSQb2GWVdtIwqS8PVMcWpTVZyCPjI0fgrLHlU7Hs0MOtsu/Yym1DX/BaUbSyBceUXLZwzbY
EY5NkP9TDkisSd7kWF1OveEV21PixDUP0EMc7Soeo2arUlQRf/DuO5tvopjnvlcUPsOVD/lftYOV
dC9sE1OXPRfD80qZYhW09/VwPRpsqRP43zPoXGisdkQhpWHXO9zncpXFVxO2Jc/s6r1CXBo6hy1t
5oLHbAiReI3gHk3DNIkKly51kyQsI+LmP7dOv2HuARRQlnYWm9NYZXCXURloBo2dFTPWdK9auWCH
cVKImdERZu0he8OoaZLEU5uDRkbwoQKwNS0xCg7JfgFpn5b8trWxnwwYsuWyF1Jj/Ia6eU8MATcH
icrnp+J3gUzf2tGe1zChEuAqE/UaLjm9rDPVjv2/NJPwY1b0SgUuM8dzLc6MgFLPvAxqrBYayR1g
DS8uNIbOqq93MdR32WTrAibhY5Ix7TdODShDS1QZIhu8A0VtEYNG8wKWL991xkXh1Aqj1kYKdU0X
k4x9LhVeOCfdRZbrZaQb+cs0iLMhJZVKPz9mAaBGWlvsS2und8pVKD3guqoaquaQcJwL1yboOx2i
iXHD7RhLrRy5kB4EtsnmnfqfJOEBKJR0rgQBkLLGp0/ojRgXkubRJyNBusq33nW/tQdumkXqDElo
6YZzNk2Bl571MSi47/bbClxRXbxRH2zdbDogAJFag5RPwkEn5+KZ+PIVYammQTg2mqWDPYDsWQ6T
MzQ6lJNdAPF1PmHggNxP0vS7VoPBgn33rOuTHRAI8c5PYMuKbxHzOzUKYBH/tD60v3qIsabHMMeD
70fpzE5nL/GvIsIQlSJwbckwau/Wo/56lL9KYhQ/OMDPW2LcyabEw+FmF8ZnLKz8uS2HcKWWJMDo
lBl4gpnEj8g/XbcxGCdIo3fOhx3ZeF0/d9eVx41AK9Evc1glAS2fbAe01QEiYbsOydnWqIPVcXMJ
xUm84c9NVnv+xzAYEp/odhmKC1k8dC8iTewoZT4eKoXZIDOLPteGgpWErxDfFaKa2ldFHWDGUC80
ZM5bxQc7XNQQ487EeZpnXPeZ1/aL/D8hYnj15EXaspCkRAJRgZRKyqKMj3MYmEbIcx2XQwJqxWuA
06Ihwrbh+CoANzlZr+m6+sdzTbhDRTLPwSuLHaZ3ZQPQ59l/QXwtHKbjrjWMo+3xZigZdRWwy77A
uXMxkhh18V1Y5Y/1RGgep0MLK5HoMkkXYmO8i8eyMviTqw5ORyZ+loUPs/KI8gBPSLNS9MnOlqyz
VPqqnszHq1GIJXy1KPI4CG6wjVErGZqd9SWBQtX+BGyCmCO8xFLpD8fROSGLzZ07c7IRxgTbohxi
dr2mIbo8Uv6i8lHGUR9IHwmmS/MXEMgfksDimtc6kEa6UMK5SWuFMv2NSEHfYP6hZRDeC6SepALw
zCDWngEyItzt6ciE8d01H70tIhSezMHAsfst4d5sNArToNJ81MKXJcFpkQzr3qeffcGni8iqTBK1
VbpC/EoZGnzvcgyxcIQBVviM4xXievHZWbB/xGtChvzlrzW/aCDXSVO1zQ9dP/mBuAW6fRYN8dlE
tuQ2eAy1XfZ8TeH2k+sx/cQPNcYlgiwmQNvRQJlr7A4zrp6FCXwY0SGPFyqWWrUkEWvzQzOmH+n5
M2NH1MxrSXc1mz6zZRo8CbLNJGPaQNYlbS4rRrmloKfAXLWnqbaqYKKVSiJOatCYOFE4UEEuQk7T
9Irgh+cvaoQg3yGCY/JEJ7SfjiWWxeBEWlKAoV9nV1xqhYmPrXbBZtLkthTvxtPVLUsCXwxyicc5
e6haRZ5tNpf9vfYSNlPRC7l6bEFymlWorSNMyemxOREDD6x2H71KtoO+ga7/Cdc1es+3nU1+HY4T
znBWM8fO6DHSUcLavwknR5FIYTE/nd88t7eiSZVEgUda1hcVLa9WPSp73ti/Mpk7M3VlfoOKnxnd
3IkgvO6FoRUeMXXd6K9p01M0f9Grn8vJvw7ZRBhLoxQJxRmdQk/zVgOaNk7AY+IsUQ81og02AKC5
v0YDPq3T12Jtwqq5uGY1BMaCatqRH1hL0nj7XrvUN6DDp7vgi8A2uN3fAFLFujgAnAsxKuaC+VhT
atWTcEMOaESsj44VpNJArJYFwK/6C8+LVmSaJL9lpbd+WuiUfncX2UV13VYAneJZrieM671jYr6p
b3E/BkTI2w4LfWNuk9aaQ2PVliFpTp9R/V2DNB1m1iUGohlquAExb8B9trSpUB6HH4lRflypfiJG
vklgK1l1RU2kvmJLbi7+iOUGBkDhIkd+4mA+rTs6ZscfjwCNMT1f0+46I0cBs3GqVVBf3wXb0shY
qlAuLl0aqaFU6c7Fy4JUZtzxZcmvvSSfuAnUqnWhk2rzCaIZ9UfSAbXgM7uZ8mz8zUFGDzX0If1S
+JumIYRJypFVENuKmmX/NTvhPLVdCqNVqBzYQCjFZUUNZdZDLogSweJJ4tC1x8OqLGTeNwSFTp1V
yvwhFr9M2FLoelcT+/LHrUmIXQn6rY0Tpgmim07jF2lylFnLm90k26lx9PRAplcnCODNm2MH3pSj
HKZmtO5rlrh794WpY9OWwTwu6q84sYonEdHuozy+IBWB0YgUrFyhiTCG3IoWD4S7N0Ajr8AS45Ih
vs9wAp/hThODahgiaUIv+3ZOHBcmvH7cWnF+3I7uw4xONNNDbg7ngiWg8wQkwnwn+A2pHXbrAgxS
ObR7XbfJMnTVI6mwripZM5woqflHPn/5OoZCgb7k34tkAvUueq6UNvJLkMLtdESZTqJa3dUVzurc
FsMikoDFjaDqJZoqzwJqpdv85oTiMlztLaEbVtDJuV3wKbEn+1/8H1p7VVqIoCqnpAPdSr8rsT7e
wQAum6gv45wQt77duUG7fmrCijeEBehzbYIb+b8ifIrLoc0CUQJgWoorILeLwmTUlkLnUoKFnfsW
lW43iZiMSSD1erNsNvFNRHT+Jzf3nk3biiULcHeDOVM2n3SiBs1iP5UXTBBcB4DKsAEmCkGyzCMH
K20dckyXazE9eIRIar7wj/SXbiWbi30PEjWu4e6kvgWOoFchWzug+sVqnXCvPRhHrwcHsGw9ddGu
9rI6il41V4AfFuM4ptkMqEZg5KqKL//JU9KpvL6vz9WtSO5uRot2liil7oCyp5f15fNLRISCQ4ze
ELrzHCv+23TZMErCqWvPDBI2QxMxTfQxElzawvbgXvsqCaTg5MvXj1O8BiRftHxit8aPcTGpdnpe
nhh/3WZxFDLU0cgEi1/JR2eDjizccad7kXXVy0ZG6/2W2S/9PGZZVdJICqecIuCUlJDBGfiTbZbn
JDC15RJz5Bl1XcFNYQndQdv//eHEr9eG8AvbKyGJ1nbw25dEKMnd50uDDo32ZhhgW+p1jCiz+aLg
RjuERK68z1zs5S3Yuhe2hbAxJNwtMMvGHF086Juc44nrpWzhgSSeFcMJjIK+icSltkh8QuJQrWfS
cCyFekTmunrEqBJQ92G6xbLqrHGnU2xOPgdGpjb6RjTwt7xWaHBOKAzbk2BDrcMNjANxUy27Hx0H
PaPDA0GHso2Y1QSjLGJlo0zeBvhtb6XgHMHmgL8okjbqLllgkevUPU4l6TZgjQIrW1X2aV2Uxw8B
Hi6jsGp79LhcKqpWGrcy9SLFDvvNRBraEMjge0V/EjbnIu4t0JNFQ7pxCc6BPkDkRp5BeAKY3x+i
Vk5Si68JRjoxvuPZ1AA08Sc9adlOk8XWnxBR6Owt0D3dmPoXS8oGFKV1F+aMgV1agVDV/l1FPBVh
89AJ6EvkT0TUPlEdzIY3ZiCHCC8DvJBYGXLeBPwHFZucboCnZv2TESC2eoy0eDDo8PNT6/L29NBT
lYnCIMIgH8WJT3HOmZMTBpvynPDqjybIsvBATgXvEARuKmSWERCDn3SuWTEevdtt8bEgfVtRGoHR
gvJWqYHz7HjMUplZty1q5asBhyQi3TUhDay5QOYIQqqXnJ+SkzyEV0mp1Z9KdNqlaVtWbiotxqoH
Igd1z1kWxx+fPVpzr+Yt8Ynja2oodKchQ6YzwcRX0EU3fTJaPubTBxUwjQ9SY6a0SHFgj9SfWcJb
Ix6I9B+A5363uLMfWAD7qjYNDc32UTr5ey+3I2U1qvedZlCyiZJ8usFfTC9/4LOUmv3o2aa+jLcA
8X63DbxGDWiwb9mdOGwqNl666yZFK+QM0XoxmQ5rq1Y+RTKbpDIyT6/611r8AnGmQHe83vqIYB6p
lOUYx9rpWqF2yiFLq7bBJS1lxpiKvKayVYWGHFT+38Ibe7dMlzxjQzVYaVIUdV0d5fTDF/1hpuyp
UpsP0qpMAZ4PogjMl3fwpD8elfXSeE8ejKfC1jxOxDwZCaZcYV7PhsEMKYeY3tuE1JG05lS3F6ui
ijxZS89FvHXVwKR0AQMSfXarqlRfWwsaqznWiau7WLcveAemGmxXuijPyLx5zpbpOUNxUFK6E4yA
XYBEArFC57HDO2UnRGvhtwyNcZjsN1hCWnSSHG0YGXxPeH1T3RqZd2CCwvMOyTKDzJ9KWmwsqowh
RDKI69AKR4GWNZH4Zk5x3LYNgxGYhz5bMWQkZ6kaTv4rlviWQeBhQLIgXxHcvoCTMQ2YWiGz8mPm
oQ2F9kQxH5Z28/WstFu2lLvbRmNsMl87qk0AEgaoFVF98DdI6TNdCR7VowLYL/C6VlesMu/S1Cxs
d52WwS/7897y3vyCvtMt4hkUeFFKcxbmAivh2Z1zSozl4oICxd3W5OUI60Lk5J5e9FjuABFax47S
uqNUuRBj+pmf7X6udQDiLoJCJCDDZfo8pkynE7YErvEmlRMz7f7IMKWSfMZR28vdJY2i7Q/JybjL
7TGm1cdqosusP2GKhjWq0uLqYy16dOhl7XvFcaXYYHRN0dRGxfI+XsZrboT8jmFL9wW+YeyNvfid
y6edfD2tCLM/fYHD+T6rQjM1Ar4BIf1QIqE4VpM73/jtSwT+9sgivjxMOcAgcDalYvdovSmd3Y7w
oBu+xhqHOj8oZlC2msm8Pr2rqXhmmVAqcNt1ItRxP0hm6WzjHi7rBPlKoq79lYKZ3xjXbdNY9o8L
8w2u6tlMZ/C8DZQa3WfzBOmzcKwWHCKNwN1DZfMLPitIueEVCH47qD9DlQ9ALDZwxLgFOsNMA0jm
JizqX9Sf9LHuVm8uklveAkHCYlqxn+aHOET9Lka6SEHIDBU8HLVpvhYvh2ojlWqX3iirfs7zyZjG
fKZTE5AdzY0SEbVvvh9E14VQtPBBiRxPMfNcxFTPxlJSadhN3CoBGa8S5JHSuO8QU+wAaE+xKnv9
s77xekxJdp8nNujQblCzzmCAG8mHU6EXHPO3PFXdom+BbrLcFbk0uVQMpL3//Zx+cz5LLaecegK9
gZgX+Q3POmXvgophL61PgLt/d80LTAZHdgn6P3o5GU7f7D6ze2eiSyXU/FYF7aTmAjZtxmVMtwEN
ogAEI+oEUbV/6RSMCGeEZOs+VAebyG+sEptWQZkHyrSVcxjfR3BJ8Sgj26Mf+ft+cUz28CO839TR
gwBgEsM4cZ2fA6zvK6omB+PiTfjn05LazNt7iUJEf6hPDZW0ASZLJIL0Sq3sdikH+tDfgEmjgdtP
M467tVYSxPBr7Fll51qPlkhVCq96+9BxZPxcAnn5MiM2MpFTimS+RHsN+g1k6q1iTBKGjbrNdI4F
2IVSzxXsFxRU70yW+vL3xN345335P4VLxSGjuQyD2kxbRRziO7ehDYbXBZjE59y/tZAlwHiDLgZq
58H4lmVJ7LXUo/0Ja78lPsbchRCkBl5wEIDJelSbLxBF9pIb3FqUm+nWKYxl+Rl/kdWRtJtlLzTv
CGB5nCMCCG6b8JY6UEXW7D5C14ibExI/cd7GGZR9bQElwo96Cm4Z5N/+0RFBgmjq4szoJHvWxqUR
mDdYwLdWKHdkqYV1p5oTEKVxjzf4+SSTgc9vA9MobDk+9MyO1rShbdeDV5mh+M+dVmpcvVE+7NTB
iKsvd9buw+mjg7CHxlJH+spV/ZX3449xMA2LOiDxAtvlzt/X1ItLko6KQ1iQJDEyuQInB6lzVrbg
xuf8DtzgLQxLaMugz9n2gueCTASVh0tdDT8cRVRhJbu0AORz2FgjHMkO/ENW67DKelea22XsZ4xY
F2GeBuj1xhRR81gWTjBR6mDVSZrNRdi1IqQ6xw8vCDpvMlePsAgF170CSu0Xu1yT4HgiiRQIrVFt
PT9pUrqLB2AYm6pgkb16VhGV/XO3I2GRPAMAFxXnKVu49fv0on+PrqfIWZ8IsYqHDFubWiry5t/C
ysnvETXvhKkC9sIn+Kz0tGKLno6YlsmPieohpygdJfn8TvZo1VXPy5LmoTuvi1NW5LDIWOlTeM4e
I5SMVFxI3WIUJn34LTnYKUmOZXA9dvLI6ElkBLkyx45QI8rW4zfYsOhx26FMgHqDnlO0zFGzhqxH
C5BvuZzIdLJB9P+CW4mCVqB9MfwqBt5o4UG3FCoYkcNfHG412s5AAWYJPekGcCI2Gl5jSRQmFKpu
8eontSEot8AkDCPXbTgvW3RKjHsPdBKDlSLd0vTUperZQFMqDuh+ofFbycNntJjq45rpTXB3ADF6
zDlIyxQgOc7YgSFxU5n5THAdhwnr7gJWMUnD8yD1xpxsmTiI5TmJ9ZYIp93rFhyzz9IXfbplP2aE
jriMyBn0TCRdKVLr+Xymc7PtjErUlyPGTyOHoTNWyDz3TN1tA0IMTJFxW3brgAG29JNJD6cyZFeF
TcLVdVx/kRU2xDdRFO1jr+/rJjo00zN/xdT0PBETL8ZqcGKmVv7lWknS1pFfpEvAqCTvfWSggWrD
Pv+kpDV7uXmyznkYO4rmUBMWRgip2LMNvze+0xdsKBv51+a/6exHHXvQxrmLhHFZvFaue/0/KrJS
nSQmw2Vc2GZ/0c4KuZUyage4AbhR5J5EChhvUnK3O3plpXV56B1OoIehd9Vw+6m2Ku+DdK1PGAUc
R27waOo57wMRmKboZ92Su34NqrAQVja7YWbw/qE6cBICiVyoFKX2+QjlTZ3W2VNPv1P16E48s4eW
z1dCkk4dsp2Z4QAQ7KDVzaHM5pfWIe8d3pJccI7WhJNlexyv+rdNJZTfbDIh75HhZLcINdMiZvxZ
KmO+M16VplrJeX0Kg0JWLk48mht2S4Fg1mR/bUaD23W459fCbk71jr9vJZTp4/hn0mRGAPaciavm
a2CU+lA8zPcYyhCqFvcAZUyAep3aMOA5t3Tby5zbbH0vELiuR+D80BWI+AdCP2KZR8c8qoc9YfDN
PxIh4FJI3xG01Da3ifk1re2kvo2TBZlGMC6qlo+dQACNbYzw2npGpCoWAzxSALI1cL4yZf8pp4NS
ct2H0ZbOty64YLLDwuRgFmk5OVBV1AtR91yS/BCw+prPi4xxkBo+rY7g4pPegh9zGpVVIM9/gpTW
k5vUT7J7JT5b1dwrMOaHOqAX8w4aybFFvzBAYxP6i1YUepZMqTM1oyDmO0BTiGN+IWUjtVdFg9w8
16p5+VZzHJPhiwqkIFcdPlhdpPnoXUvWpCgIdtJBEPggF6rZ5dTJYFwgmrg1qfBwNq6tyVWadN6c
BJ/d43/Ldp9nX4kLsby7qbY3fZ1X3ZtlFnMklzaNBmGyGIY4umWQ+oQF5pIx1YqHu4lmuMlS+583
iKvWSWczUIEo5sSPD1NcyYzMSP7wNLD0XyIpPMkzQp6KXFJiu17l+8CpLC+Qkmr7lMrA98Q7Xm1f
5oPWTaXRk7ff60yRqgD8ceBROjtS8XsTLVqdWgl8Spnn7ogQHBag5bpDvSelk7ceIVXIc+3GyilN
fY4Ixn+ozEp4Cp+xbL1+8aUQV9NAdt1YX1pQlMCrrfcrNOv0dfBM6iGuGjFcklq0oYzPXA3NJ9Fv
XRIPm2mQh3bULUeZaq2pdAqrclO2o9tQWPPBixVmxjYhxM2Fr0d3cN4oJFxl/HKxc3K6ZSg2Tabt
BiMVcTETUD1OBxJ4plpwTCUzu6rbgd5X7bw95ygCnzXEsEsxO4jxobL7Ol212SX71AuCMIaRWfNl
B2vFCUKzmL+bQciyfdbF7sJhEZn0t9Xh+3sD0j0TGYY8RNySMq9NkxbQBoarNDxZRce5cFTyngrb
WSHrUXRMX4kkLWDuML2iyl1ofkQVmgSvGfeklw9rh9781+C5nRvlb74266fhNGioo0x5R6nfXU9I
P++xFotkfIn+9ctbApKYhJWuoS8qghDXpFhu0wHaH/ozBz+yPcl1ZGwwUi3dk0SYhD7yuFyMZzFV
UT1x5/II6GtSQDpzgOFTSFkvV1PQcTEFx3O80CpufVrVFnHW6FCJYUBN1nMetmu9kbXTVThNTN3Z
ZYu58fJ3dH5Cg5xA+c0Pkabro0yzxwRZWVJkyzlaDvEQeEqtEH57DDsrv//azRTkqiA4fc6yTvnq
PNp8I1aTYYvTsUIHkCOFigfkrvlwlkDfU9feGMXV7yNl0DNpfM/x4sa4UAmt+YaHjkm0JG++dvlZ
XLnh1h3/X+R0v/3QjoqcrX7Ju7iEXgMCKaa4Rs52skVFOd++trAIPGR+C+9kEmTc8O/m7XejgyAT
udDSJ5mGbYTWO7EqPLRMg1UWlZJY6E0u9xsYloTCsMUJK/rOOcMJOnI517qpm0BOKyEWGrnhaCK8
uMTrOjYs0hEmnpjojtw3QuZRo86r/3s8TS36onoAe5/NvpZFgDyPJzHMi180+1msU/ReNQvkxwBZ
ZKnbVgx1QmF/1RNGbpNBq91iWPiFg4Px9f8Ru8qu4A3ZV2BcBTJtXcozmiSV156NSU5/4XRQwUUr
M3rbjzHu3Aa6vzrKxhS3EWkQ7pLDALgiqwVd0YkxyszN6Gakz0ATJXbhFpKz259gfUKU2AI/v/vb
fL06KhcqdPjxOT7R/0Nf6gBxkaKEdUd/hKappIp1slXssUolvFyKkTzNmeFFW9ZnaPJwl4m9t46t
FSqyitio6UIBGbab9dzqQ9Pbq8EnJu2/TD3bRFuojoNK3QXnkw2BeAof1j/+ekcFxZsu7WklMFc1
xv1Kr4txKnPyjXjfmVi91G7/llMO9zNHcwg018EIub+SR0tiE1oPvZealYODT7yQWwjcvxCqpPdK
3IgY/9KLmj83cMvp/32YyWUo2SkpNRaFkSYe0Cq9ulfGotM5LYeorBuZyKcVJU9IjSlcIUXJPxLQ
gOv2ilfUkBTWBy3Ni0Y3yVpvQfbKru0UdvzS2ZXPgBdVNDm5GrI97M1guLqSWWqtNEIho98JVfiA
NIyUiNUhCWQ8MlszauVRHG9CJn+3GOwKVXVAH68OGEmVzhqayDv7s/F1DCyWjXJBzAIWy+NwfnNK
JiRmUn1zDBuvfPeBjLP6YkazEvPb6GWhJeojm9RsVIenTUJXWLqtaG/vies+gTE+Sqv84LdD94Vx
0EXBFF0VoXZLsEnvuL8KtliBQC29fvJb3RVatvSmEhxlbVClXGQWrRyrRGJ7747kadTtQU3Ls/xt
qQJboyg1nXLuvyGv5QivYU6nllFz6yESm17VNxTZvpZXZ/VyNDr6gFfMxPEEFBo9TSdiNBZY4esN
nbD2ncNxm20SQnVIM8EmNrqBS9cf3lgflwnOj8sSy93bCikUUOVL1RpSUHDrM4CmJCzO3lBiIx8A
v1sta6q8RBalnhkN4+zI0TxTgq69b05CnLHwcbDyL0LYImbNqj8U1+xCPbQkS4aDuW3OIQA3BIvK
yVOCSCZU4KMyP1KLKQI4nPC12G4X3giDwkL4NItN1XfsDKr72M/X0/0ZQFq+jCi/KX2vGK0UN1kf
4kqn3B12YwQb5nUDKoL7w/GPHae2m8zgGIdpJF6+0/mBbbRxRn77jR8lRt3EaCI9qnv79xMtAy5g
/EZxYKM3xekFKGuLAFOvDvdOig+ROfpEydVCLM456MIXZ2LOpFabfWpTuT6YG3nrgvlPY18t0gTx
sE0XrWfnKCXSTRFm7d1hfRYqk97tlWBjOtvmBSYmKyMmG0oBlsRAjqwAmWcz7qTmBsCSZe/qelyv
FHTRiN9pBuqawahMtVscczAsZVYFcO1tMwoo1AbqCzG8D8LwAaU9kvC4d6+9Sop/osx97rTGKUCV
H/Ut+RZPlw8ZHKPJL6lDxY9wXccwDpmz3OGbBZRq+1Cgm4iES9j3xUz8ca4TAICOa0nY6VWNp0Xc
cL5ll1dXqck2MSy+VDNWe3b1XTX3sFJ3w/X/f40L4ETX1xMStgOdwRRmrYGJDaGmoBfnS0Atb0GH
7lw9MQ3AbGL1YEIG0btPPvvW2Zymaua6FhkI7FTmusvswfyc6kr2OAooWG6rpxfvUtEEGqpIXSyK
zJlx7o+PfPHsAqS0L4hp1ukFHJJIPy2nHAhj39FNP+Zt5GCMNSYgLC3iih1IvPwuSit6yqtBeg0Z
Fa3Ls035RYNCtN/zzNlwBWDPKnrP0lP/0O0mEHTJGWf9zRCps9DnDvLCbdIvVIVf4a2iB4XyiEur
hm1yGIA9hQ138sJBtJMcg6L5NXkznRKrcmwL7ZbQKv/QykWxbyN7dHBumxqYo4+rwiQjCf0A1fRy
twVHx17zUqYrgMI1grdxg0/rw2PlOqhUJdH2AwtfkSLOlCZ4grEUHX4Y9ko/Fz2+DpSP/TzNuRiM
qwtlj/xoU+hVs3BU6Tn0kyuQpX+66/CSOAMhdWilJGP7ai04+xo7FBQkgOdPYbl2DvJgOt2EEH1f
QXryVIAP1qqaQi5hT0f/t2oDikuZaidXtub11Wo/4SjIP6rKGVEo0KZ9jLuzs3aoFw1DS8K0XdIF
Qcl3OeSkPvWQFcbWBGf9PXrYWqkqgcjpDKPzkx1ggZvr47fe/x2hgISaqO63rUuywAUUy4LlI3WF
YlVt4uk4YvjocuYJ+4t0i6JF81nl1in8+CdAGsIfpdKTZsbFKXmXbd7qqgT4TNibyX1qOCTAV/ev
+RohPgxCtFdMF+72E2v2J2ZcfAUuCmN56ddtEE0ZXUF1FTvt0YK1ylzEv0JmtklHdZ0hAXq64a11
IwbNW26QH9NJ144TyhrD3Rr/uky6ud6WXAWSL+1r+7dE3UaVIb/+EthENrHNFuTfZJXYizoAzi9p
NCeFpH3j144k3mMWIZ0ChrMJ3BIA/SVFhVo6I52Jm7spkB7P7gL2m9Lx+a9U1fdTRXoR84RkxBpx
V+Ssr+g3cW3rGYvTBNJ0U0mH5i7m+L5QyYt42fjly20H0/kwRrWFyU+C5l38BrbXJHaNLhdLvF5E
JCjwA2LqSS7TiqJQFFg4F4khEOKRjX/0a1hGDsQUGgIkwEfK8jXE9OT2cjOymDpcWGMcdD3w9Dn3
lOYCEmJezKwKyQDg1HzjnEdf3uuN3VFgQgqOhqJAJJUOzlIXhi594N7s+lT1GGftJ6JuK+zPs4YK
zFBCtiXWafXo2RMuezRfshphLDSBSA9K7cM8CjhdNOMk4ZzEN4rxLrZtqIqFSp5WYNNxpUURKCCy
5uO5mbjVoSlJFI9Yvj6cVFxMQsTpv9PSOaB72AobJS1XWrto+6FQB3rs4jmFjJqM26dDNbkEFWYu
D/gfZK8wGdhUyUO0pM0YlB8bj9AtyYyoQoC0tsB9Lwbvox3AQWsZ2n+8ycyBKREs3GXCEji0eMeu
IHq5ajRpFgGog1tukwbCFIU0rHYfWSueGOLp97vF9usGSKIpFeM6EJGQd9M4zkO6xgE/zyAY87be
5u4Baghnk2NTIQyvGFU8N77WXtC6nuy8ATOp++BQsk5SPqEECbtBATTcw9ZmApOJF2p8oJ7c3qoV
bOlhQVwQXvmWTQONLbvx0cmgT1Xd8o8j4ZcrXuvTuZ16wy0pppvDip2WR2HvWi1FCen77g2ygFRI
GB5uuJrjXNufh9kB5eqjHVuJGTDX/AT62JVE9pTqnPOCa+DtTLxNYjIoHgce0FvGL+2UWuC5Cqgt
A8/H7pe6cDh2VDuA+Smrl9ILi2UIZIzQoYPF6hISddGDNRNxL5c8u9cZp5Yw2xR62yFQ/NW7OpzE
FFTx6Lc6Tqd1n96qGHD3/9Qve9kLhuVL1Z48Um0zErTk4g4QRQeNS0/WjABOjtarrBO9bzxuTczi
a6i7CWQlkyBiAA0sAJYHf5EQIEBzlZ0fSivKfOwkVYVCWl5pT7zfFH/9/G2y/8hFyJbqyi9dNzuz
3ScLoFySGXOAktN9ZJgm1FBbCXiLpd7mCKjXKXo2W5gqISNKU7ngfIioHylHxXpnh5carvwVEj3n
Yf2ScPJRMbru9B+d1ijhTMhDHikNtc/1WyP6XJosdBTNipOV4+Dtw8bO0ZhRPICrh5mLnDESxZqa
hQ54NiHRoonM2OFGZqSv48WOhGd1dlhsgt2NgaVFk8rcRYK8Tkvie7UzSFxA76vyA60KZiGkyRKp
fQXdVIMETdPRQqSPfTy5mjCygIwu7xAruLa+F+lqtyywKKkH3zxxxdoMzDf8zXTdfN62tSleZRMB
1sbrR1qzt7TMXLxKE2WI+Mn5Qmew5h4hkNnNNw59TJJtjBDu7CDiO9Bsyekzyay76fubC/XnnrDU
h/gk7zpbPmPm/ZVkWMIWR7JXo+sRflFWEialeG2FrW1K0RLb5KGdQBNOKRSQBjwPLkQIJX/f6Gba
MLM8cWRmCLw9HGouxqim4rAI04qfO7xVkXTqvA6wQgEpwo/P4POlZ3Cp0KA7CloUCeEEoKnk9wn1
HZoss7KISXu0wxIhF7KXs5gghU1zd4EJaq9J3GAv3HTP6FQqFfrDKmYcfeO3X7Ds7n70kaJ5hdf8
jao0SIFotWd+3aVVkR94DFPLK5/5jWR8ar/Ulzn4Qpr/C1/Zz1+IefSyifOzVLssjyUjzVC7CIrf
oKskOZnbUsY4YcqLroCCOqwZw+5jsm4CpFF2JOUyz/+MHzwjsnWsN22QofsKiNXMpLK1Vl7qRdeP
g0En4F/+r19MZsPIkDdu34XRF9dtWdknsxBRuUwS4U4akt4OoBtmb5VSVP5oT/UigZJJLbRV83/d
sO6NldsUXJ7mqbi27Fh7+oaWh6WROKwG21qcs9IzCoSmcwBTmHowZKJm++0sLXhifDfpmjN2Ttei
xrjRW5mwV+oq97KOVq2bBfoUjv0VUGyVw/QPiKvDrtFpYX0GouqJmuDqdrmENnFdcddPJd+Ul0nC
UYsUnM5vjrApzH9XRn6ReRQbxJOH/KdSR6NrGaZ2jTcGsOiIg/2BDoGiLrxZInZVO3mqEkkZA4/k
UyFwm6xMkdR0eDEMri+jsCDAYjw1m/T5DmLyaoDrgJz11cx8I80zITKLsprQdFJHsVUpiTmfPYZK
OpvzyD3UwA5HUzVENLm3OGx2+Jh+O7Osq82y91q+OTw+AMsRloBbt1llBt4bfwThEphTTKavOha+
1+6vdULWjDRNSFes7NHcc6e3Lxg3IPT9WVHMPbVfhMhATrp7LCY3tv3p12aXrPm33BI7NPvvPlzL
dh2uJBr7Zt4y9BW51xriII92UsKf2s36NuzYSPS0z/MzxM0txBKQH0ONCFnDNa0ETa4dmel0+oHk
xjxYAViAo9Th8Vv7tlJbaswjq4/vEtvDXNVVGOx69E2Hekp5nlbdyRJciWL8cdUfOCpJ61AEvxiG
Yn+Ul7vB5V56FkswIEdh73N4La6zDV5ZAQMMXxfGpmwNOmzJDotYxvuy9D8AA0DQCcIz2pW26k7G
Gy4+b4C3DETbgBXMdpM56Q1hysnx0sFR6+c4bnilogbomphK32WWP+ytfq6DS2VWEOoPLRVV4bO0
K1gixJjZ07Aji2uFDF1xh/QTx+hysONqxjU7213lEgdLQZbfmffFtIn7/n8Bs4yfz2UXLdyXNWUG
2YIP09iz9tkwS1a1wvc2JfqMXzYnlx0kqcnIyFo+d390UjNzwSr48Rj+DdJsgX/0ZZ/Q6PkETcId
SQhK9BEaOm4iJ+RVcsJxqpTAAuy+eIEe/5i2b4k7gkHEFr2Vk5r/ckS+mLtFFqo8f/h8cTVquA+U
U4biye201PK/8zIR4C89v2AuHcnKKNNJ9fAQ584t0A/04VjBUSP7KuYmLaX7WQp1iQwFJZiW2FX+
419tXj56L06vuO+LL+YOuSXi/Hn5ivkNxA947adbmFwfhIzoi9AKPJDGM4iwZP9i5jSWhmRZvpIb
AU8o/fzMdLs/V9zFMddxBrn+kOaAloRRnEC7BRaHi1NDvDgH/R9xAZT6JfZwZMRiy2Oq/o4ZfM+E
m8vn19StQKDxQaDpXFKB6AciWdMhlmTbnzIEHBcj1t/+H5XOj4P5M+5YPiG8JRr3dNrQKVmpbAaR
9HsSwrSf8vz8kuotxDo2ROkK36A1umc1emj11bkrbuA2Rzs4XlF1yWfoNcvfABwT5g55Lg4aSges
kYD7PD20OwcQujoEfdvHmFm5qQNtjYISLCYnFsojn/d3yqt2HadOgLuHnQCmz9coLGFOMftlBSfm
c6scXwE/QtmzlRra0EODcKmg7/ozePYYnsKzJdTFn0P1MRmzQVi639lYQnTRpRLRnjTltzX1aB9g
zWdz9fuLU+4W4T3HkrU4OwAoCcwleh20qE4tke+NeF9CksJOVLpQ4+VA8R4dNGEojhRfe/oXhkQc
8f+vWm9P7NWGpDEZwQ2LBXFqYuKroiDsQrIrlji8Id9WsgMazdyD/vuGEWEUqx/+7hXAzg0T2eaH
Cp0FoV4MeqHC5fLsnroJQLPOpHLRefZWElPtgeuFUnGRTB2WSGvBmtGkQx1/jN34MLoHMwDVlacm
09f0mNpxr7mpAHImpW89zwL6VQ7+b1paAlL2JqxGPTnSgcipB7CByUVuSOLqBqAC0SZkqVTYCvgL
UVUpfk/VJWzE9au3I2RXkhgBLMuUikeE9p1G4osDPRGPXVTeVpUQjMch9ZdC40nggEsAoUPLpRE6
41ZasCOpYEeh2sI/iBd5u2cbk7xLZrDQnmGOZ8f+LVrbZEW4Lf1ogAcYP+CBquzA21g9233B33bm
LFIlb3xmih4UMdrk4G8knYNFGBoFoskxQrcyTHV23ICEqqWKftFMdRtHrvoU3qbhuaPICFGJprxG
dEaK1OJppZh8x/ZzPo1CU5tFusSTlaZ/FzRkLgBRuWWZJMMVLXgJWcWgihxxP59k0S+IUGYeVkfk
JCmBpAUv0VkhRNh6SByRvulId2Q/mxf80vyMAMx5qOgNc88LY7sLWhgMB+f0EICg3PkF1TkaP+pn
N/tDpP8VSy5orYfAFWOzNMil8j3F+fPJh8Cc5KQiEBRIBH2+J//Bnq64s2Qz6u4nZIvSENTUCZ4+
GTWl4YdtpmlC3fM9FVS5y05aqd1hXVd8AalqxmkvUyRX5mWUvlLCAiqx4pJnvxASkVs6mgz0IfeX
IW/upp7JnFd2xxN5dhjLEJ+S9yupE0ELQM7o9osInxmKz1LtiT+Xsnkepw9GoFwUoANMzO8pqqgR
kvMoPscPXWaQvJC0KqtAq/f6DORvu/TmKs3fwpIhlZHX4Nt0HSClV3JHiuMYQK849AhrcsfEeNG1
YRnp6cvGers6zlqdZ0nCB76KDMz1fNIbv1deK2EpQ0gkykXy6pZWCMmN9ktw+8NTfYxB4OtVHT8Z
ErGZUxQFsJonBAWX7q9RhlsW+LXKQbvnuDo34U2DT1V4QxM3nxJVOz/hFuJg34n3D38gq+N0cwpV
sA2uBjmFDEv1ik8DqN+coKLQFmHnVIrUdto4KEfP5JLKE8GYogKl1ZD3vuR9KQPeRUaALfuB5ZbV
v38iAvdZIGFrX5bIFl6fwbG/L10bdL/0nLb0SFefUa/B6AXXFWGW5ZH7/4kPVvWfMG+ompDeKap9
6KoKJyaPdlhGuZJ9ZYjfAL7H9H2l91fxJCI07m06tGfXGzeCQNRkIU1bgsQuvz5AbiWjrMYiFPqX
jelQbyg2VOZiLDy0sn1JNzdU7tUjFeaYOQosOgjGrA1KTj2Dznh1Snp2YmNFkRqtf3ZUzyjg8CWL
9xtVC/+awO59DsV3lwZ00fHSMfdTyK65t00U4zJYM/5eBheysbrp/3GZZJEx3j66SIZERTjtAvgU
ebSnNoAio7H6tCQ79F7CF0EYruT/FOIurJfgDDHMCRiUDDwD5kH/7Z9lSmRCxw9F0oqMIcr4BI+4
Nwd3m0RFoEGodRMb91Qle+UMt7By6BsbxKvxK+PaDte/7+IDyXfEuW1pVPPz6YCIfwnmBkO4PPNB
ocUy5mKpVE1uO5VvHUkVN2cc5aXNy4VqRWYmvbAYiE1Fi/lUUvT2wTdXG23IoakKJ/Fpkzez7N6c
h0uRIDc1XOK17oG6Asot9z9CB6jskFtcUCh5zNpGYJucOP/TEY2eBX326pXeREvNDY5YsiD4xNmh
iWpbuSci3LXoKh2RZn2HiFduX71B4R0YZvPMmEzLwRi/a7Gwk/esDqVAJww1LajzBXZlKeAPCZmV
lnMCZHjtPk+himIkvO8grkFH1Iu9BdVl3R9MHf3VWm8qpUfqrx+UoV7GOMyLD3XTBuYmX7JzrbRN
LAYk9ucLvADxHiYoAEbobYvkiUPvhVh5OEZ/bIqhXWEi523MER5j6EKG1fOFK3BQwOc/j04OYD7q
1mwiQHOBR9/Tt7R8zOJPQ7ry+hw37oVYqkQZElzw3xRmWekJ59g5W6wCRhdKELN1LcTF3CDOEkr0
eUARrVRGqALQMjZD7lysPzecTnIcC6MnSTA5XuGN5kAxAfPYxRt7nJnNL3u9ZbPyzdl5X37oTsIs
MW5ZpSffzFA4XLYJ/BrGDp93IsTx0IALI/1NoHqSkGNu8xn1G41WBnUh/edT4flGQ5r/U4Aeiv0w
L07kj7avg2jMcIl5X1g0yp8Uq/1TwbntbrdEjkr+tB31pfd5q8qMGbrssMgc0ykAo306/stPu6Nr
PvyOErrqF4FOD171aLE82OFeJtrIzWgNg/+Eq7Onx+kcOXp7zTkFtYHwwkJOKyI93bgpJNF9L1JF
Xw608YpdNCriYf4Puqd/lK0k/lFQ1I2kTccav7MATHfkMDX4OKNPaY98ib0N0NleujLiU3B0tOt1
KkAmBEBW1HFl1VBmBFTC3l3jXUk/oKoTiY5k6KLXKmIMCYuku69Wv+8FUeP8WeKoPoyOnbzBaia0
c+rB7Jh8A4eqwpeVK+PHIyU5Po2wcZ16oxG+ynpRv90yB6Pf4jCQw2ORGlx3z+leMwOR39zyaQGt
zL7383hw084F3kVXnTf6OAEoDTnsT4m8JzFRQYzEvw512Wxugugkzu8oky4RCJEHSLwAqRy5KUSr
cdrzVCJOPs49VmDFBVX9TLW5sBpewI0mKtCuwwkyL77ybck8oa7+dIhHJznyS7HhXuCSMzk3SURm
KRhbUcqE1WwfRu5nfHLWTdxiGsS2pzvKq9EF9ih1gPq6/WAYPWwK9MyiGi/Rlg9r6VkWaqs8JFVi
DwkEVOYZPmTtnPaUiNdP+ssAI/Abs76l0WB7D9WAc4x0KAj5M1swqoTa+haakifNzzhoBylbHytA
H+NfVutyCWzaX/Q/TglVHZ1GFS5QAZyGUrbN9CSNKOMS6U0P0BL/VGnMcRA+RgZwlVxecDhOgQkR
B8WezKIvUbGMmhkFfrnsYNtuypX/rUnYzyUGExmw4iJ8b+1V5XpS9gX/yPQowp3GwLZ8thiPDXVb
9JVHWVcSqbCCu1+zyQuYQ/2mV+/Lfv0K0HiiBZMhK4sPQDpMI7/xbEcqK+eOIUGvfuxKADVZElId
B/EzRqohjOR3h9HtTS5T3jUfKQpdrwrU0BLxcOFKpTO1cKDYJesfJZhY7anH40mL/LWGuBV1eVRh
8AQTPo2IdqGi75jdBynZ2sHhF2DyIpSwYJJoT1QvJ52AzCKa807EeT6JBMd/SbUK1hy15EYihA2a
pYrmEY9b57dR9gOXJx85Mmxu3nF9+GIaEd+bto0kIW72kD5fH9XhB8w+MeIXYfcsL8Mx5oflbuqo
G1tET+lcPfcTOxGh+ZyRlMIgmNEcfPhQCQeZpviwLK45XF5SKyj5/MvUf01SvrSk6r17hGPVEACz
CBnzh91ReGC0WKnRkCFR/QoLL4jozmppDhrVqMdHxyjZmDicwgrCzjJzNYuV0MLu4U7AhpU+GIkb
nBvRkVr9GqI0Jvy+gCftaYKcQ+8FiG6547Sle331Cn0zYt7SAfXQOWg7rrtKDVQuAcAiAbmFVg4X
hD8GMX+e/r8T8C/mDYYfk7MYml/HLpAIg1iBtOoajtvHdYv2J8VhHXdPXTKonsaAWGQrJ3Us4Pys
Xmo/kPAVfXTAv3a4Y78vKUPMkNj7cLQcH2ZRJ974q9LQwT3f3Nt+BC0Z8ZH8SBfOX3Pz41O1bXHq
tjXYcvPVggz+FVejuYJnz4OIvjKzernDXs1WBMKBn9bDew7NNxlQGl4Ow7IU+4C4wfeF3J2uLpjv
iCD0HlQIxZWJL4ZsZ6mu/WySmIcpvln3L0xXAzgxlO9dAfI2NOYazw2qJGKG5cGAdEFaYNHq0k1A
VFaIBqP+fQPe5iAKpzmiRMWdRZuXAGf4wA5jITobfDDRYVXXw8PRatu1sxuwppu4qP6wxB7t11ll
KNQDOTW2aODq8RcZFst0+t1jQPkHuIt4vc79+oHBnA1e+m7X+1R3w5rV4vdmlT3oi+1Sd5LzUMiu
xQ9eC2sIQErgXdciZXhuh/BsRnY3Q2FBm3e9cRcXTA/ujXCJGIZnFf622IDc/lcj2gM8iUZgIsDM
BcTAiEZf1Q5tieG0HeBC4Jb9kYQux5dpCKzhdTqJ6yG31kjb5OM/FxmW7xdcuRgy8EE8LbIvY1aG
EfSbWmTp00xu6xTVrbFyMxhbu4yk+lkAxJkRu/yedboWUUhKP8yvktj9+wlAdXhaH9lHL715S69n
yZhczI1Ng0am+Krb5j+RAlceIhzPA05/2TG/eEXLO/aGjlR0e2Ey8Fsw8rZVXYxOSfM4A+U2rYS2
BrZ/ZJBNlLDxj+8DgjQubMXMtX3aT7vEr/z/7OfwN1+/vXVe+DYdACk68BZPznFojlIL8WYF2uQY
LEsgh57SWOEf5c6QesrMxVHqws/n7d0VUGCBTAaaNz0HhCprbRVyu/uI2r4YqyQRhQUujwS+IRBM
oB5wHtJTohPzRWV2ZLqLw0lszVbXOKLb1d0+OEA6Z5cR9UMTTOgO5EUrzonmsZOVwUiBvOqKVTff
13CQQCutVEw05v+MeogEPl2aftkjVm1TOXyfcRDQxWICXR5j2dlGDSNJNo14IetPc8MF/RezHnwA
zqXejGY2L4mODtk9qRr7mow6i98/yP0Ruc+9CfsAHjkeCSXzFkyA18pCkh7EdPklD6j/4eADvH2N
bW9aSfFmeNuqLfDCzGjlOld8P+WAJCzy5Khqkyq4Ik7rWt6RVXz/89padVbnSJNISdMhzhwY4lzj
+iFcTimhjgzDsg2KVY+9gMWKgrtvB4LwyKhld9gfGtBauShgqyfgZCGV6Z8Ea8XVtVXZC/36DBYN
Osyl+pNgiuqSVdy5VMhDBIIktXIS9zFuZ90idia93Md5Aiqez21QzZPB/gO+Aqujga3SBLe4LE0o
WNYUgiQgq7r8qn2VItcfs/kTvidlEdsR5cInmmPGDqqRf9e24180S7otef4V0A0Kv+UYB9AQPcgT
mAVzQJodYp3co+zCXEMVasXO/yYL8HC2NOu9/FmELkc5dvhFSB8Z60T6lRJAGxTH+Hw05REiHk7o
dBHu/Y/gTiJvGWoXfuH4z3MNunaArhhpGDIFsmSGxJNmCdw6cnHOFC7Q8A0mKGRNirfqdt2GqwQM
NH9uFSsUopcOTcSiWySEABJXoX/TZftbkJt45OoIcuRaD4RkT3RcFeNZQR0MfD7T/zMjxdbSEhRp
r+9RxCam2LcQbGsibVdSH7fKyesCFDbrbfC8nUeZccezosgDfDiVDSlAEj9WOnUerds+VLugrNNs
A6Q6DbRP7FqdPfNCJcQQMFHoTdcPXks7AxZsj8iooR68MmiCdGIivStetFYtc/UUQSHzTp2t8Muu
3iQ1/pyWAXuF0a/ZH3d+VwiQvdXVEodcbD1S/5UDIyI8anMX50kxTovopzzH9IwXcgG5Cuqs3/96
C3roJy1DqxZWxD5CqSjw6WDumf44LRCSZcnWdOn8z0QlgZOVkshd42tcziqLuGR3jOW6UV9vZiM2
Bu+T/x1jPBuYVIAp1+U0FOpvys5qWVQtX1KLKpSYzNjn+ZRxpSMDi8Nn+TvXjhiQ0sn6tG71wCEH
iYy5i/+zENCwrcsepgLdv0uacunqYwiu9oc7vbqs6PMXng4Sd9Y6Fpx0cIFdfvVGHVAOBiOG5fkt
7tI7lJ4zlhrMtJWlJkWW7Qz/WqIcKbDW+XoZqyAQy6ug+rLnRu4Iq2dN2GImbX6Ovc49iUdX95vg
d7zIBrcYi8W7k81CsCgqZe9kO1UdFW5oBSmOOB5UDjmG+FPddY7V4GhH9eku+OHTfLPUVWTYEhdm
+NJxAQDvP2UjDRPfZI0X7QVk/M4s/lEMsDyGXkYg0wV/DiOpbdmavwDXbU98Gym5X07wF6pDlQ8D
tZW7Q5ls8UTJ9SwiXLHD8aEh5Nzkpg13nAbZsn81xYnWOQZWNhmz6DwO3aZotBWuzAjudn1RQL1p
GV4pbWJhvs0L32Yj5hWCisU8OvbZtUBMiv+/rTcqgjqtBJkPP58L3GPkSdGTQiUWoWOwUicd2sT7
697c6w6Bjd5b8weKff3cXRwMEV/Y0LJAa7powaBY2dljmJxCHzepK+gN1J3I5oXIEOahkshuXwZT
hmrZrScu/nKIfvxh5G4OR2tgb6iVDLN4GJYDaKrGYmlCuohfFLkAszqSY2rFoX1fDdl/Yab3yUe2
InWkgzTzynXM6Z/fD53dgsA0phqGRhb91/4lFWfSZOpZ+GfhoWTtpmnfS3pPhaZHNW1rN8ySb6A/
ZThxV7t5Q6QHrsD98F/y6M87DrEXJfgmoREXUdFQ+2SoPemYu5Pn85lQIe2lAKXR6dh1ZhFCfWog
txEvD8qB2f/TiIEZXgcberjIiOkt1ieemoii54/F5O5lU2hftUefZuduX5NlwP2V6LulQtmHbr9B
7AHalzrPfPqLtBDrj1QJoA4Lr1UeY6KwnkYENRC5HsOLs8jGGIavUSVBtZuiN1z7s3kjMmj4bROo
3fgt+bT3IUsdtSj+ok7UOU3Vm1zF78CiLZ/5G6GCqHK9UrMUuc5hGi/eTuvuqpBSR7iSfvTvUaRD
CpTsPdbwc9a9FZJ5UCKmLwyouINdXqDAcpgO3yQeVDTomIxui8xXQPrhI1cYg7GqF4Ub31K0atSF
6Ecv7VoeNlbGwFKFpSclcUYWe/D02Zw1CQUMwZlY07MUoS2jbioqIBx2oIeOKy2JLGtG0IWXdMl2
9xnWM8rjqnrQzXdcVjboaGUOC7eBvIBhclLiJLtHuV4o7gh4y/e+QM4atO1qGBWGYtuXCnw/3lx5
HbOn0ioppfLykCpQGo4Hn3nCiwmagZliPb7pGUbtu62eb01x4VsyzSBahygL+qFGLLUAIPEXW883
G184V7wg06lWJU/HjfPn6tZKX0jNpwTkLyPsfFs8M805+hReOBZOTZtXx/OMeHEh2wFIloZipSnf
ymVJzMWDTxyG2VXRaGo2psn0V7eB33w0YFjVNjiX3A0RzP6rkR7N9o+AaWRu/7sh2vbtMAKS1drC
zsMcKmw/oDf+ZZkyp6wecz/woAptZ6C7eYF/S3ut/lcYmGdxVXhIGtU4TSuD1+78g3TyxM8ep8vQ
5iB3XAzzgeFWUiXfRNkgYaWhSGFFmxzMf8nlCusICoASNpzsAsRt6mRUO6BICuu5KdMw71bdePS1
hoaoIXcvx+9XRSnS4JjxxD5eRzO8kSSGDD8ffL1Fd5TKiG/KEXRwxsBrhYSgC1TIcUUFoY1uU7xs
waA8Bm5ekXg1X4VLMnL1aF+qiZnS+R30VGtdrCZq4CTJ9gGfZVrlraA5EvqPf8cwHdQmfr4mznMR
IEjvyEJj8xqIVycqwm6NQpwv1dAwyzPrVW3Biqcx773aJzi72rJameDIccB8/LJnYFrwZj3uW8dx
dorfdYWtT4ihdQ5Fhs5oluqzwMix8j3+3+fPf8Wq72cSRJ4wLoQjGV+Qp9BJWtaVW8C28sbYL2/S
SdpJ46WO502QkAh3t7g4ptxL9l2/Ermgghjkk2ncd1KZqxrpBpd1wxzZB1De2/hy/bBJFOCUr2OT
p2oDBYgTbioh7QTJEL/JB0aoGnmFA6uDAoKAzWTFW4D1mSkoQLk0GuCLJ784XRjZQfBvRg5XIn6W
cfAIAYGVVeC9vcBc1RKh45Vwu+6CWVt/Gojpqb5tiwxbTrVkLsvKyLLNMCWqJwsZ6f897Xnf8xE5
KvVB8w2BOWg2phtuK9doHISAZWCk3Wg7+eGHC87Q64Ip4S22iece61Xcu0iyKASkTPKvrRTibCVz
DyfEH/5ZWIOZDXrRRnt8oerzTVR2nFSzsFJA3Q2g9i71CH+ksLSGco4gGYrWk4dxnlk/IcZc7yL1
MFWrBdnoQLSYJo1xappZXB/F4bbl2fFrWH20dT2flE7SFVLCxzj4fxM6qTO1oNy84mc1kPOPeePv
q2H4BA2vfoQ2jG3haH0gNAR/P+kRNsDJojYbuXYGKdbO8e4LEjOwuEhDe36TKtP7EcQ/2rCZPEnn
Z9Nu28NRLmJBTnKOo5HgUCmoqBII5jFDcyqnsmLkxSabfnQpgPGgkqYet+VfLd+C4XW5O42cXZp7
xiHbVa3tUrHllbW/8UukOq2O6LYIHGUrqWEm/Ixn7JS9abtKYu67gC1I3GygaqlfKCwrFuSOHxB6
BN030IGtsHH+6Hq0PFemD3awDPmD2feo1bysMjWcFG63Uo4Nzt25TG2yC+YpML3vGq2XnUucDfa5
mQMJ4eEN0HlwToI/RpRttYB/u6Yp9zpIP4bICCk9BAqg06XBw4X5fEN3ZnV6NYmSgPcIT/z1dfAh
Ek6HyvFHvO1DCnuJZR7K5krbvQAGoAJPwNoSrJp33WZOKs48qRr7oya+MKxJeN1FbijXpvp6ObL3
fSb8djqUz5cH3nWlq0K8bD4AfwPItJMERLo2bGu716IbBOt5/6D7K2wjgE4nxLTaFdpSsei+LwSM
yOqfvjfS12u/l2Lk0GYCEE6S4qWyA5cGysvgAKRGhb80a1jIKvJwMWhraL4qiAGq/yWYn/dZ0cek
DARGirNRaBgG78wgSjh5v5YKvwxzhcNXlNkOOp73XvSjcio17qQ4VMgSsOpfe979anmwHDJgsinb
2Wtiuzlis2N8i9HE7b2YqORe33RyFVAFRlTgGQiPGbyheiaCGsTLb3yst6oSjk0KedfGxPpXUR9u
AtWX3ZoIQZgw9piSDvsMxMx04LhFwCzZ8GyVxR6oJqWq18WU5hITG5h1Mvf7LDHYDaU8/85xyybc
cm3tDuqe0TqodiaVFN7BAxP6gOExDEwIeVVMX8KMyf2VAlig6fpeIqIpJ/MFCSR749/QSNc8+9zb
KxLVzRY70dcvErsAE8WPuBLffRhbgxThBmV+udM0WeO8ka3YItQvHJ34fyiC7DV21Y3eKs+tq11e
iWtj7FuN7GFgWR+Iw+d0htcp3L9CwTYZagMiwHd/AE2E5Nuevw19+TtfabMp5wKa+9CRIHABf/5Q
EqxAEdtdG0WJJSlsAdPQYCYIlrPIIZXwxPTvfBI7fBgDqSE61okh3gluXB5tkjzi01ViFEdygAHM
LhDdVbVsZbkL4UIq+UXTQb5zA3z85aT8w/hEXfHbZXrdKhtegMG/yZsaO7sU4ZlbuzAUSX2m4Uf1
sH/Jkt2xq4Z08kPkF0wq7zpjyQL0u5nFpm2sF9Qu7gTEmN73j9wSbwKZE4KiWvKUjDqItViZ2khE
vhNxov75G5tqw4KthisnfUvu4AfqTNrnF/xwKDBd6QlJgXQyEIAnB/pTYSVQfmYcCTCJoKSviOb6
pYfiE5+WU1TNbtkg+5lHKgpx7L68scokuZANC2ogc8qa+O4fSbiXz6FgZt4QX4jnG6DGxcZiFhdu
alSPuXBlU9QZ60wRlIu7JsRU7qfrl3mUQfibs8GcsV6o3QniLCNTYDSp4pQ//XnPPGUJ7/BZqX1m
HSRz74RXlkgncO/v3H6lLaenthM5k/cpuFPqgA3puJA/erZXiLg2HZxuHQ+RwFYJl5hOfBHwAFoR
E8VvVqiInVgFqZikvcyg9k4ihGRFLdWACLG7IfIbMccTEE6/4LzosaJu3rgnpaqQ0psfX+7VKcaB
8k5bRPBKB8JqJlMG05p2O7M/Qt43wYkOKxDju338mM3s2xqupkZ0OdQO13dtU2XuebcRij5MS//Z
vGA1Hs93zRtiY/eSHgL3ApCUs8PTxRm9TMKCDlHELjpKfuc9cyUpqEZfOIztFRp/cA47g11hg2kz
ybC9HbA3cRmpWC5IQsGBSJkeoxip19LzaSqt/Yqjbno+YmemOEQQpgknpHyfIlvDVlUvYDIxaSiI
Gu5+R84ztuztlXYFpe8ytD7JdXrvul4oYruWwVb16BO75s8X6Y5+hPSj+388xQceOYKUPJeHzgU5
+wgYnZm540UUozrUd+Sqm7f8YKWsPyBpuRlnAiNVfwRiYotnnJJu9lkEayRACl/6hHDncAT66WKH
ogDSKIPw4s8yJXOdR8I5w3j7J+VXb0nhytTiOUmtxltOGSGhaaiOxYihelhg30Lw8gDOskbSy/PW
M/O+uNj580SFR/CZH59yNNLcAE0ncPXzKws1s0+eyY2XaYu9E4OJPkDTYD+ZOwEuQ1zlJhH+vQQa
1jJXMuz5JDlaGpDWg/RBdtRii3TBVjlcl7XshG7to0weda8Xec+73cRLeOfjPJoMFVUjoP2H17pt
7E1f3NmCxZqEoEwlwqGVuCuI9hj8YONKYqLx0Eg1fmozS2xQGzJB5v7yq2ZQ50PDJdD18eIGO/jY
7tiy2KPsg8KX4BNFzqhbhp07JvfpWFUeId6oRYdu9DStMQSO4TbDCNtGiqsltiYdJIrXhOF/cxhW
OflekNAhD67pH2ieaBuEIgVmg6vm9vX2AWmmkbal60kDsf5bWRU6lAnJ5k5IGFrKsufgGHjLZNgL
a1jGqQu2Bb/psW6/9l1yA8gjd/9sKqIZATBQogQlaihSQTxSg5KQAq4vFqYuM0SHq/TBCB5/uKrf
JVmxapHywDWvv3UkZvJVZAIAkgCv8NYAU1GpJLRMRWZAChRFjyG1dwTDCk86capAW1MWHmImUueT
qr7eu+PL9cnX+hYw/L5jYWps0AWguMVH7zsrbYIWwOFr/rQpveVR02rST0K3Wvbgt1/TOr2406lh
p+TSS7JTDaZOFubj0XeBl/0NGtcjBawBtMAgDOsnW2nZ4X53fG2tY9HPTbLCgKOK8gkJO4+1E03O
Rm8bNBTlQu96t+ksnEz+D9yO1SsFeJ3Z1Ci3VuCFk+USWjldAOSd5LXPJCZP5ZfxzCVftvVs1Lw6
LuymMcPqwAxtJzXJPt8zadwhgxEWqzLDAtIWOAX/ADUDIDq5+VyWvtYjpUsfD0Z9n0j7OYIgfAsK
4pQ5K64ME7wLUoHbbRqfVm0wq5VCzGCMDb3+2ezZgNFVBdoUFauKQnhKcg3pG3mBK/JONI+YHc+r
NijwI58iMF4rIZmAHczpl9ctW89nR9VYA8nv/yprifFkO8Vgu1PRBtB077npDPbVFF8uDhgU8H7e
xyt/ZPsY5PSk3v9EmM6oi2w67+srPRmDig06y2FZEA3rEgW4b9AM1etZxH6D0c7H/YZ1E14B9CJ+
ovWLHYkRBSPZhiN9H0iwaZ156zDGTtkJff8ldqFB2NHCsvv4E3jNFP9soXMnxIPM7oK3HVG+c/25
OG1DRBwAj3chdO1xRtEu1bTWiVNkhQs7JYb3Kwak+4iPmc96NVwGZNBh6RaJ68lnvjK/GkTCLjcC
UrE5Y9Fkx77FbYpC2qrU/wRQd2IB2QkgFj4BcovQnkh/LnCZ4PUrf4TPMd49G+Qg+qji8+3UVuAH
oUk2BEKx5ewvDkbTSLS1o/DolaBC9Vbq5UChDB7EFPmG5bmpC9zYLtTf/I9MfhaI0u0HH+z3fE6l
z25WGOfniEfO+WOrQ3t0r5stWF5KjPkgkR/bnHQGOn20ugtd6J5dbHOnlox1IotfU27Y8fqNCUx6
LzOZF4kns/hLCvTpcFPcl5NBpXTMlIdJL71HF5+nTL/AjjkPhVUDFnicbibOzlFvGbzzAtofoHV9
HF6EWX5fdq2MbTwVdLYHztFbpRUARtN0R9agCcpfXQ0XfD0OFiPXfwx/j83/xAftdWKfY5f6p2Xa
hxYFclGwfcUesgpMepKW03bPeltlknMjs7d/RBeR9FcQVTSplPkdeyOooRzbE+XvONt/aWTC5xpa
oijraNU6pwDFWHceweRHvI8Z+fLjTrMrHRlg+Y9cTuqdOrvUCJVh+c62nHwyeXV4W571mIVtPT4u
yVzf1nHkjzqj0OOkuO1d88O0hfJWZe+B31+Vs2dpnGtoslIS/dVty1V0la11sLxgKpOfSMXqXTII
T8Hcr1kssw1x8jb9pbgypxV6HJUlnrjKu7W8fZ8IpkwPAxVtg8IviT3MLR9aRL7Yq1tsM62PiT/j
P9sttsd78+EF7KD4KxY/xbT+5kBzWZHKZ7RTCVvFkfoQYfUEVca5BNH2+4JbbpzLi0FdFC7gabOI
jSJ0hrydCvfrdQeLEVUv9Mt6WcxW5sf+z8unnzpA6P3UCuV3eUnTlcJ4biQGuxvZAbga+rkwjcp7
ph4wCludbx0BtIc2WCKmAF1QBQ/SnMzSo3dCyDuFNomaFNP46QRbP2A4/k/V1YGFVB4hM2A0m1Fj
/0U43VPsblcu8+mWoNtPVNBK/nbYrHdYVUiTt+a2WD4tEjVuT/0wwf/dyy+4BhNsK2z2ZiVCTvBb
38g+S3/8kplB+OpodPX85F8RgrIuvkwLKrl41jQq+EMZ9M6T2LpRbuqR4aaeyIKXT6Is0cUqHqgz
qFXQtfAJMne/p/G76U/z+T/oB0cA5T64ylWqKMBj+krGJy9u92jy5OSmO/sbipWsInYQ7o/1rkRo
UFC1ictjzllcSkZLwiG/HZFJS3utMpp9V6XWzyyXNNtI+7IE6T5Q/eiJEJfT9vMyOJyxtI3sHr2k
/rZTaz+3/41ayF5cT8oAOocngi7+55Nuh/jmJr/F39yTM38iUfx63xNh4cBv/nTSfuPAU6SB07s2
I3VE1DKQ6zocSykbbIK5nph+ZIIncT1ckK3cbCYGg17xkpfLsT4MywvuM7Q7Pr9FyKaIZ9DDYhBA
zYmS9kWd4bLxuQ/DVQdIPljraQ1zeoFqVdOHyCNa2ZZYCqXzINxeOxrKI/glUsox+WOMWit/3s0S
FA0O4BBF0Gk3/K2/C8DM5fVOghB4OkKi3yxjAoMy1aN1gixcbY5xPdOD4NPWo8BVs1TAn5jPwk3d
crY0eox5oP35whHEBHmP3DaIP0Lm7jWL6M0I7ceEUFuXKVIAGuCUaIq1dgAzwPj2zwDWQwQQiCVo
VPsfVP+H8DvmwuzbvYs2RP6HY9KCgUVjd68gNxDMiSHn7q58AbdjR29/EY/pubnv7YoeZKhFY2Hh
LGZcmJ1weAGhG8WzwdP9UxNhq6dLNdDsxVAdwg4e0sscv4b4XIEIEiOHEvY8FOahCJn6RmLrdQLY
oashU8RTZePbQPI7R5StjDc2Xeu9Gfxrs1eaJ9ifAJCmuBd6zWQXsWSnHxj/OiWaftlOt6HDwDoU
GhR8oGLVshyWmjjdoArT6n9wURIpAw6htdntL95418mLmYgLM8hZobSmqnlvQignLRHmGhixP+65
LiMWRfA/EcaBs4nBEv7abTJ7XaFgvMnHBUBz4UxXz/Tjl6VV7pypp4luuCW9so8hhTpi5tKPinLw
FczGiqrX5wWheNqju4hcM98zWGiCsZXQ6x64sPqgxf9RY5wXsXHViwJ21BFm3Nw3whDbAgpgdFAK
sJacK3aBZpT7TZNFz74mvyp4uO8N23p5NsgIoZOXJFebBwIkLbYdg5Xhb222NLBOI+MaytlTNzl+
qT1r4SMJ+7ErK5+9zHC/h8DoHxsfHyzxcXcgpso+XW67d9aBHtlhVVsQ17UErqUO0qDRUTv/EHS3
u8rLhWvNbaNFzmNvshRKIluIYJtqUQCHmCb1XpHETiaNUinK2ul6HWdb5mhcdUz5AZfBz+8IhSj0
xIN60MQxyOtvmwZueyse9vwe3pC/4uWkhvFjcE14VpAEgnM8VDxwRCPlvbuwlKuM85t/cbSPS74L
BwFG/JSlidezOX3BMQpFra1C7l1nQtvt/4v53gDNaAfdMmPaawTt6DH1SHwCNVmgHxxhZX59cR8o
BONJPhsx+cr3DT2dAVin6K2DmXv+sNIuVJzXHd0T+VE61vtXq6fRSzXkBG7lV4lXGJbC5IXynYCe
MktnNbRRqhEkqEzXHK8WyEsxOaseuTBNfXOjaIhg9d2OuNhEfGwROc73yT/qIgjrHXAYXl+xBWU5
FQt5uHRT1Uv9tsEwELOIyYjVdP+iM2TgtJTUDoE8WFgZd9rcIU2UadD5E4zNn+55SWkhqVBxbsqx
SggDx2RQQEBuY8culIHcI8doI6dNCVVYOPqdg48CBRNbGfqIBOMCtxpurFDUrl5wBcZwav4hiAYo
Lmn6yJPWIzsGCEBBTNRhvva0HC9A3MfxHJJREVMdtQVPihn8e+3rtqIYygdD6Qh10DHS6DcFQJms
8+Ohb6r8oQ3oLG8Du9kOD0TEAHweBylMwFUOQ3eZ5enbf27G2XnKtKWgGFTQNFYm0/PkXZMRvX0N
GbS4Qc0ZQT/7Gx/TLeipUBWutb+7caGuKz/9tEb5x0+xvo+Vie4T+hFlK+kGfaZUUvg6EMirUSRb
E1yGulDmezXcvOv0I+9umoV7aVYHNZS4MVeaONFn07OBnSJgoIhYziz25NQNssv3HdqWT4h95PMI
w8npFHazXbFYvZFIsN5ZzBeOSR4749q2Wcg27lSBiuLumRDwLfolNR1s9RfIPsO6V4SKmVw3K2Ct
kOTyhFMcf5+k+4812GYaOwwFqEWtmLFMTMtxGozdpdpqH3IF5wyi8jFbkNaTmRLfJsSJrO1uGKbK
Xjye5/fvO4kPZNhWPMULkDdM1bUd02uS5CuEzIuelPTSgkdEuGKd1KJVuHev3IrVBHM9qTd99IOc
bLSa85/Eh6dlLMbZaa+DJ8g3ldrEUJ1PorWcT4x41kTIGQQ0O9f7PJvnKzBqjrfLYsG4g6YxCTRM
EGIsMdGdw+DNLJglsAaV/MZTeGl/ytiIsCsIecWU5SvnRCf1+XQxzVAVQMNg7W7MNZ6uR5ZZRysq
vtsPV8s1iKrPTOI0bJ9VzDyRgFrgUMmkwgQzdDxUSKe50M0ex+HYc6veHO/jVe7vvs6Zqk4nMNIU
2RFtmEcGY2mI7ZpSUSXbarzqBe6gjOQi0dHNx3PnopKp73ABEckkzwgb4q8DAkc761aj8ZkZ8iTm
kp/rruXHvmUd/ZHIcSOtxLz/r44v+q73ah3BICtEwMEaIQCW4vYrd2J3+vZTsja2g1gEx6leaqRF
qu0GcPDGBUZlN3YPJxP+6rSa1asbbKcP9BwBtPZMwsbCQvjz6ApsaaNZeOP4ORRLJsObj+E+WlNF
bamS5LYUwTp2B8fqcO3olth1MSeBFD7GuQzVK6eEw6i+qHCw54rtuwe5ryG603adbrn/V4OQJo21
rsWkNtmzCAvUhkU29KY7ir8LGVl0KRq7ji04KGDfp1aNQMQARGzkiesjX4CMR5HAXeK8dmbfoyPl
v9UYlH6kz8YpqSEI/F1kybvhSJzOUKIKuJ2lLvCXFnwhdMlnFQv1Ki7xd2eF4HAnfVx3k/UFp60Z
bclGW21CAPt19nTq/WnNhc/c7/NtqJUt/MgkuZF3sNR4Zmue0yFgtZ7tJNEqmhM5QuJCC0MsPJ8f
XOc52bf60MQm9hsEv3o8hLkC4PPs5MhQl3LrQGg/cVlwxBG10FQmARFOnJb48UDFtC+Ya5w8OCLk
47qgIkNG11WR2gSWmzaYeMUyjp1ehIcDbW1zS47QYGerhXCsNDwckR15X/aiSCDLZXWnJiAhDYbf
tSbTRdMXGWoRLalGKauQN7XFDBjUeG+LWXMnKfrduye0Nj6FNj9spjgOqg2JUeqaiaYbjivAsE7z
k35yhbU973QqTHVj3wUYcsyJAjjOJSUYHIP18Wlce1GAzBv+QJ82x6e4uiYamYrPr7IL7MOUBpW5
2I0DEpmthDOUJEl3MC/wmCCue12dkLACWWIBsIIOag+fBVRc5ACxOohtB8Mnhbbmjr1VK6FPw764
2dBViw59KlFDMWyNhoh94eZQGJbnmeSe4JnjH+lVutNNzCKPrLIau/iQtvfwXL6fLjf7aVLmslv/
a17qb6BKjWUaBF4Ud+1deFIogF3XHn55X6CGedw6R4zXNax10tW28mzGNQkJbtqVxEYnGOxVP3+A
0oROfkpwq0/C9R7mPMoA/dz7sonbt0vx53rDp8kNMMDxEQoiU0CY/ap8xcn0uys8XL49yfz/VRsF
e/vVL+T9IEB2Yg5Nt9hrszewugIeIMX4iMxcngxBHuzc2zhX91qOTyV+Ro/vzy4LX/gkj7ugYpIO
ObZkw/EhFv8vj9LCL0PIZwppjGsyYIwWmxYJkjRS2GxxmAn/dstyNQXZZUpHb3FZZa66vUzWvS9x
SIGGdPspnVGSgleAV2P8ImGKv3sPo0/ih7/walyz0nDO9+UjI3iZv9AaBNEUNFk96YO2w3Il8Br5
lLSV55LiSjAK+0sSgyEugTGpDYv9oXk7DOnX3vMDzbH07+HMj1Z1S/9TJ1lf4oFL4H8SxA+z3BqO
CsPclGWEjhXHEUYiFc09P3LMsTNjrIYF7sqDI+MPtB7BiTuwGGWk2LY92uR/K4Hs5G3229SbUMLK
hVip5RhPIyDRDu0OlKxnce3h/cp47mdsvOWKpr+ZRULtMTno7tAQZiYaTGrBRGNmd3AHTwTD87UB
GyGslTd/ep8o1kA91vVhfwAcJENUJSB6uUatc9Uc/WZHXAhJWvs8kWquHySg9BNw2NhFT4KtlGyo
Dm2j/08UqPF1oMWDDaA0YronjlT51OJLTZg4uBYd3Bu2WLHTYLvPgfFE85Pgm85qLWwYh0hNeGDv
3uh9b3f/pHzcmpmD/7ztTCOGmP2i+Fz6em6zpTePIZ81p+ESzZMJ+bvPKhS51MrBd5LpQoDl1ZQy
2x3mqjgFLwQBFqSFBDVZyGQhbfe1o1ey2wyLtfYCGEortspXd1zBj7M9/1/ttYf0Wt/ozY/vqPwG
Pkn9yAbnwA1GxyCCHjWlV8GU5co2SlfBes8nwLRupAh725qH7TBnnfQduEfRX/MO0QikogIAHdtY
VK2ptGdQsv+wj5CnMXOZS1KFg28YDBiLNQvU/O0LsprvYfs1K8jHnSpemhl0YfLH6BttsNXcLYsi
ka40CLrp5eTkTINPpDkKitPSbZF5Y2PfYZ1wIk6YmZthwwiq38WjxZSmGHnnSBYQxvpd+2tol9gw
hml2Rl3m6PZzWuQfdZr8/eGYDSWN5jD50zJChuooNe+I1Ei3wuCMMtaMsLTNPzQxPBqM2Brtvt5U
pIJ3yKe8psR8H139/agiJ7TFBrEdATEATIcx7niU3yByzXlUklEJ325fQjxfcje/+mWGi0FPEvRQ
DFeIaQWsJZfNJPaycwNakY+LUn7+2vFIXbT3/xKaN+fX8yu41jyPUP4AqilUFvAfCXPYLu7kjmHR
rhGrPSpJoECJySXLCTLdnK7agPSmQmi1QVBgKHfQjWTejrpTwwQbzBwf7Z4bdkRr3zPz6D+Fmn5R
ioDuIrZ2HWoUIxn8IYgjD+G/5JH5zm3Mvy6BRjo2AAVvMFcrWc+2tcuvZd15apdM+2NxTv1IdfrA
sFHTGsN11P6TodnEkuxkTZPtuSMLNWyblMTrPq+TPh3VqlbY4XI+uK60jDcd3EC6egW9ovef17Ij
5Aob+137CQmw9C8dFhid9XO2bOdNSLzN2inov+buDHjSzZa2ErSKlayLRmNkOIsVkF5rXIZILiyP
RwnG5R3gh9GSO1k5kKENKBvXuG76Yzy6AnNHjV9ThVG/Qd30jN9lN5zlnlkr+uVvDpZ4THHEDlK+
WzYu8d//UddMzAZVGZXS9wWG/pks2QX1jNlQaNNDoTEmX/4cFK/KZOXPa/uGHAlpy8NzWE71w5Q0
Lf1Go4SESWRp9VPm3Rb1+Y/n9zhOp11lZK4EdmgNJAF0A8ZW+uKVZBIa/v5DUGoZeu0x0WpjBP8j
tFvD7G9m3myE+8HOEuTEoQyUlzcBpQt7YYxYS5LcL0x+bZykFlZTs+6Mt6ONVn1WFgxpP5fSsDOm
8tNUYg6UJxeM9HxxAXwTP5b2U8jLKyakWgQBSAOlDQA3W7HZ6knN1KMNCRZcUa3wL6zpqFYES8Wb
CocD/trQRLKHrncMdQ1O9tCzOEXEiep/z8584y0urQzIhR4ecIwpP+P89FqoVaFyKBn7RHf+uBmu
inTnuuSoLDpWRcLDJ9Xbc3jqDiESrfQqzlxRQ5x7Cf7MtpTGtyKJEh2Ir532zFIo0045WEcCG5Ye
5aYkf5V60myupqRtIsdEkNCz8wWDVPNm9nBKfUwToLfy2JKY0rJZpIjDpUFL73nAUyZEiA7CPbLL
ugG28FX9ctMzYr2mA5U0tYtqc7bS/X0hCuuOayrsQrn4H0X0xrf3zBkBPfpjgGRHTYWcUzrEpTgm
GULTEQNLziWWr/hCJzFYaY8YmGxpT18kahlEzzi6B5uPtb4FhyOlJBFl+hPxFpZJi1GfotI/NVQH
autW2Syv2fccCsxozrrxH6I5A68HJe/lQnTj3SvyWwmV78GQlZb+Jk61uxs8/JzH1ywhD1Qf5nW1
7VaWJgQ88b5UGJX8wIdLC+hH4pTwF5g/AWd756QRopVxTEsXahUFtX14nPmEpdRaCPcflD036xhY
lgfFN3ofgckFFkcg/f1hyO+MgZVDoit/VBFy1wNL/h9QyR+8ym5AnWhi98xDDCD5rLFTOTxCfdMX
p6aR9PERkUk1bKBfP+Umqd5Tu4mNaLoEOFfSVBrszKshaCeBbPXnhTo0JGoSZg4Hj+arFk968Bvw
Z8sePsmm36Q0SeyCF/dVgMJZauvLHvxyxKACP9M1ZScaLlS6YbMLeZfPAxBFBMbYS1YCaG3Qcmew
r/PjgnUtq4QZA08dDwPbKrp1esD6RUMbLC+rQuN9ubZ29vIwe86zaRtmwnrvBWepUK9uBHJ94Mig
1z1ZZn+ldjf1VN46duKBzUb0Dt3dQ/S84Ti1MqN+3cu+7doV94S+3VoCEdjp7IEAo2gpCSNpAAmU
c7oHjRY+tpG5hvZky5KQq53pTvgIhnN/6kJwkBO3fVjCRt5Ixij7hjuCItmM0Y+LcX76BbRk68p9
HaX532Qu/iFLOgMN6q+/RyeiXRxkhMILG5tnwSSQ21kxw2c7jcm7wxxOsK13JG9A+9VMKc0hDb/o
BHQfrM9hl+iME5QVdVUO07FSp3msZJgJOneQOGgKw02TRP/hkpNnAn2jfCFlCmmKXlkBHUPir4s2
64NhHC3SXrPNVkfPp7bHkYSZKCiLOce9Lu++qiS0LC4oZqu7p5FU2w7xxbZSudK973EzjiW5FyAa
pMYEuY3yNwEbPuC8pknm48JYU7Bie7MeO80hOziVB54Fbx1p1qx1TnYRmadAUSneioJWSiv1NmJO
OWwZ+GZLd2UMxsio8HCw4rlRFsNpsTa3AZg4WjtlBwJujIhRlFFCFA7D69JiigH79+ljLDNw1/Vd
KcuXsUftXnYOlqjHlnTe4IXlO5p3h03ochgRaJRAosbmUbeKAwJ89J/Or9x86kIR9p/yoQntY6dE
L37OSWkr95eYKvDEIG/JtAT5xZywdFjF6mNM7IhXZcwmrUIT/XNm7VFhuICTN2RbdZwB09GXq7IK
Ph/H7Y6Ved+3YMEPUD5n70sWWssxyq0g40AJ+lKU0tFOqshJeHa5bJWnetuu1AnQ/peaoUMJb8NA
CUxtU6OLRNGxufe95jDsP+NiFGoOBPpwAmfX2zqATzwzoHmq3tcf0fW0YF8pX5d/EcfdKeY/6K7H
Lx7xOBXWFbfNi42YqkB9qw11HdSE0/Yit6VjdG9NT+fZiDaNdR6oWsBSV1Yuwoo3ODzE7SgiKV2k
doGSQ3PJ0GK5T9XTlbEgI/lLIi4KpuYuOZlH9xqp4Aw2zQIy/krpzoaq1rVBjydGGhwc0xJjxAhb
Dzq5mKYkgSNc/C/XF3lu2J4jn4R6uoKfhdOkSak0WC/cR/2vECpWeXjQo/bPUkoMcDYwpT5P2dC3
BTZ/4gDC/D9ExNTHB93oAkjhteJ56K948AyipCrToAkZCyL6rRQ+UsVRK8oZaNb1YOTB6UrNeiZq
oVTZabgKk4ZCLNwDvLfxIEHdooBd3tsSVYu29COlMRYgBsckyxUxivr1lPrzUW+AQL6pKb+pSrO/
qcPekIriAJZ6Xm91L403IHIJPOHqvOZHKh2d/nldDBiyb8GBVyBiXcRqRzA4EPIYNzOOxxImOMWM
8Dfln72+oaxaX3EkqwKgxtknRrtYqtvwVuN5DBWR5tVr17w1j/b4NAWgUWYIN3bFZxe4zO6sL79Z
TDAkf1/40LlL+Nt+tbbig20axScD8ZKxfjIrE1jTK/ygkMrncb8vpgoECEKD6lZ0QjM14irfPOXm
iTtjXqhLneJBlhgWioX5KRWgn1NKK8kx0nnNlphN/NuXAkDTdikRBDZJbL+GoT4M3MerRuA0RNAL
TmJ7YQhue3qeKj5xwXkwFLlhujkMY7HrBmUzCt9/IKsvkww8ayxsFVqobTY/AuQwjvJfDDv4PH7F
Lg5AWBHpUJmcJVrQSQqgsdx8UELJSGrZJ7QGdkGceoOz3/2j9WlSyGZyOMxg1ewbVfwqWzM9a/FC
B3Me1MYj6RF/Uh9d99ufhwUpsxRMbth338zLGH2ItmBQCy+qrOeGIDuehk1tbvDPdVIWsHTM5mhk
tH8qzDIZOwyytI3FKFwzKVFY3pjeaOdi9/JapQ0/I57tjmCZbYzrSTiSAOkYTZ8Kq28vSuS/fNKu
amKGsdGe6fuvEU/o0GZZBzCuI3o03BhDWgkywpVIFHJF5PDbVrQY8M1Azo5w+wUHTqLTl/YErM5h
kXrmzwYurdUti0/RVMfPBtwx6EO/rrPlJ9Lxj1XhwnlTvzo5VI/WjFu0K3z+2tU93793ONRrocoT
51tbO5BzxA4sBk7cXxa4xxKQR5DZyZHjqfHCjAgLWV28+Eel4hZa+MCnUjHs3A68floNThU8yuyh
1iH9AS2BF7jtfbba93l4uEccg3zb5frh9od4934VmCsWtFiGye0rfCA6+TS+rEEk8qtj4uMYjFrx
8mNS4qSuSkHD0G4AtWGzXrQGXTZL5tKPSkYMzqPyx4CdGk8u/cMWnWEM8ar5E7AvydeSooN/KKQd
JU5mhCD091MHV2sxlo/PTfAUQMF5l97laGA08MO8mz8t5pHxMWocyyzA/VnGlHQpPUmGsAy/RY/V
nYm8LxjGFpECbGt7DxX9VsitQ6Wt3n3W6IyZ8ogk35irswtYHYqAmRrNpibxLhyJ5MyBaqsrhUMH
je6sU9AeXT/WOJLb/to4BS+DJm4+L2OdJ17g9yziYp2zQS3z5VEO/kSSLnvYSNMNmQtwqWxy+jXE
DenyJennVyVYwiEPuvWuX/T/RYavCNTqQswtJWJIqFNbIafD7WBTJtI4J6aSQ/xMOo5jgctVhcD6
YOZux3TG3X/Z41I8RFeKJ+7FXhTlL2OurZfjwdt2qRf2doUVjLGsNrOWyzkHKtpVs65Nryr1fqHg
J6TxDgG2Gac2uzQcgXBT+t7mHtVu7g0cBlvby+J71GlFRAiZJ/czpXVB59eJ1tm0Fzx1wXSa3Agj
OGG8n1zXcRBVhPxx6GosW1P7t4JOEoYpf64ajUI1mcLJ4n6sOIicK/z419yavxPBf6uXQIdb04Rh
EIRtfeRy98c0V7HBbTJ9v/CAUvj79iBMurayl85QLxCdbLhOHh9lUqnFwrvuJQbB7gLudXq8h4et
NvyReOAEN6dmNpK2lcTdhfwdqcYY+6+Ncqf/qCrzqkewxVYop2v9s3LGcjWLoKXrfD4+iDnfoH3H
5jFNUvN/oCrKzlbGT2klF0JXACep5/4uimj+QHcfr1EMzLul3/ZbbZcIUniQf1KeFHvQiQtzwTWo
d4Phtw9JXOuUQvabg9JKJkWN+Bjjo1yChHXAXhmqr9LuYnqLyxbXTj0PM3lFbHiXEdpZraAj8F4r
iOy2qIYW1ecR1pCP1OPIR+ueJsacR76Ol/DKvwbNZZwHC9zpga+TDbl8DEqgrtY4FAGWS5Bj+YBc
m3K/ZRivriOKcvodUiJw8i82yGy3srzTXUEIzE4+ZCMfpSqX1j46/w4bfkVKc2XdBAabkloyWqc4
wm2LhPIqxru0y7C8IY32Lq/Qtv0IjmHe1nzvkpot9XjEldwuRQLwYU0ZAxMSk/P80+KRAqKbjiBF
hpHIYnVqYYVqR3WUCIjjvjZs9Oh567muFg7cH+7Rk6fQ5AiOTrX/HNpvefEYr+sSrIZiHWUjfjED
Qd19aFEhZYqX5oAGq0ktbSL3j++1FzSemSsXwjtRoB5uuoaS8nWBnq1O6jB2jWi11sl8+zq13eK7
aGTdnsxjEZMXLbN1XPJSEpN/3I4bqfq8VVSuvDwbEKWlUFhfChSRmBw69QHDZU1HVFNUMnviN4q6
4R6hHgv1YQudgxjnFX1HjEpXLsZeWd6+Tyj3aPKL4trjA1svW7NUIhBNd6tnsILOI5cZoJ/SWwDU
3cAAbFBCZ3lg2N2frC79n3Z/QnJ5LwmiwUxqxtrm8MYEs11mLfcA5fEjOIWL3o2f1cT85I2RZT1V
0bTNs0ss6ZIm0Qi21e5JOkbVvy59r/saf6I+U5Ppc1U2R/sDArOB/ueYqLJ66FsdQ9h4dXvgnrmf
5j8aMompgFIh/L2Yn2AGHlnmqXnsn/weg2AQpRzBr3ohQA689+WQWfKMk226LuDx1hG4RX1L2z9D
qngEUlc7UHpNKLc9SeQJqSOvwuc5mijN4tv8yCQ7bgcAUxkjExA5/8LzJ1HBZPzD+hcmtyDzoDE9
XzVfhAm4b4nutsZZGkAmnBeCWtf/6Hrm8itBBI/f4dHaIwa2Qu83L+V8qzoVLsuNiO/drFNic9tN
NnWaNgZWiCYbivHCRtHQX3i0Nk7hsGNMBdLAZ4SqKASUlNWFyj3eUkA5Z21ciVw3m8ZV46LM+kLx
1b9k7YhZRQLL77Q5aoy3eSFv6mrPRvL1ZSX/HG8nt43wddaK03nTC7soKId9lQRqeBK4ovg+oNAo
DHooHO6De2ZLaAnXp8H4+mftdIm20yrikLqcUXC+1RI8zbU7cAKdP7H5oBYeNCT7iJCL2SBpiceN
ikMFdwVp9dJzzTGllWAzGY6hmxHlW+Vm9OtL9HM3K4p70VAVoZSGgjFPnqa1WeEy52ozc8y/hRhT
j6Eaw/etWPhxlGFaSLGBe3M3ZvlASYwHHNbTFzngQ973C1UTRVGxyiBnk7AJGwUoXwNUJ2m671gQ
EwHQMM+KS64GBLjiTTd8LNn6TfDtkrNteaDK6wdclG/AijvxVJj2yk8+MdF4vzCbp1JuHw84y4gy
FzrXUBrJLLm8GUZziiJthqeVjGoln9Plkewog0vpE+sF0XWcNadp7ia3L7qSVnkuupnJ5pnoyYdq
+vfNUGrBnEEQ15f7PQzklmtUM63TOU47PbVAJfFJLbXfXiMpW3i+oGCt+wC1FbdfR/qXs1iyHduR
SfroRtz4MJcbC05B6X0AnIzVAdOkusYGO/SAIAwM6+HIsS1Dgsdih47IuFVyaGvCSbbM4sCHlPbF
E3o2krpbecaYm2nCasK10ToegWVIiBspeQN/zBN5RMWE+FF2wdU31WX9jZC7hLQ58QrQ1eXwj8RK
YZex4oMxKJy/O403DXhsQcK9ixplxTQNZhd0mnb/Ew3NgqcWbHykGfvy5qGMEV05npfeYbwE4pub
uq9paTBh3+i6rR9XDEAsstgrWxDnmQMVr7Vvq3uUCfAXJJ3dyccXh25yBBoYVkbNfl9gJrmzz/x0
wG3Z3vnAmVDwptEmcKrCox8HT2KVDrEQRvOzlxwQ6tvsqVQrM73kwLg2iODPp7/o9HZU+W3lnXFA
wptndU53ml09Wk9GHwfXQmuhwczx6obkoc6bOAsWiIboSdxjwGTdrF+ANN5tlqHv8Due0lqAC/Q3
mLvKrbPCZzjPvl8kf+sAoUmLtXdFS0qFnwypEJoULyjoaFx8zWWmVtdn8n7BLArgIn9Ey53ZEH8R
fnTU4up+EhkjS66d4cGrV/OsS414U32P+u330Izsx967TxUJUJ1zLW07jm/rnBEv+Ui9eg+qFiNp
OTlIvd5g6T2nuJAkGD9zCAcf1G5rnmzghkX5FtcRCsO/nVCxx3Fm8CZSYXlmFwqvEgIo5h6ZtYU5
OFxgFnSRSTXVXY4BljSMwACxaGwWcN7j4guOkYjFka6n3VYGDveyxNvBLyXo5cTyR3airxTbsgGC
e9Djgf2RQn3K8wPCCzuK3CyecuczHQzirqaf5DQ+uo28bEhnqMpWjObP39byza4E5lUbd85By3GG
r37dk6lYLuY+0A/VCq5oNLKuLrGds3s35eTTHcr26ColfhtCnDpu2jjmTqi7i19D/1wXmlWo/HZl
TpXlTLpSx1UALHsyQFg6ICy7egdQUjII1epBodhDc8aaO7Z9vdVaU0ORnpFIEhilhIPI7H+VuEU9
ZbbOEc78aRcYruR47GTE/ZFO/Itvs+ZLwnRjrLT6aVrH9wZi50iNp+ipTvXGssUgJ28fnckVhhX7
JGil3fZeVsNIoskCKbYR8pOOpx6qCCmZf/WOE8tfHnWn9R5nq7pZFb49EAdgCl0iPKsYlWhXEAsV
DKy8ZGsRXfkVD+YhRbz5BAF/LkGH82FR/sYJ3Qy/EVjNmYauDBHIUCNnlNOOli1+Zy1744uNqqi9
0rFuFj/TLDCCI9e+mCaaTjbGVykaNpsGaASr0Ul+G+Dm3IgsMmyDrq27k1C2VW6QuUUsSGNJupcw
R2vuzGTLdm6Q7b37HgdPjiy72ufobkVuxkcNcA6jBWnu12OmcBJ8mC32V3J9rJn5yw+Q7NM0wgQq
O5crDyPExfeGIC4tzLmgy71dgegPbtEmM9hsX/HIhoPkdj++ta4M59SX7PbXT8yy/Tt30JZ7UBcQ
prPLVjX4bATdVXoMvwA4/EM0WL1d3Hs5MTzv01aYGiIRXt6RanqqS3kzViM+Zh/03TXcf1rH2jz0
r3gRucj3yQPTqFZoXU/Qm0Sj4eo0iowFl+y+sTG7KsNbdUNvHUHxxjzNIpwVi7zEMXcndeoLfBmK
WxTXbGARVMAjMrN0x3a/mXJZeDpUfiaQ//qTabqsrM+DuexWlcmChA+pa/nGS+erBZN7kBT1ZJwC
GM3B1C2YG0edhFpeSDzODU5cQxc96XLMEpk3K4FOoBr8KrFkEztTsp4lR83K0EuC2K/BZpV6oz6H
NpwupDtNyPcWTAjvqQnyDC1nerDfS9A5xI6Ln34fpIbGZNEr6WwSFWnYbR8R2GvvYIcNKOE+aen7
eJRqzrhk46+uudylBEHnNG/M5Qooz7Cs3DQf1486FseYdAnT1mvxaE/pVm4G2i2EbGhWYOdJl6o+
/CnAhq+iPRfVfeYeki8l/8oiHqyuIKNu3xA85iEObjGhfjj84DgyOXybzv0W/v/f6cOZMKzO97G2
MGBSsEGmRFQh7ZkSyyyZzhCju9o0LA03Vqoy8m1qaKPnC+hYeIcSIppmrs2BuiIe4feYWKIIohlr
aL/9zdguT9GHZlxvxejBawmpDyaZjyjDrfeMypziHZujhdMG7GZyCLWbYR6aetBpVhAjRr0/mLvy
pZ63aJm216mVIxkjtn0LQXTzMN6e6mfUQIOZ75qOWg++ijXbkYgf5Vyea6mK+DayAkQJNjT++Wvr
8AmXzBUx4AR6J/IXMt+AjczvhpH4D5qE7zy/i3tFLsR0y5BDaE8CBsYblX2OBwc3PS6Ftq8UAeTa
m5tbjTa/xoJdf37P8kRyHY5MtlwDRhvGqT8j09Jv8m0FlPiBKfT9FYeSZVM/0Pdli4u0sRBSAgzB
BEl3lFRJgkfqadUmQPNloPosYUNPU2to97ZpwJxK9NISVPN8RhqjNwkQ6yH1O1bLKmiScyKjY0YJ
g3WkNn/oQoRenYc7D9aRb8eeLJ8smNTqkmyvFoEBX1xyIf1nN/dvokFWmBzEpxB1ScQTECGznR6l
3P9a33P8AupxG7dehpnBcfLia7kTQ91TkeY0CH8jYkm5ugD7UWbRUMCfXHPRVfHFc5k6l5or0Qk+
hQ1pv4TC6+jmJy/BomJpGErlwtyVRXra/Yv5vuz3tqUeSWD0PdEZtNsEZn0E/bWAw5jYXza/Wplf
g6ixTZsv/Evi32WGjEpFv2uSwGUPDp7WJ1d9vR2ZTv2AsNud9bGpVWgLhgYhOg+C8Dd88BvD4LjH
7q7OkD2WEJI2q/N03M/Y+TPi3bB+GqddSkfDeR299s/GOBKaaEyuYDZghfCFwIWDCVTEDcnGKrFy
pw3P3gAnDWEasp6vZYFA/qqeVy0qhHXCB8V9fXoVSMvU2hBQW8TI9Ate4gpjLwbjQF2OeTCEWReZ
eqfHT02cNvEKmCV0+lpQApvJBZVOcc9WXyQIQAlrWI8cH7BRrxXH3hGxkWcGIRGPx+Pet5VKMK5x
Q14snLsM1s/e8SH4JIolHLmL9InXalfJzaWI2p6irb45VOM9nTnU8OHvQxFM4qRv3vJHV0jUszqe
bXHwh2pUDLY0jhtJebg5xZQEggpiRBUGWO0ikXhAENmsPNRiMSdm6sAgBMDNJcUa26Cyhr3Zlova
vi8U6rnRuNSVhNNisb8iTm/9yLSR1fpICQq+KGMzFQG/MVgn/sM3ESrd/ObR2JErjQ3gjJH/XUgK
Sflg2/BdxwNaLzulFUy0ISkCRRc2Q7Z39gEExH2f399bj4wWAZ2QZZ5eVgZGpsOuKNwkLgpkrmt9
tO59PwsVK5BxCxUGLIDQoXp5TCIcyJv9ti1HQCcqAt4mctfBVtOSl6ZXQ0W2O9Ivu52Xl56evhab
xJ4Zthkt7tFuNItj/PMgdEWfoCKkq4t0ff8A2Bp/njnADUXuoEu8I+jnEDHlBRjjuK8PAMzbQiUH
4nc6RptyPnBC5G9Vxp+Yhy418TYdRZutApuhVIF/ODzzCN7Zkr4ZOQypatRpgF44uorL9TGo+t88
LtKZj3TlO+pRlpkxyojlkRenA7n6/UjGCXH7FxpSLd9OXxskHNAkNQ5ywQWX3rZUYVrrkWiTv922
4Yje/lK08AV2Wiqhhu6VP5SdWBR4zlxOCP3mrjsH4eY5GEM+qipCtQGxA+ACfGNb9VW/C6qHcGn9
aQSruU0lUdAubsb5Yj1i8EpEs1MTziCODdXS/x4xVil5Xn2RsXZEaHx8PMLMeWd7w6iZ4yiM574Y
OWCkG9qYK8TDttHLWl3RmPEhGJYnCQXKLGKtQHAEmTH/JAGc7jcJ2pxrXowUKyu7grCB0IME/cnR
CwPypC9FaxxHY7nWWRMhiXr+7Y+SffwMxecGd+MyKjV0l+QsmMr8zSTCufsVSgeAKnCX2gUw8mah
9DDph5rCFnIlWI+6zjkNiMQGydNToHAX9cgv+d9hInyaPlF3Sx0/UUJZypGCnOFErWofpgrpGoKd
bKNrWQ7Ow0H/Rl/UuzVA4QiJkymBxL9fQPRRLNUJFAL96Nt2TCgbfFan8ep+HV8HmmE+y9vhTRTw
etJDmf6DL138mr9iTtr2InqydeYXVAxYPIZBaqv92w01iqW4Qa5Qic0kRWsECwxJN8xBoS0KSqXQ
KJsMpuBf24BPxoGfVxvGF8qXdSseOy9f6RpIBniQGImkpCHovnlYMvXtyc4jqdUbpvhuWNKpEiok
05LAD6QkMYfhrscCwSFlSfD+0pGeVk1q9og83EF3yK3tpMesDPJWjB6XMWBTou6hSC1nNBmn/zOW
cZ5Zc2MZ6/e5F5EROHUuIWxSuoxahNu6B7nqA7hTEn0jOKdaC1QLY+SzkEayC6g+7YZp20cgKi8a
Hl7A3z7cZAIulyMUAll0WNMsGO9mBhUjgR5BRm9sDxboYAbSHSsB6260KCbtaBQjk0ygwcYURMiL
9KEym5i2heRK7g7mMtfJ4Wdc/BEoBKHKhsZQSiOVDV8qE+YDGWEcXqZ17c7wv7DURg+4UC4IKmRL
ul9isX9Iw9oeNzcE8dTPwLL+ThhhPBVgcHjqFqxoLemzj5vV5ZstehLMjf5kiI49Yas98dt2AH95
fmYQItKF54J1smLJsKfiLOGM7MvxhZWPSZ8haoD7q7OgfWAZ8Xp5K3RqUzXefYsMgkHMEm/shrGk
xBzG8o4SId1RqBG3KScJxST9spOKtCwTjyyQFowhu9urazDJol0wx5S+b4c0OTgvTJZ57gA/dKD/
p5R5+tHzGOigbVn8p3QBdjwVJrbgpIYzEKRZTMzJva8JCpg4YO7/D6WLd9i2drqdvQzBSgiNerc2
/COmjwhve4l1u5JIYh2q/vQeOGiivfQV8GwSeDUEyA9BK0Oj9e6/ggGtzu6PGVZW+Fw8xDYij5FY
/JUPuLZaqS5jtaigtu6qk0KrbTq7bc0vTppT2ikdUg36PYHd9NkiQWBigfOTD51SXo/bueFewEce
60j/AuhYYeIo1U6VQnilWhbaKFS3oLOBPLQr45zOyVt5Nv22lZmaOFddQqDWAPF6JYPGwTfullOj
VMt38nsOHMzj58FI+4EgmP4m9nl+qfw7cVrkJN1XtE8qHAOHHugqO3deZ332c707w2Ico7MiXOAw
+G4TcgrsicIS8efVSFPe+jVh5jBwG8cbnaDsiqflVbvX6kgFs6rnHOq6g1cGb4X0rxEBVOb5FUgc
QTVZerOM/rz+rlYtsX6cvbJbL8WX1WbxBVyPC1RSsM/4cYAD5RSvo44THloak7XDUurZUDi3Jgm+
4LiMaR/bQFO1rJzrkV85K2eXJMtz8SqLP+eU9dVulDtSgOHhMQjwcdhVmYvKOjTAUUxFTIevnJwp
QgCZTCBZCnw/bSbFyPXd7/eOuw5RkndGrIoURBlV1Azu3DXJbwjfqiMc1tNtOkd9KyWo1XHMscBv
pNrH0GLY5sNG1BRakgA/d8qEi16urShxCGRNrH4vpxBEWKTOyLZeKnKBpsXM5ivz4wf9BPnW0OsF
3gICztw9hwunqCO54mOdjO2XuNHfDj4u0xunSP8w5mKv74R3aX/oak8DlnICCaXRTmOk0qaCxHg5
ami3BhS5gFLfAgooxO1roMRemOqclzNLtietGnwg3OKL0HgMNiKQTz+W1AYQhp+aVaJJ6DWSuUGB
txp8plC0OPK2CTljR6AmWpF/5KvV36lY7kAJZnRHLjBpfrtHuKF62WQbPIyP0gdIyLLzVTpwJH8C
ZXM234O1DRCE3Cveel0hzYt4u353sCNieDahiWoQGYynUodUCSsm5PMIj4+FsxDbyUVXroe7zfRH
txGxhoFqRrftRuNjICRcZ9UTtwxVJl+YtTO8PevXlG6fa8PImDgEnM61kj8SHjOfQWmmHycdGlnm
AXMKEx4URX1tuH9pA5+57lqrf1/54HXdZarhpzrtP9cocJgmKJ8+YitQ7aiLydGuxch44lDIZrYL
kUPF7RjV+puR9bfFmvDMHAbfNEqHgWNvBLnXi16HTcBoLcyIcZIodz/5jlOlUtugyvUla+oExogc
h9dQa+ODwc/KjXuxcClUL0HH/h8ONzJCnxvlBZWpjYLlIMdxgMzcqxocPYI7RA9hTvTd1z+jnYm5
ugwpOEFngKTvJnjaqpUW/YPiC3/ZHEUzZsq191OdXF0nEuLXpulM4cInguwZmZF+Sd0I6od9gLvx
5UMy1nHXhl4/KLMDMs2cyhvNb54BNRCq1ZpLdKnF834b7lzoYjgZ/btUJuZvfpG8cads8d1qf1Xe
wtn5mQNHdcdZQQ4ZU4M8y/2mSslXyZaiUNzYuelRY9Nrj/ZV/riZgGzh1Cp2HasI4OaerClkA/Pc
MubOFW4J6wN9BHhxZaZwzqAFISaH9+m+0rMcbFuc+HnYwXHnFr76CNrC8M6IlnfWZ7jvDrfj89Hb
IWl6ewDaU9km94uuUt0TpAtniAmLfgQIxwLcosGznMAZzbhTQuESJYy1mXa7yVNWlacy4v+UexNb
ZuMkW7ToK3wqQ/qdxihp2jdb987sUm+UOHS/wwuq28aOdNC4igFnszx8fXgLhZ/TC4Yscs51mZqf
OlSLjp1jkqaA8gk2ZaY9ejbSM7uWQWdSPceQiIpe0BifGzcYSzxX2TvzlPwBNL8TmiM2jx37qcne
KNQJayU3qfFxHzhers2eoJlnPLgjKjBlSao8CDJyUPfw0+5RxZ2l4y9GiE5d6m1bg86rjBRekgvu
EG7QEkSxzSIT5OCU4/rfZFvIRCwrMYtinM4gXs34pT4vg8aZ+fC9BBkYL9HN9gv1eYqEQmlCe9xF
2TIHk0k5QOlBaTWMd023BKH2FzwhDTv+AThqUv90LCSnDfiv92keeyJSr7Cz5j4v5UwUAw3DUN2p
PUqf0f6DVsDzOf3cemgaSYVHAtkLgO3mGGDSRzz3kFG8+TUHcgM94cNn7Bfd0wUuwX2KyJm4P5QP
RAkY0lTGobbdCIV1h+Zk/NAZmDLgLlusjwzqEnEBWa4O4UDkFHNYH3nsRT2jh7mp2jsXTRaYd6mi
5ImKRcRcLDBkodc6tFpjbpCM99Y1jo76z7B0kKWZat69Y7biHxdE94bClFR+OZ+kPeCRJNmQ/0RB
BnngHqqfKjyVQyVJVpvpj/dx+opy2YCOmbWMquP3JRu69XGOjoY4us3naahEjongwPQNG8EZQc08
3jlOydHM6+Mru2JsK3Pv1fo/259XeCeOj8HuslC7tEEkEEAouyddSw9l7BtD8x3NJlgZaSe3t60r
XH3Wqnrq8Q3amI/7hrLZyMAulyFnDcDCyelPIVjalfWFJq2BnaYtB7Dc0BvXqNM5jpN3+mll4Hsy
R3ccAKa3PHkSwiok68UbdJmGPnxv9IGkZC9JF58Wbnep/Z10OfgaWgqwjo0KXD+71CX+DIpq5WVb
uWDSLeBp3q4ztF56YpMlMl7xiKtdfB5rOyR2wXOYlFBGHuX3GcW5FgxTqT9jUw2yU0VsjOR57fKH
P4fnqAkIcjmjQh6Vt9YBOFu4fUIQnuYTIN0qZyfZ/GJy1ixBzYxNUyiz3kNWF642AXKBmwLmRn3j
6XpKMcDxxVvms4ZF0jKzLK7iswWZT6mQK2wE3DoIS2eY42c2bEV/GND/UKhnrmVFzcwHN6muj5gS
EJ43yYi0BdescHKjwvW33RO8adif/laRtTWOoc+OtP+cHDfbOw38JCgw8dowssX2L9d8OU2Vrjfd
PLynqr/bT5LoAJFNwAMoXbkcf80wr1PbF93EIXER6ZBJQTQz+rNnyVWfe2XSKT9wonpaNnmq9BkN
UthOlg8utBbMvILJNws8CHv0JmdWEcfc4z81lr6VTkptgkC4Dz/ufzIR+/BA4sXVHq+qQf261HPB
OeSLrTnQ6GzP16bLihPSmHBngcxWDEWctvzAjcuqrIjM82SgoQ4yTCOIlP/2pSFpTVGYtm4rKiic
qFjhciT1bfx63j7yhSgbzX840d8a4g4apEh9fm7Qa6BpOP/tE2Y+UKJ27emeFpxwp0alDW/a/XAA
bml9iUhlRhJ0+HgW8V7ecruIvUAYoUZLlrVY1C1KwjRmgxjp7ePIZbDn3H/ggnHFq7qIdDstv/WZ
DKBozfZ7PqsBE49G9bLH+9ucZe0wkoMU+flRBkCF6wzoS96hQzEtTXLNaW+j31jTHwaS4wMdMcRW
JnrLiYRp2f0E63NDXrWCYYxvpB3g6m7JHyxhmaM91eA5NyYQ50e1RZQwy4OWzDYUSCylYTSnAuj9
fKXs1kG4wAuypuUd+m5Q4MuE2DV+WlA2Us/Ro5eq6sY36Brq8VMMhKuRDrG4U8N4WLJqm9Vf1a0h
LKF14B5hixT1jmM8hwyrTKoi0yncBYo5DU0IHVbrjuZYHun3AupwaFkbO12IJFjM3mAqi2oyapIK
4gLlXneVTbgIJa7u0jHhqXegAlyCI8eYTY9wB52177Txsn6VpD1od7nzd12jpaLngbN/RrVr/uUL
ZcYkrABO4itJLHhAi885KC5FUi99b8A8pRB1PGTRnvNtQMEupk1stXsgIqrGqdrPIXvCzl2J1rEj
UVIis5MoM/pnnzwrrQvvokpdFnEMmWnJd2tNk5oj/7TbnAyYWPrdaRtCCk4YyF6zvXjYBCuzy2tv
nkOK8SzJ3pluiBFhM52+fdkhIDMvin4Jan6t+RPR157rdOpMRtQw6nsBYG3eU29aKeFY8UqdGJSm
jOKC93ZeWyUcFX+4ualgNUDhPtQxf8L21D+dOlSNpKDwQMYnxqixpfKXpnUspQCwPV+sR1a1o8zp
MhaUayja4UpE8+jH0q393dMLjlpf3tnDiBCKK2V4uTiVTWfJLjnWsQwMQ0CfRRMUdWX/XLlHgOP2
Xy1cSeJZdyPkBH1EAaOjoLHh8uiaJh2CFbp6WXyaPEN/vo1Akbx/glTBWS2LDr3+A6uvHTSIE0Q3
zMso3h6k29yeU3JT28bgH2A84UXBnnQIDQYMwJw/aqqURSIZTqTSq24HT39/bxKpba/MUvYnIOjx
xSDkQDwIAWpozoQYj8v228xMpltnUeZcJWtTpdNf+hvlJxJGD/40dmnqWQCPYCCbx2HCtK49e8I/
caZIRevard1+t5QqX3XODQ7J87l0a3r2znqTv7rXyDxf8NfKx31R+q5horL/xK+efTb2GgSDk8Ak
EUBo8+TDEnujTQaJZUGUvEBBeKPDWC/+UKU9GqbJsyD/04aSWMM5pyi3Jk3hENLt/ut2sPUwOiLb
U2Qiz/UwljtuH+lKOAWqVN70vrZnUPhuVodD8OxEb1k6bvsm3F11mbvviV9DkcIgyDpnd6bqA7VN
tNXjMs0NQ+qH3Xz46uD4aSBg1NYRt2SwV7e24Vd/Ku6e6kQ35dTOPswKMP2AG9bulGao3zNuO47v
NiUOGyQFzTeaUzDr2zzBSsKGZaWl0iVgZj12rodNMmrSPN3z+Q7WYabzdN9C5FigCZzWS/YCRtYk
w7DGmivUuml1AQIlRjavifonRuvGD92ysthKv2wUpLWFsAYxpUSd7N4bY6DhGuTlQVDuVPn4DzCt
xrORGc778r1ek5gZUdBImQYIZGe6fgAEy5LLuVWYUadYq4bP0E05dgbiHw8W0AA5jKp49Jr8Rcel
tAvCqZb9Jw5mjfUfKXoLXm6X4ryWL8d+2k6H7mTriwrsDQYPAOCs/v1xNN3xXlGRDhXX9Y8VDqu6
nsxllKlImgFsAIl5X2n3GfRtLrlfM82zq0Od/L0K4AIWTPmUnWCZ+wHT108pnPGbz8Btn6z4koys
hdu//64GdT2hfhl+KdBgpimn4iiAHvHQWn6b82uQYUkTHfGT/idaKDMVkHWyFnysAwJxxxqwC58/
sqYnNBVPcnOTxzc8jGr16RZ9iAi9696cI7TZgMjuq4smuzno0sNd6xfnq5g+bV6tZTT/6NaEZpML
O6TYc+azEkxFfQZS2ru1jBFcq+UgCtfvqyRSXvyZAJLTvyHKUBJsGyvt58zkU4uaskOMrRLASrzN
jUh9/26d29sprxJCDPPIfo+S+5L9mtbu2FRIVlPZro7gxYo2507jbqeuZpXfSgC2UiiE2/iSz73n
GnAYzEKF3jnAnymptxYa66m+YurwlZNF+JnohJ3rXyziObOGWg+hqbuOw9vmZHxKVd2DfkGysVXV
uoZJt7tv4vG36/WzLKufMnmpObRcRiFP3eA9KWDHtnyB9LfKwXO4B1pZb2RLdMGQvdDx/ca6uARe
gX4vmAnCdIOANAgLD9DeJImSl61aTHyN56L6334IRvpseSCGTJ8mL8HtaIOQWpYMvF61fxMAltQX
PLeyPbtfIZSSQ7fie6bgxTnOPDLD1VhaYgkYt9fnTFg8mJJb+8Ju0K3YbQQNU4cdVj5XglvXN7Dw
9rcySte82z2iaqco2jTl9NMRR3lNm4bYG8cciuYmRRNhJj4XU0BwgnjNnNCwfhp8gcCDvLyZzNse
3wJpVlUD5GYylLmHFTyQwZcupcB+flgWBznmzeULPys8CqXIq8EbD6efoSP6/tr7f7Dtf3k1wCkg
2uK98wp/iaCEiikPigXY7TLkJKNG+0Gl4QXp8K+EtQ7PFiN2vHN7RPezD7Y9tx3FqMvJ1/j9LxHr
TTSCLb4rrr47gzZHDuU+uxcKofejzTE//s4cqh5hLqselWH71D5YCqJhyjRNgOAzVRy3VAhpfAzi
9r3FOX/G1Fdl01YC/yU01f6kL7SbWXBniPbD7z2RcWe3aIxwflC9l51vEDyVQcdzMzeP4HjCyKxE
M5C1B200oQcYYLK2QlDkx2hXPDiPGjsaBCS6w6zK3H+OdSJYNJfnImaLjTdLNLVkIIqivG3/7DVn
Z3Ruuf1MaBOJGZX9jcuuNp6oADEv205wiDHUMvIuTgiSSAQ43VBRYDkBOKwosEnCmTjDSE3DZGsw
szVyFigawBKSBKcbVTaExNVjPJf7tDCnOOxju88bVbjTSBd0ymhEwv0kU2DGZhVA5Hme2+RTdRrM
Ys/PKjJaBx+0frL8EG3or56LAsl18WQbHowmcxXNy9lsYy71zNvNt3rIqdBAAbaH5X+x8YBmTLzO
fSgcJBZeOIZyyFFrJNH3ZT88XsF7rzT2hOf6uBRejXP2mXCIfEv4TNTVFZFhJP5gTEoTnP8/js87
ClvxYE0UhjwQsDm8ji1IR2H4k6Ys8b6uQn+5PAzIpPj/L6IeHu8To295fiY6C/7Wn1lv29N1kv47
fA9P/HAxBVU3xUqIu3w/wGrdL9tJeIqZPRB55XB3J5Yc6+el17OR+jEDh+O76/87bu43AKvsF4In
apJqT/nNb3r3Vgu0WMWsBUqwNkczbBr05GHa03d8t9uHQBhoPwOBLvpbP8K1eG50GAqOrdmkCrsA
UgvaA0JG/38S1RVP3F+dQIatfSO2XErq7r/D0g5uEo02EProxJ3HjbnBTbdE8DUGHFulLr9isJ2S
uUlUx3iK5I5vpXmcB08/+qcpwkE9PuiPqV3pfh2ABcqXvjpPll58DRhRMvNm4WJ/Iw06X6qpwDve
8W5/HhcMjjPcOUiPImqAof997ZC//l9TuHKHCX63ud1qrNh03QTu2iUKMv4o/dKDdjylDEjNQfba
4y32mnbXpDa7l3IdSjMHPNZrXOSYMTKZmsD9JWm+HJ7yaDmqojCRiI1OAEsxM+cXreY49AEfIzAA
+d9wZXG30mUjGqO4sGTgAPLtmC6shVB0+s/aSmjJs7TsnNik9nfpw54Amt2WBwTtduNpjUcNMHpy
cZN5tu/nTyy1Kyry9up2BM/XlqPWITYLcZ9e0xIuzw1/Ue4gjTvqM/UgxI6Dn03qtDOlcKhRYhzO
NMEbOpetfVnuEqrkvbwOisrS1TE6nHz0/G1L9pBC6nrREvlSeuzCQzmVDQjdyqF2QE+OsAJsQgl9
dvrFk4bC1Hvy1GnoZwqf8iaYkzY1FmKrJrGD8DhdFnq5tLV3umEds6MSJY9JYB5sEF2gk6IjkSOv
qdKOo6tpWflm4XCDY75rzo3wVXImYq+WPUc4bxgznVbJ+aCt12m8HmCWWTVeUp3gFKVMii6Rm3vi
iMIQPHriUBtHvUaN1mB+yJ0u1EyVZzleLQq9iTiIjKJEZXSquCcNql6ef9vhY5igYTSHE+YV2SJp
5/5C8D59QKNAPP8k/2Nc5XyIlRVOKF+rvtIcXd7DvQ5q0vmDeO7r7XGCmvN5jwt2CySKYe0Qe7Gu
2Vf0RMTVhjFLB7PJUjsIwJV/86Hfc+IsaNQOTnrZ9ME/mgtz+qMbrBPaWOiCe+JemE1FHl/O5Gbz
DiBEm709h9PjUP5kEBqijjjM99e8rO3rPE+SzQfFqB9m+e7TD9PmjSkUpK1ZybA1O1ErTOQ4KrOw
lACwg88zQcve+TebPrL5Uxa0UQlRYp1KVS85B4AytqGLkdbuPNabIKxesvpcq6k9COCWkaoSBWSX
HqA8r2VUvVPblV2RIJrUXanz40ofEfgkCqD4bfgGMMU5kkElOjMTnQ0V5uuvLtfUHWfZiGz92bP9
qMVWfzKHlU6FEQumkMZRJVR/ICKaRRzpGf6Pi/d9MKN6qp0UUiWvsDugdSRNSgKvAgiwheNrpncV
bd/vmh4mFf6Jl3GoqtjFEcv2ltzn3PN+VjLNo94/QYDBVYib9dRi1MGV8pdYAEMzk/b8veFL7l8L
mCdtL94ejhK6ayKphYyJFOH0U/Rsl/XyJzJ8wmxt+/BVer+7xLKtuW3BB5MML1aLxY+B3qvr7CAI
BITF4t/7zU2wRufM69Z7LKCyVuCGHV5L8UQU27Bki5ykqRkA8bMZKOksXUY+6CKYQL1jOgvbH4P/
ykQGn6CN7NtaiXCq+85Gar2F/qgZ2HXf7grC/n5LmmJ777EGqtcgcD+Ox6t15utASzwu54T7wBra
d12lPM7iTr2GkJX8hv8R5JUgGN+yf1HAMskI9wEZxjjGkX/FzyVJqIX7icbxEUZ0ehzeosHWBv5e
KXKf9yIBYHAoWCEwXlsxMJ0qYgee40ETHTxb7Mmq0Ysrm5b7TEHpM9SqVROPv+gLLjs+Qn1JvS5o
sWuMk3YU5eUrnutPe11uWdo26OI5KuIUtB20vLrUc4FAJ1hdrXLaVqh3OmjswZVDpCIS80rFGHFY
yepbCjjUAOoo0OraasPxM1for8dkHe/ylierPb/4z78arummD0wg3ANmdPFa78ZFsf8+sVZuvWyo
4FNPDs17lbIORE8hxKR7IhU9rJj++UQ7YZ6zEdx2Pqw+ntPzMLib3kB/i2wyMT1Co2A5Hadu4nUU
njVhmbdPS924So2uQSKv5OUNIfwUPIGcLiCiV9e1kYo9pFAoSgjMpM4BpxQp/rgT/PZHxdllUEhw
EIlKsoeg2MZcGz5QvThGaDZ9hjOa3t3/l8T2RoG5LIrL8myl9GLYHWd3vXu0YYTPQ4d0k3GvvpPX
1zs0kg/j9dZxjmz8iTBrkyiWxZz/cm8xl2LsIw1mW2Ok83TWeoVQrUMjWfhnPnzjtL/x1swdU/3D
BQEKBrK5jayH1ZJv5AvjXqUfaDwlSlpjp1LCOhvZSKjRSa38jHWsh1D/LB6r3njsSFAobH67vJw6
BD5ZFUz8HNizwYeSNGiDjQ0JFJlsBABHkYmDGKhx9+bT9FLdrvhsTfMRXBD3E9H4kUHUS60SFjnG
9csyQlJppVWU0V30zyKxR8Au5E4EHRdehZOpV8vNfjZQL5blg4jZaEVwsErj1T3T2XvxcTF24cS0
mZB9PmCX8kGlFsrfhnI2eautoVmWwJ+B532LBZqoojKsg3RlvVwbKcXAAkI0sNwyNvCWk4T6f4aw
9Kh5oFYLqlYF8sRqW9ly0B3/htLV6bnIKZQIPmX/OxZZKwovYj4G/5OiamVri5a7gVOnLhY9atT5
U4pDsS4HYcWFuFRBPbAE/g8aLuRtA/da63eq1W9Qv/lc+3hr1+NXO1M/krywsMuYuCczUsnkiBno
CS3F13CP++1TKaNFC/STm+lRpPDVZsoTHOHreuw769M9eFOqTkcU+p1aoE9B1iEARHW8oslEE0Qq
Rj4+4ay2qI9y88UUlSoWarOG36dyeNLffTfJUohsCVWZkpjCAfG6PR+kIREVmCYX79oNyKbvgOOM
U5Q1Ol2ZJRiYABwCwCPtx+R9Rk/cmN8aJYvqDcDtR9XpV8snotAOOHwPwpKapWUVkEjUf6VDIEKc
/weboX1SwvaM6R6ld3QVWvQrih2bbrYYRnjNd671dY9C/WvSFSoGLZ5/+qJc3HeKv/nPPoJdSwPA
/QE/mZF8r4B+LZmz9LLhhrPu/CGj/AgmphSRrpeUxlO6j0hypa35oQ2uSyn26eucFDdZBp5I3zsq
HdPI7P4+XaWX0Oi8DkQXSfDQ+rlKVslT0GpoRb7GrwWXww4treSKtpCYMJ71nU9cIDVwDEkG+rhl
1twJuUxhx+jYlRRGvQkHRyRSBJP1lLKd1HmH9OcKElCP7c/WctSHlmtixi/fzFygnd/M1D0IvbWL
lY3iyoMspyJLt0YXT5apa8VByeWpoEHUcwZujBYV6FwLk6eqlcYuLrtuUVA6/0tFLr6TwxU1LQqs
dQFkrNx9TleB4JbnQbA/QNwDeMqILoiToa8lZ9uAx5zk2ICO4HdWZkO9sLMcIo8um70zqsdkdZCR
BjakEaY/Q3UxWDAKEvAQKItOS7bqrq3Nr/CKjN1vwGQxB7+IHsqg7335tAcvn+2mRY+AiUTnZclP
FeswBHxfTMQrLNab1XhVe00Yblyto0Y48UfrQ9HXjsHjhX0+WoFDgc1F4Tw8taA8rZDT1sHI2aRX
RXqqw9jwxztc5MSr7Bm75g+EUbslA3GGy7M/vHDVSXeTmhPp0V3W4s708fHKISKKmZArJ+F53tO/
161w2esWRGpHakBBSvU+vKBvGErxiCmvL8bNytwsuDGls9mvc4B0DqL1lDK2m/6FxgfBvfnZHd/9
afWjT65MKX7UskTJBcq90PtjXGFG+aPpeQxuA8bndG6+M4eHEWvYNk47MFsS0jNJIMkAIAf6fbkM
rJY5Fr5vE4M8VFUkUN2fyi4I8HhUd7p/Yk+aq3XCar42VTZ0StpIk/Z1BBhlg4ylWdP3jkIauerG
+V8GMhebh8qbsQrKOR7bM5OOgdEevDsV/tYJh4H7nXBLZ1EpJlD2UBIclKtFW7Pt04yCBSoKohk6
WlXLVA9+UgfdN9wKh442ke0ewr/+w+VrTK0UHOE0FS/I28k0U83o4qhls35blYVTa9q0UlS463ST
dMSflTV7tldSDKf0QGTrMzGlFYbAThma6M/XmuaZVxPyiVDq9CMnOCEdceL8T0XqSfrTI0Wf7hzy
GTuZ6eVDmO05gs7JdBlpf2N4PVjEAX5dhCTCc4i3E9rv+vLvlBSSKempxXAi76ayYL7iCO9W8n/O
Q+x4RcdN743ZFKp3PAwN5I9fkNA4EfNni7N2+q0FUw+V0A9v4NydjgUtitEEUrL1bRQzHCCeW98c
XA7cJRAmZMkyjvjaQJd4YDBe/Sk4+WlRdh81AHeAoNGOOQrX/c62AQC5k6T64s5zlFatFTJQ9cEk
fjcYyvH6qFsxlC4IODU4menZ52lm9qKOyqz/WDfqEXR/jQPgJ+E9kWl1dBT+pUqG2jKTSILr/eMG
Mjz2sqh89pSFXgvEUqpDheCUzlSyA5p2kywYaokXhkhaPxrXuDND4nirN2QiDf6HG0nwEG4EoX6V
4kXwEs+Ih6hC+fWiXiX+qZPJCBhCSsCrVMZmAZpaJ2x4ASkP4FbaJIVM1+QqmmXhcU3fWJXh2xv0
qCbrjZvv50/yMixxeNPKkJv4lVP/cY0kjq1NBHl9U/FpjatAtbcdG4G3HplIDgN/Cpy6zrfkodfc
5eZR48JYsVbD04/RkwahXmM7eSvKaKPU4iDYzdLq+TjnP4E6TlARj9H3Yu9RgiloSE/x2wUNj7NR
H/Y6RZSglJZXAmyhgVKWjCwgnxFRqeSL8q5k/UckZ/ZdhdyZ5UOV53mSJghyhZu5gdLhkWuMUtLO
kUW7g0lsy1GksC8YOpnA/atMHrcQZDYc9SahKZHPMW0Ir20iJWS6XU1N09q5g+dVBCxiyhOX7OU4
gvtwTS5qNCeanJnhhwRSj+AGeuKYup3kV/U2Irs/0F02kKiCh8G403iE3dziRa4pP4TG7r18xt9y
bZhE6j1z4KAUfsbEteOBWBvf/AgTYniBmn62Euf0AUDe4XmcorTplAR5GYB7fyo4iDGg2CX7uTCY
Elwx6rS3rEMljGVTnUMEEdaIXn43Vgmp6i65R8Ruk2UtLY+UoS4poseHMUy9zYRD4SYvz6gvoO1b
3WhnvJYM5LqS0Vqj1/pOl8DcQuaiEvRaHa7zfAirfVp3emj74NgAoUsSugUftWuYg6yaI7rVu4Jj
6T/qox9UA70ePxQWXdtd7lIjEDFuK2egig5RMAgARgdJ2qbwF0QCtO0jdZw0w1ZrsrdtYKF/bV5+
QLkphyI3gG+VNxR1TCDHmqOgGPJng6sCd3imMzcbXnBUNX2iKdelK4w683yZ90SmyGcqyb5xTd8i
cmFDbeTklrQ9Rhkrh8Q6MmwqJBJNzawQGwBeQUJ/VTNhi2CnLatx8CJ4tsuvZvViCczZM7e26zUR
SmDTlo3hjoy8CmK2at+uki004F+LxXTeB3jy7132gAPjPE7awt9t/F7OoCTuyLCW2v8UPSFNsCGu
EnRgIFU2stWnzcu9I87QwtJpcaPkQz1ftOlp5uJfSA+Js2DAEkyydz7YK7zhhvvBhsEJRjkJx0dQ
4qQorynYdgZqxZurJhVHOINVcO8ppSeMxr0bAlDT1QDuWR2rR3rKWEPykgSutNSD21lKPCNZ8/F+
9eVWE1V2y4GCq28K5g+ZrEdMWtUhCqyuyfQR9iLceXGJM4Gq3/wmqFwbUsUtnCWMnDadvhFvk7gx
C/iHtrbvFVefY+7pwU33vP1uRiUpZ9f5tIpZycv98+2wBYyf92YMStKRBTegeOPr1rixZ+kAjbaU
IFqPEz33UfIu7SeH3/5IEO5Zt4DpP253eehVNshteV2Eys5pz/3kngqglZHmKjdTSdh17q64kX9e
6v2lyHTnOz/LfcHz3cEVNQNMg94sUhoFmMguiYmeDn3/iKU44RRB1iaTz135kv5OUfIboapgpS0d
Z/PvtNQUbbcqIgxyzrRJBrpCkoMtwSYwgwmFah5H8eqWoEWRbTBqFHol7P+AVJOaZYAEuLig5MoQ
A5yt1ygJpHSh4JmIRH32jz41W04hFOkfzbYzYiqf56ZrTu9fH0RZ9qmTcve/V46/ykUbKHwKx2Og
y0ITB2YydUkEbhwJWT19bQpxFCdLgtFTGhjZDPSLwaM3QoR5jhpwpX2U7/hVBzbNy2gg6wLMNk4X
rhiGm2iRfEr3RvwYsqnlKmZ6ohmHx1ANyloW5oB30tNMF2VMzDPOhLbJ/sG5obbmomUnB0U3YKiw
uQxS7u8dV1PPOCX88yfvqg5rry/WCvWbTvk7mhCXfaC5sx3/MgTh4pOdyPaikm7150Tvqn4jkh/N
AaCq/SIQ25Me6ctiLdlkdX7Y/MARY5cK1mmA/TgtoT6O7GOKHmWTcYp1f48P3QOSYGSZk1X9haio
o8UNHx7gmK89JFFzYaMU5MlnfHVaufnJ1DhtEhErGajrkoZaogBo8RXpvbAz/OkhZpcmZ51hrYEN
dFJ5Wgga/BpfvGOXNVnjmPGoXTZ5wVqJYj/T+FVUHrT9B51b7CCFFvPN7yJ1AypIgE9XlNorHPkc
kFMvC1YQyNMj1FSHpZqK6ATCLXMui7CecagDSHzw0748unz76wvy1IbjDCjZoJqdB/u+Tb1ej0hx
6sI9feGzrjdYzUlnJKSb15eczuN0gz4gnEpWEG7YxGOeHpfSCs2yi8WkZ/hssOj/3ba8xdnoburm
WYL6XvWdKb6NIWcQ8I9Ny3v3Fp6UhZdVqtL/D5kcAO0+0oCagxPNhBKHhKbZaf7T+48Xks48Ao2s
CJDfruhRRPOp/dogvl8zix1MB5F+F0IVy+0SNHaNQhRwK7zRhCHs+Y8xzMbsFb4wTnjzbymVQXVw
OEux1Fi0lHTC/WhQAoCoI4AqWnJQgzNLHBCzWgwTK4craf+zR2uD82/lasptpAtJG6LVvZwd+B1P
3DauPZQSZv0UtL4FUU5cspZXqUBrpojhQSPe0jocQEPhPERA8QsdYmdIJsq/SzFxSV35f+3+hICH
q2I1gB9cCeZYRuDrs6KrzQ5sHtPxLiI10gt54iugtRV2iU+drJXZuXIBIczMi4gGIRmfeNXFxpnw
SffDlGBqivhXSv9nFKjk6nNlVhXIZNpQVdj7/8R281nMKGnvBrWlrCuOo4HYigrXLXTeO92eWh4X
X/3KL/41fbLOUA5AsK39f3BEROYoVKzw20DrJOE/1SY6IMVwlY8MN+5v0gkgth+i0qrTW4U359fl
DVHI/Jq/SfYY3uAKCclND94fT6ex345L/jT7l8XSICLpCrTEmR+BGX77bRwWEIhp/9MqGtKppzFM
4xpb5LVk02dLS19JqJCeXtF+Y4xez+NlNQnSvC8xBUlvtMatDDhsjTB+fGxkBRvF4z8/fv/pUYWu
lDI7aLTYW4RTtoqU/PzFjZh4HYJToWYs4zH6BA0l26BX6Ie/gKJunjaE2zvvfT8e8I6SxxZR4S8J
PT1huNmvjmryS2+jSylJ0DqqG4hYrgePXGlM8X6OLIhfNFox7s/Tii/eGktJ9NV1FTkyHtsUlrQs
3DLp7Oq/IXxzAOJbnQ42V9OCxrk6qIDLA/uIkQsxwy+u+Un8ctXKPEnap9k63lEFgdqsCyVJVUpR
UpKAxc+HpMQVT2Gmr+bcjVq6Avx4tS1Kdm5PL2JEO9bxSGzAHjmXs+ffJPdv3WnQ1F2LYuV6/mRf
E61q0IEgfGJeTEg3gQLbLiTq2mHigk8HBPCo77IYKmxNtw5i/7y6eVOk6XdJhLgVdK1MJDb/GQgY
PA5KdgXzn3dCxfee09GqGyYZz2ljCTII6fHu6AWc0Vkt2NXheOReAjn/1xMV0Re4sKEomxHoDkft
gM+XyxV2Gm4zwVg/HrSSHQGvNWqNHlZuUzRmU/5WJEIwjhMlvvtYw8NjfY8oL1tC1j9n6pcDhrdv
W2XB1PIdVSc6k2DklzUkf/XgDxo3f62tK/FIsRpgZxj63ODeK+VH2ZvMmx1SaJGZ5tMZJW04nVf9
6SdJLQn2CdzwSVTT5vZawK17L3wr+/9I/EvKKCd7cfflflaB5xJYvqQgDhHfdbBjQNxSelE/XoJE
4HOQHcVAUKIGwtp79tFVXi9sgewA/qAxPUY+ABunKiaEU3ujfni1LfDea660dlArbIRsoXbfpIXI
8yKZH7PrYoeMAGAC7WL9xu2Gsod7F7ahaCe66fo/SNlIx+pHime9aheEjOav0GWAMSA5w7S0IYep
sohlk2+/3aat54/nI/MTeVP3aSJ+rpB88tg8fA5owundRrrnMafhQdjFJRqQxfJpUJh9e2osxxcL
bhrU2Y1HrieJJexZF4XVszWXM3Z8leQR9CJLdVwXrppSl9IBV65rcwlccfqZU7g5vXxgdMwl8l29
1QTL6IsQIK6VMzgm1Vn2DNrj81XLvw4Ipc20821v+7ZM0UAk6Jt4m1BgqVltC7VzBnbOVeuEYOzh
MophgkzaPYurMGSyqxDWRQFcycZpinokIbjRhsNI93twrR/Z+53NuivyszWUViP9pWqc4EooCsoC
lImNhqLXF5KY37iwt1bFSLwJBS33QRTrL6gfl5pV8k762DVDDFT/KMCWUcXsj5IZgOw9zTA+Elb9
hFsodRX6vSUOrmfaLDrAdajZ8wQJZKWcIBvYqmAqToamoiT4UUZwWlVfeSQ07PoDehvTHRECPtnF
YX/fZTlC1K9knM+Nnimq6E4lDa26wUSPhwlJ/wsxquzBYnAxy3BTF9OYZPVmBKj5wV2yjVjmFBRM
uCSbL3dYg1rvwZWH0J4oGF35XpbBGAMdwU7+HnKdjsBpiICOkXdjSYRkpzqYyHsvIn8rbZUeZHlV
9WHA6Mn5RrBJq30ZY2hvI/yQswehMmr3R3gzfO+aBsw4g98R3PTLgwzH27wvBulTkBl/k0CmPJiE
M0KvnctBuLCQfiyQAbcW9rSuPAJ/v/C1MILIVTyGO9TKImEMwjKtTpsJ335LtKoxspiuRKlkyYRU
xtNGu9arjztJrbrb/NUM/oCaEHbIIM1Bc69E80PiCE/6eI8+FQdrO2NOAF3etYKW+yrFZOyMi+fH
TRwGIPxO7fqR8d+46dAyvSSWHuMV7AVBY+RUG2p+x5YGujndxXS8umRN+CXBM+JDP5U2xqDLVZRU
vFzM7q8Nn7rCzmwc9AMseKQL4kceJRBC/UmiRlX0rQI244zJULc+AuYvHuYMNGJ/a84RX20aIwwX
OP7DiEBdPOcZo7Had0L+YFDhPquF+JD2eqdHtQzd2gaLRtp+JxsQVvv58PlIMB2dhKlxNabch+1X
/+xQkUynaCb8uhS+GtVIUHGgnGrvELwWkzEqNGOzWgOINUkx6n+PQ++dOjJy1cqPsu1K9Kwg9Ixo
4mdJuw/nvn+Iqbodlp3Yhbqt1LtkokgjIskXIAuyHet6xwqQ+uHc8OD2gMOodBbAfJIyPLZ4ELlW
pSFBVtCg2cbr5IxYayvSzvnb9/p+XJLjv77exqArcD/Sy92qr5SZIXUJuea62OrmkRqEmyIBqWCt
XfXabMdUXFIna870irJI6vCC5wX04STRHNDP51IiuBLrc38jFtareO5u/B2uSH2fgXSHr3yKmsf4
12Uai363JuxwqMZ4QFoDxzYDoIJpj2kTkjbCQFzQplVHf7boSkAOrtvdU49jprWHo3TYzXC9QC3u
fYnkrXbHXfhvI2XgSScC9PDVePJtQ3j2Ua/iP3fg85y27eMTToI1hhNHx98i+tC/cFZvOIX0DL9d
DSxq8h6Fw+XE3aoBnoRoeeBYL4l7yYWB/NGjog2jchfAd//IWy3EAITKhfpuOvQeVe0+6ZG4A4iA
UgkvPxxp/EPPQBCFTz/zy8p4kxXQSnmNApW+HmZsTnAAkc9CrXtFS792xuK4mKT8iUFaooS72fHU
F9Z1K/LR9eIelCzLy2nY0ZOUVqiaQKfCTrOKjlQCnY0VwsJXNj6Bn+AjMdzduHFTrw8svCM2KqQT
JiB65ARcSeuae6j1TDESznu/BjYovlQ+uECTD+fcbziQi6j5WDGSoPpAPPRTe+wCoqFKkkGDP9Xs
T7GeGuDR5DXe8E1uLSPZe2sf2qHQ1evrRnMeg8J3I+Nu7phYeeCx1+v6RdAnNPcLF2UIxggKVVdD
PfkR/O3EqH3HCADEob2bfkIPNsOEgYUGQzzaSASm8nVW9a9izebLyepN8aPu3HVf4H7TsLVbqsK0
ElMjomfqOR6Tuf71zK0cxCmnUWsG6Z16M0c3K4Pb+OO5UI6IcAp96lUnjzjjPDRRB2syBV2l/sRi
RQ1iutBTkD6J+/Y2a+p0fgGx79HEPJ9mqek/IiDi5jQ24F3F/9vyxYRH0OFYNCpokOuXObDx49Qy
8qWwcE+B+9xBmFRzSdSYCQvgZFyj3E3RvNVHhU22khWQ7fwYul/gWQlXArt7mTRL+1QteoihHADu
dGZFjwSemgG+xa90eEGTy8St9wiDQWYuIr3yGrySwOgGLLGo5RAakFrgbjS+0UyVzuYCu9sFwgIs
qIwrUqN6DmrmkhGHqQZ3YMJsl46vlkBDzW1iOS3CZF9lC+oU6Yk70KUrpaZbd0kXT4ehs6r4oO2t
VofhfTgUaPrF7YiNSlo5IVfedG0Dk0ke2i3YO7uinj3+8F1hMHyKkNYAcySsLFphH5l0guiBc7ff
R40ZXhl5BRbNBfEeJrb9NiQAuZcnQk9je3MSXxePvy3/9ZiT/HIxOBnab4maVFbMmJpyEfMwekoL
ONhFVp7WsqDx76PMt3ApKMEt3iRlIZ3geYB9jNha5Yxu70FW5Jb642dY+Fc8th3Q+kb2koMB+tc6
or51Bm/rr3u7uGLstDPSvOGeaY9O+6bHbcro6HOQvYRshKxlLxkW8RInqmw700x+PpjUec/LN93M
DY8CorHeIeIt3ba0f7bj5bo3cg45v9ynpeMDn9/wX9PkgOq9DhbwxF9+7iBDxeKXXlU+F7FzuKwd
KUNbZV7Vm4o8avQRc+yQk9X7Cqt0xxrUnU4o8A5fPD7Q6p2JmPZ2PO1T27D4QlbQBDi2Sm16sahc
ALqXZHiBC4QmPEjpAlHlwZ6/utAiYHOhnBzTsg+bR61bVAReypzkZOrfmQbZ6jUkk9+K71HKOyN1
V8JhSC+EygJGvUk1ryAc+e+RT6nK2XSuxrD07AUfHOD/Q0KfrOeciTBGIpm8ZMkUuFHhhbebTR4g
k62RB9l1N4rRAeQRORovKzECHHhuS9109BfpLBq2E3mAfQwaSgqJDOVaov8vTYX1mFo6HtqNkySV
5jpwdBEyyYiukTCBlW/xBeg6sCWKAqXBekBJpJgfB+qTqRj3yWWXZD12MX9R407mEt0KWRByxIA1
fTq0my9Xgn8pS9tGdUo20ELRq0UsgZvXY1XJBwNSuZwBG7nD6N1P9oGK4C3bs1CYn15ZAAe/p4el
Vdbh+LmTvYTPtP4ENYdSvRsz4wtgF3fkC1BPD/mpLP0ogZmasJmBWn2vKlOuBJdg1W32m1JIJZYn
FbuK4hMiFyzhOUW7t4AOKlH8z04Rrfuw9/XObtL6JI+Elr5TcYab/JCjT8d3PPkFg3yn0aY3lJYd
krJjpgMBZAZF93wnucgfqnbp1IUr2KmKDhtmTJpO4cffnjkzCMG1R8En0hfjshnF0POsa44mOzlf
Dnk9iR/2QOzTyHSjrU0RiVXBYBKYRtGfdnU/NGldEMzMDClEst6MXE7S6v9fsBZTj9KmYxR5p/GV
AJKhBD5z34o+bUA6BQkRvQJG1np83fF/QbdjbhRkY2s6ZbKnCn0gJgti5PS8JZt6t6TegUPzUpQ3
8ubE06/Lwrs9iByvltR4JpGi02alqFY2L8eHjiiBqqBZHw5vL5n4V5pmpLk39MxMiSr9QZe1PJHH
ldBGNZnn5ouCxbtAd3fkw4gsv16ZnpPNK25WEFRAieETyVpcmeCWddP18NItNFH94Tu4AtfineJD
MEd2w0TZuvkEiQfBOIPwtiSjkfSAsB+kHq+vegtsYEzi6EFPm0bff/bGyWwkKJEBFEZq3Zh6n6dd
oYBpDTFXPVJD910Oi/zZccKaXm5tcekth87xVmpI5SHJpK9GSG52KYG1TAxPZwAneKRDog5WDJNr
nSXJghQ5LEbseL59lbRDBJbMdLgigSMdXj1Uo15/XkP7PwgsXkFKQWeILJ0bCANCcqZWOVDWffEa
vKzF7ESTrQE4YkVAev5L1mNV6twsK9JoFqQIPw2rWnopl1AUfKyxXW4sG14tRB7S93JGeMR1zEKS
XscmF15SEv8RCGhtHr7ZDJ7ulF1OaixRdnSSDEYJLfPowbZAWzH8OSd/z4FGo1rHKsWGnzGNmQdE
vv9I4kFT/MMRKFChzTSoSw0bUKGmIE+e04EQojoqiSb0LvLCoUWqcyYap9na3sg5C1xzst70f76T
tACcjgOOGCztEdfZv48yAUNl7g573r7kEl+bWxqShuTxbxWL+ctr1ScAyqsHiXVLbimiTzhC3Tst
lnXh37MY3q9RAGpmnY/NpD65D/tDNC0vGQZIh+PHy7te4CgdPr7ca+QYcgdoT8AuDZC4xulPMLJn
LXuNiwXIUasNfkriZ3O6xk0Xko3zdbX3Y7skUW1evn1sz3FEqoxu4MAloo2Ju/1ZJYU2/qMKgfh8
GpguAiIOTPaFKjhhWas6HhPspZOYCaczEbQBumzPScAC98KNl+3yjFlsevMiO5PNdLw+q8GGxSWL
h7qyvb7c5ZuJ2w9U2B6CT1/+IyV8ZtaXL+fh+wnnlj60SmzvWlXPl0Yo8qeBlQ8jxn0vT0FXSCO5
DG9ROKDxAm2QccQfBwuuoy1iWJbVnu3zA59vCcNowjBfelX3EgxJtw+hzk41iZIERNQnfhbwnhBg
6+A+Pk5rVcJuEnDICuiVIVOC6hN2kqdzjuqzwcIGlNPRvaY5LA45jqKYuhhuji0a1qQ6ttIYrxVv
Os0a7k/y7l7rIsncfO0MqwYTox2tNoSEqBQwtddrqWuGWYyEYe7MbuzaPqS3Ie3oUzSPMvzNUkb/
3pNJQR4AhHnDTDNU/QrBgzgk2Zo9FjGlqebanz7htHQgMKuBSzeoQ0fyaiy6ub201yS7jHZilAaZ
nHEvqiXZ0YXqcjNRY1eBxpabnywUKPK9B9Gn+2+N5JUoEeOytfpLn4kC4Kj8D1IVD4gNsX0N1oVP
BPa2ifr95/SbuAjHTT3BlFue0db9hlvgQOmYW3V+DDg9BDic0F8YCKcH4xZ1atCm44sW8wyD1zmB
8yeUfUfL65SrPzHzlwE00rqa+/zo0PRjsjYFUHAQVCTsWMCjZ0TzJG1Vup/otc/3tIlzrqIQtIss
aFaqU3ww2o1nRFLuDyz0nyvVmQIarnIhV0M5LDDOTtnCudlL3SHQz4ypRR6XbI32sfUsdulbZdRN
XsXVQDxWyy69G+zhj6BjEYiV1Ju6N2dIYXwvLpHnLlrNwwjmRSpzKYAmmPVM/qcSE0Vnti3fLzUw
Ra48y8AUS5o8UVQ+GIDCoNS20dJArpqj7tTnZ0Ebfgo7TmWrFEtoIyDX+kJ0NpiORHi/wylL+cQu
vdtjcYquPfVXOePyjBOlEBndh7zwEPizMDi8DjzSjCA+AyuZpPo9vJRQMEwy/cOPYnr3f9hB+bUJ
HWORbvnI0JPQs0+k2jvvd59gwwvTLIok3CtSRIbnphuUOdPY+5Ra1l2QmX/LdaBkotFu4CYfNOfb
2ASIwtDFC4ZuXf9fyaT0BGdJzKJ9FTv2deyHfCRIbrdISAtFQMbtjuOfLLw3YusA9/GXSIsl1yS/
6dn6W5Pq1TNl07ViUF6tyoZQ4WPi7Dxmi4XtmwAGexEjyoXRGUiGjeWaszZeGwKMhAfSsaXXjQkL
Wb6L7NJBlSjvajE3nDa11lgpwdLuTj0yLdcEyD7+WgF/WJ10Tve0SBlCu8YiSy2GmrrGI3NIFj71
SKoxcEGrk6T785XBnAghDaY6XctCqSPs/yTW8ABtaoCIibhjK/5FAo7h884R1bc4yg2bPIFwSzMq
B8XKvUrmwA0U3an3Rbjk2AqcKwxkURkkUCIU9caEpEUSDU/xCRqpSBfHPl4COYdfhiSBn8sbTxri
/a8bpGFR0onR1wyAVe7JNZgyNKJ2WhDVN0vCp+kdcMju8zAyI2sDntjCl/feH7QSfRsWdU1SDGns
NtZx/sU7238GDLHHlYIbDDXg8dV2ePHJWSEtZ2NqPHLiIxPht1M6ZW7Q1AN65wri41YWi6zGLasD
xqkl3/4JpMsALPMBvPr2JmvoyuZp9GqvHyiWcwA2NzZVgXoqcr00oBqCmg/DdbBcfQ9hlDHsLlJk
sHMEms5s5S1nUokNZq5eGco3ufcVAsAvJL8rfGKkn5b//fQZeEqPRG+qkYAZKwwH3ptMRtqFUo6R
xLq8snZn2tiMBwk+ZXQERIcviBTAb+wR+77xguqWpv6sLifBbzyyvsVr7mo6XvuV1ll0tsy53jdS
kLzu8qnA3Hpxtc6riAdtc7SRS3L7c+lTmETf4MruKZflAOs1LS9C1PNMZYT2b4YCxc3JGe88MU/n
zIY8puELH/0HqrEPxkYFSWILDbH0+AAiSxuqGy+P7ippM/1+bpiGJcgUu7r3jvV76YpAYiO08TO8
8ebv6e9fKElvAFTb+l2BvVU3LpTdN0+DuouPglCLdGonTnY2dUGQMhBvUXm/ThoT2V8e+UAzHWEH
fhyYdvmIlTJB5CvHjMFX622J61zf4Ypo9+8hkQFbKcX5Q+xEqKHZ+/FK64PalO9s53SGWbNieQ6y
M44GqN2AlkPTmzMY2uwP0T9N/HcGCwwcVUcZyhg0TrLQXNeZFudPsJntFlv8wLFi0QtrgGI5wCh4
tuGiqU71FWXsF7UQiur2FM/zTfuAPGytFiqtPfwf+p5UXsRK7FDg9IosgfWVWNwb2Bb2mPBx/ual
jjrMUKr2xK4wmpVnfwcwNduraeQgqaaVXQnAG079fDUuh3cgQ/V+AnEYC/dNiJMSIFhlLlO4W9JE
kmOzaTq0MwV9KjYZ0DTr8pcwOD2Su1hYqkAQMMioqMZLexD6CGEMSGIDivCxY5/Z6cRtnuQl4SuP
xJa51Sxk9zUGPBeNXwZ0FVzznwbSFRTggZ1JvoE84JhK+fsVOGhVJ8GlbaNH9wfleLV2JgUoqDIm
OcQII2Yr6lLxOdAMiQaqpPnILFYMCFNtnvlaNSpd69/VA+7ZPckz3hggjB778SIXvLCZ8MfdYFwj
U4dTMjW7Vlgbj9u3ZdUIbyoMcdrQoORBrynNQbFfES7v4/afs7XpIC620EgkmMMwrS/ZVUQFTQ8g
+5BvQ7yFT1H5R1Or+OQ6iYHwjsOiN22x07xQUD5Zp4QKYxXbreLVc1XbzHjksf6AMgQPSWkg1vW4
sv5RW2gZoEvwnKMBqvyTKOUfkb3W3VMrIXM5vWvyrGbd502t2EqhZ0gTRhsx06zfGupNJMNhCwn4
Sutcm77vwBz8/gioaOyBa0C+N8RGLTrJbnKo1KDVLa365fecbjpu3UyGXBkCi7XF44jRQru9w/h+
Rj290ZDyTCa0Kfpg/+3ninP4MUKl+1lUCTtxkt5eXKrVK063fa4iu0yJga4g/4zKWBn94AkoG/KW
b0fVsAyrDzH+boUO1SYWYCq3z8LgFYEX4k3ft/wNkKt3z7fjt8fTBzWDPX3tGOyebn5nkdvFS/Pu
qKMMzRP3hWe5RtOavjQMWpVcxBgQcDtPn1H8esxOucD4VRsSywdEpGGbfDhVUD+F8rS8v57dDazM
GE3CNjZQQMoRiu67xoknlT01ZvnbMC/8ybYUD1yugw8vgp2rwSwtKqe8t+IL0MSR2ASaBjgAZKwY
RHwrYYdc0f9m2iunN7cCK5sqeJefeKMcddqouHoRfKacMSSRIEwe8GVBD2T9bzdbYpilXW8GS4EU
IwlD373MnRosznSaLXEpwpvSx1HUVhLGzjm5Bj4MCrbinX+mlb3btgzNtAngdMmo17ZRtG9p3CiV
u52CVGmPG9G0eduS+6diNoB1gAOmp1Gx+edJFy1zR0j9BWv0QVoMrozzmuXeQe9tfmRS1s45jY3r
X2vvRoK076ZsPZ40oxNbbqxJCy55nAQ3D3+dz9XwNCcDoXQRs0DEu1796UMpalRaGgMDgsalhkQ9
fG2EF7BNuDUIgyuSf1w1Q4dQz7YQV9yyNbIlU+6RHeZAe/L9hIiIrgjfGL91HVcGl0MQ+kQWX6c2
1NBQYqRC6ZxL8Q8OFINxw+M9m9ZLiaN5zq8ZADJZrwoMH9Op0/hM2Y5a8aeawL0DZ71vOR0iu6Pc
vPKLNm0SvLKxSXPsEjZVqFSoePDOyrmAhfX/RqdndUFACViyeFzak/QwWYPkCkc06OViyoa5ebsc
ZpzR72AlX8bzybJPQ1GUDAzzOp9ZHzujA9XjsCvhnke+1vyRvlH/EUXhxiF83YJfO2Gf0lEsnA5M
ABD2Tp2eEsBlfV4QCtPhsroupMeZxEgEp2xu9/pJYurf/P7qu9WBa2qoLorhNQT/sdufEc/J+y89
pYjtDyF4jcOITn09ZZl1WI5jzunzSFUA2qVzFNyV6orJAaIIpv3dY4jTfrP2OCjxlVCie1a1DUDk
uXs2LUL1umKT9apmpSTzkA4/qAlCD6I1DOJODVq3u1jZAssBPjSNAEYyf2oxwTBZ2YYtNCL1dvQ+
9iMHyN4hSGu/OvSnlxQOXSpTaRDlrHKcIOoaPKNm9mmREA3cidTKrLJs2mXl+UTAo5YJKQnYWsde
ouCp8Ry06CcInB1uRQ2phXBZl5e83HVDjjW0OiGR8GH/i9BeaA+1/T9kkifbem3yy2M1qnxWNxp5
31MzNK9gt6b9rVFtrIOD1bGski2HhbzWwrKjt63d19vsO9P9qpsUKUMqmQ/vEPZOsFq0y2kltBRq
lKEDxXjIVU3kRdfbP6il6KP5FOxIu49eXwMDG/Nt44avHwZb+TNW9F6ZfWJApHkrLWyxkkEl0u1R
ivc+kseJ3iw5OvXfCyZEZL6m6YqZ8UXhyGTHfJOs3s9gY7JarVML3Y47g96AoDgNQ/1YMyD+DpFd
slr8aVhSgjhKu210LU0D2xHRtszGWxdfTxYlITKfOd0ecEQ6k0ejpr+Av6Fuclse19lTs5+FbRVO
bLQsOK28Pfh0+mAPQ3TF+gGEg05XW897/frWi7Gd1a8SQfCHoVfQdDQN/yEtK+sCv//bSj6s/Vin
aInW5mjFuM3ffmPMY72xkIxTM2n6AhaYHysvJ4i4o3yb3wwJCDTy44D39GCkWCe7YvweBkZvA3aU
Dvtdm+QKs8dDVQKYFcInP57HQ48TBARQVsMEQB/VPyHPpGkHCstTT7p2TyAFeTjXAjhp+KoJVtoQ
s7IYD2TJLQqnJc144Zbo6RwVFNReH7x1Z3C+IpKiB5wpnXzaNWdLZ+MvHm09M0yq7FjeIbgfVIzc
TrKG8nUSw/PhxGZMuVUclmzLwFDCF+cTwEy1dau5J7sywXQJYSWb1v5BXCvws9CUj7HC//jIEYAh
T4ll4f7khmeINrsQvbfChjC/61KaGRnjcAqjs08vWgebynilfP+BmFRzs2oTbctZ0HTZJ/3n1YIE
xNGQOl2432N8eUIKQ6oy8JU6dQrydfcXfFuRcu0sUV7L8yl0NRFjn+JppT/w7VmAALVHyfH9Ps/+
gW2EuOvFhSa0TNPW1ZMa5vsDgS2dm78gT08k8qm7GwQIwlJHANpHsvNw97pHFrFkxe8Q/PsS1C1+
qsXR43DRqBdPwzQ0DDxXfCXrWY/XLRr8fMcSXM3bGT6prPrCsBO9taNjAPa5Olx8OVc4xO1wSn5U
zjww/WXuPbYIaoLm0H2w89UJiriILXcDIfQp4pEgx16SyslJJTkLZyVKFnsFwFnUT14RQICgE/He
opuPh3u9Ic+A6H8i2EHI6RX3JY4xVlibBHRoiI3pcYCej0Utz8PC74Hpl5yIrabv7crBWa3zRlv9
sFYs3c7XOxdv2FJSs6IjRsE9Hwhg0AcEZAUpqSlmJaX+sJaLXfhuxlwjiV4eWgl8tUQ5bcU28iat
FUfACgZfgDz55cffnt6zuK1/uuVVDvtNl6jGP7+ldM4IBCmNusUANjuRN566h+dcv9d7iJil6/Cd
c01uzJF8qAfykTGFMKyZFn/n22Fn0VS6oqkoSmep4b0b/tYsuH4FYD5Nwq0NbAjZQAsPrwETA6k+
IMSDCh/0MhAVAG68FFOV8U1DIzGm/z0sP3M+gsHJPaLE5OLnoZ+OcBtqccKfG+f6tBKhRhDawKR6
9u51ep3rKwHwYW8Yqa2Z+umyiPF8ZIgRTM6vvjvT4ouz+NLcJbNb2cEYksbJMhFvFFwgfR1nJBu7
u42PiMj1NSBBGtsQHwfxRmrXnlrwqdpfNwZdrST0B+OttxE9adq079mSZ9Wq5NWYp+A6rTxLKhiE
uMxrtt5lC9OBYYU3Uh7PsaOUmn/DbgLYOPWAXSamo3/IebFD9l+XrB8+NX3GeTqtkq6E8Y2GiQ1/
jCamabILJQ+V6rckgQUwKFA1eCG909q944+Awz8pecyllyJ64sdJW//CvYzb6u2Hks+1Fqdkga4Y
W3Lr/yO5upV/kSf6VZQmARaoaFwEAQRSCBXG7FOgTN/YWoJCReESK06Kc6WFct2hUhuHET/+1PPV
US0I6Co7j3095ZcxXYEf9E5WyGpVkT/D1XC9iPtcaPNrU1c51Qgn0hU7M51bUfnq73K/MnifCTbY
AlBT/OAEEbILfw9MpPNdyNntMK50pP2lRKUT6gqQUZzzYsw7YeUHPMfHhYlM7TLgGkrBYlnXkKZ/
Acbc1/TDNG2yLmCTahuQMlkoYf0zBosWwSmfLxuFj5BrEmK8Ng1ZJ2kbArhBpBoVB64e/iwFxGNJ
O/GdYDHX7CWnn8g7uJhrAcoanMmYkGJsYReQBgpH8V76sR064yqtF4DFNzThWZogm9FRIbxLu8JZ
uS/3no4vR9ml333VQytPAaBzbArigGzlcrSbrE8z4HoUkn/AboX7Hp4XMm5VlAi+JEpT0Tuj0AX7
xOtEs6R3KBIBx7yswdBR0Uki2DSbn0xZS1+MN5YasJNzWsSY5YnjP98gSCUt6xMLiO7XZ9tNNFTS
6LkNkFBcOFSbyuURi4df/b6nH0+4ErdMoV8OW8uVuKPqxA+H9ZKHNrcyTb5PxblAb8HESxhZwukW
gEq7slFE5kIK7mmY6mjztvXZWd1mKXcc46j9mvecengzrFHNyAGEsGm20AeEIzaz9EYW6zNiwkIL
m5QcgfY+dhsE+y6iFDGACEOFnm7U3RkYIFJ/f0O4bqwe82Jn6E1bliimMBFu4LPh0q6xO2jitHHb
k0XR8OdypSUnIhE00AnLhxnfiYTF5CKf3eNaticuyY2ONJdYANY/gkLqLGa9Wx6HCDmS74NK4fR9
gdKL8KF0hyOqx7ut06EdQm3sPibxf0LfeEFllerB5WI1vOXC0eQDKCUxZvEP3b2HRk2a5eTfOWcM
KqkxoUeYflWjVxf+GTAU87h/pKno/zu00aT9kZp0Zx173t3KS3fSqhdZdaIlam8aBtC8nePEcHxi
rxycXrm5aXdM3v21SsY41d3MFGMiWIVJEdRjvpwSCfoyxRQIvH9AOyWct6mETlVLy6YoqC2bwldY
Emk8/YPhy8G53Vy6+5UFNTs9nwhCa+WKVUueXHbBPaBjQXSglhKcvrrFF/dtimIB/VtjHcEliTcc
0EzP18Q6cT+cGPBZe16jw9Hz7VQbI8cDfEcjTRvYawLN7UpuGz8pqYzZq5uOaC/QyNyzHLB+Rct+
AHatg3qubKH30MZL4KCjDDS5uIXpMzJjzKITEvUbRb3cVGl3mXUSztotSIm21JeVCYMDjEJ847Uh
CYWQiVhlU30aplbGAEIMgoVs59SXP6kt5MOBzw16AZtcUFuv1+YjooO8h+iTu4zG34oU3n/O1qKI
mSzG91u41+CElOmYAIvBc6ESFv6orPTL9eNt9xTIwfis8XRDYePi1MKtDJne6hO675SZ/sRWJKag
LIDZ+q8s5z7d180fnvNZRFyCAtMG1qsgBZOuqY13giAiGrMpcmyDKIIRAHIEGt46+8qJfdGwkBeY
nKWmmcND0WKFGFY0HUNum/JHJuBPXmMYJanYlLXxg72ZLnRomkHXujbMk8dnDieKRBYAdfCS6gK4
T8/NkcfFuB2X3E6GDJcxXMPQu0NvBFU3YfFtqvn9o0szgaRhY5iDc69iml1m/8KqwdqjrmB4SASA
4+QNySOIHlfh466hu1xjQjvVjz8UZI5K+R+V15zAsDGSbDuwNeMDWGdbnW+ioHde5rnirhG8Srcd
0qt1YyHYrryMMMkIYDhwbbtyJKndJNqYTkqkrGzlK401z3bQaw/o06FUgg5/A+gwYK7CjPjr9K2b
/hNE6oTkdxA8+vKshpq6Bg3UG25jDkfsUiFcp42EaCxYPgsaho50kwkFL4klSybT4CSc4zPSX9jG
357faIbTpEoKAKrSnjapzrRqNvcq7oYJA9In4RQAFJDKV0q32aFyWo1f7ydAlrOWoIS1qZjMKVTk
bzYx3iz80pLUG9uwUo661oIqnIcv0mfPlrYei6yc2Zv1FEFzz53pz3zaTVF+f9XESqKsjagcH3tj
H+8QUuP9SxS1YD+z5F3nap8c9/RifwQXtT3G8ImHyr98dYkPfpy4Q4pRHH7ROOt6MJ0ydeflPohz
Mxar4GISdfSr42dPp41zXqJeWeOP8JnCVZfm10DFauJ33EJJRfuq+O/pCKv0PzesLNtyMUsDDfUq
oBPBpnCMD1AwxO7mB4MeI/bAOZz6w8drneAXGLxGguJBv8IMgxklwnIRK23rdqDpJ8FA7D806YLt
zM1pz5fwFZDGA6uImUqZEVqkOI24Lp/YT4jI9VLZylZ72VMbAy5B6jVfH/Y1x4oThUI3b+SJnUf2
CpdAHhpmsmvCZVQy1t8jCSEAGUPkVxSP0S9g4FIVGpLqAH1BDft6waj2hldmK7+Mj1324XBUppo6
m6lez9fQlAwFfpoPJSm9sAYQhk6km799daKdMMoe7gyvoGiVTPpe4Ygf+A/KGwFNazdzRmiVPY2u
z3EbYBDHTqvIH+OXtXgam+xFHt99f/u5mQ2xF4oorUPNrG5dGGiIJXtcsTKM01WE/PeIOzykUELn
BFYT00AMTGN3iZnMEKou2MPpjKeLmtGCpy9Lv6WhhTvY3bU1S2jUK4D/lExkcotdOkT0ievtEg0a
o7jPUuZh6bdRpBlo+uCH2Vmlwhu/D/ngx4n0sj9M471sLsuEe3ZtLz2tN0WpEAuIOnWVc9/6l2/9
7hRoESqSOCeiGWZmHss1Jt7/x/3yINzKgLn7ycwPyto11cJ3wcESKklD965RBcsqB3jEyUafMsSU
13yuKtXJOTvwFlYQO5YUMMePNm88e3zRXt8EecWuUCifYNxXqw5fZww8NkGRP0PtvSJporg1Iq3/
TnjkT1Hf3LP42I12yv+DLGpFYzaVAQPo4cdzVdu3SFhRrrJh0lfMVsE1AKbOCoC+Cqn5eZRycpXh
YfeAX0mQQZEA2wQEbEOgp8WW2c8WCxAXh5FOQlJcqR2T0Dd1fDCH/HGvvlMj9pUAdb0oHtvx7MeJ
Uy5fLYy+0YWsoAU/Py1gm5bjUhHMDlKWvf00M6RbVLZ+xbZUR/AuXjNj87TqJdurtpQgE14gjv2g
fTofjO41zfGBaKUpVprGfWdHNK2ekuqxMytIYdCry/Y42Z4A6Mfo/jvA+8ebxUT5jO5D1ELQfDNY
p8A/z7cnTExXgKONSBGxa7pj7Isi+c2R3puOqZxiD64fxOuiZzSWD08dlEc8gMu+n3yfB4dmfdKB
cE0d5oHPxq+l9HtqO1YS4tDwiWx6fmr6NshA+R5OsReUEq4U78qSA7Fhm6qJIdQf+kSVk4MhQJm/
uI9XTe28nk/n5hJyifr+5wdsX6MBY5Z7hubOg/7MjXSblz4hHAu3BZkubHgW8Q9PCPRNxZEFZ5n3
tGyhUAyFeHE0e6JTI5rAnMAubpbE3cJTutrG6vbJFxhL9yof4PTeREZmX/5OXmrODUbSGrB+HTvU
3KOt3I0lgRSYfHQWHZsN+BD79fj98N1BEGLJ6/jURWjhtf8QYUba2Usfg42uMHLW9+XSTupY1Zh/
AajCbUwKydJx7S/T/X6JT4k6XAvsNrDFRt3JertLCsSJ3GUxTsAR1ADwV8SBcdvvfQSOA8bi5X9C
2PofKBSL6jxq3xDHoxywf7flEhBZuc7mighEbzLHVswsVfB4gD5Dq3Iey8Ef6GePQWSiNg9mOPbv
6q8euZXHHZsCZzjawOhNYKAGB+6SKsNM2ChEOY0rDml/Xbi77E2SQ2mRdn4N4kv1gpoC02auII3h
dM1Hd/NK+U4TvGtFTqxRnXCs7OwcnQ2DCWJnZ5TzrGlOQQuV9l+xtm4Ds+E8mhJ7bSAajdb7q4C4
s5WRvQDz8aQchBff4LVcxVaBLaVTLd/c5jLDVeg4/0ALb+uu38ed39VIc9geonX2Inf2YzpDzaI0
cLk5ClCI/bIcGSnnSOlofIcxVltiKHnoHEuq3BkfykycNf0PMXIQOJwEGCv9BLeb7rHzYx2k+zsx
K/3o8kMb9sODtxgkO7wVWT1NMItZMwXGaEvCLek4L5/vkp1e/LK3I2dEcSx+sdxEQLcGbQjR4XGc
tuMr4rfVzbM+xVo3ztG6Bkvin/r1SG/AqEjRdnfQ8RLIV0zFVt8/z+aJSx+i54S3l2aEhhxH8pZc
m8bBr129NsanODHbaBw4I4GA+SvwNW3i5tzQN4xCzP5t95mRGUGklVCPKYTVHLV/Nqp9hr/eWlIz
qSN9MDyi26E5UElfWCLe+17P5BwFXBcoHrZ+by3v27B3LGWVBJNrwtB2RpyJbVXjDnsUxtK8xvN0
xyEpgTt+tBClAIAHc/QbNGI8HZX341byoyfpKiEy6ewk75tZMPdgu4tZRz+AW8hEYWuvLryPGYS9
LnkL6Tmi4nYpcJysOufQpZ7YjXq8AoVwlZgPKuWwHZJIjAUxWLSceHPtTUzIi8Zvhk0rgT83KtcS
N0Ja5D+nzxo5DcJ3XlBR0zSnPu8/JL7GgkH9GDkHMJ+rrdIwnyfQqMjAXt+phfPgz4LxEnpfkBGz
xg0SQFjjFZ+T6uJlyCOgWl5rKXYVSYryeHlXAI2j5YFiWCJHThwWSixV99ubYtiqNc+TAGQ5CwOY
UQBbLwwb2uPj01Qu5sa5x0lMUeGFBTpswwUOJZ87musp4iK5GHafOYxcoUAPQnAbrZIZTgw1Dk/r
rEhEQBMPOaaee9AS0+w0wURzYu74pd4TQc5iYSCwrDKX6zKXLDUg2SBuAMUbV5uH2Q1jS6ulmxui
S0fxx2wVdmqay+/xi/G1AqSf0rwMrUOsFSZOryiNtp3iqvXRifsyYmoAtT+h5Ens6GEh+csoKs6A
xG3kOQ4ES2bFP7mmY2g7c6eWmuAGB17AwcvBNETFOxRayh+nBmTkDuFydiP/DeTFtF8PsEkwDglB
CYe6FA9gyCtWLMyu6M3zO6P9XkBtvMhULxPZBfsfNWLIl2TupgBGUi8eCiSnLSGD6LP8b+5JGc5B
Av5ClPeE9n5qcXeogD3wFlPZZPIx7aeOUQnAWPfdxxSuX+tqe4w5UTPrduws0EasA2hK+u/Jlq4w
0lR+/bITsKsorfiFXy5xmywAfp0Z6OTpmHZnlwCkb4OG8URT/2gsAYCXolxiHo28ZD8osDGq6DAj
N5FPOf6u8cLpVK0csp3HjBEoRs/mCsay2IjgYa+Tyi3J5TK0ACbThmWp+mwK13AOvRL7G4yevXBf
+qtIYlCbgD3gwull22pampl0Fze9ARMsoOxJgUS2eHW3IqqY+SJdoHDfatI+66Soj5zSmECTLX/H
tsg0VKGtxhB7M/yzq/egpfUe74/E8k9kytWHnAfGoNCbYjg3I9OacX1OuVfrTDGj6Jxjs+H8plPV
nEJPs03NSHsXSOqqyAwswflUoJeVEGtYCA3zk/H2iSBphc03boR2OICyROrfVofWrKMbUUrbSB/S
42jdguGA0anaNZD60yeNCwJc4EF6/BnKVZJ74mWrbv2KccQhSGbsHzk/CAv2GMlKFa03yaCBMye7
2C8Jk2f5q6iEo5CEH07KGCs5/TUWnpKHn8nuyxb5rxeLppeQ3iVCKSkpFRWyIkkFDkCtfZTpeHQl
5n6fgbdzJbphqOlibkMM9mxqu13TLpsY00fjtaireag8eHZ5Te4Fk8LzkUGTu97u+1dCyal6will
2BY45A2lFtpBJSjNSp2waftKDN1n+/k1TpDfB4bggCLMYnBoqW6HQRPqDuUbiH3AkbCm7J2g/wgx
cfYTFk1WhKBMwiNZwNIu/Fmhx6l8eAPOpIIlSHRxhX5I54mB4MYWlIMBPDtoFjy1grL7e5zwpFvL
Z1bucJaj3dHrEbAQnvjoTnEFhdxX5xgXID+RUgbhBoPwjFvJeZuzF9DoU+xhOt5TWbRIqZnvtJ3x
W/aEKHYv1IWefJ2I93VjT7B97fD3DSCGNXe9Tz+q639BTZPGbzxSfL6oQeh2S7LJ7d1IaPkv8ar2
SeVOO00SCqxIi6iU3aXCq0zgG2IslUtc95Dw4NaJbr74YUN7EeWRmnQvABVLBWmioH029gElVciB
hya5HOMM6G5sboEi1DYg15yWWiQsK1SVA2B/kYqctNsHLOWDMpZWXsiUFszDWyYxlwsNx7zazdmH
zKGAAsM4ZuNj2V08d1hCHJm87zZelAm+uK594JFuEBC8gf4wHPVaGty+TSVyq5BRL+ZGhz+4uEJR
hoHjUpm8YKqK6DvJUYjwW4S4RuBPzv1UZKWbvkvz1g7Iao+kHXZOxkA+VPLQwSe944oe+RQNwUU4
CvH3Cr7CA1A/lhp8/aVMCbf5GowKGp8fZmPLEQjiIO+zpG9YWsI0h7Ho0RngukKlChcF7y+x4RuL
0TXVQrJjr9sePggvRj7rM00dbxIMSLdSEVcfPITLHutc/SgBKOpQBWXd3W1hDRSKx17ceEt97vJe
uotK09IZT/ud0c6++H/lI91QbQd+ZObNtUu4kQFUWO6mikRgfutmjL8Fekyoa39VgM/tH/06TUWy
DC3UUicsJGcXQdYzEkLAHXr2TAiKukz7a2I/kECpTPMEeTR5MM9GH9hNgAQPHtRWuzuHUowsHq1Y
V7EITE1PGhw6H2BZiZfFGibgPYgmBotJuDhCmFidx0TsIGvoF+YjayI5h7hVEVvIXah6uF0EVXat
8sHR0tf5oGGhD5ELeihIGSDv/gIb/h33maynnybRPu5hx2peHqu4y2v/mOFpbq96a9jmLRqPva+k
KJZn5CDuUjolTv3G8CUuCyGg/GQ5UJedSDlDxAXnRRzkS++brQOj66hZ1XmwyLMgFO81D7w5shh5
aCovJH6zO9Xs+Gae+sUrJ9Z2JH2/fCetBnYLvSx+q+QdyvGPuAlCGe/CoYaEcmhwLlatUNqViBH1
PhPvIh9+/ZYh9nXiIbrZv58ph0L+Jf3ZvX93zoe1r+lbo11Fts3wuOa/uoMpgs8oxd5+aeLIoROT
Zmpf8gUUj+o1uxQyY0UP5Q9n22MDWCHgVgYW2t/lPNjYdurdjo/n0r2VfKnnunTS65fGpiqhd26Z
Wjt/L6lMk1w0XmdBGd/i5n/kGHI1us4Sz36VhTl8ieprGyS6OMzwi9KfFOTpikSWZ8yJVd1kRfo+
ybMyG8zvSM147J/TN+rh330T2z4Y3gzAiGxjkTBNCjhHmhaWXlSXYb9cpe6sq0aGyj1d0MBx+oXr
YmCPVbkDMKt+e+YOVMZySRLd7fozAG5d8IsGm0FvFMCYxNJyCVdP9KWaoA4P9itoODe0F6rFNlMn
ojmS2gyhyq/W6r14hX0Mcrgg2ZnHZXsnFpLTvC9oLE+MT8/i9B5ooqe54a7REnmGILK7P53q8OII
HifaEhxDnXynfpRu4nP8n+cYs7GJn5Dg078Ytrck4JBfFbMv6m4esW27uOeuP+xMylx4qv7bZ60u
87gpoPfPyE+TjaVR72XmE6QmzWKPSbkcNS7dFJuoez1QSJ2e5TmLdpNwUrFb0Uv86IBiiFFyBl78
NAF4b8dc4oKLqBPW4dksUnmWZrlcXZB0/LBsUYbA2wrmuBMd7nUao384LIOCdmq39Roq7xFnH6+A
unn/1O2aO3VoegX258oX83zdEgHJeWgFY+swpHaywLLFqLUzAN2Jg5SfJqvAsvhJQ0u0oTReNt4i
LHjSpELeJcnuBIcL9vKXLOpeWmuH1+36u7RDavIeK1E2CS8S8EjyY+XpFzHkngGhrXxP0uxTHCEx
r1TNlUyS0S3IP/lDrxWzBusVICQeroqnzY+B8Aw9nBVoiNzV4xZmd0GjeTYJ7PnLWTPjS4oikd8j
BKErYyyedFqMksUujl3MfFJJt9/UsoB/F+ddddEya62KusSHDHZ+kbqucFIXfVqS7OZQMA35bLVB
yiUoMpcVGhgwGtCzhpVOnB1qjkGg1o4AKkvIcafy5nK40WP2mzRSDhDXECMKA0MOk/hpktvQtNRA
B6dBZ8Qs/mSAE2v6XXJnU1XaiEFDNhZo9+b6icW+o/D8NG9Y9UmYPR3j4MPDJdbDBd5uEYnoY3uD
nPdixbY0sDqy82G5HYs2980PDQWiFj/YtJiZZ9EmviARbF1Dz9FslKywdVSMFL/7jsOdK4at0s6w
RxwE2mvr4R5qi1YPH5mFOXgly1dPfiRtSfHiNUAN+4jExQL7XnnCm+pCWhPy3LBLUn35yxI6Ga8d
pqLpkP2aLTJ83oYLpmq/5puUpXfwGZxIl1KPwZn7eXidMsxwbBwSqE+pipT45O9PJ7qg6k/elmcn
/su+opPlEYYpM7NdbyYQiUnZEnkZF6FEXpU1YZwnS/L4l0l4BD2JhnwH0aMteALWZ+dDOOoG42z9
n34eUd7ADwg9deloGw7IKX1d0VpZyCtQic/HVgpBC6m8+9HCfFR0aJeYK72VQjE3tycQ125p+eih
BB6lqNbrwj8Vp5rMw18jyRYkLsTLu/7gXTxJoZWI0P1nUP7y8lWaZQWlbZpGao9r66tTPdXKc/OZ
j6McMlhTB6j9DLxamxakKq2BHcA3Vp194Jy7Jrdr1LtwabPvhE4TiuAcmvgeqNCMEMOmFzkkqD+z
3lfTBuKIEgpRt5I4gRAHdnMoayPx123R8eR/8GGbV7SKkNvhkK65Y3Ip7pPUES3iJaSSKDocMr03
PhNsCMrRAsiJQ/gQ+11QjBoTuH6+c4+GcFZQt7ViFIOyInvXzsZVfx84lv8y/nFIW3c8NSUzdmVe
SsZDA0DoeD/PgSRfv8VIuSpA6wLy9Cgrx+DY4vkyhSVcxieofzgAY88AYtAFDWdTd5H4YdW5lHbQ
Bt2X3TEYFbE+wBZdz7Te2TN/iiCoTt+lNQggf3Bk88wu7n2maB+wNFDWHaYPFVn3HwXXvwlkWfIJ
li8yqe70CRm+NIAXFZfMjUmVydWa0aIVX1yNdRvmPAvFgALhmQwuGeMVsC/P/npVsvc8PE7usDrY
5+ngk67zfjrkWXE/JmncXDeFT2Z3IVuma5jkQSz9khu68duM7MXnsHGDI+tI9fPvamHU3CeNTGVX
Q8DqE7x6LEUp5babxRb8kEOi9LhoXS83orf8Fu89I7ZrLoMyexYspOTs2bKAoTAD2iNXl+hcyFb3
Ndi8/ohjhgVWBDtGz297UiW5iA59tJWhE2fbqCSLKr6TOe4vXEFpqZXFm6Ywnsv3fOjxCarvHbwg
Fzof41IPzpSvpr206wtzngDeoX/A2qrSeW4NsDp7WpT+yTnLA65qWLWELtuKHl41AJRfYQAErk31
Xv++pdnefEpj0BXI5RqKWamS6m7LFB10Qhe3OcfWLIPqnOEPr9xeBfw+ZjD1mGF6b+OevO+Wvuxh
1Kfh837wZZqUPhe8mpDENdTHCQhoeNnLmRSl8sUy2m5mCN4I3xgrCw+GkK0XOi3E+qeKS+Jsh4rh
UFL4pZAyrhCaPCwMYJ0HvKwVMBwxLIN3II1hmh19+faL2oYT6lV49A7rfsev6xohVD7GLww2+SKN
DhpmY47lXI8jKwBsP6yTvLNNGB0Xw0uVhCpoQHx8m39Q5fhOYy9aSiFDKPrXrHTsR+iPH3JOqN7s
Fy9WqWN4K5A3u73lCPizVfxlFYME0O8zjxjSGFImOb8O0mM2eBty+jepm/tyta3bXsdR+mCLZyqN
FGeXB1JE94eBhzoYtsF3vmbQJY9Nu7zzDJHkiDUv55RpNUZpPbH9pMslItvJbG/rM8Kc4Ie75w+u
JNGiaviGCmHNJHcpVwYA7BapL2dhITYVvCSVrxZ+ThjEZGdmmI8D8SIjNghaQmGlYneC304NlQ3D
SmVglithdGmTnF3MSkLgTucCzi3PNk43YimauGqoUiNoVpzUVlKj5yF/aPC06XoCq3jhJAYbH1EP
AjFmEkBFtNuZflgIcAYPm60N3MPCE9N9k1cIMdFbqfnx09d510eZ027yK2+bQveCzf7K7TTIt95g
/AJvXdxKKf5hVTsYecmP3gvW0op/wx32W/b4vlm701BVd4R7Kb1ogLr6Po4DlUA3QCkJZrv1SSjw
RX7zu6iV6cPHs8tTfnY98VLuo00ySkTsnXCWCItDK2pB0x03SeUzXxwAuzYDlS1qtkOk71cZcjJR
lY0noFN4TCoO0p2MdmRmtRyrsCx74nUZGkTsRuyW6a2dzCn3tjZDedDDSoClZICrFoNgR/yEHbfm
jsdxMsQtdHXA08/FlNp5NY0+NQx0DbR01cOE4USMRO5VplvYHXrvYO7dg1iz+vhN9tG4Yf3+Ievj
wJWN9HTXWqGgVUutYmtnv0qFcRjYYy+0lUlFDXfoXU7NYOvZF+YMEcwLoc7zOCDVBohkvwoz+di6
XHUp6o+sKE8Mt2LYWrvoH9nmqSWH9xEzomBrSkshWvWWQb1hv4cEYjr3EsBVfQ1RRQtvX549RSzU
o96eMaUAXa7yJoE9lbtgARoiS1/KyhVtrJSvR3A6wY4aVfNf38o2O7A/2wks1wW87TAEqtsQA47S
9L42+2m4o54TkLhVfNZBd0AU+cQyVpJq+QYxmZWrxYIkHBRSlfavmTHqRjH8H6R8AkTYmWOWpFyK
INa4GM6d6JHsO5fe7C1DpslmayRxpfeCGBvXXRmzWKbFwbEkjagfFBoRn9h4MMGrV/aftRaUxGHa
tsryqvRfQ6r5WtInQyMxNrqjBzb6ugnNSHqpPAUa0WHm5nHdeZWY2vsdTJXJONZS448wDGasQhWY
/W2lGF2E6F6jAZ4IJqc+KMKEtGg6oMnqbP+bwyXm9w0WrFzzRsTInZy8fUrviMm/1W6SCZtAe0ZJ
cSZbB46WLOAiZpVTcqcOjLB+CKwHkF4mvrhdPneTlAY15eOEJxJq7Qw2JB7UpGeuC7/+ZIPdRfhU
H2s+nqimlzK93JciP76Cc1dRQWqqMLf4rP9ZV0WzhmTkFQV76tk/fgHcU5upuN0XJAzfQ0Pvu4Rm
+GjbZch0S51ve5A9FQh8UKWMVXZIzT7h+/yUl7wwt4vEqN8qy4EVFznJHXPrsci9W3vn3FoXb92W
eBcCUJ4kIJ9DQB63LeZ8/tHi1JMi/nxXagsb1OwWDcrQEB+l1ZenxQ7zQ0jeb/s6wT7dYCqPJa+c
eNEw0J7CjmoqvSe1O27OGvMt1Bp/f7dd8BtapcjaWJVTZTy1mhA8emXwqHXrZ3Pk6hDcFh7Kmkj8
b8OFh3UtAoNg8I511cVwBqMgjdITZCCttDx7cZf5jDB4gFLa4/1ZA5akVuFPZ7XLcFmsqGUitVfW
k94R/EN1kbq6CiWeMZlcenfqogPi881gW0f2ws8iVnGmNVqOJ3Prs+enKkh5YoEOXKVFO1ig+EmP
Wkv5XM/E3kbrlR3nGQVTKFngakL08UJ8SQtsaPumz5ouFVeJGqQsPvKN+wCjBaMUeZ+Xa2yXxF7f
xsN7mVYhY6Fa5oZHOG+5MD+hOtvH1bgrDb3vfR5nadurn9FD9cOhpYd+SzChVVn1xeSRxgVJzyYD
x1XSM0c39QgHbdvTGL3y4HB/PyV9xdtP5mxTi2uyLnXZ0HyM+iZWBIIP2WS38IQpMf6+FHGRleja
EfhYtnhdNKYmjIhrF0V0RdxQPLj7mSONzPwy6XXo3dNHzb4ql4YyK/ju2D17j1SKsWAkJ/3XGvAr
xQscrK+3zzT+X2Vmhx4zKGTAl5nm96jkG2cNTSGOt0bdQhg81K3KbqsQ0elYsJWQFL+9SntjB+Ly
yN1R/fpclcqGgXl+DsR1u7oPojqTOpRvy3t1kGef99y5w7eRPQuBfsebeGqgZ1rxgJpI9UevCfAJ
aKrI2fCqx4e6pqY0xtM5kdSJGIMQVQJ2NY9TD3ixgPccTge1xrfODjOYRVLqoG7lBppeAA6IMAmG
/USLJN3juPreRPZXLyLiiDthKSO1iFcjEGtdVhvX4dCNXyO4JvWyNEsX+AXfnFWRDTKRAxV91Z0P
24M6QExn9lu3sT91wOh9K1ModhWQ+hDTRFsOQaBPov5vR1u3l6vU1MwZPZ8t28R9O+GVMz5hJ03x
1iYe83ecGSS42cEOH4RFW/7DM/ldylqvSoaApQfbnab95BS+fPGjUJLIlVCu+TeiSxIScyk5VQqj
/NXLcqWSjnm88M9QDMmqtS9eqsOSJLXstB+/ig2ZMI+vj2c3JN30L8c15anArg5z+r2wXvjZtl/a
Rqv32ZLGRx/Na2+yDTwA+q1XpqEEE/MKNAPj2IAEBhnOnNwUVS2UbQ4doBglylpta7YsnYZ+42Ew
v9LLQaUw+dANyabrBA+SIdF6P0m6Ffmfj8KW15KX3YGA1+CasgKxYbHCV6OByPehR/NAg65D1Yj5
J98RpRDtEUzhUuVTPnaX/znaxksO89rfjbweon78B81Frg55T7xyrNAeFBKQgPuwz346SfPd0AZJ
SjFkl1KRTEWLgHSfu7f31KfewtAsYkk3iqVuuupyhlkRiGXe9V5MFW8Dh9wpTrJ4MG14yYmaKqtc
eZeZh5MXK8BBP61/fdC/kz+uPu+xkRS6i4EoGtNgr+hucmKoLSsWaO46TcERHlI+aeesi+MShLK6
lAViWtXiBly+Y6O+WW7HjJIBiDVuybFSqr2bhsVjlOZaxKar/HsqEiOQji6vEJxoUPo3rh74qG8b
0s5GY3Id9wQoPSLSBCrkDq2z7CDtUoOswcF2abCvo+HOUuNMzmOhyCIveu2HLB5KUQi1rbfg6XWs
Ynq8QFbANJ4WfDB5VOGFjer6OEFbxQIaGkVfAWdc4ncWd9Gm6B3cDsD23JuavHmkZZpw6WRouR33
3JdBhfzozG/yzpKuegI/TA5MRHpcMI093kursl5S6klmaFUR8XtcXleYBs3dVhfT7Td1dIbArT/r
421kcmi7+aDVOSDernrRnTdbkLXcsf7T7CUjYrsf27sVw8/O7gz/xdIl02nMORmNAcHfcvyxBLvZ
Wmxct6hlpzDasyn5jiDIXDebMdjvCUERzlEX30tqy5z43FgDCR+rxhWHbFY6KkUd7P9gurbXlsA/
EHHLdCxw/2roXa+jvWbHe7CohjOO0w3KVQQqGUHlnXhEdmZVCx4dIuaXU6Tgz022v8m4aqaShBVs
u4R2WvUFbJ+Guqvw2HxTkktgrzUiKPbvu2YBrjUR/qZzDa7+o832cdUyS5BOJKgUXvL32yRns/x8
5KIP3efpg7aB4CuvQxVVerIw0UVX0qtFIKT6vbsq77jz2ufiZRnA4MJerMrh/AFM5I3wROXFfTBs
U7b7Y0HHyHdhKxFHTNcN3jRnnXNs0cROHhW0ojlA4X9IQ0ZHPEZcLq1MJA1I/RPF6uMvdKT7R07P
yHsSxHbwt8zAXaoUDfjy+7LXRq3j7n0eVM92h+rEhxSDYXozFRp152xu7kYoQvSbs5SlkRcf9r3H
UFS8NjH627QJB9kLdLOog6WA77A+9q91sp5akRo+/kETpiI4ftr8wA3bLowKqGXT6+4f3rb1zo95
pOQgAqh/2ifVmczP2yJDPvG9JrWI10uQDJqcVTU8VfGYO5bRaIv865m4xoAPjRTEpi/VXFsZ2x6X
LJlY5srZuCdniKgDHbFRjLM8PKXExE6LG9rpUjW0agP9yGr5HPGQ4+pXSS56jFF9mi4GwQ+eZswE
2xfUJozNRAZ5WBzLcR/d2UN648wq5y37jp3TjVbhBnf8oc8oJGu6DikBlJqr5734Eq00GEjSyvaf
EQvnb8ZY0w+uyuXIJTN3x5F97wt9Zbkn206XrsQcgs8/dc5ACl8CM5X9w4UYK+9kOrcsWPla+FZq
3xkmK8Q86sh9nMLguXXB668PP5XYnA0haFMkmV2HES8eto3IA8aO3HG7tJOgFA/r8EUnGHAfTORF
lsgLD5A+uceoQ5XeKl8DW+vdNh5uj/hYCX166S5AnSnnlmjnHW9MraW7lwQ4YShASmutZuBX5DbO
CrMTI21YUWHENSLiacAA1hiefJJ1ceEjHNILRoER5EDFKIBXRhfhq2qN5j+6COucE8628lxSbU8m
A2O2n34Hl12DDRWSXP4lu7jJFs3wSllwqn5xnkJiXkJEVTMmaOeWoGn+p1dEoq3kuXe7CuhdGENE
zV10kRmZHVtJ1IkcNVUr5RUdJ64p8cBLWigeG4Y9Sg2X1I83A3wg8X+Sux+CPVd8Ci+7Wtwg7Xte
hDoGpXhDmYo3iwxk4Dwj+OZzzlR3WO/O/mGJuSIlo8J4y0leQW/Hus3Ij1fVMyf9VkA4H0yV3anq
5vVlRKrgJ6j1uIo/Fi+k2RD2Cer1BRFECVVNJP44LFDiXRqAg9G7wmaZZQGRGu47cw4o2nKj+GZB
VT+w74PlFoflANF7eAmkATI6lSNzxWNxd1uYjkbIh/sRNpzRVJpLJsIwaqSxOhG9awjg1N4UVl8o
+ItyLgwlIdyMqfM6bZDI1ilQI8jsTj3bBncnwLTJbZt+EvjfwJ0XvG6w/5PWZ3xzpuF5MeUo32Uz
IXpD/Ak1U85hsdm8mIIoBX1YM3zB1a3FEMsAxkdIkFk3a10w3IBaVdYnUvqyqx27clLD+E9owLvU
RQhPKDm0qQ1rth9eSSiAzxC9WIfGHzvzpMJXiE+FHo8CLcp7ZP85+YMsmmfnIHeAKpDl5rOnN3VO
mA3uJxyuJeL9d6oU6Lhbqh8Hzcof0FAnmBpT5rAb+cNbjOOMduupJEivIZLam502O9XdKqD8Jf6U
2WZ3gkxc3NgBfnYvqGPAycORjhHKXCwSRcA6yNg+cSXKTZi8ap20+XOFtWMRQeZlqMmWZaiyGIrp
9emxDNyIv0++B/TEX6wqJVb1oWjNHzBCFjSPN+8tk067psH+r6Y9ThoQCdFS3Zo8oREb0rg/UMG9
OhNtIqc7U+euobpqDiApIpThC4cJwM8YwiRj6TaYCd+pabFuBFwt7FoaC30m2eUA/dqPRBkic+0X
9fnjVUM0OriJkbUBAT5gy5jjCydIMo193AlaQOssUH8sRcUMgPhMGZK6ZZFmkQxg2iO+oGtLa3Rq
pAU0vnL9OXYLHjQ3EqjyesIvV3NBXe8dQs1LSisO2lRFSACrpXAHnFgDw63RSGfQsWpcA5JODbOM
tXKvLhenE4ah9xiG/smcCJCe9eRm0uiuggDUUbEo6nGe68EPcbbB2HVJwiU5Eba/ojnIFXjP1k6t
F6aC7G06d6AJhznCPObMtvP0PjekhrEqYKpQTnie7Vyzg7py/+QF6DQNxlDN7McKaZpID9dxfbZw
Pe3EInhYz8ymHgT4R17+H4vzywGhM1XpXwWVmnVEwY8d6Z61z9C4+xbM6zk7icqH6ztfAi4IOxNJ
fZxR1O1aBnCGZHmmsbAJOIwVdJ86dvkcwpmoexYWm/mv1guHR0nnYVM7EcqaeV0q6r+GWWrWzCsn
z3OgGIfYN0+KjZae1fS6WnFrGVzjXMDQefPEq/wKvvcY++FBoiFxZHSMx6VjmewWOCZxnP5D3Xpy
1nxpiyDtgBkCUfrenYC1Wed1xwBDzz0L0DvX84FHMSkcaZ3U7FGIsXMpXjLRU8lQgkLIW5aM76+k
NZBahZ1HUaGP3bfncyRKXM3sUAxNqxrEZ3SaQlqvszMEhGBdM0EMIdd7zlGMbyLncmKKMoV4CWy6
TS+QHa/CYC8jlDZ2PGFiWKfvCtAjgXlhV7le4V7CcFLrj7ZpZQlvu+1MCbRvgUPKKC/mI0/yEYXe
UrZVZHnxD5lVtsUatmXCoGxiHrHZw8AqLSZ+rixWr3riEUmUIMnMWudxBrY6gTnBoGFUBEGS1FmI
HPsDCqlqPYln6hnBq5y5qSlfQZH7+YWyZkAAMapedlqGhVUJmOegRwt01jHYWo1rfBwUMFSEqW/W
oRZ8enZaFTGauwX5k03a2+GLYAhYTW9W613cf2DK+sB/JwMicYbeY2AKGzUqPS4WpmlaK28xMEwJ
C0HmBAEbRG78Cb+hReKiUmVPtrv++FvJwG2y1GpAr6LkKAiZsIxYXqzRjR+hUznLZfXI5aNtr74K
R5gEilU2wlOU+vpOvGh2mtCvWNuy5O1Bn6JJJmQVwbzsPb45JEmg+ORyORdPCy+K15s3g3ulPII4
npWaRkLtXzkAQximJ0aR0H48XT4PWh+dqLP594c850ohTDtz9/cMrRaCDfc1NWnt8cE9w7MFiHSi
FBBtnN1bu7SIuV03NfpFs+niW5h1epvvdm9baeUHugh0jPKMF2EZHz7H5JeS1vaCnQN+8Cd5ogfo
FK6yacd/+ui2Qv7WMpeHuctp8xgwc/9EAGSoMIgsnwAL/Z506E/g/yjnmBCygGdnaaFJXhlNlyB1
DPLfBb43sypEqMlmfWAd1pxH9WfxviFiknlFVmENCcJqXjMKKvqMiYVqD9I7JXW6MHHbBQqf2Hov
U7Vc710mPXlV+0GE9/elXZDiNydQYusjTD3QEJZYw+fza+tC5Wqumv0ReMsf1Anc0Wz7OI2eCatJ
WqluVtzSD9Y/ueesoesgDMxj/qBJ0NZ6qdERDm8rWjU+IsnWIKb8+6gDzBRYaSDXMIOFcgei7113
pk6B8vuS0O+Wpu96MeI9ZGhU6z7b4WWVx9yLxlBvl1CK/uaN/U9vCmKYSR2U+A+0fG6mYDT/sOIb
MuxfTiVU3MASmZdIXW0gl0IjZzxd9WjBMDTU9fQS4+vzhHW+Isxyyz+KUtJ9G/gzEf06ry2gnwXs
vdT5bLA/pJWefTcu2y2BhCIeUBEN0A9ep1iSAe6mUX/Ma7YqjPlu93ik8OGqeRvYhywvJv2vZGSI
hDuh+o7jAT+EPqMExXGQ0Q5Kk/XCeyy1W/ulFdzmqjDJr0luAWAMwzQH6lTcOOs8+vZ+NC5rBs92
YknXypdBTe3qaAON5UHOuHV8U15dh5Xtm9ZTTbTpq/4lTda+9Pz5aEV4XfnlmiJx2DuugV8om8uR
OB/Bc52eOI7vfd6P1oQeSVyYEa24Iz6hVNrMHxiZ9QGz9JXErAj7irk18w+TibffbNSBzJU1Jesu
/jXup7/rDAHb19cwDLHfOj3R4b8LGbo9gYZRecFAk+3T6BpB6Hjg3phDVIttx+snj5q/MLT5yNb0
Z7yLkxYlzdX+co9PNl6irloI3AndPfa6Wh7yQ0L+l7XnBOuKfSoVK9lX6p5BKhCJYipLB6MFzbSZ
ZaRhBmU3/Ce8o9RLmS4O2ZnNabwRCBycJZ8kSWBrMg73thCc6iIHIlt/9ue38tnwuAPhUUOELpRS
73bKjR3M9eoBX8+mBaCx+JRsqbur/HeH72N7mqQEv+SPg0RXaS4jTfzAaD9IbX8LaS+Va3YhTFF/
5Q6ImqxUAsRCe5qPwaq6vBelImk9Tpfv2kzTNRcsMvo0Sj0hcdRSjI9e+grgKH24s4/Uh7XaOXwu
R8K+egJDGgu6VFKhAVfj4Jg+Xj/fWwFdASx0rAtoH19Z+kmiuLSoCjwEWC/JI1appsx0JY3XTZ2K
udYqh84vaTZj/VS6eDX+4yezRNc8Q7tU53tRwTlMI4o0mb/b9OECRy/CV8rlRFvfFCopZCLdodtE
xNOYLLQrYhzV4jQe1LfhEqtzakoFY4bBXigiiCVHn+/SKDlxAVgeJsVRZz6rTS+KQx96qXXxGdgU
s6pEf+P95SoRt2Yv+oofwRUnEp0XFH7q+HC/rYNgFFwL6nJaGi1ghaJ5NvRQo6yvfO3I6ZEnbB0+
yY4pspftNKD02Eqb86vvER1AZIUGA2OjXAnxZomqBUMdoW/sKzBRezBKTsBIjcvD60K5ipqATaVV
BtYm2ti9tgTkZ8XAVmhpgC+xWQVPpWL5dTyNQqH17KkiznDpGjuSfgpJemDfiGKYMWmoY4fYyH9l
HZ1ZHXxVGKKD2sHOp58DLYkwE4yEhyz9Qq2g2DutzF8k/IE/XI1fpD3qdPctbSgPGjFT3MqkfyKm
2sYV039YXij8ZOSkmzFaFpEXfhtOE12oIOVAWWPV6Vzv3qKmDmNVpcA3qWd4EDOIH39zZfUstq/r
lr01Ymu8nhf/Dg9wmax8+28NQS7TPh4z2ry/5cpsIOvlSQoGJGd+gVFxQveoQx4/0FuSHA6OBv/S
D3idyLLwjJrYFmekN/rmiVu8o2OUYZbHBQU0j5LPCdbMMGfSv8GKG60KUr6ikbCa07XkP9QpazTu
Y967kueU8+Y6/lr8yWN4mgt8YqfoMdxx/Yofq5WwMru7AkjD0CaXo9hWGK1RoVkITYvLsH9WAy7v
/7CZM6YvPzz8QOwpCrcO8GY9uv/8LIaDMitzb+DU0IA56lzNl9xmil3kJsHDN5O47Eg3+h09mQ65
5srWKgLZy/1DvEMy/d4tH0lRTLp3+qeUan0i9Mphvc7Acs3EqFNYAXLhuBV5Z0CJP5h1snFvqsTW
d2jOyBS6jZd3xGn5aG0HoVLw/fzrAd7ufQXa9NLjbQw+D1JGiwUgcfWnIGxo+WHSCVI4H0lgDjT5
a+mSwFGxPwkyGfo0lKQo2hIX78v7cBMEuh7rnjxT/MqlQnkJco8vaFDRTGBr7A+7Q9O7FPYtO511
ptwx2HK1OkPD4oUr/q0uW844cgkj6D2CW2zYa32XegZixg9tn4H696MeEngEHezRnDHkfaqQW8ts
XfatB041KIxqVOSBcbSKNN6bZJttyBdIxPYUOFDkE7goM7s0vOn5d2p0DmYlJsffDAsQfD9aQA0R
Ka2Ls3isck/0yiAMuSUDUfWRGosRJ53PjXytg8GbULUgJguiKvxLkrlkqjkSEWlIK7RiY3cWfKk/
HkEGHRMGKuqk2qD8up/oK3hWTaf2lMO7C7YQNjwJTUkbop58sqUJoaZIWfaDOhQyZ6JzepTu49V5
0g7vUmrFSa30sVKJDZdywVn0LZ0/TTydifAnkUR+Eowhyfx7ZrAHS4UkvNjpn47z5PHu/SzWDX31
TeRLPcEuLKAmNy1tVSIAALEQjFNFMcEvDkUAwoBIo40dXiiQi3eMFP/MX5SRciyjkyqbQxuJIgMx
ulvlWhkAQzBnj1kewUB48E129rMqBr9oi3jyqNWFQCoUgu22en4ZRyd0cEmfIwuJ5hXOfahCALDP
BF9Kp7rOFCAT1YgHSqg8aV3cCVy0SoCqS/xAfMPe4YjXxAk/iGItd8vO942LybzhdRpeF6doOp9b
Q0pCEBxPRIV9TVYEX8v8xQEqPeFfujYfcn4Pp+gaAZzq6hcSC32hUYqzbS/KCXIwrfsIYktzIwXe
zcuNNUdocg+WTSTx/mT2V7z+bLWgFWDIxM4ytr7mrZSHu7iiJddy1bxu8EjIxNaiCRK0+QzTk9oX
THaaI2Vy7XOMvFmkAzFYPO0fpOsyqnA6kd9VAvNkgrER1fjHdTJCOBvnpNZRXk12UfSdi6f3X4Ay
1p7ltiyg15k0jtehliOAcyOBAui9jYjCKR+jdjA61CxA9z/xiokEywg3BDFEZt8rKDO8QzEd5how
FRBim9b18jeIXuiba3FiHpNYCOl0md935758o2pdAHaAPgtfjw4s+GjIHHL/vgdpsoxGUy9mjRVU
+5ah3d2f/RKh/t3D7wY9OlfJPGKnH2HoKOZsfki0QdaLDvn0lp2xUCPsK7YA1kmnZpjApDBRuGG8
5x/X+KnWZMiF25NIdgGUJbyCgY7ZlzeUW+BL/cEco8f46WJY5G8O+Nx97bhd4HLZZRjYgJMyGiUS
Not3e1MDlP1aRQAylfkyT/AvTxjI1EOPMv+UUkyFZ6OAfv3z/cU+J7dTqxH9UEv5rMlqDyv55PEM
EAlquEmElBH7OmDbfk9I7F9kNNnOcXgRGEtFo/2aM3ohQpqCj8+a82D5uP7OjEoC6va7+swEPG8z
R2kNUXo9vi2Tlsb0rDqlIHPpcuJ7eFHHcdILoGZKfq8wh1th0Iuwe6zfYqKYixwpWtErMV54SwC2
cXP/nhxctQp0bBHe5dtwRMBTfVG0Du8naPmYoIAh6GM4SKJD3di1QbEwD3tfEZfz/QnsDOwDzVLC
kN52zOmjTAfTdCib/gnzka0VzpCcbOKaOMjyVY1jPJoXZY71DxHP8KWGc/gPInT2iI1v+wViUc3A
jivJ2YJhR39OngC7lP6VA/g+t6Rq5O5Tlfcj5zcq9LQpXbCOJZ57neobqgadAgUstnVYCpUHg6K2
BfsgOOryuRlPcyk4EScGAWYdtJTJrxFAIxJ5bj7k55+F4KgFMRtWzALEu/xZDMDIk4EY/QWZre12
xg1hu75rCbQN1x2lvTTt1MmDZZkSAAi/DEKsTwzij6BSpOSzoxV28aGfmUQ/a5b4W30KXU2CAwAq
oO6U28hyVWq8vhOx15TIZyirzCkdwUaMifU8jpp8nPtOAIWIMsISbQuG8avat4oQuCyW3vr9K3uA
+nXyANzf5wtiSvqBqqr6cL9co+OVyqgAK/6aJUnJjoa7jRe64mBaPHBoNr9FtDoXEHK4MjKHH/2c
siJYXMza4R/1MX4k+KQduhryBea8mtidupV83kov7pzgVlPDNiPE5oz1burRQfUKay/W36Bzo4WZ
JPBWbQPlv7eXxmTCvIMBUvHiDwX0mS7beKIRC7F65ZRjAW/PL0lQYokOlGGHMdaFzqdBfR4FXL4x
wvECpSP7itNQxcjAzsCGmoGVRHf1J4H13Yin3uyJ9dYDylvOJqsZyIrRDVNP5/tas5g0GXAYYEQR
QrXSEdq0iGiB1uM4GW38zeYNBI7oXVOViOGtEK4DHzwwP4fVUfAOF0R0evTSVbqUxoPL3CGzoXW1
H701UPdFNIe5HJVgh5dvukGrKx7Qn57d348DdBDRI+Ths13WcI+JrHjj+2+VqKMpfuXl8JVVD2Ff
/QhSNzS//DML/fCBaNohBt+rc+MDQViRKQrPvUun8hJDREpA4LKGY8Rgcj+v85JPgpgiKshSB/k8
YI9F/8c47Jb/9ZedFXWtUnB+4OB1C+v01GlZTwgP++ksscrhgg2WBoDwWCyLunO1A7uQabBRHQa3
XWbz2FltG2lZbmj8/bhN9MyenWfpT1KzN70OTWGrAcslBh8yAHX8IW4zXs4OvwO6xWp3loQPAKDT
PViGjBiGBOXH3e6/hhKyndN5ueAupM9ZbS/gxGdUlpehyG6Gm0C+mL/HzM6LzvfDysSijNpMH652
jZViuWgItUGTsvt4+f9Jx+VUbgx+KoO/olOsR4p+B7V3WUMY3hNJUAEFqHiKJs6V9jOEP/I4BgDl
mEjDY9WYf1h+t8p6RZcyMQvw7unjCnLxt7WA2D3OueeA1fsUQY0OiENgjz05lH4tGN0REs5Iwg5n
EETG5YOoFTXnM7GTgqNSQkxUi6LM/7I50LEsrHgWCb3WxMZJt+jOZhWZdg2CaQ3N74aKBkQDiKtv
LKjgrknsEbZRyDnu2p3Kd7zJEHhLmD9YQxsie13un7RSBm1zAiNiQ4RIjMUZGec/NQyBuVINj62F
EySVvh4+n95dOcIp9b09u4CgwelGfkUBQltgqRxQ6+EIM07K+odF1kMn8pZPoFbjyyBiTTfcpCO4
LETHF+/RsreJxAuEr8yW8WLXYRRNB/hZPMCPoQLDXQ0yxwFJJPkr1HE9UNt9DSb0uy7dCC6fUyr3
qj5lHULUWAD83z6wtKa2is5V/v6R8rVGfiVkd19Szn0mq8p+pS858oIGiSjBqZQX7qpJuDaM1isq
p/Gd5+AztaMWUeQOqKKeKWMGy56Vq1tYCkkKiUaWaZ4udo0I/nPc69TGlCpBQV/s5G2qR9s1ZYKD
UoNHgJO7Wa++K0Fmg+3w+c4Y7tyxTfIZn3xDBynzBZH/BFryJyQrxFSHcgi/e+aactdUhi8ReGM6
AiKHRjibaqi+upghuToGftzGK5puQHhICx8MXRAXzaskhO+ha4xpUqUW7dGBViFodIpnuDuwhsQH
p/RGCmP7k2nqFr/iBXUSENeKOekApkCMyG9o1G3FsMmnu+S3Q0aC2jwP54amtRzQCG4ycwlPBJEE
TREQ6JoZ+L+bPtgLQPLguqcw6iUe/I/DP8lJWSf3JyRivask0y9AyrMg5ZM9GJCLrxkOgF5jIM4P
ARNjNxpzrrfin5Yqq3/cUU0sJxOkpe1LqvdtxolWBtY27Y2JHRoVTTtIb+pVtezu2zqBaCnLpFA2
jK/xyTtDb0tzSRMRd5EQQmbdcYZiKH6a4Y12tUb1by1l0Sj6I3v+rMPvncK3IL7ldaAGZ3crb89J
cUtykGR9ZFSLl1YNbir+nBfd631aL+x+vVc0S++9qPVsGJb0ZFy5upyJN1wcNRTAuOdZiwR0CpPb
hDSadYqZlVkum4TVOKquR1XJhVyvw3Y782pHDHssiS2N79vm7e0NMYXYLud36rYFZSK07cPZj69V
YRkzaagpcKg90cCtmEhRJaEnS+hkPrkDXTLdq2OMenJpd34IFkW/VY0oRttoFaUmrVFT1qp/VzLs
WwJKtnFQwXx7H1xd6UW6plUbSu/kZIYSN/Iw1LwGNThiW/T93xLDmzz+EZZyFF1kHmb4cYEDW/B4
DFSbSYyImfHelPCTfynreW876lg/Mcny5r1/hjQnoXnoKNzxX0Uo1VOZbVbdAxSolGxciV+NofBo
aer/XVjojls832u44ybabFT62oXLa3Wgl/s7gCgUUXzDUj7krkY1poFUDfNQ/AaIpHhOVBa9TiJg
NJeCqTogeTVPzlvrV7zWaNKBt3c7t2LemF0tW14SAtk+CG4lUsn4WiIz3UJcCuqYoxHswNVyY0z3
Vtb6PtE53U0MhrhHRXNnemuojMRJkBBNvZVnfV14XugZTZTEFM0a4EI3xwObXGxaBKxEV4oDf90t
PAA/pUOpHrzKjlwZW0DKN4YB+rndESKDtN0BOTdQj1CjRgaf0ecrx0IIS3YjzjjYKTu97Z6V589e
tEv/tVTUIFPYbwmjfDSa6rnks0d6dHxay3wG0hcZKbqugV3AKgJ/B1AlKSmT8/MbF5PZM39IWKLA
cr964QA/ZZ7384A9JAul3FAdMbC63RX/ysRplyPC30icVbDXGK673Utpw+1Pbv39o4G3PqolHMwV
IJ9KsgnbWd0JTvrNgOSRyQ3GLNiNoH2JraOF8LzUXPm0/kxjYDhlm23Wbnd8ZrZyj+4Akxd+DyhT
lFIHn11RSUkd19nMQQTpzqMEKdyfiPGUbI7HI1yBP+JhHctcTOaaehUKDXgYvWuWBIltAMhKYWb1
aqjtvkjtvbvRzADZOiMKxLZSvkRP/JKEG76BFqIBaSAlWNgsj974kyfsqDNvqdyMZt3dVxBZsPRn
pQOtiFXHBvFcgMIGqZg+u56dyWfFfeNiHsA7fmHe2WfzRUJ6/5cE9M87ME4AqpJsplC2N9dxmVBv
gQc4tF4vQ4jx962hQ/IKxvZfc+S1tqwD0QQHdAjeSkEHCvnGogXP5edREcQU6ni/hlG7LHVEB2rU
Gyenwnd19lgBIP7+0a7iHxQBhnt/ik2yMP7mag9IrpzNGJSNnLxnsr9KOfWeGwt8/DS/Q60+qOzp
3VlWApGCGV80BXs9UmYXTASPJ/6/thG9Hpqw8ByFINTlZqarvSWqBqvXLbdfEH5arwkN2LJrQUyY
Hm6j8ZcRcL7M0YDdmnVuKYJEnefHWk6L+qeg3QmGHX4/IRtQ4adrKPxjcnF7W9jn5/JfOZ1NXCGd
oE/j6VOg/py624tRS9DO33cIfRw03nUusSy8oWGoT6996Oaoxd56PgUB4CCoDtza8x7Me62q2m5u
RRtckUxuECIlRWyivSdKYU1vCLRKfN6rzUI9tf3AOBTy0b6Wt18JsP8zg8O9iwJ2vE0PXM1PTyKa
8oE0wg+yTNiWbHYjy0+7a4PmRDbPFPDc/a5O/30TuHJPzmGroGZaQuMrO06BDUTkCqqXeFwqcIqa
KlKI29hqW4mSiKc/C9RypjzdIB4ExeIxjbY8MCitnhREaq3zYLVDGOAyN8/vtp7b2CjUH28ylmCc
io1Yj6bJkx1Dl4BCcRjJjVztGagL74hAKbPLkYnPbnW87jb/nzEEoD65B9cNhqGets7Tr1fNHKo6
tS+xJHD3twqKArHR0ykYFoDkf+QMAjeMma0QPYtiL2QlOzhGZptIYaJGkjoRhVi6ulYJenUEdnGT
HM6WBJor3I3QwKLo/dpptOp5h6fQxIJjrQfIpV71nDUdVq2wNH21tCyxxIJDLarcR6pahAXjHl3e
yTtPUfAqlJ2bScJWVeQorLEtKUfsGwr8fNKyVZVhzBpVbgjhvlldDQByKuazMXKchfPz0KnW42C0
KADMr0vHLE1hs1/0QB57SzuoEKc54stfOj3aqHJ3LTZmTLT7mce4MGKbCyMg64wJ/tMOBzZTQUfz
vPuqlyS98LKgNMv1d9nedJnX4snd8J7qGxDJ96B2k0o8J1M+hdPgdE28wQlMjcvUKIkEygym/j0m
yqvsPU1EK20EhNEQWxKwxHBF/olfJJc6/DA3CDiqmqSIR6CWE4PIvqMZMrOQ0FDDqp9q1h4rSR0D
5I7mYNzUhPxaTbLEdBmL0ghFh5/R1rQxfInIU618XVGnt+YNCNMHaPgESae0VoJZpDw1HeQd8XV6
ki1zP3/uPPplCdZ+fSFCrpZYtKjRRNOgL7g++tPPNjbTy8pOvZNZrbhC8O3OxG9Q48iw7KzLXhhP
3D+VhDPk1TV813fXYk/NQM+9FkNBCYlIg/MneoMlkHXywM7Qy8PRjO8O8WsTSFwuSHqBEayw/R0k
FaU49jyXSogduf5quR3NVhl5qnScMQTfqN0txa+nifHPnuiszqFqx0o28OtaTsrk5sbZWnerD939
oWCdZNzWIu1/QYlAT6b3SC3+uDfjwgrSsqyRmU6IwbTW3Gnme3LyjNVdkL40KjgRyYZdtQyPedyg
uYz5haUtCObBaNFQf3mlaIHWCIvTvWIR7e/NNPqxqz/QNogdwt9pfid6xNCSn4CNxOF+4oiiUmYY
VUa+mqPn4cVrOVKgNCWI7xdjG8+S8neQ/9CWJiGlM0Ab0jDELfKzwzNCcStgYiYoZFqhAaOUZBJT
DzFNSj0fhA2MHwclIj4JJApsdWOmedVOFLOfk8kzPw1ZpCCWQVW6AHmebHFTtukDkLK3PnW8Cd08
xXiKN959aOPXqg8jQxdT9FqKg+57qhCVTmONlbThItUKs5X7heQXmgNI3NGfkB4LPLU7QJ/NMaHM
g9ulShin3wLTZsmTTk4eVZbkmRwVipDwrL2n4gCVJxKAyfngt5jwNNPX27kBON7mQOwc2HwJfXwh
5Lpw0fOEHuMEDs4aSNnOXY6R2yA+u1PI0O9Js2EP663Uw0v+4gB53oJ/a/9ftgdn+snO8bhDPyBN
es6xq1b/+WTUblzm63+13StqnoJt+pe6nvt12QtCO/LBBTp3DNLjz6AGzsH2trH8S06bghGBXflc
eCnBYeZF28keUR9MYHKQ3wQ8njweV/hNa4LopLM4zD9R05G+rJgp3ZS+ayXPRjLXZc0YHHNuHKMx
90f+7xxo1C3znKA8Cmt494XaGmsOrMY0eg/C4KHQcsnJig1ubvJ+z2cRqbZbuXTnQntAdCyvYNzz
J6OOHkThSuoqGo19tPW6CVbSshXoPJEUJEwVu5ZGTD1WcPnRnaQbv8M18l82K+EjFcgvA8M4pJ4q
n5A5PnV8gKAKJo26tG/KJfh1CrH8onaBuqTwTbdN87jdh1oRhXJtFCFevOzh+UIxvwo1Bh7GOdRU
qtsOv2IkvcH6z/nbWJ6oVH6cd0Bv+Sg60qmGOoR7LE81RrbcXVLJEh/AHTUPUWZojcbcxTS5uhwg
v4AeAPg2Ua1r81RmvK/iVdODrD8lDJd/jRY6eS+x2dwTqT84uab2FqHeXAdfZTg2LGSkNBUZ0R2f
c3EKKtlYeIRKQXuc/W5Llfd1N5qwNpWSJkGaAlymsmghh01DFJlW4jqoDm9r01yuJSqUy5XrdMQ4
MbQVbXQAKsUFCwGu+NW+wrtWX5EWEHPmvCxEevGtKScbY43hGxJowTSXwcCmU9tj2d3Al29fMGp1
te6dq7a99xjiHMqiFPDepPzMLFw6Wx1hxa2ANZn3S+wEpgMuhHd6li17fy2lCOdPkZYIJJVJw3us
GviET73LFxlyJkjHCr8nq6QvWBe47h3qLV86vTOPYQ2Jri32qUzoykgoF98nVIWzvDjpEr2SqrRR
REcSjVlQGwDopYF/S8lvQUCxQGGrZxlxPdzrhN+JIXcN7FkzXO7aPVhe9pvhKUxNbHtyKqutnenG
AnKPgi3vLPUtGdJ6xMF9kgAndNE1WMzSoJAMRfj5JSV4xOFvTKMQtrdPRMAm5fdBM9cTX9HxRZOb
3yyNbvpkC9uynD1X7giEah74f/vG+EYdfU8HGYC6n/1z5AdZnmK/eyhCCFtasUMCP5Mk8V/2mclD
vIxYhQIP15mngOAHnFEG1OnXZmsFvyxMPUYPAF4d7HZu1XXZAXhuQY9KtFOj61mbxJiDmn4+wHPN
SmI/03oCNWHwWM8byzoMADPXJDdBDgwapvo2e1JYlSStmn7jz77PKn/mnwQ03G/bPDRnmnXNlK42
/LqvvgtUAZQaUtRC4ZM8F5BLMgZOhLmQObZ5tvjdtUNhLRzdBy5hkaXNqab3DeQ7f1XyrsDf17km
Ei91a/pwMlZgksBJ36SExof4KIeqC4CjDnXwi0We9ppzMWD4e14T4dcZSAUIjYuvA0LIcH9iUD2I
A07lBjiNv6i0zHgpFJW6abGkfuNNv9/7fkoaYz4TlZw72GCIlHEqT+R8bASwsDouSRWV6Oknb/Uo
NPemhal8IMYGc2kcf9G6bpccz3VX4+bdbWI59UI8q1Sy2YAZ2mrUhFp6qj7m+dF4RODBfWcIxdQ+
kNYK0Eioix+RliEph97gJ0gIaH13pW/kPQs5gzQmw4efh5Sc6XWCY5n+ihbHNU+OtkKL3bPoAL1G
ImhnjDcevGipwBFBPR0nXIUCbNJDEycIbldTNXwELesRjtQTNMyjCGd+k71iNiaT3YYTVoyRoZN9
8xXjH63ok3tIfOrq8s8cC9ZY5NVaZMMqe0DRBhyLqUTP4z385RLfyei02ZAQzhGCinePsKLzAOfG
7nSRGYNENJ3myFG5M0EmabFNpVBZPOhVpX3wFMl+KDJvJhLknmdZeahZYWsBtt/zH404FDO+RIv5
Og3kZuKdDY1Y7kUDGhow1axjNvqQ6Vla4f3t3WKkndOdCxdK3yG/WIW81W4SFLY3iSfAhmkY1HX5
U+uA4GqAlt4L4QAHdd2T7PCIXKGseSCBehkuIPSC0SdC1GhM64aS12mS+Q/R7+4pLJxZinKJ/np2
lvA0LfUqJ4m8nt/xbLGBOJ/w0kRC0/xbLTexAkg6amGWB4Bk3SW/5EnEj1NAxHC4h1YqZe4CkdoJ
mH48z6nxVrW9FGQ2ATA5l3cU2jl/OtuwICH90Ng3f/gPlhs94LqIUn7p5a80neMUEr8DH118qKId
W5rk3aRSK/bvG7OyYJxTZXNnXvL+Y4Rod3Sy7zs4G/hKzBYjsgzyGghf5tHnNXD25WXOZ8g6UjJ+
5fszBJVwKzFqeqb4n6AFMqGZUudnLtwgGBkD4ANlW0SVBNh4Zs84+dxX5iSTJzaNiEZmFWDQix3v
hX+RSh5L16ecGNnNEHmMjWNbQlWw1VsJx5iGPkoXKm9nClZ+lBvcxmiPWH24Bx3Dg8jqA2jzgazu
tDRcLVR40v3+V89g1rv1OzWU23bf2279CDLR5moErNHeVFIq2k2ioqOTp6VBTTBVP1/v+fOUEqYM
FGSOpcWXpYbjkYyaQFOdCpkl5vEu7u6bAoM8YWtaw0olxR4vbpXceaQKSU+8dWEqKNHvTsmmlfYO
g/I7/pMUZRSgAHTiAeMUsSziVeCbn56sqoEAn1izsgfWJWa2vl8z6Lbay/CROro+XCK4dlLpHHgU
UD2Fiyfc+KT3uscn5JsM21Zd5ES0kh2gT9fhNKDSQJfk2bqLZw4MJu17szAl/O1R/BFrMQaDpMxQ
f7G24VfLFb+ln/gEzquv90gCfMBwfBQh8Ti/S1JoPxkuvP5Znq8xKUtkK1gq1JGqD5vQQ9LHWm/6
FqjF0FLFGPqTOSur/AwtY/OR3wIgoCNwRJUaguS/DzujMNAC1AhlV12O8aFS0lVnRo4eOXeblwWE
maDW0j/Y8adXNAAVzAWbpXMBVDAr/ydZpYiEAUYch+PS6phzeATzlDeKY8JTYVmbafcojDc4KZin
zVjOvyl5D/99UuzRsmdyULQM4hJj8UanFMSgubBAYYdIedidLhOt8TsYEEsMl9vZCyf7Kp9BoKe0
T8oITlzPpu0SxQhzXLopl4nbCuUM3GtQXG5Rw/aIOYaZHqew3X7NfIndIsxiCvOC6XKu3/yA8hck
so5MC4O/2zSG2u2aKuJvBq2L9bqt6XDUD3YiIJu8oDXd0V221t8OkQyi++8RabB5CZCAdzG+HNdo
t4+lOXwJrKKMDpTIoIWZTog63dhsr8xR6QMiIZi/2/FJSboeeBev1S9Qlc94hycNnuy0BfVf0OWg
phIgtuRdJbU+1GYhNYg9uEIsKq5JcTonexPHiED1dbZZV0VdKSKGVutRuwvAIrCLsbD8hptnbgiL
Xi6PAQ/GfxLD3WoR21R+lBYnB50fWEMw+8D9kZu6sVKc6bR22bQ41F78giMFGf+037FlbPGcKlWT
KzfqWedlDlwSRoCfaVgeHTzv78CQ4EbrTmfoRqM7pIq7u0aoAwIvlPNkaRPXa9Veg05Fbb9eIgfd
t7Kd+hJfSlm0X5pI0ZY9CJzbV7dOhB6T4VYuO4L2auJKkCFtTmpHwtEwosCubZ16T3bgaHgJiQkt
Y/db5EOigtD5xzYt1JtObamGfjHUKiiWhWMba420rua1RhY0BLCgAaIwFIjVAFRQBhgOni1uTsh9
20VecBJVviJhH+Mm18MwH/N0I0gv9oaKaa6BrUBi5g/en8dCWK+ryvQIQ3E/MxXV9KdLiuk/7vi2
0pDiKD7HF7q19bxrRkjoBwKJ/0WuBTf61mdf+8S0zmXCFSMKrdpqXnKygltG3ygM4peokjZbVn8K
3tH1wq4JEbL7QAQm/lGdyRT6r87ayrwIEm38C/jGuugdnUoEGjOLGRSJlox2yGAcpGaTdJXUhofn
voDR3oLpAtcZEO3LuAjWNqfiXlt6T6Uwfo7WOgR+M6tEVyfIY9zQnvJqC/E6cJCp9ccmTbrPENGw
78T6N5Nhg2dZ6M1WLjrcG7adObERBQKkb740du61IaAO/uzy5Wb8sIYFUATJMTJJaYXGa3vUsZVQ
Io3oe5bVRkegB0J6grbGBY0ZAljBUIL/82kICb7X3omYL5Jgxw1RNMrrAbac/0Sl9uHBKP0P9udo
poyBJin/FZv1NIuwfYSCWhiKiPLaGO4KzqDvcePCVoXxJMnD554rLWJdWmqKOmavCpmKWWrbEjLZ
wH3z6+WWZfSeROnUxGcUSLCfn5Rp6arG14Mo7cXOkNzuV34ACX6ZabNALNJl+WKXtvlEnDpFgGBQ
EkPEwmb3W72NnlO20MvWs58PHlaHEV2Ak6hhoYPmMJuaF4b+nw2wtu5ghjhhu+ifRtrr/ELmsMLQ
dZPrgOCFPFcomwPunnkRNHBjOjRFMGEcKlDCB5H1HqDZhotmUVyb57TPv9AXEmoD9LGfYIVc2x9i
7cEraICDX0tcB2Ucu+pxKqRNNoHK12KElqo+eAc/g1y6Flt1j4vf2ZtJRT9PFLfonDLW2kqHW84u
7HMj9kN/SZUeSTNtd2/xEw32hbtKKd+0sei+5CPYQTLaTnMdZX13I/jZiIwATwma00AdRLhOvQSV
/RvLcVMrwTDUNsQLeaXT01NxnJTx2noE5zuFOVl84E8SLqyvsx/Mbo0pVVC5fAEhi97oErbWiFNY
RocZV2f0NstcVUCWZXmjoI4PIg50zParAIGlHwToCPCq3vAib8DWsX5nmLFHMgxX9kpoWRdgvQ6e
CtVsskbwg3liUDUMn2Njt6SK1TXbIKRzdE9FEZj6ZUxAZv7/HPCXLMyqm3usYdbIMC6yRvJMrwB5
obmO/Ul+o+kAj0eCJ3uOa0zuW66sC10+QjptHiY3FLpQA6QmwTLCy79CF9lCd5KeCy85pRqw0uk3
UtllOz5vknTKjeAsXI5KW38+vjJgU6/CcLZipkm1B1TltfpDoSUF0GBn9fiB7NTp4BKh2KlbHR94
YPWOkPQbH+snC2C84U5mZzzJhwGGXNPwdYJ9VNTjhcgXb4Zyj47RxPqZcCh8hAQMnZ5LoXuz9k2e
y8RlZdNdyxCNHtq9GGo07YaERNKIOvjw+BW89RIcTRFanKqdApJfwRZhFYX/aSek3sri1zXA5kBQ
Hi6AzN7TiFzhkE1nolBHOBaZZyriUKLMBEbpvExD8Jkx2IyzHuVOP4DxIAUYAZYkE/qRQ6F4KWfM
Z9V3RugLeNuusK0Mo2/hH/pla+5sh3psSaffiF89AJQ4F9mXTZ4YmpFfPhcVWA/tTZ7gOkbEbg+a
mUhJh1VK3hkj2TkYJoopX9uUCfqghe3bFZTQFM77w0V/V2yK+9jDy5eMOX5eWPgDnBu31WD0/5Wm
4CMeyH1qESrpTucu356UQhqQ/jKq1QTER3PObCdMffTrif/7TDxwbJu5mYYkPOMi8kWrhzkgMplR
F58qBkvw32QLPGqmqTdc329e4PRwandAK8PKPomj8W7UpUTDAAsj0u1IyeqKwCTObixltb0/aj06
vSLlK5Pm1OAZ6lSK7GVqA+1i3hmxPjAYA4qtOO6f7/aZf3CSm1Y1xTz26/19AbF6hxO4zVm35Zc6
XPFwnHy/ikjhxLSuBpElSeJmh/C/ZPTMVdHy9MVQdSae7xtgvdMOTH8+Vw7tRJsz6+2kSfGkQ8VJ
EW1N5Uhyxduqh4DvDvVpZkQIzK6fwADl7Lt/oo1MoPCYVJCmCbI5olEJrYW0AQf1wVZJ9ONu8d+j
96AGao+mC+rPB68mijAoDLhIJbo67QcOsxH/st6qUUnAlGM74G+Bcupe5WMY+mkfhT3J0u/zVKcl
9+Yml4DYeKsa1MhgyA8fmscJt3ejZ7GnRxm0AKLuLGLRGRqXIXQi18eX3XHZrqEpf2VvleX7Y8nx
lCuD4evcrahu6lO0iX/3W+83p5FOkajWJk9LyCHDHbM+I4JJr9p+5VLsqY4jc2oENsWmO/ZY22aC
LeVk+uR5MyzwJ1Dhx1hYY0X43iHTaC6zOMo4LlNm/r0B08GZhm0wLgGT/UHKz4eFHlk8w4GksKyx
E8QPli5tzuE5Rd+Q8xI4jLRFoXLixKsACNnsC6gVDfVO5t1omj0B56eYkHmigvG48tumlrcEmbSv
Q59CvUnXGXFWogaqDesVtLsbRdES3VvdWf2vKGJaX70ASsY/mbCbXXXJ+2fgj/aCW7FmRFwpdykE
9tRzr3udWpNhtf3w/Xgq170jo97HupYOVNF+w0hdlU28EadfO9C0AvHPsm0S4g3EHNVWCICDB2ZD
tYRgg6oGaQjki/pwNl3xe4yKa/fU7eHXwH6P0VNfojv2jS+5lJzXMX/4jLOxkLPtMP4lQvebFZVD
eh5Hyd4Xb5QjoPxomRmFNzMu5JEEuMbOhCpbPZJD3wW8PIwcb6FiEMS92sXSWMPl8P0kxPDHN5c+
FRVd7p4hMKtRV90HNm6yR3BzWGc6Ktsv0TkazoLURP001H8A0crke+lT+p8gExCFZC7ySvhcU863
WiMeK3nYokQ+ZwZYxBzbT5TggMCCKUSXsc3e2HIdy7pLxTAdYDggTWuEfkRu/fPd3ttcYgPSOPDl
D24C8Xa0xM/OetLkE61HNP874nuYzOAvOUf4X2pWAmxu+PvhfvbSsAdZbGVhrLH39xerwLun6gy/
Qac18grp3kkAc+PNH1sH5+g5BDhaNIlh0RhQhReZVq8wE9BxIejiHUXvE1kqOJetJ3tabbqjX46+
e3shjyOR9KQ4/jYb7f3whjum0iKx3we3nZETKqyyUZ5SAc6Je984LKVkvPduVb35IzJdiEeI7wRd
zZsc/oSyu13jAsgcXmQawHlTKwesVQZ9wSgfGx497/T1/gRZG5uG9x1aXRXvnVPVMIAGy2GBU7Ae
0Q6PoM8NBXHmK9y8FH2ePnOmSCnzTZMxJvo4w7GvWQ3C02H7S7wSjRSShXSf/ZmjLxXOqo7TjEbe
2WoR3yQaa4Ql9AEMhdRXYOjtlxjcunr++Vdx+Y05hVmdYlg6lDqexW54UEJ6YL/RP4RlkE/HVYYl
FYL9eymqmxvFXO/JW6NU/9i6fU96pkouBLzQpJe3Gl+80n+P8PipIWjUvkMqIDxWorL30ZFuLE9S
R4BlwwtXjZSx8Je+98t10EP+ncNiTkn7CDCzzKvl8Il/EtVK2g5nRp0ET/L50OlVMq94O7kb0uXZ
pkB5SHTYpXexn0LqTl8cJdBGdp1+y82qfqNMCntnPFwEB5GZwilWB+SX5Q6rLhWPiqwVAyTW8eqW
h4JbxP/ENTtGIa/HnkSIuZqQ7aLNyLbgghoKmLuiNMbDSdZkB0+apeduTbQrtZNriDzFL/LZACwS
BEOhqWfidmFQW3gzCa8a4fv8C701oNHpsk/tVLfQC+AwdJ2dx7FTYAw/Q1/goLB5xiZvXnatqvp5
j4cBIFX7QXd8xPBizRyH2bFwFKuAebBkJRmaCEgWA9KPatPM1XxEqSL1s8+zoTPFU1+pMp0vsl+6
f8x6XZ7ivufiGD9LH9UOj4pgIerva1o0K8cFlNsAkqdk5MluJvHVqsN0BaTboP0W/rbstB7nI6H1
Nh9yq6LZ6ee1BQl2bOBx2Jwz6KoUIkm4O++YYzA9fMDUK1ekIWKF94x/qZQLQHpRV7nXXyPd/Xu4
l79toJ1mXbHfFF81oIlsOSMIO4q2dGJFXnnrN6iLkwcerDH5jr9fwg3VfDqX8Vb/UxviCYewXHkl
qXxORTds9WtuLCBNvS4nK1tzncSZGeBz4gJ+WvFpulgTq+l8FLngmAWlkw6zGsqEmw9f/npx0Zmu
dv7TEwYVp4su2CRuDe1P/ryS6q0Z7evM7g6Jgi5IvSMA2kfc9fyu26uMxu3hn2wlW9OHP7TfouJV
CD+gbZTdTZD/Xm6+k7ep7QylOSGuZpdOPVdyyL57zG2C0cpjrmdA/Awl+zyJI+qhemoFLHmNzUT+
setIevrd+67xldof2svdj2P3hwYt23FBCTeYVFfDFP3KnaatUxDQBZ8qW9LiZ8KyJF7KK7Qow9NH
yTBAJJvsOMsBj3FXFOzsNE8F3ErR/K2nqIiU3wSpq37Y4Eh2z+UhGBXnwhhx7JS/Op70rOSya0U8
FT67bsQiux8XO0e85MyZqMuFTYNudqDplZ7AOTHGo6dB7B4GBi7wk6uFhLCH6BPjhrs4KJTv56q+
MAmTm8C7uPTUUhStMgYnJRUCKnx4yoeBk6jmQTEsvVbsvNbBlRYuMkoOyPgT9Q5j/+3kq4z1bL4H
w6+mnVcjM463Y6hr7nPcwIi96An68xNixDPjLX/Zf1abMkm/iKajnYu7BKhBZW3OpgdTq/nOXsdU
lf6dwdBqDVZxlmQm7gQp6SjF/Lu22mkUvJTz7EkbuWEXqtRphB48E45DzVkUKzXeYRpHcGOaQCoB
lnwN1A5ktoWlRuQcjjAsAWgtOha/tqWAghaF8zxqsU9ZzVQQC384o6j4ZvZVGX0As9yvFZfCx6YD
VTh75rH0j+4ZPVPzVV5XaqZRyX1V/Uj5psg/TCh9dTdtBcTdT0fkoCmdE3nrjwjHVvTEjBp0bI3m
b9RERrJlOBJP+BFyQxb2bM2QKdIbsjlNaR3ziHjFy4ZjA4seKsi6TiTVhVNj7tM4FldsF2utNeLW
4s1RM1FDBAQm3BGwEcqbyTp9R+t6qapqTO4dv0GnnZnPKjTprFxwFApxxCPnCFuJ26DJRNH4PaBi
72V8eSCvdTNyMHFLJnrV4O6RTiYyRzGxvoNqlvpZxxVD921PqZcThso0+UwZJK9wzsRaJoTCwQKe
fSWt7qX3ov7kaHfe8oTrLIMPVlIClYY2tIS/AV1ETMs5EmY0lW+wfxjE4WUmC6IX6SZ8249kwLqY
MxGYXUTXlqoqDc7KFz6wjZZysh8EEjhk9xuXL13O8mOvV6wLybCjDFMPv6MjY/gQ6pmgCt7j2xdW
sG8IR+sPvwPsCggWJaAe6s3irr8C/n1oS/wXy9FhoDGU330AtraF1t5g/G4DTyN8kNBU+VMzoHgX
3XWDN+66oq5DA0ewW2xLP2lqlMZaWxVA8ZqoHDOaQCog0+uhHXIgHyMEwowxhEzuKEYgtUTfXdbX
W6G+a82YTqN0oiLk+IfYnMPhujxBA56lC9r9afkarKT0zCCRAaL9EwkuYy1SkKQQGB8wbYBaukI7
vg9fJE/0pvagIYr4PV/RIvxTWPrLCDV2OzJYHf5vUJc4rxDMVGS6wIGcmwgOK2r5PkI6a9zcSZIT
v1Kyx9W8Wby/CsM1Dd29klf4vUkVcMmm+60xF/y/DCNPU3D5k1bDPPQABgquECPzK6nVDBBXMxul
Te9qOPFMIA9ZjzSV2HG+1T2vwCl+1r9Em2lzGexq/F90UZgIhxaOr+npfU7ieHEDlzfO6jT5iylc
jZWh32s2SZiUqedBsxiLSfbNboaif4PCtGH3YGFhn5473MfplW5iDuyJPBbp1A2TIUtU76rbs/NK
zuAKaLW2O/t6oxdgarnNgk5MiZvcPDrzJ4BIJV+nfhOgGTE7FXFNkAWAxi74Cj+AQsufZn9C2fg3
DJ6c5HjIdX4N94ykWaev9Gp2GqWl8XtXtd+NFcW9DX0Bsfwtr60bk1lpZyN3nukrAAsBQzq+PbyF
QGA44P+c3atBN1WxUk4AX5AlRmFukt1wqSKUw8YJfvhy/QTKG6TEXebELHSPjrcKPXVTBnMovvn/
pQ5JU0/CaQNGuL1IYvyWpJyORq4L/du+NiyIcSK5QrrRjgHrQIqF/mGaLFgwLbAZWo2UkVEISFkJ
P8c5Vl6InYLADwF5agxHpDsxm5I4GhwaPyVd7+9J5hVYBB5jTCpStqjzVCL6u9Js5moprEph6WUy
tsAiYEO1WbV1R97ukFBWi02dPOsAyTMWLYIjNoWbhrHWGDwmYr5DXyytcJckpl2MIIqo7ip+ejX1
6KiWpmRr+YHd516pCVXTHOndqhBl7cNVaOPtudyhmc9lOieyTSOYoVaZ0igX/pW7QE6Q5KjtQhaf
mN9ZH4onGxPKSDhFg7jMF2sTZBtmALwo0JinkGPBZMVmEANPDv6QcCsuYn4fL6JOeiXAUgmqRGS4
EiOYcpjMtm7FF+2TF4bDUcXknjGk+7E05ORAU6RgLK0UBEMWd5XD1j1phT8yNMEUwOFAQxUpgGZs
Ufr8bU7/IzyE5K1i5+z1o3AuhEGgaaa/vF1EpIZZWzM9EckOFShCinH3n0r7rheX/PGATBhRauff
Fy8iK6yqfdrKshcbJjP9SWTc4rb/GIR6A6rfAPAp/8dWoQlD81fuIiYR/iljZKgHfXBj2Yz2/DZm
t4r4xs5l+hmehyTsRWGJ9QyKeNmTJnS15IUzzK9+MfX3JxBzQ/tM9Hu+baPVCMmxqAITi1MpoW02
fvYzxQ+QFST8e01AT0fTmdBSNB5jDEmVvKT1XXDkY/H8BnR4eITRh2ITfvxkLZaMLfY75g4IeN7t
SN9E0RtOukr+yYeURIN92lsxkc7qnY5A0ILz3BxNV0qyHPQfHdUF7+OJOhJ61IkJkTbdBU+n52fg
/FbHQZUUs/KXSe5ZMgbfQyWlX50PJtYLG4sIv6Jx+ht1bwiu4BUcOnUjPwbo73jd4mc+6kvYnFr6
YD3e3RoWwHF+axWoP1Szmo6AGGVhApjPSIvSVO2kMhS7+GOFeZea4oTysR57Z8W8j8s3ohz35Mas
TtMxZu/10Ss5VCJ7iIgC3MlboieTPnSaKtg26jjUh6rsDjAb9aR7BabioThBUTWT2+HhvRJjmdw9
mzjqQJoe3KrdPdkx9FOASV7s5WSFS65lzpSyC2LutU6o6t/qI4tBDKMryFIv4PGS2nG8CaJx4S02
tPr9wCZI/25uZY7NvHsk/CsjcSGs4BPjV7gBqQNv3rol1XrTS/wHRI89d0RGs8mg2Vr4UgmOQCKW
cOIxf4XV0ZpD7BGH+V+J53usGmq/StuZYeoc7fYCGCP/G6wyuZx3MSzdvlurUNWRLmKJ3fr3JPcv
9YaaDsbBH1vBbHn267UHxxpDi1oGYNesNbdxhwDxUZnlhxZtgt94iQOXRfXmNRNQYWSUFl/LcTU5
nKSqyt1pR4pwPNprqv8Jk0FzndJPM8vlYnbHEAFQNxnHqlr6RAXwbx7y1AE2QN45YH/dnVxAu0qk
sFCetvrB6cAIDQJdk/PZ0BPSMxMsK/kzJpuhbPtqZILzCaK7ulyeDXf4rNPfE/ag7rwniKjWdYBl
giMULFbFm4sVUccuPDE/6Er1E4vhbud0HKHbz7VgQnn10cFE1ajbGKjGauE/6wysLInUI1IgsPFj
71HiaPugdcZXNDJMY2TVk3gFdBHoctZR/6IhOujvd0kba5R8owCEF7D/jGB2606XgaXgNks2AilY
KUYD6s/BRbNfeaUBmbWhmORBA34wQPvMkzekFTgXnusR2V8Ris+5/xbCqUgGDLruZPA5RuAZ1Thu
BSBV9k6EKiQnEhUeJ4FcF5PvUS6f6PwS+YxMoZrlRKnDCheotEXptKgGQw02szZ0oh+MtCt2A7HU
+DAz2w0pYlos32gCX4Q75P53A9qd4+gs7QIq5XfRA4+sHLNu1a55j3OfHRouYCkn4UA5fdDDBjeq
53BsIGmCy4lE8EPYYiLVFqyCx7j/l2WLIDkc48Lf45Av/761FAcsK4hHQxaAvbC0IGv7x4PUNVUR
Cnz3TJPfsyUaL9kYiPpo/AEX9Ar6K8Dr3y4Om7Sad3Vi1GqzE+c0rEYnZqDJMofj5JUJ3iwspS/j
C0gcWFu3gxR7J+RHtnRUf8xdLdn1pgoA85Wd1Qpv/ATqQu6DsfvCdqBEuOZVTsNm9J6IEgzF0/Ci
tjwOgAvvo5IqqdTcE0Fl8kfQqqWJvlOycnFqm8q3PitrIFzm6pT54VPHVs3N4dide/TYFVz1aHjW
fQsdtYIWD7R8vyiZkVxxR8a95s2uKnb1KMF7I+36JGXn1QmI6bY+wjr3IGQ6QxwEG4iTEAi8dcB+
nyP9HzFm5pvkePOEfPMVYB76dsOKlM/ATMmIMuC/sPtDE+n6Aqv93bt6Q/Iz+Yj9rf0dluh5ZUdR
7M2nP3/WpY1oDviInnEucQYH7clDSl7h4PCn02IWx2FIgfMlSuNIwxcQxIDeE2/RWAJHHIF59HhJ
MPGQXFCCTiQDO1VNtsDz8519wGvmh7PYHhRoqWKAYRbT0rQ6uOG1CEy26XJ9tL17kKjssP2YUaYf
8qIrzC9l9cf0Tn88RfM/JsRI7U/HjtX4+RRGa3lHtpDMzVFcrEnYIP4OzGrSiDhsxYEOOWc51mvO
Li0D74UMnbpOpRSH7rljaS2Vp/fE3u4g3Blb3GMwBqutBblGRXfqJiGGTr5HURKV2Jnugip9o2aj
ZDR/8tnmxSudmt7c5w8YKIjhWYFPmx364vs63ANF1GMM465b6dcBmwme3Oer+nHiOxrKltGiRg/j
l9GsMPqKZ5osHznR9VlAz8AgsB01HQCfDC6vAkZrE4WT2VvHUJu3lWmOtZ0EPD3Bdxi3dF36vfN7
B71H4XDw5yqAhmFG0RyNvZkrmLgqJbzhUQeBx/X8axvTy8GSAMXGHOBbM6kSnKQZBTrPZ0fRxh/5
sFN1f9OxzN5L65tSVu7ShBNNW9NvWR16tjReog3d3629Q/795BDfj4ecyUzidu0DKyYXR8zUhfls
dVJUjbVKd6YpkkSL0bYVM0jWB9uyZTD/0MlnGt5eJoYQvh0hX4rOaA4VBCx2yOPnbAJCuRCUzII9
PGE2Jej4no8zd3JtbZf3POo4RNMMrraFpbAJ1EG+xVrt3N70vqHGKJzC+eBew2axQzNlWzqKkQTb
aVI5BFDk6NE9HpqG5+35eoJQKQpZBSriBicg7sKSjb3ep75488WYThm33jN4NJYa44+EZR0mOyFS
60qes7hSzo9bOvXymajs/D8BZU8EfNaC2tl3hDRHxNPK5VHgHHbOlIfSgKQWupAE/vgXlAjehmWY
1sP3fV5CplwqICSvbKikvmlO+vpJPSXsgdmbXZFXE9mvNhMi2ECPdGlaVwlZsWkL4VVaTeK0JmQD
J+VxRRSMMY4ngyoFiPLA1u36pM1k02GUa7rftZE6BpJtJwmb5KN2FmxTg/pFLTA0Z56lfqWyWG+v
gk5JrGcsQLhLqcwP319ylhSKOly2vApeRQLNeG+DLjxXvi6lAVprB4R6P3IDUzhgo0hwVPxqtMh1
n1vZB2utxUMbywupiYP4B1jA70oiR73N57xvx5TIkxastu37tPioTtJ75hFITNtV+hjAmF0StppF
9tJ/GKbCeGSJgxOPGnhxv3h43SWN1Gazqwz6r1bY93iw1XII5nwT//oUxpIiLNqXu1owjULpmJxM
9gbJmt0iL2L73pQ4cSIM6GZU5rlMoVwfJswhOaDlZ59vuhy6N/zHK+7LVU7vkXmdm07QV5mvzJSD
VF5h35+lg6IWaqf8I+S9OlUcyngCqiOyw7XI4uFfAgSJ/PafpI1Pmh82eyglX3hNQINNVgDYkN/Z
7y0mJY91GfN5x2Gq2+e4ZIwvVAVE/qJORjcTHhoczp5Lb6UTSkzDIHG8YTJA86UkGaa0LKlZZQXe
WiytVlKpGlnnbp6KLyD6Pl3QkAnD39r7CqwTXS5E0xo25pUTLyeSKmX0W3gozNgW+d3megzdnCuo
/UIw5RQNmHBnuvcapugSE8XqbdLJnSAGlvfW/CxUXtA7AJXowb79Xz1k7nPSOaqCIEoBNv7W6jZh
HtsrwD17keHqKBrS3MZdJ9d9BQxuAtjBBb6CmhC3Cwv5LCL+xK3mXcqLCGAECoI1A86oJSHxVO7U
FS3eb10xGaHpB3KxgsDGGLG+DIPJwUQl78as8SA5ntFHndWcZYkpd/AdMTBfmkxgMW6w/cvkfQMi
N3xllWsl6Eqzti6qn8P6SPoUwcLHswI+j3qznBwULy1Li9SXI2gXyLnoGji97b5WHMkFjTEDB+rP
NLKuF4ei0qAOM/QzTMRTNZfhZBujyvhpRSU9qLISDTgtO64i04KlI3d2ePvrpme3jlonI87Toc+I
Mv8X2SKAKoMUz6wf+krL2xOP7LHH5WDQ8QaJHsrjXjqNSyY3819VpFkH3Shaxc/GSCvS71kLijZp
zEMsNHfvgmr9c5Zsjys7WlZfDoW7Pcf7rKFgfug+XvP1EkKjHRrFwW4QdPjTrvs6jrtvYuzTm5ZM
NBoZEJjU1zcF3gifUUwNqiHdsNUxmjyVe3E7atoZK5911ph7ZNflh5w7BJHKTro09VD7PrR9a4qi
IghNoUqXySoWcDZ2zaNssj6VqNLS01BYHBdSqP0p31prW7PwcCVrV0A47aE3uHqTd1ZlVZPeN76B
/v9BS8VGtx3fNAdiuyuBRJuP83UxWXaRy5SbC+jFnoimi1E7/QzKgK2V2RU017dkDOl+Lw0MjYp+
YaAdCmY1G+jijIGxqTgRMKJ2FqoeI6bXmkFGjOdePkX+NYt9Ze1eLKh8xZ6R79J0zV+B4GbHpLvm
TEdf842eDAeYrV2P41g2FFQpE7trQlqFsv/Pxe1cH7y0SUYUfcv0Lopcn7g2MmfJp5Yw3ZMqZfMu
XdrCBqsS28zLO9vLcyPDGi/HlMl/EPs/IPOmOeTgdn/dRvhNR+74PiZovR/mTwh6B9f7EMj0h8n8
ALSuhICx1wv/v5bZrSad9RPiK3lNEzZN5cPwD7xYBUfBvcZIGJvba/+8MInrFmV+RU/expwLhOdA
HC57Q7FqYo1VmywEsMT0ErYrqTl3hO0zDA8ZxwZ9MZ98Sum6d/RfFe5MEoXeUW4X72Mwyu6ddKLZ
hkwjBa4wAIeMLfpXCGLA9uoxd+3KplullJgc76rY7UJZwnAMIo5zaey7OMX4+iDbug3Lm0J/vo9M
uPhVjWcHdNwVJMGVHeXZAtAKRnXviSWqcxuKIcS07aDXxmhQdqztu+siQrr3KbYU4nkrJB/y/4Yt
h9xlmsp0aiyN1MTt8citsg7G5juckJJ//IyPDK0l7UwdRILBbZVHY391gb+SGpxjdpQa/19mgUwU
PfpSZbrVCcMJbNQYZGZI4bASm5glctBDMDctbdG1Zl8j68GsQD3m5XbI9x8Csq85lzbx7z16p2XX
SwU+fJ/aexMFjQXkbuDYHALImtGC4l6BcZ7NbGlDWvNrlyzrh1g0me4Fcg/1lkvSGmgsEzobrjHt
djCJoIatSNOB534QXhRtf6tQDYwSbQeAqmg3RszcrVA86jepjxLFlmUEA6Z6kaeC2zXAd4xgE95k
m11yN9au4doDPd7quaaNFyQIegX/LBzGtZpkRNDvi5WrhNZztyWEbo2W0MJxZr8N8Nu+5SjvUX3X
u/wrB61zfkstX9TLkO2LnvHAFpi+LxB3QBhjjMuWj4M98mB/wacj3RDNVLA+GEHSTmXauFlEcB0o
K+YPVXZMemL86bpYM7cz9VCDsa6/RDGCn3StNwE8XJKMAOH0845adsfXwVmOiFY6+ltrKcuw9oG4
q4iZQiWknD+nI+K+kJ2CHObq9CNrkpnU6V1fF3DFJi7Xp9JXhEpjkCbLqXpA9jR9X5gHjsQ9pyOb
n6yPFxdel1qnBGL5ChlRxht3su1KUM2NtkSV3mWyF46HnlRmYcayMwZBDML8R6gYAEZGSf/N1ab0
UGUpZhowH1SfQnCy60xIy40GrEY7t11ZELjsPQM0ECvRLG6oDx4BsffI8+uBJCWWNXTbaJzbTb9S
SLpKBAt1MPco0yHrP8Mr8cSSG9NataEO4QmSdeDQ9KXfmcIPyxQjxegpY35/wEyr7ymNvUNhQkp/
loK+skmvgx1HPbvuQEMj6/3J3xOCKfU9cFNGKzSRyvC0zaof8vTKCsQbWlTOoDlc/76+pxqAc3Rg
hW4/KZQ8D7OM+m07KCxFymUlntHmBR8Kw2khAaGGe8uUXDbE9o15EppEoVh3rsTDUp0JZkfEHIYl
VamCjs0/uaEzggVzuS4xDRTOsLCyjEjm+i71/gPMA2iXcidDbghDQuduPkV07r3hGlOl4zTsgCdr
r78JrmOyh2EHGD6TcTdXI7z1WQaScfjS7hfnBLDlN2BmRHAiYpetwFUqPAQqKaTjvzZk+BY9Y/2T
rw7kKthChtqhwyBFv5p/Iyd1KMexCFb1CgS3k9W+ZLYUkFK2J9cG5tv4vCg/+HYBA5bBdx8jMcT+
qEWiCMlUJoQw4SuJ6zJUCYrYJzg8hOBt5VsOv3Z77UU0DflpNLPUC80qjBDYBL5t5gbwjZYW91X3
9ueZ8y4L50BUS6k4GSvL9ayV3G8OahEafS5GQnamqA2wz8aKmpou7479T5A4PnGdkyNOyRpmVTHQ
mI4Kn+Lag08fzdD3Vyq8zYQWccOGpHZq2S/v0XG2451LSFPKERIwJct6MG7peQEzdUN/iq3QJTWK
otenUeTDFO7ViqOpDy4wNPj3sryObVqRk2m+9vqPmCpQaABqBVFfyh4HSbQSgUcQ5jD9RcFkT5qN
H2VePm2+aH/cki4+K+9BASC1CdBLxFvXTt5bpfHMBUVE1GI8pfWFuaHShkdsc3eRF7loMwaX5m8+
/Ng+SfNVOiKbxOpQeiNk43W00JVPddve2+vMariVDgZPHigUNyolNJaOWw2/3f+h8HW3dGyTbHve
XCMGv2tUbYxbPJjZn86/9dk9Fr3ebhxLg9RG9q9xXnDE8fd6yYeZitWv4J9hzGgLQK2x0ub7fPvF
2suSJsh9irf1x6HLJG6lNihdEaPgr0ruJ1CWM7IE93QTAp1yCOFslqbzehFuxXUgnUAgN0Dc+n9k
cC5N+r24pcasdahwiFDLlFoRswJtSHfZI0N0iO/rhjSru4ZbZn384xTRqcvVmzqrIdkNpFcF3wVZ
jzkRDV42cfqVSk/VGbWFknmtZYGe8D6Hqez0o44Hxu4PV0PUS4+0MZvCqP9UlXPvrlgGYlB30/Mi
Nirv0XUe20gygWqPCxQc8ZNmJ7ZdPfZsBW9wQx+4Pr/SpKytoEhn4U5lCbof37slql0GH5PHC111
jE4TgSQ59OlDFbQ0R1v208b4u6y7KRkBBJlyA88qIDDBFx5mDc3vt4RblB3fhbrqm08BkFYqojfX
oS6NO21ThOtMRh6ppmRf1UDTu7vc887m2PVIo9MwCfpkTZ+1j2f1d5zSPL6HdLe3B4IZ7I50P20/
pUVCMjDOQyrESZ3zia8yjXRkg41qTxtvkQBzFTknKt9wgAJj0HhTqi55rDwOccl3rwThKS5aHQe0
kruhAmYiiHGl9+G4Gdoiy36Qn9uiqQkevqHoep6L5MYEGeR2g7DBwJcAjm9JFzBr877YQB+0scdv
zEYjrpDneUJyI9cuoCO7cL3KdFE5LQAnp/wJ4UUKFPzmKMT1o1VfCLRDeoCDn/BPhjAceiRNMwhv
Elvfl/YUvCo5d/tC7CLTrvWribZTUVaD7X3sgtQfbKcVg1sYVXyEoEnuv9J23H21MHZ7VRgji7jl
wKAwR8tMZpBPiYGxUtWRRbABVcx01KHMlRw6PihyIj+nzv2rC1+ycZI/oNkZBPo0eyJhl0HMWruc
df58tyIIQpd0wS3iKyFxJjm7ACxYZX9c0WP34EvIFHXPdjyqIaN9JyU+0UGWVzr8rjddUfTeou7d
Mnt1YRYmSQD5ks1jXAeFs7LmqDFxtSXa7T5MFwRuuxHsd66Ubv5Int4g1JNhEA9uhf9rW2M8D3DS
mz20qpQjOITjuENEVchHlYBHPYkWAqGUKo8nr96HfuDOAL5KmyADYaxBDATUutfsV8f2I3vUJD2t
MTcU3VQbRzMloN6nmVzSLc2sWd7NfZ+u8p7t2cpMgxf5AvpUqOiUi6sxSe8yk8lyfkrwtIt/m0UK
ZuNcQ6owff+Qi58yzrIBeqAh1Lzqrm0lZ2KsKRpmfDHZpjQ4XUGJfJSQvXA26ekCZqMnfuSCsODO
vmMhCkBU80X0jl4DrLv6Irex/1PwO7vNc+Xx+ADCzKIXvxk5ulsBDuDB81mxYemU7izk8+Yu5uco
IbOlfU38LL2a3FdYjNsewrQKyJBMOIlQttMlnoEugddt5lKADX5JVhXam8liXPDhG7wEj+itQGc1
y6j3XlGYm7WEbrCbKkbE7Dfs/usn90Cj7s9u4vt4xEmO96Cb2UfaBqjfaoZ2DTX78lfGKE7BsnUN
bwqbRe1tj2lZ+878T/X8qvF1PVKOLP+VBZAi7fzpT0utookncsvpLKvUsQZKcWGujNse/RNAZFSr
nzxFQwXOBwX1Ek3qeRSGB2OSjA6VLYinsb/EH2KUfLIVo3UHeoOxK4L7VOMWzR6hXFSiPjOzBaXF
x04Uq68wmMt7ghpkWZKGfqQxjKjUNedMJEzS8xVfb97fvNuyOlj1up/zY7GI906ab3EN+6GtrzHG
plJnpelaczpOl68CBDVCKmwCAV3+t/DBdmPTLKC3hIhEqEfTGp6oNZ0drTM4XnGe1qh96oxJXJqQ
4DsRoaj9E7tsnnOW/zXePuzHVvy3A9RdDn6ewT7NJUkgbHuPkJFoHlHcnu+94CruqTwsVTyCslLy
9Jd/4x2oQf/l8+diUJdEoMpln4pnArKIM02czTmlMbDLLVvDQNfxnvP5KqaYpNof5AP23wjz8wwv
2AcIKrJk4sUVZwgrURHItbZORyNitcGeJIltdHhGCEREN7s1vULJ60hQgpiR5ncysVQ6i2VBgKUE
wzF/S5gBHyP9RmL7GKeEBxGZsc+lkuRz65P+Q1gn2iFP/7jhnUQakWWySAcjQyva0o/9/qunC6jb
OhX9SPFdX0sKswHo6QcVhpH/etUbSemVkuBkI7SmhQZDdhj1MEq0vI+2fRBfyV8WcOVTx46E78fy
cQHbtpHfCY9tNJEeKN2Y0M5jYhFJCusutsvur+ia2MWH1G338HOnz577YdsrYT13WzSf8V8/RlJv
W75RXkFPvg4XTHzsuyLqqJyhc33EJy0CQueLrmHWx9LJNxW7qzRpP+fLf2tNtow2cmsSI4kYWBdu
Zt+wjWLProwJZ2/5QzlxJmmwS5HXXaig0UoxI7FEV10VI9wUeHaEUyAq1AP68/tCVVP6rO1qXWH3
qneGMxQ/G3SUl55Kwv7huSxJg9N7ekytT6W+RJe0EZhTy7phpyODCnRXigG8GfT1YfJkUZdRLLfs
Yu57+FTMjY1+PLXUCN9Kqq3Q2VjWNka0P7V0K2aMAehu1JZZLr1LysD89Slt/eYlLFN87FQwzAsi
h7HcGv4bz17fJmJfj6zsd5ZfoHrw9UsXOc5T7gNGgX/k7ljFsBxMW4OlfxEYq441aJt1OD4XJ54B
m+WpoyQNxB54WM/55ATxc1VNqcQvpdV8TWXuwXyxTzXm02cpsvCI4xIO712lzVzzUcqC8tCuzTFB
0wDilLFUyaPp6UNdW35PB7txES5j2hS9hi+V+H6MkwQ3DrYBYe7yZBNf+F0kI/e7CQJMD9X+m/Be
O/FOmJggJe7eeQEkIs5s+/nbYvYBERqWOTi4F4x6/ROGAXV+54QCwM6FqgRUHfTZdhnESFnqMGx1
1VVJIEA5A3bBSYdPPu88f2Ge8uqIqk7dtCjHK6ur77ss2mO+CcEI+s1rqfOXWk82HU/UkJ0g4wZB
hY28o1xALB9mJdndk6kLJ8dEwMdfQz+OLTS8FSM2AXG5xunWtwNGOCe+tJA8su5Q/ygNEIYodbzx
rDFMU1jzeNo5Qs0zaVYL7t1Cu1Jmm4C/sPmtCLFuKPPxVGFT/Mc79URSapkRexKy4hnGB3ZZU4ks
DqtQ40Tk7xK6CeJs8rImHGBi3SlDGNn5wACcWFsD9LjJV/jkO7RHsdRnRAYkarYvyNXUBDriqzq2
0mwADNa5yokgZH2rYKnqg4vSadjFuB1iO3Imatk5CG+8bUgDOIpXTNxHfQBSEt6ZfgL18Q94xGYZ
PmOoXBBSFKq5S5ncTA6HOTH//zoH5/nfl5Me7LVLyJB5qNDpewye2l8K7o5V54u+UBZ7gzbat0X+
zRQzHYDTKdPsL1aArjMLcWs3sxDzqs+OgHvmLTyOsv7sYK1VixJ7Cqa+wtmDimYKo+faA+m6bWdf
/jsOativ1Yygbmz+iLU20+AlmYFtuL7M1jRwahdyAYAAdkiEGynVnSo0YpEviwKIcwtfLbLSPxaO
GBSduqZCKUwwTdR2V6hPLtZQzEhlAbowp5+PCrqE6v+RcmmqSQLXryfMRFsU7+/NCw5UTfeT+1CF
8eJD7gCh2BJ0hLZP5VKcwsZLh92ElKKe0tuzBnV38YNk+HLRuT8jp9u01MULXP4KL6cVl7EglDPS
GMe0K1mnQWaRElu7HpgiCeSrMyFmrV48DI9MkgxhR2WA2glbZhgvvHqEpMhoG6CnKH0ieXtciEBm
l5G8Rjwzwu4U2mUa+yBD0r0QJbO5AcWuD+P8RldgXNrmtbyZ+KJ8T0D1UsgSChUfJBrD66ZbijUj
LCsSRFDzjQga/QmI88vrl5jHhMwmIXQ20Iwg8depF2bEdgNMfJVmeEFDoskxwCfLnOQBeAW5bn/L
iL6WI27iEfoBL/gnv6WUJR69GyJSrB/IGi37LJGgC8vIl68MafQTKHSxuno8RifAZIJCySYtcjd4
HVdgiFQbZUDPQdUPVKc7vCWY5CNcQE7QVRyTqa2v5i3SLARuaiS2jmXEJ7LEjSjHxkyVM7fbwKqp
X0aK4L0+e515pd6SNSIP0PWexhlpWFA/vgrwzjQuWeHzeQv6xirNoMFOvmpYeptMhk/whYDr9zwL
Y00RY9VgnyE7srlhLEeW4q0/lMqPuP/ZhSiWfzf1KUC4sDeT98lV+/AC88W4DMFxjGlQ+yq0cnZU
WqgOCIZhuEpWRHrAZeQ/rqrk7D56tb7TakhIue9U8ZFWxved65iJej6K4gj7LXipmHP8lm0OkVPf
/NYH4gc4c4Pcdec5AC5nv+OV+WU9JSawyBulbKGPvoOpBVq6fBMd30Oets679+D/goJVwkqVXxcq
OB+yITEtOejF9mcXQatZgS1E6gLfQOsOx5WCRf7EPXGQSRZvy2+k0Qf/IVQkE7nPg8TJfgXMthkg
R7lzr0T+XSP5K8c0fXC2/sH5zQlXAwjH9Q3Zyd/6ma4eL8fvw8MzEuecS1G5UDDgYR0ZgTqc3lES
ZTnve33B8wa83x09UDSBYwBM9nGuzsPYII84NWUoEY+YevRB1GUkU350chSYmrvX3WD0m19n1GZw
05uMYa8g7QUZ5RDcZxluUFV26cdU478BD/12J9LgAbd6Wh7TvXwYcv2xBnhWmuq4qtgatuImUHcA
s8xJmLD5t0TEDnAU/bK3NLIKqvQamya7M+nzUX1k2MEYpIgdR/zysgBjso2d43arzryjxWRA5Zu5
UqUANJ8ikicviIMb1a4+5ITd7vTehepU42CXkoKquqc8jxX9pvGJXjGMvyNfYs50QFGJpxH8Hm7e
j4riuqDQBRnvF6CWZexFBjV5s0YESnAr4cKbBoOYlmF0Rk4+BLWEuVwVtPSWMOdvHVGqRfcGMIBX
I2DuL38UGuoL2IOsJi16GV3wqfUVozsIlOXdOdfLhNik9ARm1bJxebFRcQOXQWCltOxu4jaQ9nMW
JTPdooGUfT4PsX71pE+UcIKgXz9HNm3GPWVA4Wz5xqdh0/93K6kELOYxExDAh6lh0xajO05Srh2d
bPwB2uyv26X8ac7y7FDuoREewYyzh3oEpA+rYXCnOhonwvGnTeR257VW7/Qp6MUji6J1VHzT5oo6
RNUyBtvZLnqDSCqmw4pzkat6Dkeqwz0WEWTLF7A1fj2//m6IBww49T/DiolijhM0k/Vt6hhOrU0M
KW+S5+HR7NodTTEaKGw7G3sBd/sbspVN2u8yi7dZpISKBv9z1k5QEkCXA3cCg6OU9BHSH1CMZrXy
Kk+NeKo99UQjZ0aJ6Ahp+3/ngh6tIt3RKrTxDIFBwzaJR2WjUuvJvL/pyyY+oPEl4BRnnLYl4+A6
2o2OHjfgmSPKEkS08lXnVbMKVe5g1nxJn1+Xl4y/3eLiVFcI/nyaVs2yNsI5RWUMoPAQTYRi7h8d
efW/J6VlD7ooBlUU1WW6DPre4ZfI6JjaCH7A0amne9BAQKaBbCf02YlsfP+20oDUO7Zln39aSnul
xxbIT1QFrsQLdWkzbFhpymqvaeSbTMat8u9K0QUXPTLStxrKIvY53bQaZhJD2Yz+QbMdvmPmeWEt
3OmvJT/N8aFe92twp8GawGtOio/CbV3QoGpNqEHzdttSUMKbn+B6A3MszSosK48JxuR5VDFNh6zO
WFsuLKllGMH3osdkGyzVMq/+gYLm19CdaMypuSmhNLIqtlPVjH9MdFnIla3JConEs5P1LJjeKfeR
WZhlT2xQmBYPVlCTqZ0nlnsVwichIUSJ1oQrpbKUyHwJ7qv1hXjIb0VskPqqkVYZ2fR7IpEjE32E
CNAIhA9Bs89xAU9uzqbqD7PVBz+kDu1jHAIOfqCtJcnFuAuKimR+5DaJOlqWyH1zzkJlcWtS9Sy+
c6dCUcwBBszGZMOp5b0d11osZsDZuZqaWjXt1TVkbQSidKYaX8/5NY9Fx7yXX3Y7+rPTY9xYwTIc
+69QPc5FXOZaUw/0Z+aRUlPvJY6WqRJNEraARYl0sQ6p8aN9o2gA/GFY/KQDcemVLHTMe7F24G4A
sHTNMHlmMe/nFgWbQx2xqsgrIk+gQCZ4m4Zf/PU40BjbfXuh+3ntxAvwUuuL3vk8ixw0Zs06/+yW
wC32NI06i++JeVktQtXFGuArvWjiIUe9jW5JvUaOWc2pO8s7O9RVvGZ+sURg6vmpjBzjfPXnzYi/
5pd84oyLvij16EqUiAoKeofHOZF9ke06XFaHAC4vWG1PA9aHx9gSr6X4oZu/4/zry7LOuV4zGBvf
2Ou9j1sCBEQ0FBzPKmLFcaZbbQ8WLwaFKA8+JdjtKeMiYPFLJ9oUZWnsZC2vz2apnxnNFYs3gxex
H5WMhBZlqDRWpfxp12rsYDhotSMehPki1EjUKffsr/QEgQIR4jVHByfnNmrL9dxZYa7WRnXCkN1f
bTz0PhfzQgvBPPpBWpKk959Q8au9eeOlukPqzbtyjJe7KSjcI8Md2HqS2sxwb1zG9BqfDjzr61Qp
BYb+xy7VL5i1wj1pjI+RARHCevRvTuyuX8hBEq+mNB+vShfvmuz7LyapGLQ7ctYqKICZih48j8Ct
naKgmxkuU4AWKuV7GFdAGN200NmJnmiAY37RJmtIbLA30kPnrdWYoAsR/LpkaQNk8nJA8Rq70LjW
FpcctC/l4T/L9XsnY8LU7pzZSvBtqRVmOTjZj3AcQ9eoYbibgMYaNJPNvYyC20uBi+kvXwhqIlza
uV1vhVUWXGMOAMe4KObQpG7nDtPfSXOhH6OAI7B30buZ9aPY4eDbDQYE3ZOYN31lBzCsGsx1QGk3
d16i0y+hEMMQL00y7ALPy0sxD/1XBlEJQTrYnehCpG0SFBQNx+q7jPywdxeYNVgPXUx25+0BIQhm
DlaQSyX3ZrMxivNm4QdyY8l71uWfPOaVEBkl6YG0KkQrhmHIzVpCwWeurtLOs2fj5QJ+k80Rowwf
sa2qDPo6Ki+ke7+UD2P5vVFNCUmYCVfs5fStEbcKBZnlHmKP4ejTJjh0RhtCdzsmytEcVjcoNiDu
8FovCMk1gy6stG1RUL5jL6oEOd39GQpi751UuIZpPUUkU9V/Z5127nx0mXNG61h2eHCnQITyDOtR
Wz1t9PjyVxjeosFfk5gavpR7+1iKyaftew31wi86DPRYc3xmGbApL6ORP5cGDfiOXDMc7rrf6/YT
nzZHAiUFcO7YF7HeGdmMyqiszXyAd9gMfjXrBZ/uBC60OAn7DOEGKxDC+V9D4AmXUxdKd+ciZAsb
nB4qXO2itF/r6Q7duIzTSSFq4LMBiNalap0fr9bR1PM7uhvjhif9bs9oz7m20RVwSXLC+6G0ATJe
G//0zGclxIr914Tz5jKhDu+RAa/7VJoyG+5nEW3pU+Hu3vRAY58MRzXEDSRQvveXH4UhsibTvYv/
oBX20AlvlO6rqIohmpVYd123NjrD4BjRpc2hp96NsUHWQOXlV3KaOPXeI33aIaYeFTQe/DkU1/ZV
E25cxvkrjSt9EhZThHE6Sf6F+7LT5ZkpfGks5i/gbAp2QaXoJBbgmy10FtrNZGiIoc8V8FKpTIhg
ooRQmB31x5M5uLNWwdRs1liAdbW0yp0Qcv70LBfykjujAREguDbEvJAKw5bulLWM1+IFOSvT3OR5
U6ob7ow9fT33zO+O0OVZg1IfujQrPPlUiiQiqQjV22SUMYaMLkGYDjTZ3PdPn/oVGutKlMGMP+8V
yhiYuuNq9FE8M21HxtkBiFNazoj/rzFR3Fk4fwpVMd9GQ1EOzxLpHhvO1CJpFSIOLK8qf++2sXAB
8i+pIwAS2SVMmZavT9EZFUuJ8PLNHtp4HUwfrjvC/zQEu76Zt/O/Ro9bICBp+AGyibjo831qqMox
ooEMJAVuw6Z71S2guifJ4O/p+SMk2JDi6GhkX+IEXmlsiXwbHGRoCtKvquyk5oibta9x7crd+A+e
Th67E+WF+it94gha0ioQ0Ekmh/hQ3tCK8D2vg4tkVawq57TZTkT3u78kVia+XThZMP6E3b8NzdTY
2u4XzJCJftQi3Ytm6RWpHw/sFvTKJCa2TljLgZb+Mm9XfQoaws694ApqLQOu2Y67wIadN9usVaqL
D0UsHWLMrMMvwV51BSpLDjwCbLoeGPaYghFSOIz2u4tVF1kwh2C9WJznqgZiwEsTvbdbib7IMwIg
wZgqAMZWI9RkgNNY5IBZtKm69AydpUjNIxgjSEC8c8uhzqC8Xv8KndjVUr+uXL7a96twVwNGJ18V
QFCm2NLS2CuW9MtEjOtpJLFhrIAoZ4modlZIgJCqYNhfclQ57qaiG5RyxeATU2gvAUbgqrMDwPi6
D597cCLGiL+hZTfBvEkBH+nDX+y096oYHjiEj9RQW8/Ehhigh5oDROEFKNmdTNf68r1YOYU34XWq
iCn07pFaDiauS4+gqZ6mcIBw2cDhol1l/VYLx+RsAemOtIrXfmfLGm7pp3yETMDF97uUOewLDNQr
U62lu/nPH9hTd6BawxthIOP7iX4Ec1fkwr2DX8INJ6TlHzyujENOesj1J1zQTgZb/cGVrW0gikHG
wuPHM9uMLLNsphBtk7IAIb5+zXmueFHIfD4hjlZGJ8oM6ubuArlj6IsSjkCDMKsbu/IwPtbAPtZL
kvs1460G8ZizMf/+6W+gP387xBI41SovOz1/hDkAS1WNa0dwzTOpp5JO8Q4KpqztqADE0ki6VTx+
eZ3rveqBD/U3VjJ46Syhj9JUsxVuWXo1kX0QttfyGHP4org95WWr3C8j2huorVL2lLRfFR/UVa6L
5uKa6n1PRtJDHlZhbtBmQdovtTpVrN1u9z69I5mQGo0R8al5fBPc+dHqbc5sjTwX/xiF+U+eJnMT
UiuSGm0c/bLGJBbT/lSrpH2fLZEohpHu6+1AARpxu/sk6Cf/WkLHeE98oT9iow5IOeFOA6kytOpc
wjS9xd1CvwYw0wKRSeuXTpgsO6XEZTVR+yYsS1EHRfYrTbPVht9oonRtcHlS7WJ73usVGzq4i50T
8Enw2U3n9hYCjjjLbILoutupz9MOGBZcXtzhPq0FtBldly2UBD9c8vyfDPGSFbdD0YG8d5fAvQyd
OnW49XaGHv30m4fcfSvmMT7yIrzDBIZvfjiHaUkkAA0Zr2P4PgRZa7vXbH3hPpqnOKLnMmt9YrJZ
buA6nKg6e3fQ++rmcKcny3YBzcKfHNXBiuVmMLvgARV2BJcjVbAknIFGy55lCcjKoxLGiQqgBPDJ
8hNn+FErKgZrRrXXYT9MtQ4v6jM4EnY+clKS1yUy7kVROhLhYGm7gejRwC10RdQoexvAif4ZnNCs
40ZTOCflQXRMAFLy+43vcIV9AhTUUuMQjAdGE2ZjQoHLZaTtQ6Nqk+LcISw/nzCmqZ+lNY5LdRCb
duY4xtP1CGqLSN6klsTPhOprBTv97l/g8jtErgFUA1DByp6DaT2xE6qnnYHD4crMX02L/+ZI7QwC
OOnlPAzuVjnHvFtTVX0hhRjlta84S8TG97b1UtHHGqjCfZvS2CWVW6x3XCoPjtg8DdKtRe6wWSp6
UZVaMHQV69vKLQsI8p1lJhWP25kRUd/gJTzXaJALyzmJEyCy39lPfbtDxXCgEyL1bAE9Efquh/ik
lwHPwvyv0dKACpP0dvjn/xqpU2iQxwBMdIqM9NxRl1DkImEKqmXNG9B37EZZywEnXhw6LveS8Exv
2MkqekPitS9kSWKIGogIrZpuY/TGNN02UrUbwxAckZ/0L6X6WZ/DU89CTy5Jnvm7xqMz1N7tPyBO
NcXJkkvTXhOv4kMYyZP9Rm1OLnci/gXxcmpy89OjP1ViBsIuOa8TWHEzMRxg6ekHHsMKlUY2AUGU
ogsEqMIeTs61wFM0U8lYK+zlrsEpUDWCZ2++Vmw7n08vjgj8I8C7L10EGg58bHZwfpbIrR5qJ4oo
/+C8IBeonBF9UvChj/vizC2kG+AbSdI+GjMmf1Wk2bkaJuu7+M5FaahaMEbO3njkg3QXJEaAHp8E
Qmh4mTBbMML4I/U9GvG1VKfZHq0//QNh3jLIFL/xU4O9iM56/AHIuu9rHbRLQC8iiPVV/3gYDN4r
NXbn+bkMZNUaeLO5DDjrUW1TLH78yLzJxt/QBImDxpTgqHNQbaqJpnz8ZQoD0JVZJr3zdB3EgtYC
dFRlaMpTcDV9eulW94rzs8iOalcokYmPOXGhLuRnsHVP1X5SYAtQalzfwAJ5GTaWtE+i8AIEHpjg
swT8OECJ+YAlI2xdDBNgJ/Ul8E5tW3MeAyRglsX+249uvklb/SP/OWusxvVxO/pfQJg91EPbh3vy
V1HjCzSAPDA7sycUlS+EN7n8dSsnwwU9JzPMg6BhF7z4AMQuZmUAFwzHf6XQTakdZ1/gUhpPUCmF
Bdi8lnblxgBHA94pjdAEuHsNhOFLM5ZblZ38ennR+FyJYbH5VWL4DJIPAyBPAv8GZaw4IT7OtWel
9uUrLaKTxYTalvFqj7QZNAERh4DwhmG/umf5XoxZG//BDu80DNRrDWUr0Wto39fQRi0Rot3oz7A2
1Rj34Azt9s0uSD8N8TGFSgWr7xqYV7QwPCvOLPYE6lCFoXE0kkzR8pHoScsjzqQAIuhFZu+W5XbW
3dS0rpdbtctuOOZl7JtdIwmFGfP2PQ775pnSfcui+50t+CEFJdttnA6KqksZbXgGklqMrh8KnyY+
pkRPFhQLnAOEysPfDlxiF9yiObQIxAGSuyUYB3QS00JTS4GJIgUbpMZNtcaKALWWfdxy62OXnOjR
1X1HqU5orocZsUo/xd4enqvOcBQ5l9XeICvzEaGTbyhYJA6E6AfVgMHJNJqbxFnQUvLBsvy2T0nk
hNa9ajwWJlCNqaXR05QfrjWJoEnTdzsrxBFy1v0HMYO4vrcIAIUPd+gGy7zKpmTqJSrWeYhRDegq
u7wYojFdH8YGbK6DNCUvO8kgBGhnC7RzJ+qrswy/IrP07xtsTU9Zkt6J1BvKfGsrgZCb8s7lhrHp
r6crWx7Ele6Q7I+tbTnXwJMhgt2hovoE350EjzYXXD8xcTYLDokv8Q3vA5cpQxIU2O+VSdSfRXSF
hjoSbQI8oS4+ZdxcvcSQe1X/HMuKmNPrpATsvxUfp0ms15rNm4ZDTGmlxwAYWvgy3PZ4JPD4HO94
bMgM+hQH9UNcipofW5FhlV3gYD1NFyvBhvg7WHVNaPgkOHpT6dX3GBnlDhXAgWqPKd4723FoJQgJ
q58rwsI7pyaQNi/5+i4vIhDfZ50LTjZkaq0ac+ZpKAYULrOeDH5bLHooqCWv2DmaQCGGmwVPWg2q
PTqppHHw8m6KOahVZvZW1yOfjxzAlqS6iia71mpCbjfaRJLk0ZiYkfXidzJ40EYABiLHCDEodd1X
e20yYuwfGW5gRDSVkNb0xvL4A5y32E8tKkC5VyavEfK15EZsZx4hg4W4cMj+VqCOfHtxf6c+BQyE
whvAWh0Jd8BtXABuiBNWsi8WRXQaF8PW72Hi4gxJddx3LtU+AWjZk5sx/6u9vw4V14pU20B0bu/H
1QP24gorMdkdedAMWpP4xAuP0TEM6iictkvP/M0tYcE5m7CPMGp7iw3GvhaJF9c8TRdJC6Rl8xyC
DrNwBnYFuyFppq+Pvv4rBLmLzBKGlRnbgrCB5HKHLPjEVoZLO2bOcgcTpaqXpDLk8aghHxMj754M
fp97axFfHxsIfSppoPc93OYtCkWI8XxjGVBBzFcBqUN0Uo2FhWgVi6bh2RZTXGhINOFrNoO3AYIH
IDuA4KtDlVUPNajkgT2FjLdoymvMAqHy5XvF2S4Ndy0gFKZD9rXApTClB+oeGC0pYq8LiV5LZ+8O
eOJ5DR7ehO/JpfqMuHiyjFkSOsRPFte0hEZo30PWyPpeyp08tl/7NDkRZ+zQ+dVI2GRCxMUcsVSF
HIftDWbOw/1Tat6Y12qxdoMMpFF95NJXf3oJvFcbrtcawRQr8pH2VnyUZIrRO3v+kfAFdEOT12TC
C0cmR5Pl52tMgzx1shSFNu+gdgBvXg1stehzBXQccQReO7rUGfL0jKWggwB+MS08zS2kKpZ6mdkU
23GHnRchAQoz3K9DoFnAouNfcHexayPjovDrDvvdZ8Ki/uj0oSTo09qcOj6zPoSW4Ct3Rqqs1AlK
LdDyTVPbt2PieSWw9Rei/AAoCxDKZcj7FEzz/pZay6O4igVwDnFiXzptZpZikk4Vye+OjFOB+++j
Mx4J2kcoh7mdW2A9s4TUJfLedQwXtaOdsWBSh2G8J+gvslFVOXl1fdeega0y6mwQ/YzBx2k40ZIF
Mfoj3/RzVN/9VhP8s7jBGbiQb+W8/8lo/Xz9yNNOaIbMejkCcExG3CrRNphuGqM/7m5eVHev0XWe
oJb1a33iFRLXgISRdsYVQ9o0MPh3v/H2m4AApWTppuDP1vuZT84Y9yLa0XjnmB5QSMV8KGxjTiwa
I8nME4mZMJ1rrePdcV9ExEiJw+HwMhqpzb7VUVVKbs4Ef6F9aHQ7QxDYt6GEG/t2LOukLi3kLE1t
HHeIUFOcliLWg+15KdQqBzO+W9xLVmuG+b/KVMQNM7ebbvvXpVIm6WJKAjhw3qvpZdVLopi5k5a+
UILT8bWv/9YVw0X5iF1WSk6j2BojVVyL2q/6+iyTHhCQWlfHv3oEP+bQA3h//UwN8qKn1WQfxxXm
grvSE57A3INP8SvhW/VgT0jWuFIzq4kok3yrHLglzevHs9+0ispXgsc0j3UPTbxa1VFvgreis/ri
qlyw15Vh4s6PT7QDL8vbUIia77kdiaMnIpGDRYUspimDKhn+w1h5SutQq7Yo5oim1MvOJalo5rxC
UlEgJ6iFwj3PhDgosCkLsPseYimKVnD9RCX/O+E9xq4+qrLxwxZzl9hQz62DV464ADbR+Tit0N8N
JdJMAzY/hnBeuIDTuZGmuzTF8SA40qdhiJCaDEIS+GaKwgVdd8qOKdzuyyM62iZt5Z4t3sL8pM1f
PIsWdlL0ihFWr3I08WTU8UjSAfG4YIZwiFUwICW4ggAQy8yQEUkqQAfvYTBWzzyIaXTofvkaKiSr
ifIy49sEhZJoMVrEgPy0qR17hBpHc1nZsn8p3KjWtU9tEgMxgtEYib7xHvJ4+aLJXi3e9prQcDrY
c0du8DtG/1gBk7pX40BjRxFbAC5mvKEz1hNqmjCG3ttKCfx8VCSBX3NKsbcGkpYUfxBkk72je1UZ
Ow5izMwsfTLsZJnWTcd6x5zlRHgoVIaxlM+Z79RQZ8YSZk0tXYsrQlSTy7zCpVOu/PxxVMGN1T7Q
LlCH6sZ407AifFZ0Cc4phcimm1/WHWJ1mRJI7CP+OiF9xMTzNgu1plnv7mIDnyZFkSQlYM+SuWjo
D1gS9f66S24XGg6az+7a5U9dj++/+659VZVt4HKzFmplCqQRKqtq/gDe0R+NQi1Akp5FJETFmstc
IxGNontplNQuWwu722FUU3NgsuAGi3UZ3CbsEQfv4/hIly/Tm2co/r0Hbd4Rub1YsvGPy42HM0pQ
s1Kc8fver3CU6GsEn04IgvjZY5u2eczE/Tq67BoBX6psnjwmpZoEmDSd8dCG8ERK3VVuypdzYgcw
dw8SJ8FsaRoQOQtiqSQrnzpeHIXzM2LmmsCl2rmQnGV7/MzW33Svc2DOo/9Mf19fNIu02dsN4YYB
JG9kZexdZ8KX8jpl3x8mr4T2wMUQckKxd0Zhv5agCyjz9N3Ex7mHs5E3Ef9zr/RARPvuOuVnRaBf
xNZhhlXMOwpMZxxD6sTiYV7gymS8jfGyzpxn2BjRlzTN4nXMu7RIiD46riheiXcI/6K/U3i37JL7
iPeOW34HWuf9Nkru8AM/ZYZ7v8ZzUu2kyTaBNRU6hV+i604UYQPqV+3AFwiXzLPMS+sAmAU/JrL6
vCCXzynZ1MbELL/nHI8+QF7ZJr6LwUs2PO805Ec1HCRoumO0M+Lc44h6yOxzwdqz6pnYHEAMoNrz
F558lUQibmrHqxMHYY/c62gSwFWD6wJr5ct3b/TkRbUjqXO3QOb8KYvblmFIE6AZSIhfR/UQCDss
GhEgVAP8D0lZJEtCOTgrGIdPPS65ypXLgVXQ0Vm4fg1akc/6LF5r6rWRl+Wzz5vjeYFNZOQeQBAB
lu8qzpYVQxfPrkYg3Z7jSDvTIucda7Os5EqOPv27gdF0Xap7PRHjxdG/c+vTkSTlo0QQKmxgGXTL
D8l4EgLF6imuqWnDEgbvtc50TyToIbv9COmC6sWxuMOMbL14u7MyQin/UdqyhR+JjyNELXltlczJ
cS0iznvISaUgnnoC1Qx+kVJhK/lQB2itzJKEnvB9+bbeqN4v2cjear2wJx0Jq0xYDy4y4s05wj7R
XaQYNyZAkJvdE+6M0JRT0WFTBiKndhWUX9XhHsyaVZX6g7rvO9tdms4z6nQHwj7kDs2IbaH0vSPn
BsjyU44el24Zh31nFUAK1TxQZ1u7Wb0ewoX8S2AZqfEBCxUPjT2eKAnjHm8JbT2+yPAUhfq1JboG
5QftIaT8CRTOlGNeBE2TB4TjSNw3JogmJTeMQpnx0VINMfAeT7aMNGO5AL3aiiIFNluRbsCEHfIe
0LwWxVeh1QOwM7Zo+FkUFNwtjjJZAt+XV2Xpocvgpau0s35dFZiTJmbtVctPF1oM6aJRr8tiZstQ
H1mqfGEV4aSdm7T2dRETRaz4Nd+qZh0zuu4PPLwPyLf+I0In8cuO1oXHJWDoBowDxCbiyfWiXadU
uVdSIbz1MYyJICXdBd+2qoAepOnqR06VIAzsdRvrgx7NZWGE/ylOEUg4uXTGi6wUxOl/E6H5Znbh
8Ym0SBZ92dlIZ72MgYRIDZdW9XtRRfxjk1cwG9nD/TeV7Iyk0+H5u96m5RTCruLnppx8WigYQCrN
p6cdm6tuLhq7pqvnh8KWu76t3lOVtkHgKywQVyIdEQCkOe5j5zt7iYj9yGdqZNgBczaAvAsizO3n
CCtRflnIsVn7f9LtStVnav7fTaSKPG3mXDoMPvdbGBylgNdLi8HSMkqNemXS0YF5qtmBN10DDQSd
nSyXHLMswGQv6pjhME5RfY6xp+Txtz+V3deJHPBWcM46KgddINRIH/Tw7v4jIQ7jaFwq6/QKtJkL
WEOYYLWEg/xoATa8PCnvbOJNrkNnRWaPFvAWOMkML955r7Ht/W5ARSqGG66sjBKkb6X24zz+b07D
OpTaV9zYYapXSj3rlOgbd+snnSHquUewUIKCssARgjEjrAW18lpc9ifG5w5yYH6wYbVPmVkkzIhn
gHsP/+41TN8H9pHIykeBJR8esh5NQEAyfQoCwkWWFRqhJeq3F51OhDCqj+BU6+6cJIA82uoNV/M2
15F6XJMayV2DbV84be6CmlvA1b1rvCA4cdESs8ZtqvbDlzQtZYhJqELpQN0GP1tggVkMFPrGH1Us
6N3mTxqB7w5+5nK1xzSCSbEHmLxHoz/dLARwKczG3vQLGsXGfFUnE3lmY4YXCUWvxp20ZDofbBPX
1oEV2WrYY8NyGwYCBecCW3tCq/6k/biecoDnk7ly4kyjuB150JQrbBerSNKzPCQgmgTkIGp7hDYX
9HERvCpycHymtWSD5sh2tBN5tosGpXsE91tYIjMCYrdn3ywuwM0ZPbJsHRIwl8LPld6973rpvWvn
70EiP/dTzchTZEK2kbflksdB/sflzzaCZJmOu0wfgar/TOg6kLi8io9dueJO8bLH7v/ERFGHQ/wv
StenMlDc8fZKIpI4PIJOPtauZCcmH3BUAfv1PjF4OBoy4X5JE12Aeqi96tV2j/gL/YnOPHWIHcBv
8CFmnUb3xCuz1ZxKfkXLKw3iztgtdSOEpVJYaGrr4/OP4JZGDnC4lG26zB6U82mn8g5+i+nYrMYl
svPLwCj2hssCY/kJ2Vj62ODr/uEJogZmeTj+OPETgcyj0h6fPJPWVm8cpFiqZYhs11R+ekEqYrNT
4Rc5p2q0JaoFLOM/m3ScvAFRz4xp7vIzxl8y49S7+ZjIYS6WR8ND+HZsxjvoo/C2M2wNHbw7WOZW
bgxAp4K0llzYHvOUHPNCYVGOCtjTr1f7FKGgU85QklnsJckCtNJbFlESzpGoucZt3A8cVtmkcD2P
rFNybLtSGvE71fD6pt+nUbEI1PPQVahxmk/RC2bFzgpGLwt8tZ9pqpg19nwvLpqFFXAqDY/q17IG
hrz4Eg5SYijIwYJ51ZMWOcZMggsBu2Qtlkkm2td35U8NuszIfiWXswrdSaacU7G37zn4ZD/CD5Pp
76fC+38QZU2thIxv8jPNF81R3iOhgZENMfuQRmG5JSXQFoGmuQ1zx99/sjBEG59QbfRuS0q3Kpaw
OHwo4weoOyiTyfcZv6aRQIV9ynqLFM0xaSKbDcVW2gLJoEMMa0zCRANt7ZPdLxhX9sqonAFebdD4
2qvKlKPoe36YEHc72uD4nXYxZv1hyl5mPIX4u9puJIvrxios12Cl22bPmc1A5CExdikOx1aM+cMa
cVF2enXUvq74XKsdkorYj4RkVWqGuDKs/UbJ3ns57O2WHcJt2GHXxFmmlHrQTYi6pgoSSplTYZA1
jeexzet+8XVbLh5rY/5wjI+aFcgxm3/S3oqi3R2Y6HPeURn9S9VsIrpKW9ddNOfdC/yPVMqLIS1p
EIFgukbYIehINQqdtmACKOUo968/h9j1dl4tn+G1Mxeu+O/2+coaB5xyeEPtN5LHsJl+6nZjHFhl
ythKGa0su7kfUWp852bupyRoNeIpjZ5pnHZNWyPYN06cpHGnMKkQ/Ku1+wEF96dBUa5BEoT9sk4f
8dxjJjx5fjq78NybdNd+IJ4Qo0S5SxsX0h0i+5A55dTd06oSFk/4ru3qCvIDZdXBjeUrbdANpK6m
yZh7eoBy2G3T+S5yQ6KbMBgKVc+QqdI+iYjGHVu9B9rq4HDrPfpHU4gYx1qVxQ9YzyXAds0Bl4xo
jc87hS6E6X5U/tdIbkNAgPShRuQC4e1+CKAHLIdtualQ6/6m0pNy9V8F0w+KOp5vGqrmWV77ZLst
V9m+HP8PW4lTb4xyoJ7PGHyMIFisVpIT0qTpP3UUcAz05PsBL6D0gO3dCx5hBExKNOS2b+EPG0mS
MxrwVFyoKkwa7Y/8N9A0ol6WeWqIFjrKTkVb/utJ7ADCMQQxClekMzW1TP32uOOG7t9MoaHdRksy
0Kq9d0Nn3NofZ5CwyRHulAA/oNiujtAL9BYB7Lk4x24ekAjUFEqEQ3uFra0KSCibRQJUEmyL3DqV
HIbR4FwiGjcr/a3PqYZH1GGJ/yKU7MqiVR4286T6c3IB1OeDM/wmh7sDE57Vy1V/yzqbVCrhEaky
LdZRGnOnIXYiTc8mNYHCsDiKk8hk8w1/3CM96Fp6/kUJxRmpzPOvIr36DVsJmHVVO8zjYL+ihspD
UzrhHB3fwL+WP+0hVE5LOOoL0KeTpk0GfyPlv4xznMa5nkHwJ5inrB/8Q8E+xWJDPFurZpk9TZnL
GRoSmDysB30P4Dp4nUF+Zc7PShJsk0oeMNYwwhCKjiLCemDMfWK0JM+6TkQYlZXdFOKSreZq+QN/
BAcXksy4lDvdg32grPn0X4+u6pD5f9QHzUMgzJUumM8Vtvu81sXfCqNGSTQGrW7lfbDExB8+hnDs
rBA+ZaeJFR+UzDaEN19wyVOEfyIu/bMpXCVu+xZ6D2cDuFfwQkJD0SlWypi/aDoLyVMylyTEwK9Z
vmyd9uCsUoOD1+U7P49a/BSxqwScUMo23AoQP8yeCZPQgEatc7vkcf4Cj176cEXM6U4nhBeKAPQy
GTbQDwE9X0oZtLNTHRvXAHf3Af1VYN+qtF6VV3jZPK18RJZc/MMsWzsPteZ5CTb0v54qdMetcFnh
H3p17fGmsXMzFaLJ11iLYYIrClZenIpVOJfxG9bLC0umgfV+/c9+6O1m44Mp5H6SRLIO2m30LQhj
f2xfg7zhYZL8a9rutZ/9QHYLExSZxdjxkNJ3/317Bz6EQ++ZNJjdQ4tySPZGaCvwz7fDT3qE8ZUs
Kn6DYnzBmqAVUTzMrLG8Z/g0quN6AS94Y02mC0jt6lPJC0iqljmJj6zU6hEEpYxGv27ZiYE7iaFe
s/WVP88Gs/fQrGlM83GftMbFiNhAMT4IUNPZpM/Kk3O0HwjxDqbGT9IFIsSm3nk0xDm3Mr5CtFOk
4W910vz7U/GW43vRibJhEAMtZDwzrKQH7WG4cyD5+JOpfmxYETa5K3JibeXWvIThpksgj8nhyjtr
acPtpfd18YzHnB8rWau1M5le/JClMW4bZE/jCbLTFGsEtx87Ao9G6/rw3zOI7BTJ1MMtvSYiKhTG
nS3aHnOAkrLVWqnSEYPsQSO9GppcaSRld8g5r81vi+Z8KgRH0gYmDSWDZVH4zkvnBItSicnko8tJ
tAcxpGR0imdEONtZgie7uI1jpxl+IAaT8oL+yO7F2Mu68tBgjPpegeuAFIPp7nLKUnn+16O8fv/V
mB92s5XKnUKxq+eJy+ZrVWUqrpPCXDQHsiROtbaswBUV7Xuo03wWAWpjlTvf1Sg26TPxUEA6aYW2
K1lppYXL09I0zr4md+Yh79ufwHi2WFcJNS6+/7cXkJtDYyBfSqwdi6pFkE+403g9OsX1a302hh3X
KMD66i8AtLGBWawCZJALq4Mm/SiPs0VfwgvdA1ZFY3VJ1xw+4C8NseQ/aB+oVlXlXVMTSXLbGFMD
rO23B720BAgYmLg0DGkm5YebzKvQ+DSmpiGzmp1hzNA3rpAyiU/sJmgDbXWW7BKpLClIIKWmCYzF
fJYfoWhQeneX3cMiTUocSwyoosfBgGzp8UyQjpEBLES9cMjFpoDs2MxzFJAlv5yTO8Kk3wlTs7LT
hzTPCIICMBy+SoercPbPKqfdeIRu5MNsSr38bA3sdrj72GtAuZBtaQq4AxczVyrbwNbvIcxlabJd
pwdB3vuP0bS0+KtINQ33XQacHQCylQHAyOQTCqhcbBN4HwxS00ZAWV3z9c0f7Ui7LBGF0UTdtvNw
ZAO8GidMKigtefC6ZFpnQOIp4PiIB9pGzG80mf0jdGsCxvChd910WdI7OMx+65YRX1t60wDDHL3P
9UrFkseepF26KRWVNFqw+vPp4X0fnAs7nLX+Z10IdHMuN44tAaZCrvI2P910Nz/x5LdVu+bYNEJl
8GyjF+/NyK/gi6Y+Mem7eipW1ce8yFdUlclX5jN2f8tziMmyuayP7v0mBr701yaGE3GwFfi536n9
SDP2YO6jLGXXZjnSYp3meILYfYy7lTrMSzn96OQJE+zvLB0JC/+hDf4xuV4NIsmZVUiKPHh9B4R9
rcfJlPHjX0ge3pACHEOb26B/r3WtdH0VF2NuKkIleEhwsbEFdtq3k0xSm3BC9/h2aILWoMEnLOEC
PT0yJwzr+sGNdBtRmv88dkoty94eiRlAGL+MxgcOqfAJ7pW5UAS9zA6e//sBPvNvS7sHp7HAvfw1
A7pVDHcn8E4lDjl2gVDyvJ6jslOpvfYCsQ46LFxc+iDTF8lfA8dukAiT5TIyhd1QDYIoM19f/BVe
2qaWkbSwSfbI1W4d2atG2afXigml9iySJqlppLeax/TW+7KIRuOvj08xTeaNArH/QCKm736HDWsb
U8MgHn0hVE+/6ERbnPHGfA0i51wtvbp+x/sdzasjz6ibKJ45eDmOtTLuOPpXPB47JlRAcBF9RQn0
gGr7lrP1WJsBOKZARbyAcaODlYEyfkhzPzq9iA2wWlHBwRvqyshvRqRQybwc7cf25u/RJSpLlOmh
CP8WO8GdOLDQ6ElfbhdOhWvOtJCBhaUrsj7PH3F7JXzP8r387oMBmaEfl/mKaVnnCbIOKbnM2+xD
CnKng/TXww/yLIFOXYsEuVk43kckiBbhUxv0SXZsGaS9dMZdE5UF3FN1V2c1TNXYHPcx739xMzLc
fLAOBldbSHINbhnkLE1ObW5QTRlXN+7EUizAUHaNY24pFnHpeCA8DEro2InElLDRgv7HgvukZxAQ
VwJhlq/jVP0xzi+No2wA26tjEPv4Pmxic96VXRitcOFmvPENmQ1N235YRQi4yRY9maED5J34mTmG
eo43XV2+Fl0sA9xuIQnjGprXD7orzb/wWdwmp2bXcFFFM1yrIeA6ZE2MGDtdj2ALC9psEQH6Zkkk
ygTkYKOTJi4vT4U76zbV6VSjGtPeiaDtOB1I4P0sGMVHpYpBoPWMESG5SNvM8XFwWUzWAsAd2YfE
F1nxth1ZEX+sLj96aF6Vf5B6dac/yuM3IdFf4K6LpgXKlxp1Yo8pgH30YNnueBPIJ0YCstWAkB1o
gqO6RbXECtbCPSoPCCraMP9oR8C3sJzgnhYl+ctkjKG1rPbbKJYe144tLQb5j3Yarha8CHFzc5WT
gBhvPwkTavjFAvBzroF8PfFdywmS/rCjZ7rXik7fAgtCS0nTyzOTqdavHrUOqTdYi/k/wh32aKez
1DQFbEhs36CAqfYXbKXN7e/ct+/eDtiPiJkkv0gvT4+Q1JbNhyBmGTJCBbm+xWYn4V0/k5sC8PaI
UWcCPEQmrBU9uW8TeFbPp4MYQlx3Tc+9cF9MXMeSkq1u0NlgFiGwEWlzGC5FkuHKcasS5EZWdH7j
mJsmBCm5ORWo8tCKy4aOJtnoLFk5FvNbOrQSWUqRUx7IahNY/Zln9XCnqppA/QQJf3vJht8MMulh
nNsuatqp4eDPP2bSQ7rnLHIc8XPEQZsye7XFcCO4Nd5YmISWtSvMfGMJuSiJr3hFCw1uicRaxxD8
Vq7q4Whau5m6ha28FEr72OzOU0SYx6Rf2mZh6XsJquObGoXf3VHsUTwQKG3mp8oR7VFIAYZjOoJI
E7155tNyR1efTBmaR0GKy8bzYLwU2/XD0XUpaxWAePn0NtxS4mWZVeLoep3kYwBHuBNLsqIPWFrB
DrTmkPCgPZz7a6EnQl8jQFY0CV4ZYtrCqmTNo9LxlCVDlciMSMusx/iJGQOHgci2aLj+YLRKwEp9
HrpneeMQ7k/L3wufF531/zq6DdAAUQy1PVWZHG6E4LBejJQ/ZwS7ZEClD/qGEguPPs+2hcxPIKFN
sbZG8GumhFQkCkkx3sYwW8I9JzQer5qjn/uM4UPwvbMu7SPJNqU0YgxayW7c5aoqfY/AIxscyH3n
hA0fcPy6YewhzBNs4pjZ9UhtewUxY/RRaeQeKjRAcBqQDCsHSIZ6LEKYRvJRGhD0yDCrN3iBR9fJ
GBs9KULfcqNlt65HcjII0reK+4NjRNY+Ey2NT1vvcB9/uwZFIjuHBR/rbQ7fCq4iXktHQ0bTXp1/
7H6p9v8wyRz8Xa5gmgTe9SW6Pgsnbe/ShOWi8ClhzxsnTUhaiMEvXdeiGmreFQ6Ps8kQ0fTeeGAW
fvI8u7rPs0QTBHsrqiQdPNT6hOagqm9xQkSBX43RQWerlbmC7/xF+4MrFkLOcWy5iGKbXwOJ+Vo5
Gc/dWzHd5epAxAM4vz1sSOq12NhkB8ukISloZ7t7EFzWdKPkbDBxGW1Ap9jpWFHAAXJCqfbExjJC
H5Y/4d4kJzI1gPEZmJN2cRFZxm0FH+ZODiXH//hMWODYYp2OgPg9KtkAMM+tB7AVgYdjMjqICT7M
ubHQCt3JYzxdxHpDxTjvXsmXRUj8PQr4/2aEaK44gNk62E1R3m6ZeVw7UnRXF2REvLjcn0u9E+L/
lVHhFzngr+0QrPA4X9tvhL2heq96rhGkaH4o0vL6ovuPGY63CYqxdX4COqFlbO9NxTAHMYtO4TdE
G9p6h/iyy/TwUCQBIl1qfYI1Usni3sTQoj4dBz4hGPVAitvqlzU5Kincrne/dYLI8s+nwSLr8Q4i
0TKbZvrPkZaZnYAigmo4jSzxH+6KR9bcxhFkCHWPLAhFKt+QnQ/D6mLWAmoaQzpqUmtWmTMOExRi
msTOMag2WUUGD0tm9ihxpU9YCf+yy8gYyMlmQWyhxm5aqZOHcFIdNlLtZlx13uldDm28pWPZlyGt
dQD7843ZhpuuKP7vLUtxVHfQvKFO/JpHZAMkjPvad6EMqVqLm/I7Al9E0T0F1toRU15te1M5cgIW
k5iV+z4LxOTNX9A91mA7CGKosDT1FsamctG9TOEMdy5PBOhtyusF9NgVcaN5D+Nf3+zvXTxuF/5C
kcBNE0ZVaXxiS/yU2LYsfi4rs//HoRwkHi8mJAg5AV8sGpXe8IKZqvee9bMmARSh7wWIFx5YM4N3
KCwqjSPZNw7omw4S0dZpkIF11CvUEhI22fadZ3iaqDVhBaEBAmEe3k9qEM/hjcGI3MN2BAFqFlru
+anG+SWd+VDpnAziEjWVZUqmDJRdlZWJ5swn9450ebMBaS7rsAMkbTbyA20U3vwgJiie4ONVJzuX
sXxfItZ8YR0yYVGjQvO2mxWdAJt7SKTIbFDVLiXacD3sHNM4hNk5LvSHSkInsz31GFXfUeOyA2/7
BsqXrYG/Hdatg+wldGdr+tsWYV1pCsulVGNMHYyzCdVGb1k1kLwA2xP7yEG8tUj+ta3C5vd18/BA
L2NVAF4gEBlvLuiCz3KJ2wcDK2Ys1jNTs5vp/CtH9qhgXSXsPZQI4pXwWrCN76CvAfmmQh9DladV
EFyx1VRDHSSH2zQdBCWiGN0lbenYNxfvCsqIk+QlD2iyiuODfpQiAOrs5mwoa+xodd/aAMX7dEv9
tgHh625b+mWiEEcoP00CDsNNOaXwLOG9G0zBAMX5XnUdUVtqOk/pJJVx1ukeR54Vi4R3rWsyUyHJ
D88/yRjxtQYfZpLaIaFEaiIdJamtOGreEB+RvbPjgkDCWWKCCGAAhGN+krdilw+l+aQXxoSR456U
/MWFiq9kLiaPsmiUE4l7jjN3aJr3OXVIo35BJudWFTPZsxwrHFKqPO5b+EdRIZQDrY/aCN/2Xis9
VwGHNq98WR5XpB6+dKhCrtbyS1FoNadQSDKmyktXpOUER7paV9vnatlzblyrFHakWV9/CxqMW1FZ
AxRhsK+kcXxz0LyS/H60LqgIsL1t/XJCld3QQPoGvLYeze0epGYS9S1I26mc02zVgh5XXfcYxU2c
xoBRP8gdkzXrfqdkUut6+7K3ad+Q8Ub8wvNEVCju3uzHGE3hiSyMpnfKGYCD/ETvSSvDle7qSmg6
HhHRUFLl++UvDddyEEitqlsJYMbyDPXoswvJ5qpPxwTfRKcH09EkmwLt79PAhdTIzfiMcXUcXArj
ffTqTe9LEISjBcu/TNtCp5v6/+U5WFPWP3qXwAFBxD8DKsP1xreUMIPrZuECcWJrA5+T7dLzu3lC
oA4w/az4Sx1Ci5uFXqbnuM/RB17eLw3PgpK7wj/V52EkZG5qSWp2cBD8btFu6bs5FIbI5hhqZj5h
NImff9B+i8fC2ZubPjRlOt47/lL2YQXlpdoYALMuIP5Q/rCOUikzP/Ih5gS1KSX9nit/zde0blya
0xQAgEVJEwl9M9+4EX7vzO3y0dB//4PdI7O1IUNpveMJVvNAV0vYTwDDQ0TXtEB9QWkIP4TgdTWa
7W2EuURBZaHzhrfNzEQijrt4XAWHb2whHhKWtTvflh4aLBdcwkuwcRibzgfrwytUIVPAQT5cBx74
lj11M+fo4UUCduC76LIIvpqcT6j/vha1Nc3C18819Vaq5tx2eg55eW3H/7t0/s5W0YILz/khlTsE
htY+sgqTGDp8Gs88mV6uxH/ta7x8Xel++RFLpjTsMA+lc2ar2jVkL7K3+MeRfwu2OZapG+4YDBz4
Q+hmUwhA352fQmZYQmWY+ATUOqfiYRg37hKnUOxpCu29wzBfrZRk+90P963bWFFMtQt4I3m6fQF2
42BYL03YJ8ZhLSK1fDalcrxY0tUvcFrnP/ClotmLIdm1tpdjBeH9b4lYzk57Ll6T8mpqcaNe++TV
n73W5SPtiILkNgh4zy8vt+RMaNRYzDGjHsO9wwtbvofCH/wmkH8a8+t8tvsn6ClGhfWv5aIlu29Z
Jd7pDfwWx8MGGiSwAz7IoOyNC4AWjo7nvyYGLVIIE655fqIa2AvmBnJ3NbDqOn3gwrRZNmL03wjW
+bYlhhHNGPwr20EwvIWlYqYHJoOD/UnLe4IOkGb0nlz9+aQoHWPJy9olMHHbVcl/jVjR1Vsrc3Fy
EaFN+GYpIDflKkYyg8bJFjAuILLQnZhn2UijQq7s+aRDetHHZEjTnZrKn/R6D/VGcCdqw1FMRMMW
/wWtzCUattGzX1uOsrhPTdkufy6MhPXgvfMdJ2HwwQHIA2OLNdu/ltx5pDdb0LsDIsDt3RilCTRn
aYT03qLTMxPWDtkfIIb9qIcMGluL2k47/AIxWlJC9HwnOwWQkfphRdoHbu3+o4Zw4Jq5BwinPtLi
StwehBPnfhfs88l6TtJIspnXmM3Z/3vUdw7jNklE8m2Q/rQr1Du9gcXWaK+ER5wUhVQZgkS92USs
sg/1uDKrIM9IBIuLGOsq0QCEDec/yELMyy7VRBBZCDviy9xTJSOjabNzeHE9y7zm12+25jI5fwwj
fjXFgv5tPvYjfsKhOMjgkFTKQZsJWxKT4gLYxqMDzcxbi4FWsW8FS3cGIjH6EiSlXQxT9bgMDicV
pOBv15q11gutL1EkgUSBXOuATqyHaEFjy9DhZOkjlGT3g3Mf/un69ahnmCM4FxpLBDAhckY6a8XO
+bfNA0JVt5bvAMq1HaMIaKFzA2Ee6G3cjTO4Cs4zeOl3+RHkrbNsKN/1zbx7lpe4aCU8t1to4cnN
RZ4qJoLINJt/+7Q36HKgcW3ruoQBRifwL0ednjB7C8GREv+dcJ8ykfeZiDrm4cUmg8as5QOnF0of
JHGs1KB38axinPkFZm5RzGq1Df47aVaestVpi2MwirDVzjg4gQQMvuiufk58aISYfcFtAH72QAST
wmjWmg9twws/5U3OhUikE58ZylqXl1f5k9GIoDH1Eu/vqr3oVfZGGXO9BhFXMOvGbX5dK7gPw2HM
UfhwvrWyXYeU36QNzSPwFfLbLnaNucEhj7S43TOqMQ3gF0ID/8s89d8qCMleX8luD0peE2BD4iRC
hO6axmVkT9FBeicuM3/sLyfJ9HTFMIOAQWi8mzbcQogEo9ypNU+iG41iwbEoT4gth19HVaFdFBYv
WjiOBvxmY9C8h7T9xALEsqy80onR5TJ9CiccQNKyUbL1TKRRxQJ6hPu+BP6dvhl1x+bi2uWl63t8
tJrYY7CblXiQmj34GVupClsqh8WmUwPPWYbWkJuihyuOxoE4jI8qv+N/U8zqO/tXNXoKWeJCJJgE
1bvfx00/PkjghkfeGVkC73zR27NKMAPgGTwIgnurBS6Zq8Xc8cIjXCUraWzRnfVeFHx0tNxB3xnY
R4PE+ZvMAaGW/HsXIBpUwKmVglyORU2rKMJIokYxuxA7yU6h8fL/O226RXat5Be7luoY4I+0/pVI
8Bd7zMZJqMKsaZ20ckcHu5H+o7b9sRUDkQ1Zopk5YVZKogpvBsXvg31YG9jvO/PouQj25Kw+pYg9
4VuXHo909spJfz9Iy7wR/8Z7vcHO+LAff9GQ0Fgza7RjDLkbmoF+gVYY2z4SzJ3f98O1OLzLstTk
RQK/0GUKSdcPmi9a8uyWgq6AHz2fbYQqbP90d6ux+/vI62SFMUXTu+1/PLQhKwIPgZjfzNgiwzqP
FmLlNHhKxdVKnMHwaObjFSU5iJaqa2UQHXxe4nJtYWPgI42vt6egiRoPfgtTv5DUF0eIBnGoMJY2
dHkR33cnGrJziD/3zDU82dTgJxV6SJiV29ypsAhP3o9EuE7PKEaYijHcycH7H461GSpfXwvPH0yd
eB35WBrdHika3MtPFr4AmekuhUHlyQFmI3lZWiIqWT6zVWP72RwsU2nQMBLtMWvsR+6KdANvuFun
S/N85BMhAuuzU2FamPEBPHGLYX1y4W99qMuPfqP6jqAlm98KxEwx05kWfZsQtdjWT57Vc+tK4Xhj
Fi91Ep8BPkg0ye+sbNa4ps0fXvQ5ZhJ6EcsY73rBC83lkNaSmkSs3PgBbZ4eOcAcexYvyzypy73z
k9DpNnNNE+nMrExs760Zlj04f2y01KS7aeio1wjkng8VvNVlx3pmexytJlx0/ohzsoLKkjEaji4a
dljlHADPh9zstD8/UjD5vOYbEP0HebubM8Uq/5ns4uyqeQ0/Lp9CjAMdbZSrq20GBIYpekWRXYQX
+FW2pufvkntV8Fh9QpOivb+2Rar7A5iVHdEmi2J8sTnTreDlpTRZwF+cgSo0UzSZiYAJgORpEfQW
Gcm0C2ogfSt5bf9uDrqc7lZG7aclxpbMlGjmARWda3GQ0q1IeUi6ENmWsif//gjeJOdHIYpwjvcd
w/UMz3RIFRGXYJ1uAYsfj65QY5qfq9x5tI6WrVL5wbv8Ig/ERvSUNULzu0SOzLoyE2hk8hnbPGUL
NJT7NPf6N5RX67nkuOnxZyQFQS8mO/dzVGoDny2sF3xt07G4WUXXAkp9HT3pwAbu9W9DY9YYhnxC
DREKN54F7nzqqDxYBEUEhqU/PzUE6uQy7HEimZtEFcYzkiRpo9Q4lDbPFfijR9nV8vWSn6Kirs9Z
rwfKDOfCvdnTaUIzskiGLeMhai2Ss+wl7T1747ILkYHIQbptzi6F2bMRejHzCTNPOxzXrHbOxACw
ne9Z71ipojiEZyDUWAAg1MdShnuxh4ahadJluBPl66p+dsGsNHH4g0DiTd2P5w4Noc1d3plXpKmM
fFK4dhesuJQUVMFYhEJQzYePeAcItnn5tgZMh/HLLddRErCPvtbiFNf9b5kM9UZZAl1xxtMqBlxH
RbLCNu2cFs9rhDhigZF9b1XxeGdyCJ0HYx/CVJmfvlX9wKufJ5sYjcKnloOBnHFg8vV5CPFXUbfy
SHkFaIwhXW8O6OHS44Elhfq1Jn2cX3BRASK7OOV1RHmWSuyQakAbpy359jJT32QyjY6tMMCs0AG0
x+9w2CHJJZkqnf99Ek6nfTcDmGX8sih0sw9NLGQ96BasbJ9k1bF0amgfFwp81nXe9f6sBS4ih8UZ
+wWH+E8v/WVkTLko7ezGGqU2J7BU/7DR3vDuVQiHpxMkbfzq+pvVBAnhuk9NFzoM0AVValB/Rzgt
2CTeGaw/GL3cQbADAXyeQvK6bDEwHdnUvmftCqj3D3ZPXHEvUfwC80CQHyRmuzjLDkGgXuDWh9bm
r8GEASMrEa1QcAE5w5lqjBnPYqI0Yu6Ykkrvh365/+6e7gzrXroz07Bg5wvTeO0vUxt+wy9LL81b
u5+7JcT6yZsY5DrN4XI6nPvGLreHpm+6btFzxjNyanjCXZUmRDALH3FIKg4pHK10Q1ONYctB2AlF
Djr8j/ifwyODNVWZ1ElgCAOqgwtkC/HUoinf8rV1vYHtbjKW1PGJ9hwM7qVrOMIiUvhzQM5aGtlC
15E7ChXu+jkqmXIepOIpqF9kYQszBIrSIFPfZmPsSqSZc4jiZQyWk/dFrAYWJjJlFxCUk2fA77rU
VNdAf3kPX3ljkjkZflE8hMctjFhXh/0L4IDeO7a79txcCptkUQPt5n41BXRpzjgQ7qL8IJ5hSBCS
kdg1qyNQjIRB4oerMgomK/fx1rMC21DDPSX8hdxym1W2hJLyAWQu+TOlx9gYIgSDjzHdC9KIaKxS
GeOrDqjxkTFjKDXaef7GIKGiHcX4EHKtvscqfkBdWz2rhCeo54Rw6avhNvlAr5j7upkDBqj2iRPD
9sstqzp7aDbYIOE+CeL5qQpV1Znt/uUVex54ASSORhYvKdZ7w01TlMDuA0fMegCTT6gPU4M+SoCX
8kvvOmFiyNDipulHlfEAMl6EN7mdQuSWeSK+HC6rvI8rGRkYbViZBsOTRIDW1KX3jg6RYnx4XccZ
X+CgovO7FhzLc1ddGJeCB+i/nvlCnbB+XuH00sUit2Smc5Fds7AkmqPo4WC+FY6Nx0HCsRT3YhpN
vwsd2QoaZZIhsueR29lRMCxVK3SoJ+2xru/hiWPSdOsSEnHKH7JJIZged12xDE+lqISDmTPv7CR9
TMD6CXAGTHM8NV8JfetspiAZiyrP28shbDqtyIuaclhKOsFwb+eiW1GAfa9LBdV62KN5VBweGK+c
J6hJVTjrUbJHQDiRsiRl41apiEkClcJcVsTI3ZUcWldIwlkWn63pw7lAhfD+R6RQLwgZkGNmov8A
+sCuqQGVEY7yzbzfkOWgoVNFMlV/P5WQADg6to5CcYCk1xHQb0LRBbbtG+XKszVS5juL34cKbf9y
3ejE98g4+ocBJH7LtonKeu15PbzDQSpOfW9khMU3Dm3pmckOgXqrl1eP6MmZyAeBtmAxq/8yCWnD
t3bRvxoSNkaj7/yQGjH6SP5HyNH+4CSeEl2ZBXGp/6jQWDsLTHeO8sdouXVX/TjTpqZBDPNk+vtl
fxCtTNR+z4s12ehV83tiyIS3VE9ElX8z9ncGnP5iqwvGPOrrlhcqClvY+RjKrAK3j74ttTxvpG7+
D8ew1hL/C1qOvp2+36dA/sCMyY5JqxwZvoKN9C/GjqYEkw42FSCBgA5Q0RT8v3oOw/GaxlkAVyWl
Wfd4tLaYM9vYLd3b1jlnV0tPPLuh2HWD6oyWuWjWwGKRv/+eufu43GT8z/X/KOfxA2ADbXyxV6x7
H1XWKOYthgAR4zygFJu88wqNKb5QuYD+U6FPhnOPyW2cIbYUE2095hpGrmjHJxhy9FhzcoYC9779
g1LA8obPorTIZXDRpv/KlT89SykeHPX1HsfmJrMhKU4xYvTiBCsLH9VSPx+ZDkDmfX49mVrc6mQs
lp8XkMVWN9f6sP1PjwLfJYZ6zE6kca0xSnoR2+sCZiXf0dzCSvzGBAXioL2rVtZOptFLRnLs4ghT
xG5xaWEA31bCUWhWxOO/ENeHKoyiQzxVGx4iZVUW2bkqL8qPnNvqlAT+YesqRof8VzOKPUGYINA0
uYltymCqXbfhKNS3H4O3t5p+OboDuZsuA8cdmQuUfRUq9hxrLPtA7eE++4FRwp9Sv5rluPOYBi+i
4Muxe4KnDA4Z0AB1sBM3u5FQUdu2penlsKJGFkQuH2nwLva5p72scuXTf1y5ULPtjKVwkD7aY5Fx
VxdwwmTLs2ETqOr4UVXbUQo9igaaVrmdlKQa9B39Xopw+yLVl+F9fA+HTJ/dFg6p65OpbLyV7b1b
YLrnSUBjqJhQwDF/kzkblNhIZC29/nmQNAiTKWU0/zDlO9ILbFUeW18pLZn68c2n3R0YjPxiIrPv
PT1e4CyM0mJGXMBMdTifhpb12PZ9oYlmRby8JuTAZluGcIXZ5/LwnatM61ioBvaf7Sp4Bna1KJoT
DEfgBvzBc29BjyN2+BKNfwescLbL5DN7oy3SBvhcqfm/tKNfj2DmBJ6lEkuRTWtp9/fW2PbDiT2l
Xyny+dGuCR8x7Z+L+iPbhxjXdrvLN+15hSF5ljIcFs+3aDQ+uw1E3ElkprqqjEcdHO7Qfcey1hth
4njZxldX4mMdmOLFZ5kGLq4N4mK+rvuTPQZ7ti6FljSqtnra9wbmdTNHJU0CI8CMdLii5lgKs1iZ
ZIG7hnNLQr/O72rYv3zOYzGGOUP8LNGSfIUhJ+H8aZnHjXFx4ORKNUwfnnD1wRhM0xAcH5BWk6IX
VRdSLQaG3ha2TbechSKAq7cc2N4BTUEYqMPQhXLn06aVrAX2w5EZmclAw/LZYc4vYtVm5yvb1l4p
6FaylWSzey85IZjy+X18ZorXRrZW4CfiYS0DraoqnXfkqe8w8CEW6R1PMCJxaOE2YJYXRXYERTzF
UmyluPoi0UjscFY1sP4zNb9dEaTUEUaaGpKAUTp9ZCioMJpTuuBn+f66Zq98+GsxymUH3dMYbt5q
Hl7FdV5uIuxEVlTnET46t1boJ+mSlyuhWhtyBSt+wvVOSzEpO9TYPDoOB14/zK69HxNeE/dlgiMd
C+GSWlM7b34547UEWvTgPEw9JG5YVzT0GXEW2i7/H+DfCleslhX1HyJF5nmIKKHwJ/jLKSokHjQ5
3O12iF3WannfSI8R4gLsLqDiNAUHO2z4KBlr4zHnkfIeybfcQ1LD0SgdJw55yVYDmQYovz1QuL6x
O8UlrClZ8JB4HGQN2RN8bbk5wKUgnErU8igOKfuPyutHSYCAofeGwGr6PlEkZED+ZxJuj+Pw3m7s
6DrAao4j3BVfuCYZSP376lJKQb0QFW3VqVOby2ngTBvalFh51y1a02bcbvkoJeyzQsbogwZKmJm5
i2am0bvzL+1Q6TosTe4Fkr1/EvKh103BBAPiUbzg/qW+Jgy5SHva1CzPlX3OfQOqJ9sz2K8ZwVD0
+vEFPAxkjU99ktdgXfQCi+6XH+FqShBLk858SItPgEh94Qyjx8QQRnO5rq5csc0ycvu9L8q/FcSQ
Q1DwYSD3xAzPgjFcT12JivRQm7RWc24rEG5q6oyztIOdvvccraihIssP9XyJOeYr7nB8m02uBOXa
Ex3/g5Rc36QmOcQHfC6C02W9vpXYdZP0zkqng/aY9ImX5CQvgf4nKg7f5EnBzx9QNkSN5cTKsBav
r/HtMhXTrs6P1V9o/iuzq0EvKXsKtiYzBshS7MPRKfgooUM+n9fuO2/0T+QwPYgjCTPn7VTwHESb
p3TfBCttCjEI2VnebY4nbmODhNv3qmkDojWj3BIXPSm4zDnFeZeNLrFyl6gbHQIKoUBD9e6geTtU
slMQWblBBDSb/roSVqB36ipxNak0Zmi47BtkczLF0gpPJ3AlOFcE4EgKG+ij8GkKWC+3w8JULgaz
Q7oZerZn7T9yJ+1165S4/ZxbdbeDcRED/RjpyJuDlLcBbjzRSKuhHxfJhKUwpMHnz2/9N6dDFDga
V8TTNjUTgwoGSarzbd4xDCpd/J8FJHM5pipLkqaZFTBsd413BPELqsr1cKgdgzbfUhPGK0VIjhIG
TUQVjHt4l+zhu725U09sveuXaPjShys/sKRBSx6gRSUDHNuUehpR8h58GM57BV005ixesdWzjxaU
MEVDXbCNwjTbHyKzKCj0JlgZnJYcB7VMcOPzTjhifHPkcXkvSGZhLMh4BBRRf81o/PGBSSs/+xPm
6jSKC+yGz/38mwItHE1RjkGjiOTFqOxYRCDTULhBRf9rS3WHwti5MB8aaVZeYH3PowYIrurAJHUC
CG0FZz06aquHUm1P4Dy0dYtQSr0+sQFO/ZJTzB880BeJRqeCqeMVRs2vzXyyTDo2gRw7j1ZqVOom
XFJkKruFQkF632KEAdb0z8WRYZzkZbxasgYT+TlPZ9Ux7l6SLy4aIDs++3QTEdbH1BxLQ86TrC48
z+abHrdPzVJLoATnsS/Heqiz3MLPzkb4XvWaL/B2nEhy0k+a0hu2c3VexDzJWAHRLuv9RafQhebB
AFRm0W01K4j273b1j+lg6G6I109R2EFeujeastKwZI9WdiCnVtmJ8VQXRVEgEZLQe7FqKr4clL3E
y3dMetcKSTrHiG1YZzG87EZUnacKxRujJDvZzDytS83ed3/X5L/OugKvCwroZl5s3xuxV2Cl9+SI
MxeDCWaQPlKrC6WTTR3MIuIpyBMUx4DSQURX0LDMkML9JAH17A7AzkXOozwCZ9F55M1vde1mVVRq
lvEg2wTs+l/ioVfW0VeUSaZ4q5iThohwFoyms5Y10/zZL1CGAXlN9PYLpuzkrG02EFPgNPejTNDW
lr0U43cJo3Aiv4K3qssToVJR9u9eJwpgpkQ4g6a84e+pjYx1OoRz9peU0vS7UsKX+7kZMvsJWrOW
cTKLN4Rb30nCJreqEqx08dPczuahLvG+1ItSKKIKcxjbJEgWYGDbBCTju4RHaehZd2ZnWrOzumF7
I5nOZLZWE+sMI0BI87UF7BkmLfXYZc4hHd7AL0UNXOpzUicUfgNAIerZ4rg0tAwvH09nSldt2T/A
vLc+v0tYUyjs8F05o64U/66tOgfJKcf/LZsp/RtjXRPLvjgyc9f9UW3bEMSJYyD6yXNt7RzRcyRu
waVyRcucc/rjEZiCAl//Bf6/60Mv3h0i9eJ6HeRrT0DnpFZeDjTnwuTqSawHcbDuEoJaFQl1SHUL
RRqdE+8o2slnwqpdNhva3JIBj6LFvmiopVGNZsLX28O09OqXlKoU2pBxngcYJFkRy0Hf/gGQGj00
mcjsyHbBOdivcm9B9hGeGqd/rUK1Jp02YV6J4DfJcScMnMWt3/UrNViA7gqZDYwZjrU1Cn3k2C/1
+57VnzySuvPm8z203I7gFBChRpuZxJYUNUi+yoLoh+Do0+h7QMS6CDkyIXl9XrvXTWeo+xN3lUoS
FDbc+IHcivDUtJy1e7kkxLQtsCKJeOsD49w3sIJD7WfylAOwkVo/C5oWAQ54LrH3KjmUFPxpY8/N
BK+sSBJOnBC3P5UD1xnX2k3jT0oUYrZdGKFad+qxbyy7LTZfDRuqMOQVMloxqphIUNR6M99GQfGE
YR1PDE6HtwrrMFP2wY2E1+UNRg/6EPzJS+zdaupwSmQ2+EmGfY5UXCwcTFlzBD1W0NUDtEc3W4NB
rNzZQXqTb74r7yxZuPQLgXtP3jkP7MjA8rn3qhzhGL6UxcIs4L8AXb8BJI4+s5gys9NWNTj/gjOM
h1jt1JdeW5Io/3CO/93ZfACMh306GpnTHylPOTkQA5n2SUBeMHDH1Q4xRPs22L8Iicv0z/JfMxvt
pHpPdXaTBIEr7EDX4gQ2ozpI2NzO8wWh0kZCnnjByBbh4oW/LlMfJyPihPShdLvqPuVMCqkrh6Ks
13qccbUZFTlVRm8GTlOtzH2LMCX3jTAfJkd6kSJS+2rvRZkSBlHQGjL6XfLM43Lq4mI168mEGC+a
MvUE2FEv8tQXcwGaP7heaHirTQgAYHtGXnT+sANb8Eyn338INXFaW62y3SUtlaxKSZcQIB1QkY4q
wkVGHdylMITSMek5I2p8fYZA9ivMdwNU7YABltSYMUvdMjJB6fhJyE3OVJMzf9/1ivRVCml+PrVd
g0CmrXgJ2IEYvfvTQUbY8OSpPFcVLUpoQrtF86EPegOpkXZgoPPqtvHdFAjhYghBTY1tmKFlqoZA
3+9tIV0ap6uTJpLUUQyypxUS8CgByzuGGkWHj5Uy6UFK5vi9Et0lWuPkx5G8YzXX1bJ7BkNh1Q2f
pc0MDiMN7nNTwn0qz8qh+EJccGv/4v4ojd2oI2FBF7YRuW4pkCTUnGQ/XvHMauKdpyUUh6SqncWW
g4+PVT8xHRP9Ss0Tk07ebl/rN9rNo7uSaoxDdbyqxhc2Cz+pvndIhKKAtO2XcqgwCe4/d+D9stRU
ZEtmk2pDCIDxQImi0F8XiWrzHh2rIsWClbrqm0A1Vzj8G9WiF2WviSUY91UWORYZbonC5q7MlxGo
GAAfWyKqxinTz+8NrXqcXwP6ckdWlMf9uz2MnJoEFeY47ordxPPbh0NtruDxWdzb7igREL0kh+cc
4RGRVxxgagA0ebPQ9bFAzh0PPBA1+SzQ3qnQdq+ed7PHv1YppAkN7xllvREn6hJdLmZG5GFATkj9
ufQaaFfghuDW22yO+coFdBryWzgDY4qZIf9u0+s7Z2BylQ0JSY20ShYvuAwfPsYhQZIbMXnELwo2
ye2j4VA4pxj0XVjnC4MrPoCpyhYn9X6JMSXNq6EOcGOZqXNTKAjSdl++ldHCz/I7SOn8lpU6q1+H
vt4Zs9d5iUZy17nXhnD/oqO7TJMY3Sq2XDVkj8d4dPZAPq6FchhPQSYNmlehPnhGKy94kookyvFG
7REWGwm8lO5tD1aI303VDHXKIWdVXrZvoXNXFXMTUSO/P1rPyuF6tTxQh66OZRa1uXrErno2fpNh
+TsHS3uLY0Sm4sFc0e9Ph6vustzdiRg6pRmQ0gNTvKiV9fLHlOO2jJeghALUcm3iNmk04JzeCEKX
p8VyG/VtGYF6lr6zKeX2/rZqDC7Hw4eVPdJylLwNJXRt5aUpLyFZxxiIYtHGAw2LVuxYHh7UKHun
ESlDJkOBRHk4mhtfDJTC1gYoo5YeqlnWm5CLEdkpnz2UEnQ+ZMjtzYtFUmYII75DlqQ2NXhxjGZk
VIWtfbMVKXnUC+yhkPdkZ+PSzErteuxDPgRi38xgxnyHbM+MbrSZ+Guw97MZesCTvB6d9r+gvJ+T
ikBaMv+lFwea2Tq16bj2UoxZkWF5wlXRR1yelMAQmd4QZDYyr74J9jbZrvB0jUpOpz04OHPguEVc
EeDf3QuiuYA6bPIT+YHwK/CAhEH+9xpiWTLIN4FHzHocmK1W5QHmpGCorwClxZU94sRUAO6H3us9
lVq37bTy9zkYPsaVm1JTTeXJ/iMgTLVBJY6ws/sFulLfIa0CjiFbOJ3Z/hsBEvuaoFYuUlGaoKAH
eXSInadmXA+aLCVPPTCSH1au+KnBupmcjoxro8n8JrW4lnRNlGsj48aEG1WBIaDs/fSANA+AKs0I
K2V/smxbvv7tCune1UZ1wCZ+MIxx388qHFamPKx1xuXUX6ICRbp42IJyBfSbi/8bs0gRIlfniyr9
MigZP2axFe5+3EESAvC67Aee9wL3S7LUXrN+hGVQxHb/q7RMpdr47/r0/geE9NA6XeBG4ITsP3fT
FXI5s34fDZMauG77oVStwf1HyxvuFfKJLkH6Ng8xl2aSuQpYJ6PKocim6T9DIwHdHST8HNWwwwMS
/+LBXSLhALd0MhYpd0IPGVbLFkCJC17jFlbhKNFJ5f4jQx9KqjoRzc8fMvEf3rtTkwnMKiOMr171
M8OuCC/B2p19BkH3g5aOnr9LBDhHPSCxIAdZRZp47bhdq8NKrGqRf2TGhYoYqbnWEm0/IeMFXK+d
CYcmV4nWsGFJH5JbszKPc9IVweHIscyzBLgv/4dnQIh6yQrMvKLTvZ8VVxuVBzpUkTuj9MJyMR1M
MmBfNGZCr/XfzCCy+EQdMe5WMx+rKiYuyHyp6QYhwVvf6UZSVzLngNTAgxUAhMrHyr/ppd1USn4B
nj8PUNwEgcB2r5J8F0d8Y09xF5A1uM9ubtvDA3EyzwWgge0LXi8WFyNSTAaqYmv8tA+VX7Pms7j9
47IRPfRrpqSZt9gGWpZj1JFyfbFXob8yTfGN2NRaRo5Bayghz+Gfy0/ddPMAaOEgU/DsBvhqvaHM
v/KEaS9hRUabq5EH138bIY5kFHj28f9JKCqP0//b2BSghz2zW5s1oW1oqzCoNC0T8MyWU5VJ3fC6
JogVI53q/ZwFlhJ2HN9nBLW2PKKRInq6TXvzgNFQYWPkm6+ytuy+nMEs8hRz9dXQHlykTYP+PZXA
kDxNnkGisqX7HAXevgCEfdllcUBZjlX0b6oOsyo4+AvqXtT5Sgh4KorSjA4G1KB793T+87x2nQgQ
fTTZJ4uI2JxUN9PfAYTLUtxk5mhlx4EYcCV6w5d+mYB7EahIqejqyIPg31itW8HGW+jrq/cf6oKf
PUPI+ZwZannsNK0pMkWjh+QFH3NRU/dIJk/F39kqM74dCpPjQZ0pucnV8kt3QWELNidwoLgf/0t0
hlQlK01bKf0Mf4QcKYhzuymltXuuJ8IGcbCdOdC2MKv+q67iMlUF0/ymhfawROun+O4VCfqxdc2K
Rtxe03cd6+tlXrIOkLV5kfEulrABaVjFuB/IKGRxKIQeNTyGyNakfgcBIv9oRJK/s5IXPuRGgvJn
zzu0ZgETCr7rgbrjMmWLuEe9BSsruiMUicapd8cqQSoU484YBWuafuV1pE0OjEaYpsO8BTvpiMFT
GUAmTrTKjzw7eAFZFesey+sbe4GfXO5pTKMmrs+4rtTWkVEdu7kZVHgmFS0Rk9v9Z+alq0efZ8BO
cgDxawoM8AswKC/P9CvSebeEupVvnu5zfxYmJ95vyZ7Yt8S/O0lDvVFYwwLCbeYeb8FqBJMMJntt
qUqCLbznXOOVE5r/0OsKjNHm1GfJDm8hOukku6frm7ZACQ7jlJXBjEzyCksbj9nRM+UMZC5+ypJm
aP9RQred6WmoCY3rISIupTAnpQWMS/kfajrpZnbNDSal5wpU6rnY9gJABx4muPY+NtCOXeO3YUjz
p5a7IBl49fYd+OmN3eAAMHLef+VPackRAkME5DmWnUTBeML50xP6BYFNxPgVcGrkO/OK7xMIJJC/
l0JYs+f+MhchOKB4h2y10Pvl9upzGdo8+kCrobQ5jX6Ihd6yydoKbMncEoSF/2bEBEZLYy9Fdmbw
kF8QL4Ac1ASx0EzPzsKqe2KmzUMM9wEQXiwLkCYuwqaF0lD3fs9Zi4NTRrc8DCvoKXqzFowstDni
panIcy0/frfglfSsR5iphRW9g0Hvwc4gMvEcjYqjwPn8+RJpF9Xk1JU5I5etuiZh+wDIzx/CGBWI
9etmPd9IOB3pHohk8bIDqjtS5hSAcaoaOgYR8kqwmfnXGIdXYjWUDkkiOOByTAQyC2+NZrPT8CxV
xNQEajavJ86RQ+Wg4r3tDh/TyHVIMnlfX4UOvTr3ZUBw6mD2DEO/Eq+8k5/y/2VCGl9L55K7ycvT
+QorAPa+MylwRIyfvPtRFcnJukpTU2pi19U7wA1dPIVW2n9wuSBypE/CHv/rIsmQK9XrKCbWbyfS
cWzasIYmwjyl1B1HqVz8L3nPh3VWzySmXfKWSB8p5Bl+/2cq6+saVnUl7jkX4CfU3TG0IDJnpIXW
h/A2hPKHIT4Bj/RfMGffpE+vuN8AHcTu/LPdACjZ1UFJzeEKYW5uX8t2SKYZTcOxsS5tO4TCBjTV
ZIlTk+R0g9EurrqM+py9rV7BvGSftwtSEbFO+jC/w2LAZfmUKUyPta/QtYN3caNySg/DEao9XxS6
5ENQlsTk9TiZRx2j1oIhGHezG9KIE3uHj8vaSy084nKRDjZNMWKWoSgfxLrnhFprPpHV1402yAo9
Esd8ulx7mQlt9lesi2iavKku0fH6Y9mn1St6F8MXPbRfQcbcDXrELavKKeYm0XBHGklz12z9H6zy
0v9Mvx2SztfPX2uKCG+11Xr4MP1w6FK3/8y40aLGy5Ah2JE7ZqsYNhAmdUv8HXskHJxlaVhTNKWC
Qpe7E9qh+H55ljbKOCVp//+ghhWvhPp8Vs3AO8mJ/CFYSpJUjtJx43bKLxW27NWkIIKWXw5ySM08
XdNq9p5ipGYiMHZ41JBfMrhRGyCWlUPzDGFkEECenUdx8ZShUtMrfMqoK7dHPXlxcrEw2vjRv8xW
rbl8hn8SgfPYVeTyorwUvikw20JpAUzTKUEp8MHyX92VmUVXrJp3hkHegsbA+UzwOB/janUZOm+m
/8N6NqL8RSWpSCyrcuBJq+hsVmbUYieLh+wR2qsc8zjbEAqviUxEJq1KiViMp6wb/2WFFfTPNpuQ
Bxk1Tc5+6nBjM86nLGzjTVPWrpukNnZmes0dy8t/7yeQomeOhifYK0LlbgsZLuTxiLwQoKgO7xqK
LZ+mGNl6aH/HVaYsLAxnOZPT80p9NJKomz/tNZCia3NuKmR1xSkblzoS1lljAYYt+jkxH3sjXoKa
aeOn364Y0yLcUBF5O3mm043HFaMbGw9Mi4fsFu1Zry0PEGTfzILDgO7ytC0gCIUzCj66m8hJdtWN
F7aHxgvQRGTNCxDoEvg5Gdtd8hPdH/sRq7VrGt2Byps1TYdy7w4MTIbGzDp6cLQoyu55UxTNdvRx
l2PL/FOQGYlvqQeMBQY+Xh/6UDuy0lc+t8a5oe9qO27GS8S/VqaTMYowES8CtMr+EVpebHCoD2pq
nQJS3amyea593mVEYJgNdoUYR/pABQauIkY33+X4l1bIA0s0NWmHq1spkfUp/mnu5c8InUyzE82X
dl+gwZwUL6e4QNrLroI5LdXMe/Cknd53fWGMIWMj24MgqkMrGIaFpn9c++51cVVHkXG59omu7st+
rmvXhD7qXJ72iK+1x0+GF/xT9p2pJgSmS8y17oybByRDFoeTVVFDu0G2OB8/TMhJhcnvin+NEF8w
JE1NrXYwiLS3WhjD7aBNHftJzkqgszwSTiyu3kSe0bxptQR1wZB3UUi/bYXts6zrI5KajyjR348/
ZK5YfFsYCIylNeRAWtnwRrhJk+gsxAbkT1ABewVtFGPhKlDwj6KNefNKcNG3mn1knHARYTFVQ7XR
/jN7UBC2C1Z9JnplXQCXWSIsGlAUHjd7FvmjTl3H4tDjaHRBQk/eVznebHVMGd28UEqIPdWmPtFF
l6u6WoyovX3Z4Sqsji2wqbFZTwsDowePAMXVVU219Uez21tcvy2faHl46nIrK7uZL5SlPvw3rVmM
7sUmhPKgpWL5pY71vKRzrsQB+gZecNZwm7+1FzLwXncMJmN+ogi2gDDf6VXiz1P03+Fp1jIZchJZ
NGuXMcfMHut0MqXjfq+mlrkJZ0oIVgJg20/liJVKNDPEcVur3IquozKfEm0M0WwN637AT91xzryd
L/6ekOz145EDc460wtLvAdZAHBIgS3SwCS6OYB6//Z88SoyjW/NWifacb7lc5DLov5PX8VcHtivG
pQeg4qH18Iphrp5uDyAsfHIW/tht7qzH5ZtqkBnrdHQfsN6DRhDQZcfO0/b6JPakqy2H8L7lZsbR
TTWs5P/ZIbtTJt4dQNEtUay8HE8IHti4vb+/vuf4RSTC4+01Y9ej8LsqG5QLLXnzBggs3mtrMio2
9ZnXbMrGZZPfxASGI1k/8h+twexCQaJwvsEYGPEkPF2rpvnrYToYcmABciGuCS0Ggn9w4RSuLI/C
Sbjs7tfOFyvWjZU+klP8wi5bry358MBwbuNNn0aBsuYKtzRsTpp9mTfhV+uMhRuzwP0RAXXt1tCI
mWoL1wdvmvPJnvWvS54fbBc0R7f/c+wxgG7HyOWgdlPL7WY4NX9cuBFQbtH2x46/WGx4G0+jkCla
6wmbFefH+YYtZCxNfV5yOgCXlbqcOrT1rPKbGTPMV8Ev9VOf6Yqtx54rfiRq3JShzjxbMX8ylpko
cWwcumzx8HN0Tt8m3GQn9IgbvDkQtolSAHJScNXcBYd7RS1MS9s0VCn6535NFFANpaeFcPdVxR5e
Vb7D2EVEKM3bDsVz7pjswH9HIxVU8gH1m36GLOCqUiSpsiK97xDLD6Xe+MV1Mwgo5BfLpxf4OdsK
1Egel0VZoYfdRlp2b6zlIteh3GEijvQexYZswu7Db9p+PEOkKq96kTfAiG7ruwuWypBOzxfrRrNa
Tk/Euw1KdmYTzPgeklIkr5quSH/15na+b/ryBjuFEfRmMTyd4TCctEXi+UOX2RDIUe6UpaoE4OgI
LYH7gr00iz8tpVXzAqZxcVKc35s3vBxeTggdvnDlHPGQEt5KVrvAEy98cwyQW20VrEyHMvQcgTw3
yWk/+0EmIGwKPrWivykI4BwFPxuypbTG7JBX+RVbGpHnsOQvHFankcuTLUNyckPybog771HOACYA
fNIeCos7wMRVpMZ3lo+CeSu8XSfVIu5Y3s8kQktJLEdhtZDlBGHYN3iLfC5HvDIiLe6eJdVaTIg5
/HFHAviq78seBv7pH0e1/JQcbmO5Ww6GEwuRHET4vpHK/c1mNT7VeWWxuBPGi4zVtJtoMgiOafzv
o5zsdM3j3eu8+H+M/FN1j4dD/bLOoxOXUQF0dIWtCVOJ1JttQBtqpbcgMs8ZDD29JRTT+EM7GdD2
wWJTfUYyKGn+IR4mflfynNkreG4cAy8dmU620Z1i850Y6CRzgMQBnMQGNT9LYhmo2KydjVgq4IKn
EPIsKp/Xp6RSEJnjRpbGRFnnQAO0MexjFD8VItRCVj+qNrMQD+tEvVUXuPMxv2z3xi9qiqhICT3V
OfSPdgEZ8yGp/kLToMEmN1niygseN8wlxuOULH6YfldnPitdej0OJttT8x/91absWCyQ3qCFC8Zm
PVAtGzQhditX9Espcrhid1LJfFp41yk1GDTvNXBjoPxeLMBTmuDKwLqHOQ58JotcDp0LHpe4x4xi
wi3Tz1+DWMgRY0+Or0+Y8vvt0PJBQfhbn3l5mgTR4EV7Vj6FpM+I8+BO2x+o8ZEiDh6gXIBcKjV9
l5sfrbPW4ASXE+ZxAxbOHSqlBHUSz5qxxcKnbNU8td4KHizWI+661RaZGc9rkfUQqGiXZmEtvjMj
2gLOYnK0sW4PVINquBd/ACIUPqoBtBzyn1PNSy10exmww8rjIipBBtfa7FvYQx3LCgtH+IJ5ZaGz
EGf0FH/gxEv/geA1GyzmTl5oSMNMJAzuadVqFLiqYFjUiM0OjkB0gqBrG5VUsvhuZiwt1BJY/Y6/
/cQRroQZv526kpziRmrCuzR1CYbDL9Eo/JkVt3aIHokxYalGFb6Jn3l/JG94RcWAgfIqwkqn3zvL
uMINRzGoy5Am8gISh+KuY0Ps2OSfjOr24N8Lg2z52YALmgiqcBBbmzk/3CDHlodytcE6wJEM6YVM
TFy+53w/SeIWoChtcuxVvatEbRoH2CXSghSd1TrXOuvGZzdoJrY/Aiiu6sF5hT5Ft5qtn6iUUs3z
fmrJvEvRYVelDMwt65Vu8Tlg7CjhHKUTQuFkNOuGcXZz+eqmIJIlXmJ+DTS453iIPVbyRH1icA4d
7oBjJLPuRU5oiaN1MKlTUEVhexNVXoD5KbM/KBuCos76muK/CUOwpIoRfKovzpiqarhwHxi/WHqU
29rWK3j22K17Na4EbeUQMZSYybEZCL+yNyMs16LduX3Gtd60siGbEfsOZbV4KL/qhQ+zt2pTZHnV
iDJ2QTND69KrwMsFwh6aS534wnoirCdg2k2Fxs++Q/XGNi4t3Ff41xF4oPnosKrxd2VyPnUJt70v
BmVIqPj1RpUUoKeFfV3z5knfizQTrAQLozMjMU75jW9dpaFvXjw+kl1ytYfb2HiVGx++fDxRWP+G
JpeIgozmmmvGMBjE/osQZJ90y40yBCFzBS1dLMdBdH0chRM5JT+8ISMTqUepef2N1zyRrtWro+E8
Xiy/bl/iov7SgjLydY+ef5RZwf9uprbtZSoyQSztz/j6Ix+iizxErH/q16MjggDec4pa6WFjy5vh
SZQPeHqR6VSuc6n1KCM8CYgVRt9HHLAZbp87CZ1RvUYgvb1JjTGPFDspTFFjFAoM+D8KtmyC0d9M
dTKHpQAdWfTzoJ0wNHld+bVnxYvv00Pi+DVtW6uKfeaXFnUEGzi5i4AJkuFu+/okj/Rro/b4NNo5
9xFwVVWs83Mgr+kDJwcoNBjJ6Wv+U+t+ITkMYdFIvsgO8DjhkMId+9HrCkhn8KFEGu+j5pE0ovF5
lBaEU/JRM4sYU91FRy2MCpGaqn8l/NVBaOpm3IBhvbw9BL/zXK8hAdeMfephaqazud8K5KflHNTE
uAmEkJkY4O0UTzj9hA9lSFhkB9FLLEUuJ04QFFPB21FUDYruk69NOIjW6WRtuFIS9qyHBM02AGhA
UyNSGAGuF5IGGKubD+g51FK3DPUa/rCEX6BwyShGG944scenQw3XWTVKdoeog3FQmEA+Bty9vAMs
7Xva87C/1ABhn2ZTzhiiUMrQ0WlUpSKRrJEGKuI9tcOiGYMrGwItHZ6xghN0B8YxjB4Hyo/9NpXv
yLpHEUGxY2v3P4Bdb45Llz3Ameer/MTJQ6bPXs2zuxZ4Ms3VI/2+df7gDVBBSHXhgy9LVHyZxdNr
0BN/rLcnw8FdLyYgy2lroyJ0SNrUq0fXC6JnH6crKT1/Sv0Js7z9A0vmsONo7hQbfX1z9bvfoMO9
SwmH8BP3UZWhAkuVAsymtbmPDBFX0LPJx7ZHrSpuw5erpLrNBqssfvq1mqTZx5ZlIjmeVft5EnFu
v3PBdRKQ+aGRbKsCrc8XpBShiKb/ZEKf1oZdGY6WiA2dPkWJVuacmHfW18OnpTsxERLmXIblxMk/
cypeoagpepqK4jWGB9jHfRVKZ2pc31i8ioyxIgk1IKhuESRS3LFFtfR+uEYcyFAB9Jq7q0wGBzov
4CyDnDzmITkox8V4tiVeGlitIDmQvfq4Yv6rBeFiKuPx+AYGvoc5ROEhYUKDqzKkSCxCRpIDu3bq
95gcdtZeYBB8h50Afnsm/YwU6HQpjgd1w07jzCRZ7EkUkrGQUqVo177SEG+j2paa20w7PycksA35
RT758+n2eUGOz5i9AdAq5hnDgvaNnapHGnL6nbDDOTG7/tcp2diJexgvDOxvGUiePfW7CxchECGE
sRPQ5/XwUoaMpiSg4zLZZ7AUrqpfRShpJ2Z3VHmT0L4B+2EGDiIf8TIDHRh0Hfcu+lT3z2X13+Ya
QrbIrcGoL92GW5PWasbW1I81OyWcQ4RE5JycZGJsRK47JQfsKNItNbTZazOSw6zKZVgufL27jbBZ
tVTQ0An3RSNemhC76UCs89aylHBKbuh3AGXyHHpaT9dm9aV8H7oU27GDe5I1Dp6yHODClLcWRd20
aUgGsqLm2NzlU1uknxgvBVeUlfB01WvCXYNbyBR7wjCgH/xMnLgGLBxw03YpbTiDHElIGfn/lqy4
qarsoKiFaX41v625DTnvnfOsq6rDBXvi/JaF4pxX64tSH/7Oe3wGAH93V/2GGkCKBqM2x925EoKC
D2RpPTiHqi0xOZy2rl2f0rZXFE0U9QnErIexa7TF3JDXbsAj3ypzW6J9WcSpxBT9MKS5TjXa9eRO
XkRkl/4FvNpEXJOr8FCRptfa4JKOiViUFm/9C5qGYtFFUbzkNfXqKi3rIyFPZatoxKBORDwGB/Qw
aheZ+J88GOZoiMynjtBeIw8mTYBknBNy9C5cCyTcw4q9Ab82OVZPScc1aE5zFrmY7TrdjunTIz+0
YMyHAPmd6jji/0dlsT7V3NLtYRaIEwu6IcBQCwC2OUkPcOB2PrzWkpNbHnoXTuGnSa+8bS9XfuFq
aw7VQBtfO6kX51+ErsAcMKBM5PA7DRf0dCYjDBlpie9TQNgimXEp4qZ1nq0M+MbGqwiwZuoNx+sy
QEzSx5wUJPCix8eankXkPsSG8iCuSI0kRIQAwNgpGUv5F8WrIMD0IssVUTUyrV+lUigEEiJ7w28r
4s3tYvL5E6jqxBh93BKkjt2QJkUS39lf9HjWaJIikGzus1zekar2Pfjc/17QWms4iNO3563ws4TO
nPcak+dguA3g5jo/lAUVF0cghm0RhGHkxMy4hf3/BDMclMe+O0FRsLDg7mU94KmDMeJ0Xcb3s5tQ
stRhmG4N8B/eub916GFgacwWKdPjd5avgYAp1+IVZ7wGZWw0jdvAhX27vFiT++qVFtEEj8PUXk06
6J8q3YGC3ZHiDH/7MdzPmUWWLr/npZpgXf2gCECZHDw+Xou+srTaE5d/jjBNwl/6mjVZNxBZyVDg
Tu4GDFYAroKIIfD3nnzSKrcuYQnHs1nnd0SFzXjn36XbzGUNaXmYZLe0iZeyuClySxr3imBAVtQO
XRKJ8C3TrESo65Y6sGNCDV6xzHL28VY2WZ6qipw9KY1lTIDgm3a2rvGL1Bo/q8Llx//ZJCffWy4/
C68F66avVykHakroQVfSq1dJdetJIZZtXpsrrKQ83ZKLzMu0Ri+xIBn3d+5RaLdV9/we11XZTJ2K
cV9DgnF0jWVVSS4UUSlJJpSOBFpYF2DXz7PlMkKv6EPnpMNZVZln8fqGX2KoUIR17vt742o7ruAd
lsV0mfUndchUiVrkmNG2JYbxZ39cAlOCV+msN38c0g4l417ASqICn9zyDezVxfsSpDQ2SVjovuu6
dOU0KTI+AQZzUdkFGhJ9IH1TagARBt5tSv/IJZl396qZlUAmj/9j7eo8AIOTSheYII/Eb4D9hV2E
EBm/1/nigeeUBxxxez6BeKo0fQUPd17d4wE1nMd5i+MP49BQSqitNoIT9Ci8oPwOEuK9d5nFg0QO
SAMndnOmBGYXGqbSi3jWfsxxc6B08/L1mohl33gp6kWA028kmxjO+vQXWaxtIwcxOO594aI6zQ4y
218Hwf2LtnO43/IywpBHjqHgta9Y8L6x0C4LppJj9xzr51dZ6Mw/n8HOfoAgeYHVtKjTGRnvYbV+
cJAhs6TWVsc6E0tynhp8PdpB//OHeFBAhdeTJjT/gj9ZDpkS6mRGQrvzWSioh7B5MFl5kQoD9K/w
DgecfIGMaFEGD7yFhDN+PMZQwbfT/eZx1PKPH8DMf+W9ndgg6DDclTihQAPRp9+b2fIK4E/NW+/n
Un5NzDf7XLQ8YaulzgOACG8YMJbk2rOmTxfkahWVwV8UmXNzJQXZyUb0Ft8pRuYVPYjTuC2sKqOr
cupjj9VFFSeTCDlKWlldfBqwtNkF2YqzsxOGGbbcja7cBrbZxZCjNpPLr21WuqeavtQ0IgbmLleG
DtfVFZ9Pb5ikqspOZb2Vvl6XiaCiREbCB+huy3/RbA9wWWGq+5XuR7szvOWs9rpOzE0Y65cNL69t
+eGZ9/YT7PqbXAU4R0QK6u+C3xhn38rcJ9r7HknhmxbZlLajTTYO2Y0xEtVrJB3RewXngrwd/l9g
8xEPQ5ONc6uaLVS4lB+AX6aRYsm1YZIgzkdi4z/IPDfsiXgYwgfXrPJD0rLlHJUwK+ttKMRchJEV
41p3jURRNRQl+ikSNL4P+oQ89bQKjvqFCkpKgxbAvRKtJ9DE+BVALXn9AMLo2Zo9mxGgLUfK2NJu
2pKVHcd1BMFJsGyoL3/7YqM+dUNVNzGLW1BDGkEhDH2z5Qo9OnqzUJsFfz7JLrb/MSS3cWLW9s3R
Dc4nx+g3AB4BVdgeEITdUtoAbr2TSscER+yn5TXejrkd/xTwLKTWiaHtoRMaQYBlSeOklHM1Wugu
ZFUbnn/cDfoKGE93Qi0bf4ju4MK1dPKzdy5UDzzyl+QGDcISEQyL0PhnK9xpNRtE5vbLQVP9jZlu
bHWKh3CV9mQK8Qcz1Yv23AYj7cMUctk/7jBt2Y4wVxFkFZgDRw+mh5bg3fdD2X07SYgI7S7AEjUR
ArNSwEUnMRLQQhRssq16Xeb8dcyUA5VvAck34eXsndM2PqvUKXWPaJontXNfc7tUhGlmXGDq19m4
qW02N5XtZS++dxyrtNbvuu0cZ5IoUdlDWHaEGUTxX4vaCSyAOZpky1Qr2ZXDGq+Rar/rRqO058cy
a6hkz0CJ4WnaXf7pCWdHaE2ZkqaiKrxvcMmmNZK40lrUVheipSzJH6Ltz8mpK/OXTpXJyijTqakG
esxTEBVOkU06vaO8nnF+rCgi8uUVOjqUYWVTGT/jSocRsCsWGEDtCKioooqz4XT897I8jgKOor8I
sbpZj1fOAphFfJdXThmgFeLLOjgbA/6MlOWOGriP0d4NjS0fIhVMbjgOoHWs2MFrJMjAsAmDa2OD
kjgvp0SHHof/fzXa5sJxssDrSBTeIpbkLMFwidB6VFf86AprOXruEoItEV3bhixThNd24Hq5KXjl
ga8Kt0ee1qJIVeBzzs0Ikqunbt7WYuCulOxIHr1uCwwopTMkSVNdlv709Il4RIOhWdjIP5+xMKwu
DPwyjiD6q5ckMhH0xHpR1pnxFX5UnwuyvTbyxHh9U56TC+hIPhXoqSk/sJOInm7Sx26s7/uxec1b
gk5+47o/XVpTLuzjztL6GeuqX/rEHHPsOiJ1Doq4yWVzXog8hpIhsis6/zZCmlLD2fzpiu5dBJW1
zb730QxykBDKKQ45YF7UbiPLVAYBOzvEBn8ee5NNwExVm8nuTfO+WVNmVa4NfK3+M+kNeLxjqrj6
gipqYIIyrEf06qI13yo5A63xvpcA/9DCQW2JzBdh6Nh2wKu36RBorX1Y9BCWY66Dh1hW2cm/vE+G
jvlURrhMz1BiKzQBc6ByVpceFgjwdMSUkPjCnpjCmkXEcW/IeFSj+w1P722jLee+rrpesI9ATkGX
yExd9RaHHBzdlJd0n04S3pkG9vl6p8CFg3fww8jQt8SEaIKI+CGUFFXEmEy4MuZZ2BcNlax26bTq
/QyLjI0YwjLBSvE2/2hGj/rnyvoJiuUAaByPBpGQnkscbZYAbtN2330STQeoI7Z0w5mIWWRNBXRY
687Yj2CXQvL33Of5YKdn1lyf+XLs2VSgwJh+4s8OsuR6jIOSj0V/rTl6zA+eyW+xhBit/SOhTuFD
GZ+5781AFoPAYt6KKU7IhDE5vxAli10loYCa2IIs3Fj116eA83GOdPPXnR3xkD/eNY36j+Wldt0h
nEyNS+uT202yBs/BJ3AsDS6E4dGBtS6i6HMzAi7RsncDJorChGuTasYVdizFUk4oQCfVHHinPXGE
0orbVfwEO+h1xLx9dGQq0XSxzd/+rSHlRDp6zjS0WTQypjw4dQ0qoycPc3mXaID3/5a2qTOBjfXe
YdX6LN5G7s3hx5fyhNBJUC+uQTE77rfSkz10vSMYYqgHUmMLXFkmvybQlSxrC+FLvE3j5Uz6x235
W+TMYnsHPmbtt1/fxdjalBlKF85ndxy3KW05hbtzUtG8Pxt9W4h6TUeBbxzY2eufnhG0sKKZi4M5
bPfbJ2WJ5NpfhblA/Px/EIUGAiSV7cs7/Pz1avPaQJ5422sDcV0laA83WJF0G70NX7pb6yhlgH7M
oOx67JRamT6osQrIfvcZnbeDDS7GQiEKWG8cZwwvXQ0c+uy56nPVPLKgh5GUDcyhg8oSO8AqsL8T
9AJZaSSIJPRNRGx+yk/5hccst6BO7QGiClNSZQJf+vKLzKeAiwkAGgeVCqda1+PyF8HXlyuhsE2L
6b2N3ZDPVjZQQmBVzXIkX0TCSse2fR/DJibPVRhAi1NEJWNv1hncPzgQkcGb0GHkkJ3vR92hIfTM
ixYvRni0N3/3mZasP08njxPFpNa3vRQvltTitHsBgFJ5P06BdNxc305dM0d5McxlWl4Rb/7JbZP7
CdX9cuBC0VUGQ3O8mbmLkwi7Jo+TgUV65aIDzbjEEI+i/qMvc9LJYdUjGmXFGNHITE6WrdYHNGuL
fjyEBbnsbFT4z1KKJ/MHXZ8LBZ9v6SVJHSzHeJJ4HzWr1Dae0YpfU1/zKklz8+n1RuJTBR20wIIP
zVaNdboZ4EVrNydBej5Pphfw0qUFfZGG/Bwespni7Y2kCu1afvFHNyF1UisXOsRuGBxPTz4jgkRZ
SQZKPHIns+P6/skSbYJg89syLLxBrlEfaUv9X9W4lQFnXU3V7ahRAlWksAR78YnsIe2xBHXXYWb+
lPdqjMUMMviQBSzG5w9T8pLjkEjEN8n2ry8s47yMWaW7nS58lC6ZsixYk5T4V35JKfW5h0fbEKSM
GKQcH7hKhLRzBcfqaa15SgzlllMqUWzUpASWemfgyo6fBGbUilOyAtejPU0MMRklMZd+8IkGY/Tq
nZmdSQE5TIwOve/SZSzZQb5fkpVnc2QPgBSAGSQQgsfrmr7NCHKDAU6BSiBv3ZGwG2Wdwam6MPpq
+xqAngqWgeIZYDjiXFdC3D7mKLWEkn97AqsZTslC6dSHuN/t8SMYH2Shb79LQbbwYhcznD+OAy6R
X/JG6bZQwxuI6CFE+3n6sSyWbocrSNIzlMBWcSAUvo4w1AKqZ4n6p5Sjv7Tk+DI1RST1N2mCfGib
wryM/aJ+L5cr00Akyo4RJAzxWmpuGMBGYOVJTxxZ09HVAkZkxTHoGwuK11Z/Lxvhl+jAFu5LSY2T
cI+5srS4WEPtrd2Xi9BZsVZT4n7iQfFgsW2KRAmRGuPOcaeuUX8+wmV1pp9KYoHPA0B1+EgMt7bj
StFvRFLGJUftL0oZuup/HeDPTzO1jzeGwEJGCJSyi7CfzdRhdZBsd7PwFYcFKUWHMvEXMI7p6kT7
sY6Rg7/MOj1xgsL0QPs+1Mj6V3EdmYqaSGQaGvNvGL8nvmxX8cHT56bH9gwdRUuiCxDTLCefYg3e
Biyfsq+42gopZJCbeydNsWT2ndcXNIRY/Vz7bv8l3CVgoWJwMvcY3k/wfwnoN0zvgFxskzKq5JhG
YfB+5MJGyVQFX4HmYYOj07vCtKVylpwLhucvSPbXsqoHgIRRhDzFg9rYp4H8ZJ1OXziYYxb4W92w
+cl+o3Xk1PBxwjR2P+yhXuPyz/PFodaYWb9LRjxkJacOHbeePvAEQ2RTWFomD7sAaTkjoqd3eo/x
xqd7zUXkcrpnjrfvG6Evltfzs9gQ5+aDDOh02D0d8gjVQTIP7K5XaD1DNM/aL9bCYTKvvjIBQBKZ
gwvZpT209jf/gN9FVcD4FfSpeQQYXMQvPqQ70JAYZm+jDs32yL/j2ifgOuGDWCDXTBgC1nV3fFEj
zihHMCLmyT98THSWKKV0X1ThXILsgGffpdRY7KmchuFFIuOymqAvsGPk2NHgBNueGU9wtji7KmBw
i5u8ism8XqaYkfiQY2iuclTmzStxox0uYbD89ws6ZSOH0Mqxcj2EcwASaMF9Ff7OyLBJIi+kyhWQ
9Kln1c0soz4oa8OvrGm1fMtKn9+NJ2Nt5zHW+PLJxcN3gp/vI0ijAWVb1sC0gHxxpw03dF5V7wkw
EtZO0DXQ8U5L4xCuSMc9u2TgOMHQiRkE6g1+fw/ykcz58DTticHi1GfnVXlQ6FdOkyT+gGhCwlHS
fxxOZaJ0y7U/oAP2ntSZjfDUxq5gbt2/27T/FsHmTEFVZp5aRYbUidRFJChuBcOi5u0cGe7qnpNI
1pc7x80qLIeWaw+k+MtAAuC3Npw1pk8Wo8mxNybeU7mSQCu5JlLWlmoaYRYdO9wlKuxSndUknmKi
CqeZchB4Co5NouOZWRy53Yec+tF4JGJHWuES7LSkkzj89IiQFLphBvAtLyfbrgLJfhFq+uj4yGd2
Ss+HQ3RU9BpQWOXuEzJ/Gk6Ena2djbf/jst+GptBcAn+BSCTFqcwjHGtSQ/klYo/3H18drW4knQo
tLcbDgFi/nDoJGMmnU50pZRW3RUiGDOb9xRL4KGwVMD8dL53OiFzgoNOunLZ4pkhgngO62mADbhw
QJzfQktWISUjkylVtz5MY0c/6mpV2wuud/Zj7TXc8PfisC+zg8dS/1Dou2VlxWbDNSjjxd8lIpwO
ZGRxV5Ww02q2P/F3BRTfa+vQzsMRwoXYuGjYhfWjdCpdoQK/3o2rlFclvSFPDyqifuzKnsHp6mnV
gROQ9CxCv4DEb5zgUm3DxapLLpO0SlUoIv4yBFZpoHj9TTb/CmKaIDh3FqZs0wsAS3VVmyqna01S
z9uBnHbp/QBwTweX/sr2okQ6T4Eqkf1FDOOCsKIs7w5pN/3N7oK0xB0DZDXRXv4SgizD/rM0yv/q
I3KqZEjJUmzeMjtiULXhVfcBEvLfMRFapUKb3/vjfOFrOMZ1inXtHYW7UBOa67WGYXuaGNct7lST
xrSDiEI/jl5qrZ9yChcrygQgXLtTZFoqF1yhvLnN+nj/EhoirWnCKmNW9Pvu65W2MVhBluckOktq
xXOkGSXRslmaUEBMADMIRExRuuWzpNhEgEPLnMWD8WaALfVy/SHg5PbRiwx57P0TC3UyC1qsvRqR
8JQ9i9rjoHWpqeR/BipeKfrKCF66uLAaZ0T7l00eXdMIkpqFA7ybi/BwiplxTAb/FuhTc7pxM00V
3F9FiNWhP8lgwbz3PPHnkQ+tEoxMBhxX9BBFXHTBEk6MvMUwn3JhOsThpv/OTNyQWXc2L8hZAF7b
8K7X1mw0hZbMbd8Qm2U58TdI91+YMazx34vSYqMr/lw+NcpqJGk29RtNxpMxTLZDQnbrkEbEFs2b
IGHFoPJWobjZ4DlJfcQYg2EQziKGP7YemgESR+CflJYk+gn5pTR/zIqcVG1UvGpjx22o4dwXlvua
vxNfIarAD56wiX89m8R3fQpTxwdLUiVPoi/7sX/jyTM5xOhQlkvUtXEnAQzqpyQOCbYK8Ua2GbjT
3rMyUYhk4OICPZOLpDqXYln3Y2ouG7lGiPOhbwz75VOin8Za+f8A5u+pWaeik+9LmSHWA78hZTLV
44YlhBkKETN6I1eUk0Bzi6LaVj8Y7eWNMH4Vme0hFP6rN/iSihbTjntjTNHP+qULBL1NwTXCo560
ftWW4v4i1dfjLIZ+DluBIRlV+Fq4QeRooVSDiqmWmmjDJ2UYrkvYC6Ch9+XJCA5hSm4cNXG+5+yT
arC3QafeRsKw9MuPjlCNMvkgOv1OT5EqTdRgl8J6GKLaa0JodsUXkyqFCeMF/DUl5UzlbC77opnp
nz0EKqpN7IuNEFRUltySh6iBVGHiCoK/Ev/3DdMSo0hjaZpH322iTQHYISKtEocAKve92rIEKESg
AV2JD4hawsy5VZfq7eQFcwCj9T5KQuqklt+x0ylx8kJ05zkZ7mlmGTEnZ6F9aOOirYa37n4Ff1zk
jHjmEvexOKgVm3yqJRluxqgc3svHQgA2NiXQbcuAqiWtHdRIkXbzDadnVxV9zqm1dF7zHc9d79js
UBJTuc1c3OaQ+Kn/tUfpUu9vGVO5r0M5dseiL5upFLXt9FywYXK9BPgsLw6nHiJHWtRkLa7cLJFt
/TTIth64tdnWyZTcLO+cxn3DbDkvMS1/LkvoMl9ftPXyLHATB55SNyxcwyXELQyqvwFJ1WVWLIo9
E+EuJmSm0TuCXWimg6RsZolaVxyaHSg784pGWj6gyEz3z8xpMujhLSmEkLJ1xDnmXNlRDsfJ7sLr
UyQR7uaS868S11CKPNMN2Okf2zs7S9DQiJ2BzqIkIn9s0QySsXfEwKNg97xxNwN5V8JzxxegC74L
JgDodI569w6N0qy0vIv49brAMsvwGZmg1fH+VTJV//Fik/aj0oPLhJxgDTOfi6syvf1GMVgbkfCA
MC5fE+W36yfw7JSU6ThTLGMKAfO0Oe+GQPpxbntjV5CcKwq0YK5gd9yhRxPWncPnQG4+ytFywVD3
4zCoxY6OGQaisXfuBZnOZ64eXFS5Ph6ASoQLTFeZziLscP69xSm9wwpcu7rKXJGpiUKjhwbKZecD
4lhaftPIPNjGK4VX/8/odF2FMjY7n88eDPkTTQHiVaEpGqoCYGuRrJ838ikEFrbjnRavU43WytWP
O1AcBqkjY2BtLrqcCOJCsiunwLgekN4Jtawdwad9QZFUolfCxyONX5sh05+b6WIrzPJaXDJ5um3q
ozIM6FGUN91oRdwQDdJbk7o31tnbwR4znrgHnFYmowkvPEfe6/70R3XhkC3mCcPUXukBJKzhDhx9
1DnGmurSo+ilnq+h21yv1/3myCHS5OBdK8mTWGz9SwDnVm3MlV8VSA3lDF3Eqz7TlrdiDgjJMrlZ
8tA29YNYdoC4qTdx0xwZAfEiSABA0RC96OhOIDexJwt2oaKsnfDohexjphj0mdf0SIVxo+xFEx07
+XZpOPYAQbi0OERk4mvncFSoJ6U7A4IxoVy2dY8iAuVGox7njNCNcia8Vu5dSc0AbBKMKl4TloaA
qB5876nbYewadCxAWD7anIRLqE1S81Qu6GJNZl//7igZ1DeybG++iCISeNi7baigr0+lXxB6UYcr
1rHuzZ7x8e2QJTfkR3d3rE+4G62JNgoe8ppOV0SfFJC4ICH0za/KcwVHn2b7/DG7/+caYj97Mamz
TZZ6VoHHYqsWPGbeVo9qen30bI0Yuk/FG6w48JHGnQH6ZkkxfMFU99k3VpCzdF2gGs1wHzyjmhzb
GSKYK+MiNEfR6QcaOiZndM2W6FCKpAuHGoihjECl1eVyLD6c3R7pZbbWqE7GrWwCI4Ujn/a5rRa6
L5KhSt1CTwh7XZvZN5/A8wncd1XZeBMqFEBBOESgzrlTarHYSlvXzkxM6PqemEo/rjM/JCRW3I34
MUXnQjefWjALGSgr+PCsXc1/eeMZW4hS5V7O9XIzgxoqCGaUu4ugaVTaGFzJP/Nb288CZnQFroma
XhkgR6eiQxz7vVE4cTZYO2+Oe8WZsbFrd/c32ESnnIENckNdz0AsfnbYq4qAf0XwFrjhMJiR30JL
QmtovdICBGK6rxq78Y5pISYNTZ8zvFySYsStcoBuo687u5DqZmMnttV9GxBm2rJImE81CJZmwEvr
hH8wRDcQPC5D8US6J1Uq40Tibm4VRkX+t+SbwA/OdFW7w9S6PQPpg0fi6Z9tpmIwUYrLy3fn5Hde
Fhbwy49FvZ5NPtCY6btW92eE0pca4i3GbL1Sx0yGgPA+MCYTS3f5vIzOO8mCnxDPyW1blVxDb//i
BImA3rG6Yt57RCIRcAjRmwTsiHkFRy9vgU2WBDs6C2qpt28AKkCm8O0Qs+3XkiI/ZsPtFxutxa3h
aQEZta58GEo/ykxBx/1IoDFzilT8wsKEks8m8bz4Cf7447n/wmVNAs6qjHG5OcwxnOeAFfz+GoZs
w7yHiMftlRjPdhdS5UxAsIISilfLzyaNUV20BC2bY0TYVDpbe9YGBPywfA6lq5P0Rki3vja4nqKu
WVz3dbVgglMxYZtdFLw59e5HJ6VsmtlL55SX7ZlNufVCjED5fmpL3TWCJodOUQSiOAuoqwvqeO0B
R69lIQ2z+8jAlsTtjFnzntEiFQJqkUUt1hyc8r4aidE0Vq4NW45YUmk1HbsVMbxPsSZbhv66GMZE
AQmd5dCkVyXSrywG872Am4wK5r5f2zD0KZU9AQzqKzOBXRze1+125nF5oMmeBY6Tu1gWQ0hWmIj7
/iPOZD564aQkZOgccdbcctlFlrWQCDDcid+dUcfQj/VAXwptxcs0CiSUZVoEROhY9R3eLTmJe640
WgIjmxM6JPw1pWHSggLr3kasSVMebeRGs5zMFwr2AOwN8fcwDu+Z/RnZJbb4LQs9v8TizTkJ1vLh
GFQdtFaTxR6GfA/F6XGi2YdxoNUOsnpfNYimyb4qYPEKlonoStGvX1pJ5uQTFnCWO1mcQvXE5SYu
M3ZUEmGcmBMDKSbgbR2VcSLcEsp8CfgksmXvn5uvabgFWz//oobpqbx/oZM60B+0tclTZ8Q4zT9W
P4c87Kd3J+yK3ciySjWXa0rhmBUxSsNzKRaxtb1FmARp3QxvxAPczpxcgPMReXkxr/Zg7tTdHgO6
393Ud3VcNH8pIPRRVcyrIdmUQviaIj5QbZfvDKZlA7fAkwJk8uU8WZ2t32w1f7lS88oC1Bl0x2No
zqzf4ou5ez/QJ/2fKI7YdaN6+UJVA57oUGRjpuaNjdw6y0Tbm615Bzg5SHbg4/Agl/YntoWxVJfb
BS7G0CRmi0RB7WxFNzLPUTnRv/rzOqDNuEBp7KRd9uYQxdatnvb2M/k89chPcKYqyun7+wjyE/hT
qpmIFTOARVkxISGpcAC4BM4RfEAlw62EaKsMLAem3QQ7u2H0odzCjA15ZxGHYhlRoxxNZmaEJV0e
ajGhgBsM7eWdSOo7UV0NlDzU5CzrN/uswKzvKwZWodRIVGcjq0Hn+rIreXLQUHQcruNqfTjzJu5h
GO2iOf/tbaRXcB06ohsMZqrKPjgoWQIqC7P6XAkaE0m+Gj+ys1YJn/TW40Nh5VtCPLJrJO8e523T
8wVbjWgBrotrL468uECV5dtssZBNLSIjvCbDjBuZPBVYjxfFozzFhuhBfWpZGRtwpzjWyAzKH2Wp
I+ZHeFGQsYV7AxEa9sMRsyYRJizp/IirJL7jpbku2rR5eMeL6gbv/eU47KJhjsNPAUTvBL3Ljgva
SXOgSbp8be5cwhTBVsneoSeLrfFPV5Zx5V8qYYwRHLMoJUseOYT2ekWvt2LR7AMO+xZ8Ez+sUkUp
vylBUOtmd/YxZ5gWH5jGIJvfaSkSI7qPK0ShlVLlQoFs+Ly1QnJezAnL7bKTFG5G5LTTw8/yWTaS
f7aeed+Kli1fTbJaRg1DT85hLw0oT1hBVnkiByNb8A7Szj6cBM73Ldon0dbb9+O9xFYDLFWKcAsG
ZO24yqSbQRggwlqi5qWYticbC+CTi2SqCnuCqnqSoaPjG1XgViK3w9B2ZL9iOG+CT49gjG4H4k9/
y9WQi3iU167sBuPWWNcWPz9VC5inPC5F4quMV0KW3PPXXwHPq/iMp7a0TKhjSbzv5Jt67FxWxaJf
OjORjP7lkc9rNUhvNXmjryCwdEFzsvszjBgTOFz90PHAcuHrwjDzoP207ZOv0ZnCa3mbpG2Yh5hB
KpKyDvv6RgpH8zn5l1BS/if8qw616Wq2v7lSjDFNh97gwUJp0Gp/3Q/YRNQJ7Y6w8/A79xF+K2jE
6Jcirukjj86o1E/g2Y+tWq+Kc/q9oaJPdUjzEQG6Fxa2EEvXlVFg2z3KtaKNFdohlZyuTrUVVWZp
1WuwD4qtHEqyjDQyoYeEHiV7uz01p98vhONazB/NHWhU6t3snAKl7zuRHnvzoTkaKfmhjcGxSg/H
systAOGPa+X40Nrfzh8hZVhJ0AQfSZ4yqUzfF4/SCOTI5hDVkdC4BYTJDz8CTs4LxWKxTQCHAL9/
wOF58mB9xHvlPIzLG43URQq/vxStYqjL3HaPYHMGqPrYwisgFtvEM2nn8PXERNCsSiQq4vBKalBU
XevdxNoyNPR/JNfdCPe5KWdA5QYCOJymZFVk6jXKZzkhjBCmosEIaWWNGMcqq1aPQmNTrUYZWfmU
JAZgZD8JwlKH9/9GFDkntWg+4b/b+QKQaXdTseVcmIR6xy56aRb6QWvriOpF8vHVhcNLdOHXPg3Q
msknfnn4mLvLkGauNkcH+SGEEByMn1sSXG+MkV5wucu1gZZkM6MLLVTIQEFzdYre6T4rWYq3KYdp
jkbzUibfUodIdnezC/QLveEKV7fP54gGLZJ4uNqSFSJWhqX9/x7YJq1kjfaadzr5N0Uc4fj7Gw8z
EcyvTpOgDkR6y/kWVd9leKgZel+QGtxzdlzgj6EY2LwpgPzeNkGrJTwMb58y7/uM4PY/qQMxegTL
Uc8bSEgPhsskoi2G7BhVsFmKVKlk7RlfhJYGlVOW68y9teue7CXmcKJngIOYzp6izAtM+ZDoi7cs
+xCCS4IK7qOUAg56TUJicT5nj6Rzl9LsT9vJyqY6waQFnQAewWIRnrHGiG1i8hhBm35etmjLQunU
3ePE5d/opGPyhf8s7601KPvtP0uPDftTYUIjji0T7y23QZCRSSaEnKcT62+a2lWQgorcwCjDsTWf
2gW9sx02xCZd53ns00lQbFKW0JVEHZ2LNbU8+z5+ARkBtpFhR4Sai2sPd1G4j+m10SxvObuIabdD
l9vjCjM2g/JW0HvaeThlFOcgLs3UqRJrStcM+ck6tU+VtY3lhOQUXuih7owsA2Da2TlV4Ii1lPQr
+Rm/eiaD32l9UcuPs00N/ocdrRE7Nq6LLEwB7ppRrh7KcNA5MrAkkMUaqE+XPaMAlJOBtMY6yisk
KczOmquy6TamJQRO6iZwFuMyU7oOgdrjzw2ppKi+LFfe+b3iFzN5kpoy+254KsFmsAHJ8ONmstoZ
uwVWLSiDvvcEbk7loDp1EAqdDNhxuQDcgPquDC1vhpqH4Oyu+NMt6Wpnkhd87DL4lBTLXOzXk9oW
nlJSGRc4XrgVW4x7hGakB8YB2RsCHWqN0pOqiiYQtOb7Hrf4GbbPPBJGEQ1Fv6ylmAYsVNCh1B2C
f9Jrt7lgPLsaoTpF9SfuqnGxBWxT2hC3C8BUon0uyeFIAXaqJmhfhYIAqoDcB01THVcoaPCkEPvK
qcfoUZOspk4OVCyfzKgdzEbe/zwoBGj+tEOUh3chhFv7W4KkFVFB56abEqT+VFxTNeNsEHOA9VjH
vNb2SvS40fftLRr7aGDh7d5/Ty51omvNVS/kUlXhI2/9RyJeB4v14OhTwiQA9wMx0PS8nFAILmnt
k1Hr7Oa+6XMBkxcB1RfXjV/+BuxiRDRGm2STtmI5N7rfHEi6Qy870VoFtsyOpRsPKeaE0qXrATmw
SSBUksoE5hxOMHwbBa8/1NqJW9XFmYSx3YEGNTD84tvOFN8yWSv1s/Dg4ObrxxaOZ1jRSHVqj783
lUmCijSclotZfdL9Gvc0Gvp5EWwhUlGIiulYH4ZGwljvzXjVJ9nmnHUjchLiKeaOClccCTstq3xG
AsoEWFn04HGuHUVzvFN/aBjtvNjBnNk2W1+LoZBzTLtjt1Tp8dzRARqbKipbM9ef1jEldDBAdcxq
BYpVYyCLW8LJT4FOhDwUL8kjFGJE3QuVKnTj6uci83/mNufB0C+UIJY2zBFnGsDAcpKqEmdjyQRL
sIzsGcn0I7KAThzjl6ZYRfX8arCeKepurEDYujkTg+HbnI+q3fSQslsawFojy1lWw2YDU4k+beB8
Mic5fUtyITVsHTdZq1fJxymYV8CyuurE5U3lQ2HQNS4cX4QTpb7wG/1zoGi0CZlW2rLTB46reZeA
NTKWvjw7YNC3QIaHkSBDmrH9gHiA9s4eZYzNsDry3F3htQPprY8HZ6QoPomhUowtMY9JdNjDvybU
jBwowQ1Y3iHc0eZncs/LunLEe7Pl5JPJ28zyU/KM1ud3akjW9z6fQbpoOoerUS1LZ/HKmD8rG49Z
5D6NjvLGuzrXB0/MkJYKXqMu3t0FTySyZIWiybrIxwOQWB3tGN7gIOnnLeZPjBmN3C9bvL+sMB48
H3qHHMY18M7uhJPPtNQ+znq/JWAopqmCoWBC6o54LKnYCEVGquDwadyPaJot+QOmYPbz0jRJ6dB/
KG9rCl0Xc0p6KpLAcsuv9nXd4q6d3SHxjaFO2N6TIBFHIHjSE1Ard3r60tHXAxjPsYo8UXXg6FlD
qHxWaYDY3CSdFJGPZ6YTFa/1KsKLn6drL8srrylt9xF/jA3cRarWSLa2sVLZRT44oj9lgnyASnG0
IVmSLsyTI2V1T/1VpSznAhB6vQKpazWYCAhnS1oRg/+tqHx90olFOScJaDQ0CmbC2u65G8fwnIfz
OZQccrSWVsfMpot34cTYmCdoi1b+wegvoKVSSW9W1bnBTYlHS2g47+rR3SyQFFc8uTKELI/0zL0C
XAFc4cx17VX+9rR9iTBQbGe+Yek9FH7xJUkNkwZW22+w6zgXZZCwh4Je1L188LamFDsve4ImXgas
shtkub9qbfiAMRzrVTP6tpCvpPmS5aBqtP8f7nmv2yugZlsy1FF/F0/TidF8AsIysWtSBu2if0kA
Q5Sw69KNU8D70tIUPIIJ5lIIbSgawuR238HRipab1jaTYiKQ0Y4DkjhJvdWB4mzdVCE5uLEFIYxf
fRvcT/uDEuCVCrC4M7PctxfvmM3AaMRhuq6TNw2GSI9wbuj6tZa5eIGTJ8YC7iP6nWtmogubnula
P9WxKc3WxJj2D7eksMx2fdIKjnPDgYW0Xkz1FqMyiw/JBZP9A8bSXSfVJ3290vd9wsZx4f0sCu1p
1zenCORgdKgb6b8RcC9snzOee2OQzo47r+X8EL4M1ms+kBkI61MjOQPzviV7hswW5R/+LHHfz5N1
q8A1WKFYc++ST9EdNbR2Ik0Cu5xkx0Z2Tq+Q/8F22uSjq7igPRZFBv4GHy0T/k2UzyJtZDygScEv
i35Jxwz6HaWPAdq7ELEpUM+Toq/WFJTaolo6ZfFrPjTven+vdYbCDkFLgYEs1NpFlePg0NBnsV5p
QlURe6dU8x0YjP1cr9rWby8xgH4rVCIZb9f29sSYBPWXKyfsxzFmRWwLzKh1rsmdmUar5JYfx7kA
Yqxtc4xVLxex5yKuyeDK/psRlQz2I1QbSid1pXPtcq9VEuRLhtHoQqGD55hIn3y1LCdICBGBc6lI
ul8oPxDm6G3V2LU5Nm/puMHO4zDyNwfv5ORg/a/LZascJFTlvP1QXmHjtptt+e+cijuoSLLCkYbe
qTF0CC75K/uCgGrfGWDrAMO0iX9RJFx9mUuXSXQp1FfnsQeNvSHTNlpuwOk+G9lfDiaq5vpnlwpX
rcQDr7bTj1Nyq9N76bSij+VVDW5STUqYsgYNxKrkQWF70flUnKRNjI/xdoz6lRuBRh37pcd76iL6
qYPdFybbA3aXgSjUvaQJxbUUAnfhEVffFIh0Y44s37BZHzmEe1AP4p6WIYoKTj8T9nc1Igv5G/Ys
KtWqnOOU50GQy/15KUIPW7stdZebVHMQJR8cMc5NPPySUlQxO7IhSlLKzyhtxSQC6Je3ufEYvcn1
BFUlwsP85v2Peld50ziXnVnZYAt+bW0/Z6TJuzhDHM0NYZ3nmf3bIzUXMFtOlATX+khXhzF1KYDA
0gpJVCpae+LFlVncQVqbMzMeQJxXwAd7eKgbQw1o1JKxbU1B6Y0EN5VX/yadl3OaBSWMfySJb/i4
8ZV3tW9+1rMKhgYDYOiL6uYZ1PC9flgpF0MYSxwPlmJXud2PXJ5WamDuY0FRNMLJAhU96P32uuRN
12qjHsqNCGSFbXKQ4NR0JO/W64GtomxLYiTZTH0oOQEAhEP4vRWdkVdvwXUdb+zSnk4SyWpEFQvf
rdzxy2yKWbdn9KxhAJ2YhTCLtKIn+PDmUSZPNLVGPuSikVMHTanvWztm4kXhfqeaN7RNLgqU2wlP
+8rM2aSILRiY1V518+RB8bj1AxD3cw7DK2b6z1g0HaGHxuYbvmdbwykoBkB5AIJl4e56DTf3u+SC
S5J6TE/xnM0Ww0lAONsOoiFsaXjcHM8GE01f7POa0x8Pu51NVxvguybUkOGigVsnQ2Lc1+NPeohE
jqAPdamUN1jexZ1ao8uC78by/R+jaYTA7UbiOI2R+nctLtoUFQolVyIY3ucXhfoOkDzJtoKIEzTW
qP/3Byip/h+hSva1AYsvuv3vQwbUX8ma6dqPZaSPE4MiZKaqX0aO2jGMpTTNF3QVSUS0D2N/oWQH
1CKkP+EVpZb9Cu8wsPKjfeUJ6BhurkjGukOsaQwErIg29JnDjB1EzPCRPXD15R/uOZBn9lRBgoYu
kmWmwuFtyLAbQpYqOhm9lLtwBn4KI2e/xr7NLALDqJ8s9TGy2pRyiqcnTUcaCQ6VvV50R6LmKs+3
STZk4tjBgFfaSZ4/UtjREVZjYjvo9knlHZWie2hmQW4mAmz76tWFSfdIDlBEPsTldaJD+OyQaYYK
sRnh4gtnIIPZRMwKUzlS1uTnLEZ51zgjP0c5oavmHNK2BEcVWlHOfrZ7QEUBCoWLVTx1CirzFPAV
p9wJMkJHDmOshz59UcYzYmxAyB+r5l0KZMV+cLQEDrYuai8zhhZENqeaOY1a+AvDf8EUVIJ4fc6F
aDPM4tLh47i53k7X+JXxJIfQkVW3b3sVDOoa2o1vrNYNELtv4Hr6tnmMA324vq2XFf7dGlSfuqi3
vP5jmOannw6ew/CeYcibpOjmzaSXRuvtxI9ai2sFHGiLUns9Ko6A0gsmmsfDHVCoydSWXdWtp+Yt
h1vfGgQuH6eTSCnyJAtzD1bkSYfmBwa/F/Yc2ugloD2P4SMgBR2lPCoICNbkXQLYww1FzH9+cZGD
QLhSshiSkzdlyP4HiQmXYN9/T9HtTl11HG3Q4MtDxXG51cfBFPAka2XatF8sW0DrJU5rfHe4xxSr
9zCwNRz5xzvURwORtIIYXLZ3B30KTsbUOV6gY/JgRm2WLo4OVenQqcZiphGpD25GzILp60LHVRHG
NcOT7z2VWdC76+Cw0KNZkikwwp+zlp8hWFlvaC0aTuGCT3vIMyuPkUpIql6rIwS2aulwDSYvjnsL
HYU3Bv47nTZqyck4O2XUyv6xfvpdEsfq3cXXeU2n6gmINUE95GlayNo9K6nehEFFVvMcdT2tS4h1
23rASlo0X4Orv9HRRQ1CT/PuPYCvDPJND9+v7/o+dgmRd3mjly7CHC8SxrZ9Y68AqtOtZjlsovDj
04RPtjXpo1OY2pjpZ2iBdCsUS9hLQ3GXrf6HjeZNErb9nAVH1EDlOeGpxEm2303eisDjPVRn/QCX
s58Q+ybUCUv5e8yBiD6IEbKO44zR6M53XfD7U52up24ZYpLvzyS85+O7YntJyu4lFwfhAwC73eJM
hT5JFkw5zoJEshSwtu369EkBa2RTxHl0OoF4C9Z+IBqYIdFG8bMFFrA0zYRG6de0dMDH/IzpOHo4
dVM+QuUJrP0i2fblh8P8xZjuiG0MIIyj9x+UHsQhCc/FwifKtToUpLdTsP+C/VFFW4O3l8r/ZcBf
S1TeA7LbyoF8duU1g7V37pROn6J3TqgmCMpn4XyHeR1RiVg6PXP4UcSlZ0RLtXFFgzgBfJFXBj9C
HFotFo6kOflneVKLgNzTe1heXgcCCyktQ4QJ3GGlEPMGW3i1XU5/rk0OqKBMmVCVjWW+PTEISflr
8QyGmzv+1hZUmwBOj9O8w0UhIenmDH6tDKbFIroH49RaAZPXBebhdJTpRdK7RcXg0xWPT/dsKKFC
3bI3jRXGzl19vY7Cam+JZwHKEf7gifhxmrEyaGxrS5y0bYiq0+BHHc4bdvINdyVWJ4OCXhPp2tfa
3hnW4fUEyEriV2WWxRdS0utK4Z5GHMzy5kaIYUWBtljRT/ciBBrIaQsKvhzSB/T5bEhFHrFkL4HV
dVmJphUKc2MGoLVPUIIdSy30xutRIkNeIQcuMeVLhzb90F7lHfATU5FoM+kk2w2drp4zo0xG2B/W
A+UUjuJjRHD6S/jrgde9oWpwXs8iMPNDFOcF9tngNGUsrBH3R5wA6mw/9t7rZbe2OEQxeCAmMlUO
3Ym+23T6cqO5l/+47iITdTzbSkNIFLjD6dVv0QgcAFzmz6UAxhj5SccX1RiUs9rTmKrvHDI23tMh
eCtaycVyiLf5bfh8Gkx4vL7XI2tFV/pc1OZmUxZqKfF9SdI+MTsJB+J3mDnHhDdkG/7BEjxz8BCW
SuSA4XCcYn4CmFR+8Xq08L0TJ+CQVcI1J/fANiLYUBUSyUJZ5v4T4PeAB+9bd/4i0xz+CUGklXxi
nLALXXr6Ag3W/UDBUKExrL24vT4Z/APklTGlivfdEfaaPkog44rjqm1AjE+6nba4CHdCENYgdMnI
BMHK9mhF1NGiCXWmTF83ddVkwzVvoB9p/o97Bo8u9BpFc967/kjDYl/PiZ851OMrXkgjc7jUL0LM
OU3Ywfnd1C3bYbVcjS5aua5UyWE22b6/DsKfvEkQI4665DeT7IyvoZLfBteci0ZSLuCNKu3Rx5He
DTUnOLUB8lZWqjmAlDXIXm5lGmxfTDob49pPOI0qisr5BagGDshr+QI4YWZzE0l3kmQLyzkEjlcK
qZ4AHmOFTMCuD/PyswXW226CUYD34l8ul2WQZ312kVZYlx6ICRQLAmLNpirGLRKTxeUCc8Nju8VC
nOgXTvyG/rj/N7faynFT80G8oEPhlspjPO6L7Y3A+zOjHLWt1l1jRhq74hy+jnHmp7e0higMVvKY
KgMnd2aLirWU8SwxVGB/JhxksyVwXgjLoj/gdWo2jcnvo74xCSZqMKKlGiFWqjwf4+B8sZnPE+eR
rFdYfWpejHKpqkR9YnZQo70tBnUWDAJyqOTqB2qy/FWwecZUp4iCR8RJYDlri4qIZ0oT2J3vwRWa
LxCTUNQ4bw7/V1So5MEjGNl32vXIOKN22wmoPF+8a4PcvgpNw4jt9ZgBeXij1LEUJylMWZCU6hSu
mIZImqw8e8bznD2MgvcJHTFsoQipO9buDpkdVqtoFdBhktT1Ny21BBtFwM0LEcvMIgi3AEtwCDZm
JR946WoDhsGO9pg6rb6O1zMBN+VCMp9mM2qqCxLheGEDVcxhjuqaHgB67s93zgzUfEvbwlYXt1WC
7jqAT/3l9HKm0+rN4NwXUnNCvhDXp+l9lyLbD20wvKx+gnRfA+GGVRQuH93yIXudwdoO8grWygTH
YLuGyK1x1QhB/2DCTy7Zltqq2WFtQ6xZjWlRaXttbAnLyhYe/6vTjpmxryhhwi7BPQIQ+qhMsAQ1
Ag8weKEdIYumnzj/O+XSN3ETYo5gtgFwDJ8xZcPE33AILsRwPhKQ9ds8RrTXTt/kSEeS1OiFonOW
udWRgyd6Hu+cTfpV8h39oQUOEY4a3y8KTth4DEfrS+kANScHFZaRk56XMBqshS7e4eYpKxNB1FIz
yBmEtsuhI53mGjghkrrhrvi6YWDIuUWoIQCwNgiRNlwWHaeFp/UChz4FYosoiNesO7uusi722qzz
zJo3gfPItjgmgyuiBCLZNy0GqTYZOLVTG5Lb3Er9Z0rvotxpghXnOccUtv5S0H2R3h49XJ1CUnHr
kLPU624KorvUBM9nevLUxNhJDbX5OPtHXiAclA3m5Erbg3/T6PXuaZXsnO/eZR4R9QrD7S/h0KHT
2aEEBif5hx3xS2e3gEBSmUxAVoskhemCBZbbPECDR3S1XyKFWa9E5M9C2T+hIQZae6mo3EeIq6oV
N8srnWPoeFbRn3f8GKyMVGiXwtlk1XnGF/DVQZBf674GlmkpUMORN4/rcFL6jhgNzg821eANdByQ
Esp8Y7B+Vt9lW+m5ZtigknIjbeYZjaoQMS2VIxn/KEWhgfzEX15KfmlZD33zENYyj+xF4WAeU4+J
egS+dC5VUjlQU6997Qun+isyeqUYN8AA+hIZYD1vbZJbIh5CaTpZdPZq73Ygqor/lb0sZX1UqrNN
uagZaltrjDkgjH1w1fLMoBSCe0muKS6kH7Ey4rmbrLCF5UqAR2isuvo8kS17yb/PnSctV/WuF35k
enpEoFZ9Vl6pLJ/7BVke0vz78TPFRECJQkSLPeRZakNbAlQCd+Zrdg5uH/HCmuHCL1D3FxZoDnn5
574xCcdeJLCpCBcHPrZ6EZSb9uRZFjr4nGcfcdcX+R2r20q+ssEG0SrPyOXax0Z/Ca2fS0BvfZF2
s3fQkgimlL25hi93JLO5O9m+4s2e8rSbs2xQ/pk2f44KQt3JZvRn6KNjWKYejKqweIpmuvGC3o7k
DWatKa5AAq7kBo/x38mJ1eNrK64vJ7pgB7Maq+64uRbfuw+rv9tOk5+h2hOCJaRt8o0oQkPNVThT
jKf5RYMwA58lazAeaX9L70J4Yyj+T24To2wVSpisfj0UHREubhCIFn4+QuQNL3fdHxTDOlIxVw8d
AbtDkNgW2KiH2cu5jn9vk1e/h/lBrxonzUhmqoiyTjDZKXVQ6srSlERC5Y5J/esmOKqlzn5bNCQK
CzRB8docg0nU66qqul7NyUy0sxU4JiTdrTj7aDyykc2ips59RdFZ7YW/xszku0+7RX+qzwg/NJW3
P2Ul4w+lpdfN8tQRsNI07GVXuTKJFF7nxdijBsEDw7FW/vuC6YpcB1OntZMfl3pgShY2LlJb7yhD
lMH7hUKKtvtuOHuU1xH01hl32ePbrQuaTsBWuy06HAPbs4I6o778UFleM+mV+jmOCf8gBLd9s4k5
EcSNPB78VV70YR+v2osEYv5iGPrihkzLvS6lT6PjUQM5x9vr9eyjv+0wVkMozhp4bli86PTHh+tH
oz0cyD+b+McgE2qi+tZ9agmE28Io+CxC+rF5Kcfj616B1+eLkJV+K0Ni/3sgV9J/ndB1zPVoiywN
OXarzhy4WCItdCzREAhg0iymCqD42xipY4eE3vQB/1+R9s/EDvB34Q1Ew+9z5yAiHqcFAtJTxYyN
bQBxAfH5VtuVNmOW4MkkzCUBGB1K6ALLWqkEt7bekEFlCZKVlhjB783hg2XUBvwD8KT7E+gSg5hg
W5A2H906jYJvqVcm+E5FLLRNo+avnui+L9Cf2FixfA4MNL1ILEng0V1HeHvqM774xZovdU3mfpSu
AERQ2lUiTQeotR9avVBSsE6K+MRMNdMLOfu4LIcpaC1M0cKWuNCi5QBVr/F5zHshde185cP8+Zzy
jwCja353yboWjUGxvejv00PcSvhiRZgl1sAwxQ2Tp9A6lLssiedhffQBpTnjpKOp4Es8vbPIcHZv
nkLqzvlMetG4GHEoIGhdhcC8QzVKx6RiP04MkjZpDwH5tuTDYtpSM8my6maHQL6VYtaZTl2jjleQ
MisGng9AN3RZbSfhp/9cfo7gxiwSunyMEli369AJfj+ijjDnvYuV0FZhRBymatSlZrJ+lpVgJqFo
vTP9gAFy2Znpsu9bNouQC72ou3rOinBQ67P8UJ+9VlxpIAT7r/AgHcreaTDrryaChXzMBphNMovu
KG8gD7Rr5k0XPFAuMBN9EWzlLQvxOjpzcGGfAxd5BQ5Hxt0rNgrXy21govBScmF0KAQCliEfriav
ZMd0+KYL4GVY5UEZkKg5RAAy+YRbJdkglyWYI+X7ZRLRaUjd5xjgMiyLuu9GIdlM76XPEf5jMcnw
WBFcayBN3SOAzilzBmM1SE4Sk4N5aJe/JyI7NeWvRFWqyEnGcglJHv06c9bpX/yQlZ/YEHN/hCsR
1iharOpzGi9sznl4EmZAvcPAI+zTX08wpDfYTz0Yp6ruBXw1hsRssqaL9FZnX1w5vzwboLhxOl3G
WcWptrXGAs8oxRoUwlTSSQoiUCmqMjm5kEV8KG4pQ3Ut4WNdgXkFgRkyk/N2H4zyYROuZr+27VfT
doh3A8D85l5TYpXCzKVvtHHgP4/c2FzUDaFhnKj29Gdysw6B1nR2NVuD27IugYZJoHglSOfDcibC
qOyUr5OUnIvtVfWMdd0Hm9G7JNTKnfTcFL388iwfl0s93aJrfnDq1xutwJjJ3w3tBv0nj4UfNTtw
+9PqMB3hzfS0puV4ELtQKcFG9Gk2lqkafKT0pLJFJDdpZL9MHVs9D3XwtslX785AKNClpc/Hy4ot
KNo67TysSYzTTcUPuGIpFFpcj3qsyhdGjx99bPPnlzHKTnN18I+SzsYIpNHJ8TrgTBEMYjcJM6sZ
e8/s2KP2CU1lKvsLvtmtsdCSwaLJCFLNav526FU2gSgvvc4f2OQTthLPXxT7w/IcEuJkho2ASopO
06kGe7U4C6TOP4vtaYhUt2UQ8HXOnG2ZlP3/AN+orf15wUHVoDBQMd1IF/g9GPIM063Ohh1dhagw
2eCAKX93o8HHTQVHuIfeI4HlV25KItGuv/PmYo5c7PzMqagSpwBH1gGlU7mGn9OotbdJ/yfbTmsa
chFx2VCZApj/dpPmXtcQdbymPfFCRlIDWRkMh2d9J7FvbW+aXl1xIjyWgrSiAi+IACEj58LkLoIl
TQXkAN3B8E6bfoCmksY/zR5JzxYLCUMMJkv949gIaQcgIBG2elL08WwQsO7O8fYVbeDnmsG+7Q/j
3j/A9cfkL+N9RZ+K7GAIfasoTjMdRRtF/DepJK/82OzKRW4AHVJIBomoPyZLQLTmBhgBuXKI5OYh
/DrP/RGBHzVURJdoPAL4CBkLDoqrxgaHvSgUIViEeIg8/RiI0L5aNi9ZIWGNqK2uaI73lGxGPw0y
4gvW7I1UmnjmvYR+X2p/uKpF2wnCNro7TEJbliaF1xnITxKMWp0N6s4SlcywRe3yIohhJo6wG3SF
NhHedIGiA+iaSNzYhXjmtksyAxDyVuy1hwdKh6NeC4/b3qjVQ71edN1Ekxf/k0QOJ5JtvknPQ30f
cqcTHcmtxwrI2ys+ZktzA/lExpUz9Z2MHdCi/zoeVSBRrJT85QLygBpH3fRdlFfW2FCtpoHB44f9
w/dxGGLWaODD261vd52o42F2v/CcwqaXEk7oWL65Z3tLBTi4XiqxRoGPNUt73GcJQmuIuy+FjSnZ
WtIExtgEW4MCtGj8q+GETkKX484gM6jq5CCeW2+2EJjWtPWF98/Ett+qT+TPyH040UpopFaMK0qR
3orQZO0TsFDZTLwvA/3VZTHT+GpQDqZ+Rehv5oy/UzFY720qNHho1jYT/4Af6Q+TvqpsfxXeepaC
eudjAdmuukQgI/BhaOwEQ3RApac6jZ0CEeOsnjjwjeSDi0W4EgsY43U38TQJ+hxLu8d8MJC4t4qY
prPaO1Xonbj12gIBs9S2Hb8NyCeD2ysSahCbLXtNXcjBMcFivt9MH1aPFFuJpPcEMvX1wJaM8x0W
UPVQLyKxxT97+BPX5J963TN0d3WRDpit8PS3/eVHLlkJRnR31YVZpQ6YJ+aNtRF71mYnsXknKhz9
NyPj724MI3rSKcBpgrgprJJg4FjoLfK9d8cYsyK7P0yyHmJ1gaCWPVVaTiOrPi1HPCHpNTiUvOEl
NzNhIZhp6SShhbN3k8idcZyanH1yhzLZov7JK+lnEqV/RYnQze/oSJGBV92E9mY5i0Hn9csPVC+0
p2HrUl5HeI7cfAc6EPGrl5CQzx8OPxfnLKo3SUCbSvJ9yxLbeiyaLGc905ceeVYmLzE5lMzLR3EA
C02eSvR/CGprLKv6xl8F1lN3uzVvnEClvShTkctJ+Haw+kVIUTlSsvCdwpMQHHTMecFY8rCfFviP
f6FWNLbVOFDyGSppQCG9xKue0sbdOEFEaqsB9l2+Gnb8XeXLdc5FNLvPAG5hWMYy3Wv7bFcDoFnH
bcTA7/zEHTP0jsquh09eiYjg+LlQBeSw7FaDJOQw387cVws9sTdM5jJ9BlZeinOWFIsRTx7X2uSJ
x8uB/OVISV2UNm5IVsFTbvl/l4VbDuj8iPIH1nNhwNTtoc1NCm4wENVa6jRBGS5bS7njWwydXmU7
E2KvgvYTcJW/N8MkMZLEwUaeTzHDUEXlUKIyGyy19aqsCyi7tqaKw9NayFP3fBqDYZt5+c2z8Aqx
4jrv0HHJ+8g/ienU2JMTm+Z4DTGK5hdOhi5+IAseZe+NSRBR/G8BSR/ktqF6aGzMA3tCz63o8AcR
pzjvMDtNWQpjjgMAEclg6W5IaOpuOdnwnm9fUp2uzqcrw5QFhH0gRmqxhWpBuP2OaIxgbFvJyFTE
zFFRAOmRIemFHJN/Aj3KQSAgovHUj4Voa7H7y8lZStvS82s5XpyoHSm9AHWHOW9BGzUc7opYZqEW
GvYliODj56IHBMmHKZela7dhgaHiLIn/povLbeaYDDHhgbE1X+CDC08TeuCWz8tvAgzoQWzBFqtV
cFv3stDT4Nl5uUqODakgMJeXmXLfSQw5K/fvgp1+wennfO5LmyBZ5GGrE6FsBYVQX6ADvzw5V9Sh
5gK66bpVKVr8uHnrinJ8w4aVUS2cUH58134bScNC5ggzI3mNLb2ASFzSWVwigX6l9L/fj5KxOZc1
rvZoies+hkEPklx6BtF8XaF3nNzZd22E4u+2QxZZ4QaV4H6U7wjp5aGwVdYI5OlakTNPHdn4BNb9
Okvzy0mb/lbeSI7aSfg8kDs/gPB1CIFTGinpd1EzHyE7IbVmy7fyz498TYeJW5kuIvRXdMWniX7e
XUbkIl75+m25Q6tm79gnuxLYZV2X5HVyNo5U/mJjhbl8PnFLZ2QrXG4NVVkIzCpVX2LOiUa49o7e
tfY9dcXjmBEWlyKEQBwDtVR1rH6BY9P0YK7IJPjxwpL5nujNgVTPfreW0IaZ8yPPz+qfL5aTRn2T
in4s66GrPVi725dzIZuIQ0EFLG4vq1Uu4fMxLbe4Ryv78mpJAxyX9ghgs4fHXEd/qRGAcgNyJW5L
sygBVln8Y9VpoAs04dH9zThTsfo9r7UIHFN+xMv+6F8VxrOsRtA+qr9SqXC9KFF3r8VPVQ2OLG2y
+Edm0wyxdG72JK2WfajLV4Tn3ZZeb2po5bZHuXf0+fHoWcNNxm+t1J0xWGdGxjO1r18R2afrrOzi
KVDQv1j0o06HJsmL8KbTLfcwP7SD+EcCJojT65saDvQ0d3VEPi00FwzUhvJ/4dMjHbTSkILvFTiy
7VMidxhgX2wTzHob7xSTbjH2zeJxRRihmveWkpDA9A1o1OCOrQlDz26m7/au8IDUBMy7pGMlIvW3
RMPlXkIBYqYV6W3g8vnsYhjdxolyB8MGUcq6pyYYbVn+Z8cv3cTyfLUZiZy2i1h7GmtIOHOzh/fD
FYCbzZCS/d2Jv1pzVN/m8/ra5ry/yarlYUK3JzUYKD0uKsBXv4Hu4iAbBsrPii2qxBU6/tIDKxQ9
DDgAKdqg2j2lGeQqchvqnZRr1hworyPc9RgeeBXG0ujtu1ZVY5qK6iYOgkVDxSXlRSpnZF5e7hjd
3ktlvDVjpbYOT/BkfNu5BXXW7dOzb+LeV6KVs/0lWFdkvDdMEcyzcmkOYT4yxOY+lLd1xZPIEOBH
LFnCiZR2hcT7ebGQQbDwTnqwTrVdtH2ulDLj62kYFu4MM6hBJXJi5WXVaQ0h2JeKYTqezK/F0E0n
OWZ+cBMzTX2NsKaOZ2ndP8R9J0+TjbyX5pTuYle9vQDr0YQDa5ctgItScHFWgLV/AKtw2KrnacLU
pRt2FWFYug+zLkceE+U7qvEJpmOaAQuYwsm6rQOFW/cR2SoiPSqm2aoRk/AKhzhkRjpji8JKilyr
JTrCcGobqk+QKJZf1t5GL+w+0jIgOgMV8PJ8FtnRiJagr3dr3lIWRPapW4H6xKaC/JwsPwvAv9n/
142vHqWC5XPk4eNo7drCOX4bVOyb0xfWJBOp/o6AUojO4fwzZWpGCzdqA9yY0NKLmPCQ3BF+agBg
r0+zTLls7m4TdOatlp/bTsrpLe2GHBtTiO8GJJGlT1OYf5PZ33iHEit3si+MPzojFWz8si2NAcZI
sB2jpJDAiYnaWHX/2YXnaDYwu/KhrX2NdcyE+uteLRuJ0xPSTjANu5ItckeKX8Lt3Ibp/xRrhfaM
7+aZNdfgrBWlHE190MxrR1nOLhZSbb73JGi3UL90spHaapfo7bMLjQAsIJeMzNp3XRTB7ugkvhzb
kr18RQxGwfVZNQ0MGPSe4KoGDYYq4vGicRfIkQGHuNzoh4zu+6LS6tFXMu8NrqXufi7Mxj+OEf10
Ht9s2rFHO/701V0RtGK1WURvdo1mVxhW2E7COpSFVk2Tderu7Wvpr+B9YuCCHJdyKhfG5W4ZtcCT
NxbX8RdakCe8mSRRXV61ta3s9IaFBf+ril2bd9BI/rDdUMy4cZ3KWE/lQujd9nRrMfGhGrbf7kU6
BkiNpxCvCvWDsaEQOPtQ0CfRh2qpeINB5ouZO50z1fObshPi0Wcx9w2uP268rs437kb8YwwAfFfQ
cb5Ik0IrQ0Ad+OH0he0iozkgO8jR8516895a8JMUJFZAhXT7sflNiYMfRvt0U2Tw0tFdRJsT0v+f
fW3XUOdmm1EUoF1pXI/lqa/Vz/Q1R6dO4nDzgbXw0n1EZ1a7r5yAy18bMqvdYR5Ec2i/IVIV2teX
sRmGsW1XNTso9GidG+FeRaWEiM26lHhz3brTFh4P+CIheikw8b0yj2NOWSMDHD5SfOXi9AL7wZa7
LLynCWK0PMR0kzPQGCE403wM7lKwzrYk0/0l1qszqK1k07e0FpGkhCGnMh7/N3WmbGF3dgtlxJpG
TYIWZEYrDWyLCPwqq+Fo7dkAcV+pjsOJ9IADlv+y6wvXdghXM74iW4fdWzBSZkejJLYLdY8ZudM6
EAUn+uNrJYWroAPzUIsUQdEWLHCkJFuX9yqRh8rdE0z1YRva+X6dDFum/7XGBj67IyJ9wDDvi1bK
yBNDogbUC/JCwb5J6rEJCRL5PLYYSOCjEVrWRRDBon6Se5GzcP7DRqmTrju+6KV4yazGgaZfsLU5
TBNz8DK6C9TtmhoD9WTOpFIWeQL5eo5kWMDCR8mgVsrtMtNdxl6OcERcYEu3AVmTkGOmSP6WxPN/
/y/KKF1DrcVJy8N+mggJWMIhoFTGm011kBDQJn6EkUcBKAdXw7Xo/S3b+rsogdZohtZT+hAY2dMe
IcdX+yRREVkVRo/G5UTJ7mUqPBH4D6SpLPyYWOV1O6Ft8GyCZmLtMxU3Xvv5B1zEYgWbbn2FpbjP
BUaSERPMbHlqKb2ndNWdsuCrbC5htccfbV/RxJ1Mi2x/QdPkG8JxpkT22Ai1ZpeqYEJL2vUJziIu
b01wuat0QagHfom4ZI5sMAHHd+1g4FhEOZ4M+xw0HlKEu+YAy8XLlMviBIdXNwLCW8WSENzKEMzy
6v6ldScow9tuYnHPN2dVHaCjrmNSFHGUpVntgi4G42PjuBcUWCz1h3+bOVfbnjBgbPQNQ1JdvPC4
K3f3P1CXiMIa/fcTkHFX93z+5/UU5ZAAPCjqvkRtq5+6TzJF/HNOCgs3o1s6ign/7Vr3cVBxelG8
AZWBYhjrcvawyY5KnP7h1h/Y3Es1mnMLJe0NCVa9NKpcY9jLrC2T99WgwI6iIK3eTTr5JdGrjllW
ORowMZ2jCnpK/4sMvW6jmVCIj96cEhHwfSUx60TTc+uZvHuLmj2flIMpA0ZOxY8hGyNopJ9vDoGx
i+Y9Q8Ltb8bsU3o039Uj2I7XgKtFxRqNSch0S1yYmi3MgsyRm1cQLq6b+HdG+If2V+2hLRubV5Mw
1SFVHKvskM1oTWC/k1yCERPQqlr/7fDjzk9nQX/BI1fpWcfvHw8AEaE+GKzhqXhY76tbli56fap4
Po+qy0o3S63VO8rWFqjvilQ1/m8j8EfM30L0kZdB2grxbN3TBGXzo+3cDDWZzxfqXpxNuNhLIpLY
RjqnwrL22t+whwYUE3u8DMFKxqUgC8zVKfgot+rF+uQ++4rulo4XJLTUJQsvo5zVNtnmllSS70RY
qmQtBkimGVAbTgRhb1l7vjH+Sq3kCvKAmHeAtDpURz/x1sZYznUX199UtJjK/BZ+qLOftlJIex5B
L5Fv06ZcP4UmhMQPvYek44Pfu8mY1kx99NUgA2qxsfWD4hsRRbUYgeoDdLdNdGx/d+vQgzcvcvEQ
NsPyQ7v3f/y/BYBqi8bJs1mArYYddx0faQF9ttLS3cSAUuEQv2gzy1OKUHFwEuS3LuwFS/xrXRGM
RZU3BWTSK8f+n5HEkxkECUIrvqVh5Q2zBB0su+lZDOaEvGFzchqwS/BPz0pqdG++nzL0MUp8iiGF
wxmY558Mv3EWpOMq2+N1eFVOIyWWfhuFEnIiaPWauGIDd3MdZhy5+pA3JMbsS0BwasdfKI5tEO6s
Bm23PFyAXrEaMe+sK7ASGVHPIfkXLpCuzyieALu+yHpjq3HEbdj9s4aOBtYov3vwpj0toz9trsPt
fkKfgpLDN3sQX2r4ImEehQsINUHtFvsW+jOd8ST04xQXYg+Hi6lXTKQBrLPlP9K+/w8bPHmYCm07
feYZYJerh4w+9qfd7G9pIQHE4D/ysaX3kYk0EtWa5spWAXDLckyXI6hNfHV2dnsCS1P57uzb5loF
iPxuBgqZ3NsTXgf29zwvW47E29vuICdOhWNxVFsX08R4j2ismOhlrFK+5mXIYVJ+QUI3Qy4gk3+x
6KuZttuaZ5tX6beTWCsCczeVu5zm3SLrNr3RMoEQ51VG8DaRmXUkCSwUElljh3iDxfc7Wy/USD4N
Wmbw2nzROSN7B/cQvIQ7PxoM9Xv0zBVpin2izEx99Syy5jkK5MbNukui5CJoLFV76BrMLqE+SKwp
SX1fvnTQ/5CldEWluHWAKe8h9aJ2dMX4wTXFtmrWQ8D+FdNvycoU9bi2LpTq9hIui3SOzQJNEgaS
Zb7dgVSRO7N0DG4UJff0mvfqsw8PmuiC7gRWNCArEi1t4TaKutgnbbb9+dDdNhyqP1gKzpqLbpwM
EiwTQ9TPzdF6bHsdmFgBSTMMMWMLk7BvseLmk0USRIqWI2zcjAAPPxjfUeWt8a9NcBbUhLpAQNDX
dAQR2h0SDxzvIp3ny0uj7FJySXlEJbT/Bfcgk+xJDmOaYDuKB/9+01EcvAxftahLeCwTy3YPvuA7
5Bbcu0VdBqym25VvF0Me9I1/XmdgiIGS5iolVpF1VmpYdBn6s+sbFIINBK8H5EaejFnCgk7DI0yf
+DEfQy+wpsrwnJpoWYIsK61GIzLV6hDZt9cbLFzAkYl2OIObPs01aA6GnmXeE5XlKRPc7znbWJTM
GfTCIOLkKQByg4XRJ81ThjMg6Ze4KO+rSUUbhC8Jgzxoo5mT0Dx6AqvBXY/0DeMPD7tPiqM4cild
aRawPuZho6Criq+qWk4+FRbFUlBjs2FschWbV3+GuH5+LFNGZPlFftFcjML9Lnh5+xXks6Tv+p0U
xm/tzt/Jxd4TYU2raXwJsREQ97slA8o9jig3KbK+4rYzYeBuX3RKPC+6quFu6ehdT7ggpg5yDyhB
dS2Wu2v7c2IvYNMgZg71FfbcRMPyBFHbh6ZehlB3isGM6P0aw3OjORYIcccVkqTmS5G/c3YdIEA4
NG+2HwsLE25VlQn7ERoQC9DQj75Q24CjlJhY8U0hjUGF4zUQDuPYaqIWV4TDkuwssAWJpWB/4/ZY
8ajSkwCemdNmwTgPmtMwrrBMHmo+g0wvTZN8b0CIwFO6sapNzSU2XECqyTB0zy0vgGx8Oq20xriT
+7V97HPwQ6Y1WHQKrnXuEKPd1tEcikhXgWdXl5SbQsE/PsWQ6C1TekrJfTUCMrDmuNINZ6WhGQMm
gAlHVPHesxScTkOBjAfJOE6VzLI0t6oka2JXFFDrUeCQXFtpqi/EveguS7cjbpCNmnd/uYAPgrEy
iniycws5TwXWlG6Zfvo9gnEvrQoMLvayMwU9k/kJ++ulaLcgQCGxm2nl5uR69Tfoes2yfRw8DAXn
9eP+dTZTdaC/+1B97POYqFpUe3lEByihI5D3fUD5515KiHxQe6QHXM2I7NNCwLKfRIlzds363IDp
swRN7vfVGb22b9oxGY34iGStC6ZPOCnAn90FVuTEfm3EPNeIwW1A6IVnuJVSVZniG5vCKsQFN9T3
vFytaU7yM7dYzx2YuYyqMLOlGeuIuvt/B/V9ebqyuz3MYS6hbdZsUPcPVhUhK+Tt27EP6vq4lI2P
TPVhSd/RXySrWpmuna9qs6gDj4YY4mE8GZda0Bn88LDYiZZKL36++JjY8x2Z4E5myQ0cA9SE9zCf
YsnX0awLQYYJr4FmOORBe3ajW6Dz5/h+WnNvL6rI+fKEC5c6GF1ovI2t8bPqh0kbeAOHIS/m4e8A
rkUhfXR+7qmRrgipuAn9g7V+7xyrXlJv11l1EXiNoTHV2/xRQxHnhUlSwDAnfR2d7I6AldoTmDS9
0/FXR6iNHwfvP2kxOozeRT+TyT2kUwuiCPdBtmXFqYNA792NwZZALf6YAoHJaId0dJaq+lPUbzBt
EOuyRWXRDn47lDQB6C+uQZ3qcmD+ezyOBk8uonUykBzEHlK/zUsXc/c9Q0nmRxKaqrKI9UgRFmGW
DEsFMB3pk9wXGo00ofOYLCeeHwDfuC2k437TJR0z0KjXQIyMCEgeOSV+KzYw1kUe+Slni/WNIW7i
MK72TlqUwsCofRkyJXR6zoUSxd3exP1nlRFiK23XXmhf/O6n7kwyzsrzipkfo9/K24YViI6jH2Df
W+3hrwtYkHzyv6LShfRKHIRlvFgpuEc49qvuhvfJ+bJSOv/CJsWYOZsJvnNpnMB1f1Ff49x+5koY
fssmWDJnpE0EV5tS3kQL5ZmugocKmGHv3UO6wk4wba4nKub9H3n0NUFh0lhjCvQEB+0CiN+w82mO
7dGyJmWCuizJOwncDRDI7S54ln0Ia4Osxat/45JPrHJfVCVW2hu3Qnk3kIqQCEfIayXYo/vbPbHm
0m/VYkNa3vbDQb0YVH6vdZ+fU/P1i2KDCh0Virdf7Tx5vjSDRSMo1VUJEsA5i4v2/yJ7kIb7EeM4
GcBRxzeU58NTg8kt+Ynux7hxgpNSn5xbzMosFWqzTi3f3BblRtaOgm1zdd8zRHdY/v+im9V9LZ9w
RCnuN2tjLptbgU0otdJMgs9N9dtxfwURiJhSBWldZEjn+i5A58Yz769meNk87qIwm+aFHwo/aota
s6LR8Yl5knR3fRemaNZ1cKwcq4XA5hsv+RBIho/sXX17bHUtBryGxUD+e9cD+5DHBM7xWPceya9z
2KOqWYxhZWCoxX/X+5v6o4/21F2pR/sPZzlhAJRDcN2b741SULMkb7AW2hWyCWONw5MunBrUFeZQ
ojig5KMlDLXQk9l3UkjpjZTiWIHkPMhXwzCwm0oVB1mvFSUiyPAsFpM4w3k0IABzZXBbjnHoXXyh
I/FhfB5KRcVUohNXEWMiqsH5jrq4uK6g6UnpPSEaVCd9Jv5YsneXMPsCZbT8HKRs8SUlmLlvu+Ob
3IH9jA6jGmp67LoCByk7FHKDTCWBV9SKt5Ixy5JvvON48uoUQi2MKf3/xVYR16iE9ycOh1NmUd3f
z5UVEs0OfS29G3W+iz5eSTbhEEIu0v/AVd2XMsm1KSdL6zbcf6gNe47OWK/lccUWmfjhoXs4Da3t
t8/FRRPJ14SZ9bxmTNAlmfIHY7oNxtpTSD0TltgVDc9qHOYwQdZe9dyTT+9scCJCPyjdqjj+vX4a
BGatv23/7/rTiyN2Bo+ednewYugsZD5jaPUmxsueOR5WKhsJkKWxGhNpFuuoDDALRM7K2dDPe+eY
4LzNTt4tw6r0QkPnjf35AJX3S3GJUlQ6zDMmnsVlaqGQBXfbfujcXU2kwJ7q97KAXLekefRMr57T
+4nPlfg6XjJvPHoNHXvVrItjgTN93M1EkvlFPnwLfL+hzH6IItJMI7lSmhbV6q6bSDuQlohCP5ou
zC+lZyp6QXJjZLj05bmfOgGoc0ck6CghtjDL7ViCcsfB4k4V86aJT6RxLpk8a2IZAGHsb9R+ZGc9
Lyg0YuYQ7f0i/M8s5+2MLyj6cv2R7ROuYcWhc1dRqODxpNQ0H2iKUiEXQdyXz9UgmRaPe2PIVLVa
4huZvN8GccMSxUjA7iUnkoq9uyl5xwwkdQGg/Ys8htDmnlUT7MnniNWNsb1Q0nA3Kbpg03xCVI+P
OhaTq1f78adbcWZ9Lo0smFqEdboWFogqAvYysR1T39kFZpt8L+ZWuUf17gUDOOg06RDUcQkf+Nno
RryPaMDlNv3Wo2m5uBebZOB948G/pIytW4NKfFYu8vObZV7Ksjf5GXpXQnNgUiZTdcNpJxxmUPPu
MUBQXc/3D8irnkYKQ1jSaBjIC7dX05QOey9njFn117+T+o6vdfr8H9t2PeMh49NWEgrNPlBYm2Ak
b9zlUjpOs3ykY8GQ9YvlFXe19PJQAHuKqZsGoFyTPDJzwTYTwO3Z0tYXam3YvP5nkVmP73a8+I6u
CQpF5Qspk82oy4VtTkQaPdlf52nwi0j4BsYNUJO5FhfoSRJJ98w2CEDwCODv8vHmnxg8Ly1bWK/G
ZQEhLcYIdW4kcrPtY/EJESXjxhqojJUr+t8VAKM/qdP+5VwObe7a06e8K0AahC0if2/0q86SbJv5
TzuP4HyZxd2fud390Fotr0lhK5qcnkRbxOWQl3jx2g0IxCdf4nGIMYnsQe/+Eo7Olv5DxslJEXZb
15uBdwX8ufh66TUyFnywCQIIBO1Xn6jiEX9NGtfz4F5hlIiWbD3v6E5YBYnTTZWGfYkPEZYjCKTW
OdCxbyRivuH2ZmGaGlOreQJC5JNh9vkuxhE4DV16m5Xt5Snl71AqRjda/QFbDF07u5c8O/AAHLkn
y6mR4Y3Or+jddXvRYN5bOxMU+8dXODKZdJ/0yNmLGKi9lQViZTkq/tuXPe9yaLIujabgWGxJVvxX
M9Atm1JK9xuIWNZpveYBk5dF00TmoPFPLZF0Tk7aZWFkUH+YbeQZQSef1yfYb0IJ3R4PSpJUWMpL
5yS8fuika7eaWRyyiJIjTVnaqZaUV8wazOFBTlDSyoy7oAZXXX1E2R9EN3TVQUus4OP6aguGWQAK
BXWWuROyR3EqO1U/06yjreQn5yeDvVzT2+KybpZ1arbTWcF7RPv2ZqDwWKjT3Zlb0PMUEubLb/U5
dzHOeTl9Xhcq3hJNOrb9jl4+EApKZKdavckK4q3zi3lVXujATcp4P4WOGq11ZhdRkP/ts92RElw3
TmG/xclQb3ttKtPW45ybV/nr2x4PwtvwL1GemPEcDKauX8jyekWWT+rVKk32D5pA6iICP7rbj7Ne
jk6LXwYw+a7EA5P8NPNyHavN6msDyvsTLywd4NxDOlxbQhVk5EBIBKfaZtaw3Rul93ulnYTO8IIM
7s3pKpZUgSOxm7bOmbl1Y0I+N2FK3dYCNK1rjpUQrh74Wz7WXo6ja+N6ZSbQC4hlLnR4IC1OYxeJ
ijShmAUbgO3xSXsgQ1AehZfU94h5bTtVM87nkztTA5QL7HbJovuJ9yGibuu2238o944o0Z0gGcRK
8Wnv9WNatdYoEW+z4U1REUjRYPJ/+HuMk1qaEVUWYaB4u8uS4JK0rEAbbZ0MxFW5oOmS1HyYoR46
IELXa51p9dWFeuUscl/aevJvpmhrIIwLEUOYNbqqCq4AAs8I1WcKMQD+vRDfN1St5a6oUWqrahcg
ucqt6uDOPCj86nMJ/97dSLIhWUhTwbkxDOBkJkOItE2YdNaGrLxUQOpYrsCpcITQWpOI3xwxWrVX
7Nmxig1DzoIqHc9b6azoXydc4vobJ6vII7v2UYO3bCCQa6cDX9iZByFsrLqE/7Sbp3ugb3FqvMaA
qPDAq7lcmpYLKgK4AzVBLpbPMoI1O2zVeW2x0hl15g28Ujvy3akMFABMMuSxVpxk71jQwdeqA5vf
dPGHcQbb2D0kLmNXh82PG5hb/ztwt3yeU5jTikkL5p0fOlQAGwEy2rwVcY5uTI2vNdH/mktUexT6
Wubh7QXBb6n+Amy4zPFc39j0iSfbT9RdUSmh6e5tfiUzFtc/G9aZH4X4egHOPNlxSo0ZAC2a9r33
444EuIuLo/8mirIo3alqHgsOT1XHEaz/fCLF489o5+KbEoXcq6KNW6h+mfIyIsG4y4SlYU2fIcA6
1wUJ9hDf1th3BHvb2DBpy7B1bbJ4eK/RuDO6LiAbg9K9hzL+GXrkRLRFfV//sRqeY3UKDLWG3S6I
ac9uIm5AwCWrHqBwffHIc5Q7Yj8A0HulC56jzuosEGqlNQHr7ElPNZZANNOfJnjB2QXi7CLUuOzA
mWD/hebRgSe6mfAStSuB8j2J1atliuhcRYUxJ964Wohv74Vn5A+ciBGEanyt+b67HoKLFPwRXSll
VDgNOZb4crmUm9P+BvrHcc/GDfRORqFuOqaZ7VXasTO5I/WKsNlFWrsWMqwqVS+rdvxY/lZmDPAo
xgX2r36WdECetu5KQY5EFF5PPYSqgM1JGueSiIgQZgbLpZoogM2KO34x7hqhhoydU4p/isjm8L/a
6KqePh9DvmsYULrRc8zRdo15IImXfpkw5StDox8A7G10jpoQ/NM5V+8VTagiuC8CWDOPTLEr828o
QCARe+BpUN9Hrt6WKnWhWs86nu2lg8gxJxhQILYkzD0KlBBgk7Y2pAoPm1mGeM0bPm5sGdcHzcFU
88eC7slncsg/n/vZgBteWqwRW3240loHXd0X/UGD21XvYzAJ/OMrHIkHeI4XsCs3k1pdI3+gijeU
7RtXH1sobW5gnTGORBSNZ3210RsrzrbbPmq4k2W6H2Y2/jNQ/cnJUMLNKMnqTnnk0NSCj92/96LJ
IVNHbMbn+fIjQrP3p7dB5v3oHKa23wTE4D3ob4QZU5MLu1xB7zi5pEY8eQt4Yd5rvZAE/vomG4M8
uZSY6OX5NW4DGeb48SKpiITidAYG9lDVEpfinRNKJ7ZxG+JHPNTvzHE2eeBY1yEnnugr4p8jPDcX
qgYSH5O/ZMWeVAT/33K2LjNJhjKu7MZzzeU6udUpz6CFf7Q0fhU2ngZxzxfD1eOFrUXJFZbJC49p
x7N7vvQNKUq/SUDaOSHL6HgjsYcBNeCMgGybnxS8uFjzUs7G1XSq4nGP3ePfGj4tmRAorjm7RPPn
tFGLRoE2enA+gtTZeJqfb2lsBQe+kKyoj3MwChePcCz9vYcv36WeslNqksWaUCLV7gwf389CKyDN
2bbuVlrB8sGWSZEyiR2ylF7lPBYLZwFhbE+3XTQ3PLqJEJ1iMqU3dxPmuorfae/ryOVIb2smpvJi
kA15PcnsB2o95K6tNUnCAqzct7KtZzl7L8+3ebpKBwIjHKNvB+W2UlBRPX92JHPdnQ3M7ysZCNqh
F/MBqAc8AK69VfHFK3Gmo5zJEnOlVeShgJrnp+pvLDAzpln3Bk32EPbhBll/UiRWQ40V2AoiQ8eJ
CYhW/e/CStdgIV3BlSJCpZHNRjf3ymla0xiPgntW18w8FEVX9ROXCBZh3MHlMSmlRlIalhFINR7D
lYFSBfU49ZbNTEB6szUp2Y14zVCE5rhTS26EiQ4z0xuN7/vnqjwvKzIi+nJ1ezInc3ci/Ed0kZnO
i8R7AFxYImUWD47n6FfthTpeFDuw9JlnmVjxUZlLpJvjWKjB9je/ii3OcW61QglHs+V1P5EwpYUv
3dOJV50EN8QKf1OVH5eOhYurD7nKaFJEQrPpD+kDPm/rSllEx2aDiVIXo8O9i3+iVRdq2hAqtrvS
i0wfAjtb8BeouNrqPug7ICtuH4BujXlrvRhbb59bnqi4UWxA42iwItcr1wxyMOQmahedEna5V/eG
QIF2FSovOzqa35jZ3cLiaeTMxrQInyfNIJWXEBImdoLcbp6K1ODCNyQ88Z2b2+pcPVwDoiPuGKG/
UGdCW2wIhZVfvLlgOQh3vsZ15CFqiJ+6m4CAKSHBN+rtevv+ARx5WCcBULEdgUz7zFymXDrC5F6X
FRd6emGdR2vnDfi0lEZ0DvDo+AuOKR6k+X4+1T32FxZNFvIl7c727DhnSg0dhLoxinViqyFawo0I
I3C/0iPLGrSUKdqKfm2JoBLlL2CjW0Knv3llc5bXWwM73FXk5xmr2mRtSn4MvAA4jo4prp2q/XNZ
SmUPaz8ZG77fyOW55priWJ24rE1Symg9ve2q4RDzOBP7CDDR2Hp5dOCj+uOtNhft7ZoN7tNER8yU
0aZHX3k727ruejTYwNbR+FPCN1PtHteuPJJSOpec7brAELeR2bL7uTyp3r345jur5MdmrXqvNBiL
tqMHEeKkyo/LnFtT/vj0xCRDJB++S0zI266d+jdDbFhzzlGLMOWE/4XkD9Qqx+TlqmWU5el3d5VY
KMY8UEe+I+jMe2mcvj2jrP4xrpc9/PJywnF2P77UzlMHuMk9076290ENivleF+MP1SaHjnqSwO5X
bHwJSEZsJGLRHF+AySjetnZl5i+18K0CaPG9Wd/THE1zyWr0QmwOWqy+ntegtIDNA+kelYI1TRsG
1XZr4KpI3+tLgy1qs8ilbFEAiOk43nzEWVjY/7N7uoQfjt9ssAnpYRjAE/Yb8kdEbBj2ZMdmRhhX
mN6jePNfegjYAL9PzlXHGdUHf+pC+q6JnW6pm/dl9cWTvEk86kuey8z+nyJjkEXL/3WU2zRoU9Jt
gLW7ky3aXiTfiPnIoZIQ0SNOxBwEkktt1Xmm+SDiesJU0kkIa/jMw5Uc8H+qLHdHzpzFDFhJDxPg
1TwSIA/W4Gg6EAHhdJ9nYvoGHk6q852cTqpJvwBO/jHIfM6bMulhinc8HmHZivK7Z0aPUzpvFdlH
RjnYtdg99xK27AAMxZPkKmNMsRrrd+qbFa3JubG7gO5ktkI7VrGRIuNgH2nqmlX1Hj3wPFNgxzCX
EtEVWuFqJNQMDF60OaZV6WwD63hfgc8hL+5qIpSQWVG1sxh9XHm5nbkSZErjtGmETFVES9XRl6iN
hvOTMQ1zqOup/3m0D1PyWU5SqXCjQ4FbK60mYhtWRe/WabMRRQ1m/BynDr1CNw0n2jNvXBsIpAP3
S+/g4yOzgc1uVgnSe7F0zbx7HOGy94L+MIxJl1YzNM/VGSKEejbWw9AcnxOPWdPoyeLVwc8T8xIN
vJbOfs6jZucF7hmG5VoPl0c+SooLfuet3mf3R3WZujFJ42ZsMhk9HCrADRAMMlcjIbqOAsdEp3wo
ZothZxC70jySXEV/w8LCnjTSID6tlOPwGzs9e5ArIYoe8O3fcQ+VZwkDmlDiTZF9SWSwX47mr2gC
LZk1q6gxoLxyTxjw+KLcCuMQ1Bxpa+jTZZG0ijtp4MaYH/jaSNqKCC36v0pkNvnjj4nejiBbU3m6
IiZQhMB5MWdLd5STHGHinxy6LCJXmCOaII/ykAwd1IZgKi8cods+ru62M0LxqV/i3hWNUGc/A3nc
2F3KBR1nDUeaPLK/wP46+DCdnvs+D+A4P56qC/Aq89PVjTzg6Vqcp6K2X5Ok2ds4kY63VoXPlxov
aCiVP+WTnd7m2SAvqEYUFvoHC4XGzjJgztvwW3mBip7fTIz399F18LfKLi301iUz95O8sNXa7FSA
vPBVpI2jy7wDBnVbUU0mJnmEdqahCFv4WZjCBRfPh/sJMZVi3S3Z2gQ729r/OihpJHTUfPgmCIb2
D9LTXZsBkTVm2dAYNbhgT3LYqCWXwLl/0DZhjQgRCRAemXkO7BS/ZSpry3B5uioDgivAfK38xx2b
Sdwk9YGsEdAL53XfZyc7KK+IFHBqV3evenZnV1IXn6nSfbSdpXoICEmcQW4XVcqHwMl8QB4qMrjm
6LJMlk3T1hwL/OxakYXSQQlsZJLPLQiewAiOOONunYyoa2B5FoOf3FPe632cTDm6Bdrh83XpMq/g
OHTalNuZHwFDeXPL0DaVxWeoVp4E8lLuGrmUmY9JXdyUGnyK4RZTTxHI3LFedtKvFJakwiBQ14pu
dntNnUa0vaQMkT4gLznb8k0dRCnXxfo8/Tn2ucc6kmpU49+OkgqQJ/GAC87XU5CdDjZtJQqh+MN5
kHHdqVK8bS7WjRSesBND3uVg7Wu4YN8X/CRcMfdQ1oJhpbzMPwv6qhInyWkTuJum0RjACLX/YHD0
1vJuJzpEc0OcvnT2mP+NcS35ttXG2S973NbWkiF/sVlv6lGVfrHIifwUoOn7xgwwLuB5RHNsmC2L
mCKh+tikGk4p/eXylCqBGjEUSDmFm5YAAfouZRmGCMvfoe3XUBfCKf9Sd2AhQXuo+1ti0Ty20tC+
9GoXFrTAjsr4QwlcgsP0v/4hz1r+EHVrQXPh9M4TnLpQy9tYEtFFJpDXQPV130QL+rAsT5C225xe
HQort64WX539I3zWv9GXUgs0c9PeJ2tcoOKpSbYlrNOd/rnFaWs24uR//iSgqwiX0Mm6s010JVT3
K+XdvtJsVCQfrO3LuVHLZRkuzmCbkbguT9qVyiyRY20PzYBKFw+juBZ5XDuSozmPY819LDovYTF8
VTppc5aEFtnqIpnqZyBWEMOF0Y1PUXQsHQoRgIaqy54bCDco2098aB1sfjXFwGZYkAcsjhm3HWp1
ZivvFuIWB/5U4HVh+KetORZajP8w6VsHheSr0G3BOyEappfX4zIC+D3B61OYB/NF829A+Gw6kfpV
R3kDzenJRX5f8KydqjxWiO4YMKvw+bwa7ycFeIIG/ahqxRePa7fbcLvInkvIvbeW5XPhnKoOPtN2
jCFVbEWLZNqWpuSoZV09rLdFCR1Lo7MiSC5RZaLfd2uANUo9K6HIGdx0CDuOuG9PpRTLy8oZcTIn
ChUEaLRTQeRI0/7TAxSFdOc+WUjG9DFFjVsMnXFXQObsaJbCwgFS390doSU/2GsdSC34q0+ipsFw
/gpppXistPpsTV/hFilEc/Hbd4HWKnN0hebmC/ff/uWfcwLLwBhoMwBRCAACFukbseNhoZJr0kxT
f09LeFqszn8ovldgzDRR9IpnDyI0VdW+VlwAT7lTHVPkvIl1Myfi185YQnDLp+B5BNt1wp0bxEI4
4DY9avChF50cedS7Gf61tOj9uVYDAJ6Arb+wHsai4ivsxc68Mm6ViLWN5sfMNCNwh/WS4rSjyF6V
4RXiiRoYB25rBthEwMduP4rPqHov2kczTrM2cOxVOPXwWEa5cpt/3C3MYGI94rm7V7thLnVc3p33
4noTWigXmi2LEkMv+SyY8aq5pH1yilcvuX9763ZaxvV1clR8oL35pvDjG8mB3WOOUcKtmhh9I5i8
0nso/lpSu9Unj8APTUChvVpIDleDA1LZ1Y8HjlzRQ/kYvMmfm4iIQUof7q7OP0jKwqJEFwDamuOi
OehOPgPFJJGHBBhqvP/Ip8JSS0l6H54cIGQEDZgByiYWLSg8F6JDpKvPM9khdWw4mEi5t1m5IJkP
yAX7TFhM38TTDqhUftMIQ7HcbNkJLkIVYZWjEd7dp2OXqdf19+dAydYWBWnVwP6NN64vP9JppfSN
W5+O13+Fb3diUQ78H5Hr0HPG6DMVagNWO0N5e/fpQ7e8MeBurpRTV2djOitGrUW8+vgExU03S1zk
k0f3uRAvt9WRa/FxJ4E670tK3JT6wqY0ZQc3g5FV4+iIy88wxqg9KKP3bI+oTH74vGJwP+levveg
X3LKW/Bp8vxPqF16onWR0EL8ajYV9jCUClhQJmapfwmARevbTOdHGUoWCrI2O3h86f2ESHEAZdWZ
pG9R09ta9HgqfC+ZssNRwFCAkI78oA+W3wed1UguFJw/3P+OSgbAMrMAsxQIPPY1Ozqk+tJy9pvI
51Jbo5CmKuLB3i3VPxa2Irkjlv4fPJqNFvykCbzW0zEjyW0UfZA69IGdrVhLDp1ILorhr/hl0chb
b/0SYcJZ8gxg+ZpFJNU+U5vujP2wIs/N0AmyWFDvAe9oCjj51uzwtpMfCOT9n+ZRy6R26Offp41a
obawQ/trzX96lbe1cRFQHdxPt6g526KoP7GW5PcymWRSL6miWMvJ4/KQAUqI0GQIMtfO/znLx7bh
8ap3kBOJyitD7W2wEa03CnRItabzDN7I6pN78BUk3pCEXssIGq1GSIZMFSfKIWHv5Si/2H4tzqYE
eDplP4MGHUCRLMP/jvqo6cJYqi4SmLd7+Qq4gnPf+o0vDnXHIFKJ1xnRgadOpdrn4393O2pSm1wl
rRNT2fcKja7lUgFl1eulrKaBUfbEovpPoIgCsbz3msUJfpYCWwZDPO0gDRGe4KEOcljZIyiNDZSG
j2N3Ucv+Gfes74MKCX6MeRrP9QiTiea20EqIIRcD+1lupwG6+FRsrQkecGMPd1C0E7kmzGd4uWZf
uhRif3txLpsNqE4s5iAj80WkBHvqYbYxfV8FQZ35CQB79PiDp8oStyr2WSHQCuPzcJEwU29U5HB1
+wFDO88ttGbTKiaFrzBYP9K4vArzUVqQ5CjTMj+tOVAaJwVTchubQB+QMdfqVRFp7MtJGAou/qPV
XfRbeX2A+1Q1Rr3O2Y/cFefSVH7cqqdOwiT1AbgQbB6UZTIBDoZn+dlOvqXHAvc938PLsngBgVBi
ekZDRw98f95yUiPnzZlXNrtiZj+1Tjv734m2V65EGeSHtfs7J7fSJWeRnbYOT9EsKxSBv8k0vqON
75NCYCt4j8jaUo9GumOZU1jeVyb+HJWcsoOzcIBYqen1a4C1/gCupVq5lB9vmjXI1NVqYQIOxGAM
bK+SQdLKUvfhIID0beKNREzGN1gUk0Qh+2z/wPoYNvD/ADnKBMDmF7gUPamPoaL71uKprZIlBscg
I6y+qHx9H8Eb5wrpZg4qlnGxfMVsgPbSoJWgsrSTolT4Mx65oeYpw1+rifMKKmyoMHh0snIkka8k
tZvev1gvb/FDQ+xvbpHi2bncjSiwlUrbazWThR0KdsYkIy66k7wCV0M1bIbkNAnIkeo+F9fgmuEV
GSaS0E6ar1DeVjLWtf3hlmfy9eqPLSWuyEolmlvdcntmLfbAV1Szq5DgSknYt3ztLQ8Nb0qW6uzz
tOLnQe3+plWsQrjryGFeBM86o/axbQLE5JjsIqe/Jz949oKRxBTA00dJ+EUXTI/vWsN2rywWmCWP
fyJNcLLfMWmx0GNOsFBMPG50Yz0N6BFQAMC+hzRodR8zq3GI39P1drm6ujeTFhwyhMH5S20fnFSs
DoH9Zf/wapa27IA6SZIflf0VKP4/feNJ09BERhxPSNLk149NqkIohQYcvV54wSBpZtLsMQ8WhaZc
UYIVp9IJ/h1+e+ZsSX8UezcjlhP3mNGpoh9N4ldaWT9yykuFhtpsxNC6T1Suzez3W9T5kcuJsc7X
INaW4GZ8UB/smDsMFUzTXgXC7oxAhFfUCdEZ4q+zA+NDC+0iSyz8WGlacQOkKhdRLAKZh9AxmLgJ
p902ZkiNdAaFvYHlqcf5nnEj16Avilelc9+RpUTY5xlxDRZlYfvnurXnh4NrAMt37YGwFpGb9+vz
0kZFuQurDCX/CG3dZ6evmt2wncYCrSybp41XBzj0icpZbNvWouzS+8OjBBy1WPMEs0L4RSe49Fiw
6HooINW4FIrcUhZ1X93CsWbLZJpMk7onN71OgoLCpBK2N/s7KIKXCbiehtoN2W90ngLqHeMaNXwG
wzYrwqQ68b9bBc0+eQ2eQbb/kT8+MM4tdX264U5EmBngV3RvyVeSST9pj1Rij846O45A4VwGYxkw
k9btibfFqb01qASZ4XswOOSjNCvBtC1k2gTcK6Q5rF4LnobjzEvkt6iLADEE8LBtsYDIQSSHSeWL
241ZBuU9dozxDIfizHFPmC76muwxbjTRYTb3+vSJPKa2qUqT32gJCFRo+SBu5VNm7nmzB1mj7VRf
DRT37V8qTuwN8hzt/eP2MPgUdkYe15IoJvBm0qr8XnauYjjzkVvFEw2nY3/YCrsq8vZH8/pCgYLK
s4xaQPVvCbdOOdAfH48ZoqxoUbzjieWANyhzWd1YMM9C/llZIXO4IU1KJ/zG+TyYtu1MLMBkn3tW
cVgWo6UysNw+0oz0xqOm2E0BEAfg1xUkqqlrZeDFQbEyTWwSrwHipUIFjht7zDdnmXyvkJcPTS2F
rsa3udTCdeA0346nlLpyfVdpkBM9Z0gi1q3tqVfEGdEh5u8oS6XDIIBxsdhn4mOpOjdl7HjRdl7n
XLsyNa7PhOTjflnuIrvu1mieFtHupsSco2ohTrnxczqEpSBW8y2mcZUPp8721FnVdJ3r8gi5vPkj
/puDE6ijFSSWhOC9lhRmH3WvY/MLVBln2rEa7105eOT46ZGjUnr75No4/2Ezf/ofzl1dvgucRFm6
Y1rCgbp+wCTTLvDDrSCDkUg/vyf+gwSeSBJCQFxoqc7KnX9kru/rLdVLrY+x8q4lRl/Bv7gNDP0G
OlT82B6GKJJtwyPikftBQZq7q/cTJtK+fjpaER9EAzE7CCi3b0EHdqutJ0yYAQfhffWVrLF9apaT
umrWUXylFZNF60MavKuW3Ez+XtiQrOxx+u8yBQeYbOFvxhlMTOMvK/cRmNQvADioll9alUun7L18
b1Uv8xJzCf7IeaJjl0ppVY1W2mc5OLkIhiJ8e4VrKIUrI4+sBIbNqCGZ3eB2PNqHDrI2/baiShVM
xZ/Rr0V/Xd86XCW8J8I84E3vcq9TXSUQkaOMctOQnrSnyM0w95KKEI4alVf/lH+ttgMSeJ8s/iNN
o6LhA80dk0yL+apSvf1FtnhVJ0HEwTeQM3tCgolCzFCMM3AXa/4HYmFzmcL1+cHIkIp0IyFKWxd7
KvqJZcR9kTVcxspX3/66zzhPwzbVF7Fc5Sxo9fXftSSvy0qN6yAIKouJZSqotGZpYkBSaM+ItkoI
wEzKc/J3hZjmfEWux5TlVxRU/ttfZi7aBf7C637mZ/fypsUzTt6fpANjTVfds5Lt4y91vOOhIjdg
ib8RHdcMOqwWUo5iSwplU1CAh70pFKO1wjMYcpYxLXi0TsFcEB6TBdsTtrEk1J9EMtwpRO3Xbsd4
w0pxi5dk58wO7V7ZFe26yhX1QBJXXwJWu8losTKVJyRnQ2izEnsnhUlqmNg8boCcEmAfgFlab4B0
KN9zcLKMZUUdcRUQU5mVFWUWLnODiEY6OsZXHyZ+2hqmfDwLsPlfPvrndNCDAiYT76RQpF8Hv3H0
233WnXgzHr5W+cTN+QXSmVXQr2BQyN6JpeX++am6BHEjdm2FAkUpAJA6xdHXWUyZHjeQADtw1NFV
sfL3sKxemYEgEl89DwGuaCTau5l1s59fT0Kv0YMCXueB6ZWm/I3zp645U43Qf89TH41WGDQBeIBD
0cc4h2K0TuEt1sqpTTMe2VJWWS9VFZ3WgIPsCtIxGZm9jMRqSnlsUIde0aVAR2b1/ECobPJCBxhj
lgYibFh7rA5R1w5rJtoEtfDgIsSpKjPwSwBVICmXHCG0J/agdvw1Ah7midVZAYAnugZOArDn9dGF
+3ofGw6OD1V5XQ4l0G8zNvRWOLkiJxgL6X8OiTxyPAuZkogOYIh8oje7V8crZ4cHHOA2eoj4McO0
c2GTBckXqCPVxNFVBek/ypC18pk8vLms+6TL84Oz76T/2SmcHnEAEemWmMieiFzlAZxvbe1mKpHv
tK7kPV2Zf+ArQ6lXLAj2099kxW4rEBHRdNNCw8YdQYbWmIqlgQgb0JDbttXQGxRhHorhNO0XiXnU
ng4LPLpTRpPBCRlWGSE5bCZOzPz0GnQLu91rqWRGrn2BwWW+RMPNIRtvdtQCsIpHGKj6a4KofFF7
OFfFWcEUVJNt5hoRBXzjkqgn+mngHtSgKFZN9Dz1LWgMxjyM71LfAWxKlDmq7WwktApS4K2x7qIe
Y/BPFsU6CKN04U/o2qkbJD4HcolkZlmJxFBPfGkCIeGAaTK3ngbLwYy0bXUmn53wiAPJI3A7uVlf
a/LHadbqzGmhwsIruzaNT6WnEftOzdYAX0rteuWiCvFBXvOi4h53E+a5oZBlKqUhKhrHUmYgvnpK
6yZrjyDXEVIFoceVswV4l+4P3+e+6C3vVS6HXKx99nbXZUDvi3uPr9fuu/v8RFkiV3Nr68p7lLJj
PatvdOhokFPOrkek8KbcKSCVCwGMT9gounxmWqmdIQU6HPmuvO4+I/UZLaAN6Y340zFr+kSO7WDA
Tka8wSomgqji2ZF2lWnbdnTwPwQ05SM2v4sOQkOzA15yNZmI0EBCZCIJdJUzkwHc3h5bSI9aMqZa
vQc72//TfiAc6QJf6kBwyK5dWfpi91XC4HL+Xq2sbgh4wy0t/yLtbFw0VjWBoRAaZwPCi2ccKfMF
9ZZNwln9e795egtkDkyLWvCvkSpNm2o7Y2trL8flvSeMxT4Kpkd7JtIm99wkm+diIdZqFgWj++km
s8x9CxslT+ejInUVDO9cTIZDUeMhrVHh11gpaABOXdSzPoFdcywmtVkVsIv1CcG38DTUCjJD8jvd
dcJ62hqQBXQemMtSnNM3pKyEdMzngtnThMw2jzKFLWOVf0kEr18zlOnQ7NO6bUGbprf44TG2ljzI
aFm0qS7RvPMF1mwC6fd0S4j0rAsPuPO0/PD0fajkFN6yVw3ukacxJBEw0IkLlrIkgNAfvkT7YmG0
3CBv63e1x/JP0bDPwjWOx+6iTaA+o9CBKC1o7waLiKiSubdxYRIc8Kv/dBPCjV+KUJxvvNCPn29Q
pnnOFFXumjproYeaynML5M6za/2H/QqmXh/UnbrpjDUKtxv1xxmRek1IVtLpDOaMvhupPtl4/GjV
/ZPqyD45x/hL9IqJRYy9tOfLxDTw1DNv4TS+I/RStSYDBf357En8hMV344fEUN3PqYiGgWSYTODG
dhAbHDQPg0+VLHIMjV5FljzDQiVis/uZDfiB/LiRNOJHxvkkxTe3dVdwk6O6GSK/XIgfvrx+Xfcv
KyesvkQs/ZPPlIMBKAhsqkJ9Lng/6lxnbS+8+bfwr+rrfjshCWs3IGpy2el7P82NQNGvMOUAv7bT
ogpznnmU5GyPSzpqQZWYJTwV7jMqXWX1Rch2Ji0wZ+1XmPzudZzzN8x+y44/dNiAtDbC1Ir9KZwn
uXlFsSLW9pxkFj9IitD74wN7j4XjJylOiZ48FzNff/bmWOSPJC9a+S3x8wzrX/zsUDx3K6rLFJK4
WuMcvVg+RZH/DhAqNIyM8avhpqeNff3TULt9usn1UHBQvHyTDvb/hsUlXSKGJaJ8dgTUQFMPUPC5
iJSCdUPRsR9ybXYpnZoEcALVhqPr5pDV6cgCmsGgaoyqE8sfeBSyc7RMs7m+9euRD5jkfrRnrLWp
eP8W36k4kcZ3hz9WSO2l0aUxrE2zOL2MWE3wRu1TnNLcl2HEXujHUiQ2/MRjMaJUub97u3CatQyQ
Jf0mv63l2z+s7TzSHfmN8dKQvO9Lv8TVpP0gB1FnsKLJpI0dozIL/vF/yg6pNTpi/I1p8HwQUuGq
5GwxQ9zUl4yDMLs/bA+74U9Zs+R13Ci7W95LSwZ33VnBZnvqA4qeRwqbllTwVW84uV6L9wGKVr9w
Qgmb3iquczF9MVsjtSBPij7xm/Tcm3g/jdJtEMDmumgFf6ZxSf8q4sxG6Bx+IWs5k6pzXqZY0j7+
8yLqV6fg2sxGkIUz7QL1HYL2n0emX057IsoHzUmRK4RYq2mI3srB6VxhofwW4V7sVa2wDQIlUe8u
5rtfJbbEtZloeqKxZn/qj/EkUiUZRt5oIHcvcn7FFiYixawBnTkIM0MWdwyfg8zGcBi5OxfkOJzD
npUBTWldH2HniVcJBcJcZsLEdJ+2aFcDFYG3DuWW46G/cbQTQdUBWt8W2iBilKRCs4PBv3bTbzhQ
9rhBKyOGXmOzAswJiENLvrAaBXC84c56sR0UPm7Rz1PSl6B1WWv+4F+eXChqgQ7NFUqqu9bFglC0
WsNtJjtJY+jjYFtrr8mDO4X53zMrHTZneG2q+JegdKuvKtTqtKh2KAeQ6OU5l6Xrk2TMId3Qh4VS
e2+jUgZtgh3+HJKrsBfxdct81sVzrPHpNzqmXSW26xPKREDZ8J3P6KXxP4JLPWe5MfEze5wlmPc8
LVE6natOdwaWnuuzyBi0D9S1IZZkFe8IaCayjG+C9mxk0Xxx8H+4CxUntLWIF6890+Kyx+0p8zq8
TebYdGBdza88t/Yi0WDjyXAJxViok/nYnEXx26hm6jDiFKIjis+HPZ7Hb9ubVYZLOcX7FISwW6x0
UAiHAokLUgqqxckHj9XfBYdoG7EY8R9CIofVx3Ns0Q0y7co4A249t8Q4zpzKBm8KgCnRRIPt3Hw3
XOaaqZMVLau70ry2HES1syFDlRvXdD7P2hV2NhVVAx7CwVzlVBP3ZKjPDJGe163GZqrnvWxsNMHb
reCnuvtBlqUZUth7ebQ7eK5L0fPGPi1+5ec8rgyurJ+zn49z5+ZVr+VgSiGjS0ViPC00nLmdI4Zc
ASBAZ0umydGDsjvnuRJNjqrQm9IzC07gYwCDDO3CXljK4VmJG2Q7NKT0nbtdy75K29UnqEDTL+ib
KUJl0vWKVwMM4t20Thv1HUp2K6VfFcRZGW7Pb7TiWrsBcIZFF+wGevCfG+zdbCTEYKF/h6b4RNj1
/8f4I7/Sa4oHrQslP+58qS7PFEqgLuUyJYJqwoM7hZDG8dz3ws5G51QOgZBVF33PoR6VPWVk+BVH
PLUhSlv5blfqjZ7wXv6yGbZZG/ZiGPJePPhYmqMwyfbqyZnZwt4J+mL3ojKagWdhwuiZdsmVzslI
YI894xenng919q/+W4ITIBgu9ae0kzD8f16paE2GUsYVsGqV1azSl+bowZBZ1PM8xS2O+E4BM3xD
95GDMOAwTL8t41Ce12ibHh6nuMdmCS0RBtPzrPoYKK4k+4ywZRGwt5rMboKCjCWJZLpK7q67wMrs
qlugbIS6sCB1wjTP+xrnBRMsUsfmBqvMQF+m2Y840zfTWhc8uV00acThSmzxtgIKLMlNTnvjvhV/
AKyQtmTIRfzCzt37nijxYypMq/OEE14ynEbtpxeMXXllLw0W9wZRpLB8o7JA/gx/HdsUDz97mnPz
knF7U/jr2tALP+taSpBciEvli048k5QyklFmVlqML92tEa9Dgej1SJadLjXzP7roHKbi2M+cHK9X
quUxSxPaSfSn9uNAZ7NoBIt50D7HZl4cTYN5vCGbSija3CqzFVMVhd7FErWdXi0B5TjXGrsmoHpa
jh05vwXhaHeJLE+sJI41dcl+kFmo2oGdzy24KRJ/BlksWG6xRfEmHue2h/zgXuYoc9AUtwio7fBC
oUgmA+HaSHMCjhVeXFYUQQIwjqroECGBiXP1sgqMIQkUz8fu1bcydBNQ87i0fM2yMAnIUdDCKFmN
6W6jGe5DtoIzZKIkxG9XvWgJ3UslE3He40ZgashU2bSmrZFtn7FmP/ndQO+NDnaWNXltOX4EimfE
l5RApUBvdXjfPpYh87Yi5jT2ePldE42MRj1KiEWkmuwEPfYu5JMVkk9T/Ne80wuz1MJ/CqYkt1zF
+k/FfKIn84w2jUXC5HOXA/Mso3iWBD0UEQFIv4CT3+kJ0syeeHmtK9CiOceDUkBCBaBQylw2LfjG
fk9hYkEuWLGWH9D30/ojbQXUcCat81JRgsNNud6O9VR5Q46dFVFuKt41qQAmbCnPHXR0jrZMbrsT
wOwRADa4N3nsd3mDfSz0kt5JABcyH/sNetD1A9AKytR7PQj7Eat03uNZmzWUt7oHG7hhU6KDTsQ+
k8aECHbNoHPjODRmwqjryGu3jPVHdSbZ5hLs3D8whAmXNb3QrV6iz7uJmYVuG/s4KZjzDcx6SXhX
TmfO+0MQviVKiy2FGECYBgag/iQOEjJzPk5a98gdsiq8iwgjv6mcQPsYMZzZqNmfAlRVK/sWGzW4
jhnJQ9yYd+uVlQp1qbRaTNNVNpeAMgLVDbX+Ndiy9uGLwxRLGXzO+JIffygyOILRp6sL8SERCmY9
7sMhWQvk7WWjq1PXbIf8etnY3cEcK12FB7sLAtsDGtGXh/C+aJi0cYGGx388A83uW4lxbMoI/akZ
npOofiTqkDPuXH1eD21v/8A7RKcdoif2mf/L6pfw2vYb2Q/lpmvpj8woI9AX/p7xKAdtUacVLqKb
emWg6te0nzCysw54kDaZsd43CN1cYO4xXPwsG48FU6zOy2yXoZzrFTIRMFvbLGkh5fL1WDIB7lGf
uWmz0Ldc1EtjDfNbKIZOAefE8c2F2dEs6704WDcNUJo2g/cMt5zK8BPYBjt504Vtl4EDAEnkF8vV
q7Fm1Ojsp/LYv54GOS6GOIHSP1uW6jbnJeP53RLLNWFAkH5/mpXSwpPVCySphD8F25mDAlAzOViM
nci+pSdKnKca2eTmFXWvn0TZxu0jbeNqT4GlJPWQ0h4ZumYns1Njnz5jesfCk67XfSQc9RtCBNlC
eTs8ufpJ5dNCCwxNBrrzKMOJw822BRTztmOKQbWjcWOkQ1WF3ZfgZ6PG3fFWtE3gPZxOH4ZANzie
hRyyC1PpJiIOj/1l4URM8lgtQPkb+9RTlDSdNodydxUVUhhPk9O4O04JVDqUpu+T1LVHTJ6b3x0H
WMvQs+nc7p/F1yOc9X2N2GStQxVL5zJ6Tq+M4dAIGgu9SG4eLvcZCRY1/H2kWgCp6oxfnagwm7x9
Tjnoc958/QQAL3McgDFSbBytSQLVML/RcEd3wOzra8GMj+19kb+MOSath8oQH2o1aGPSCj7dWU+A
UW2NL5Ad9FdmLXSO40yg7X1FS55nTsJaCoMesRfEF8xm0xR2vA55ba4nyzYjzlKnCkhqpZSoVfg+
LPHhswqjaXL/19PqQ1dQ7QO4/DuyJmKrwu/ikxhLoCpvIFWdMH5RJJvQ7/gndAfDC1b+38dyV9/A
XarjqVdkEn9KBG61ZKyge1QWVMLSC0lPo3/qyyLcbIJIsoZTD4d+8mPjAl9V/lcsTm2l4YESxAfh
mB1y/xMKuih1k3Z/XCmJSWmn6BmPnu97oFKU/0Lv4tOJRtr4kyU2vdMwuHVirWZfHf30R06bhB8v
wpRWRqAIET04HGyip+4S87hRzcB/mX6PsQT5/TKHWR0UOAJeUQAI8nFzXkTXdTOQnCsxQwFTIYUS
KGi1WnPwlXrkvMAkxPlY5v92jjk/eWJxLn9uFXOn9luEh+sBEw2ygi5BKCrchhgfsfy0gKA76NfF
+aXXoM9UfiCXlm7qmczoPSSmYkxfWMRiergs0Cz2Z+iupoZazXfyhFiAGHIzwXKu1XeCLwfX20yO
oKRyRc9UhLzOpV6ggCYVz3blx1Mr4VqQteMIezaTPeQg6H1qciAHMiYf8Re1BbBbuNOenYGe7iR8
Tz/yoLPuiwBzUwI9pJYM5jguiumrKYgQNWRIjpal4y0U03mBV8QJP2V75+BzmmwgECoRbW7kf9kH
Uq6Z46SZsyUC0Vr4klHCsyoaBDU6kCCdFKe8ifeF7rhzOu/Qt6ZkJxQni5e21ywBVRKGRC3S55W1
SwT1XmC536xjeI41ZD/WrOirU6B8RDgZRhl+BD9VdxBb5EEXapzcGYmw0BHOuPqgCveii9Bmk6o7
iM7DUI2d9z/ryLh+zoixslgIPP9vX9SN5ubtjyfvQGPw1rnKG5L23LDd76pqLe5QgyoVuLX49sRZ
+lHk+kfMNnfoo6T7Q34nGQFLwllC+GxEywRUwfil68NeYNiagCDDke7Wh7DnOgSkSR79qxv79hme
dBU6GctP0LG1GtP+U4n5Cnu47C+7D85tJySJVbHl4Ws4PwTmigFoNkEz509GxJAVIgHx0Hs2rqXN
JGt0TI93gihogdVUN/PL0JTOBCzz7A50v6gkE4m5Hg2GlIExZ56P32qBdNxoGAazYZcRFxy7h00M
ycdmVkMPTKT/CmsUyf4fO3Zg+uLC2ZaahZOuHgb4AwCexlJ51B1zDA70N9H4nOSjxIF5IRAcFJs1
et6Ub9wwaklnUn4qdhYstihKLTz2ecAClKSCrEfBbNXaKKV4FZ/AxY8zEntdYkEPTshOk3JX3Ri9
lGYyWyBSvFzeckYI0H60pH4mmT6qJMEdy4BAEMZaCAlbSEb4NE4BpRibQCnHgzRfZVRyEq0hXhcq
arZL+Jesw7PmN2wIn1kLB8RLtLvis4XO2qXcmPEVB17WTS+bBqyvZDUxfkf9+97Ymx8maxt96Zl3
muiqfT0YirLNHv+Z9dBPgQj3smV5xDxbBl5esZleQ96xjnb3AcBl9Xh0EQ+AzMGIhSkupP1YetJB
LlPy2W3KlqalV1N9hnDlqCpm2eClI6PmUWkxOYlAz7W40ItjqFsltZN1fvdFiUPNoD13bb2w4LW/
FDdN1/iUVlmxEH/kevrRbxyp89MZehDRYRhoHVYm1SHMC2eHYn8ABW08xsy90ihGvWn+QOU317YH
UeBE98rOJLM5xYlUdAJIKnj1IER/qWYFT3l67ys8MBvMX2qmtryeAOV5cNrN2uUJWPaSXmcswNXD
AQ7tmKCrdzM2uoZK4fGYgZDAjEDFt4UocWrnuGV3BSCqzOoGC/2g2mT3PnlG7FyUwwky0GDtqrmt
XKijCuwH3IFjc+ftjDPDzewzq5UoNPJLbKSMXbuUB1hQs3YWhGVQ9D7WEdWVGWxFvG4OgIErQo4h
BL0/y0uBV494qD5LMGMLzS+Ci/GhLLqzWJ2P6WWXyXFdaCoxzKi/+2morQNy3UAHkiLwxD+2uu7H
hZ9LDtimL1LgdCds+lmzYcAE2ipIrSyvYAf4VO7LuavwOb/9/7dsnCrM5GYBi4L2sZTg1/tQhd3w
4krgK2v2N3i0Ub10b7YseBls6ANHSlRlqBMFhlfW2FHJmqvzHgW8I8Lbz5fkOCmEgWXGvDQ9ARZk
Iw5DFKx26X0zQPrQZoRkjIEUtLyMAalpzyTXdet+hMvtH8DpArfjfiLRDB+gUerWi2n/XVuBCL5m
AQ0okNuMhgFkSY9oHfz5d48zt7EPnGYcxNveS9dO0AsssjP3VtELwNuBl56hS/iqmdRx7omVv4H5
bDIo3T4F/xMgPOKHXKW2XgNz8xBMtO9l+gpoBs9dNgDK1gumwY1T9AmUCWgq3xT5DWPUG+CM28JT
bTQHe4RPzTk2LbBAuDaJJHKnoU8RF9cLNV5I1DUFQE5K2N6O1nmyWdNSXo9E3taZmDLchJMhSYtk
3V7Q8Oc+bkHX5x0Yjo9UIpXuH9PTMy7Zwgysazs1h30vR/j7AkRAio4y4az9WnQ1GDV7ZihEN2RB
kzlgNbWSVNelLZlgrMmJ1LgDrZZ2IiPW424rr8ViMMbzJ1Kyi6ipc2yx13JHF+4f1Rq9CLwlPL1v
GSWmLi6UZ+4aLS1RZEUF76FcbsGlXFm37LWk/OlymacUf1w06SMgRXDKtZ8uPI1It0PSg6dJtB0w
zhM1BAaEEfgtob1y9mMOoa7mIl6xyL4IyhcK4yJ1KUM74LrYRQDnN2WxKb5yg6CwGxYCJgUjQP68
+MLwb4ybBVFNWwPTWtqgUYwlx56K1G9mAnVC48E+663MTURXkstTU9QqQz31AxiWkhZerGhx/SZQ
PyODy++8sZTQIOBEu67QTSeCCpIAnzVX/w+ikSSM/c6lQ0oMuIBMTI0nDm6mOOyu4c+tg+pVyMKn
MKD3Wq+k3cPbcNvl3uEwFTAOVZJtstO/93EBD6yBzY44dR5CqiqLren+1d2j18fLmQd46xAAd/p6
ou7WWRYog/MWj1n7PvNt+RBFfIkDzSZWSFT6FRmnAi4TAjX8GsU/lQ8g95/inz9OF4OYXOcXXYhd
jcq0g74cPfM3rbr2zNKwjYaOFfvIQE9f+wtOPL6RBSiZ+iMQvwN+zas8XLZNysWIfzJKgUmi1VxB
VMohg6sJj7J5xeWYA6ekTAtDoEjgIrdSRGngm3UAb2gZalQoLf7ms7ztqkfeVrmSp3L6Ofl380Ne
i5P9FHsRpBO9hhixuR5nuIFrP1yx4BOjYRctnuZT39Ml8KqiiisUgi53UeKNyxh9tEHgewmb4hKW
lABFEOsLmdCNs5Vf9a16vAYmajuEyhfYZqUPi3PEHIQVxTKqxL/LHpqNxC3BJ3KbU8lCEIPVpdo6
TZWyWO7m8ckqKghf6fkp6XNXdehx42/N0hELxdtUT5H2EHoNYpTnTuiQJcKAzqjy5irmGVmXS6AU
zFm5auN2HwQSTiI67mc1OGsl4rlo/UQgfWJ3wY3maKx93lp1o1pcoPgwnB+I/p/3H73iO3q4O5oO
A54wCNtV6rAyvyOzZsb8d69kiKqctEiXUsGOsSHYaOdiBkAQReUJkJTINniEFhuMsuiAOdBRjDYC
UNzWo0kyjIgOCTH1qUeKYGoTUMim/km56KpZBCjoIahVy5oEdF+jHfX27rz0yT2+i0XwzgoFun9g
K3pMWhDxILfGeszC/R8QjdCWsL7NvEzO3NTohm6LibyZvlinOm+ZAqxvfVJK6BCkWCOhW64VeJHl
oylcGXLgZ9ZQc6E9sQrna35J9hyqvnoOpSFZIiN2+Xr+1wTr14Vyu5bzcFsKYfHSbfkrD+D+hDGH
B+zL7xDucXqSyJ7coZmIkpXvYC3qDne6X48TmIHJlqgnew7P5qFFUZ6RmBv14oOgDwouWHV9FQOb
Wek0iOirnBUsiF3kLNua0sYk2cJmTeEj3offyvnbalyuuaoKIeqppk6zfWph4/RAI0kLf/yA174G
4COJJWMUCbfRLuD4HeKWbQiViYw50y1+RqYKPmyiwTtreR0UAxYSeAlCPC53qPLdt1dtrhZRQFTi
C8zmt81un8TeZzbX05yNdG721G4u5SGbxbQG9Eztqcg3qaqzyCFyJPpXuzOHGyJHT9nMjxzZv0Ve
grfqj6iAZuLTve2bamnV2uEpZEljAfbhz3Tn1jNrayeoSxjkqHDod8NmO+yTlv8Ohk+Plhhn+41P
GdWoW2kfRQ7AaqyqVdCVn/KegoAXQOUcq+ikVOfFUjz16wJRy7qV9R0Lv4mps9D5wSGDJI513g9B
VV9FHnR1OJQDVPux52iOXTuiIrcRR0wrDcE7X1aDcProtO9FOpRlUJ1piENoRhJ/D0tsbZCU2yRh
5yBVct2hYmAi+ZVNarY1fRW6popzUj0uoV4y1ivTe34HHmPA/xC3NPhNW93goSbhHXVdV7uekpe6
U+NPqT0FEx3I5vqFEcDr7HPlBSyHeVnCicQUgjH3hXgAfUGkJttEWZ0BURiJKYp/+C3WMPL6hFIa
LkYWFRvhJnaYYhMjE68jN/QvEMlKq33qsgqeYR22KGPQvvXs+wmV8R8CJvrKd8TZYBfqwRbdWSMy
tCh+n5K2QFiHTp6FqXfIP0cx17NgINU3aERZyz9MNTBRnRE+oaJmGIaAzx2UnDU0WB3acGibJ8C6
dQWS6pgx3HbJtuv4aBFGztWkCWnz+QSXyH1SdYo0Pj5ZP+ajKQHgCOrfU/6+6cJ+Rbk+gkB8QBcA
zbZPWbUOuOIsvN2nO1QjQiUBAjC4wUCEEcZrf6LSnsk8hSafr9AX1/eZyQWgedVDlqNSmYmQQG3M
V0i4pozNXnM2Sw5ANih44dGWJpiuV7zJrE8A5Sx2Hc6PsQ87iLEwPEUoZ4BqU6ggPHzaO9gfIHUy
O/kkZyR8G3kpAg0HKM8PS3LReyjTA15CQuZn1uwUjTkxdl9x3Qdq8h8IqtxZygoOb3mFoXM/8So7
fu2c1PbFL7XfokO5b5Ovm8HsOSa9DS7Z9bBTQt21ZQXWJiQGOYQc+EYDWKaiD6AJMqFTmGZJFbEg
BgrJCsxK+TpJ+aPMUrHvmwj0wwOzJnGYNxBQkYb3XJeOqpAhDBWhXJ036woS9PWdVEsVhT7EiwlV
/14qEGe3sb8LGU7g8l7YcnbLoEINvw/fR1IPVrbfIMhrQ1TH3YkrrDrdxnjMDtn7b5tPCO0bfgad
VwwHof5lsu/K8LHU1IEo7dpzxAnoqq19LvFV9hnPccM3YNLA3OYIAYyqgw4aDGlco3wsvMLRaeBW
5d4QjP4WS1XgNTDGugnZ4xQIdasw9Yvk9HiGSmSSo/r5Yb96RIOpFNaiErEvOsw8MKvXBRcDgN9r
JzqnMaN874eQWlVROtow4kvHI5O3filqylaw14wJVcO/fYs4l27HdRnFBDDmIEEJUatHXY+l/XQB
Ihh+XdPqhSfp/oCAZ14ABIS5UQOfZTgxTQ35kurLLXF2Dd04qB4vqjMmUElVyC1dByGWhV/tWXqU
SXLIPmbyhlMWZHXsP1UkzlsNIv4GyiNgPPZ1gP0vWKr9TgzmhRN4554qxoTP5yLJxxScN2t3eTMp
KVf9iSE4Zkkn4zIizloyXELb95pRkbm0Q70WzCm8YOt/ImIvYrketHSU+Bph7aIKK7k65YJNo285
PWETw2v8Lr3Z18iq11IMTPgOXZr+k45gsc+Khg9UsKausVA+njAtwnlSZWZ3tQd0ARWppP0eamFK
VFliFWvyYU7/q57WRcOCEo5ud3UbihOHaObDCIvMP9VmOvPdZBNEa2gRb/XDXMFSB3P7ut+AiFBf
FnYv33BGmXYWC13vrcSqJHQc/d4k5eimaR5wtIX0y6arYR+2Oc6CiMA2Obg+DFQJ34+NN+PHMjFn
0C1tl2udI56qBT3DUOTmaQvTeLxqpF1/qJaPXa5WDnTdtWTNWqPgtixnzTTfq+905Vmbdb7gEmCi
98yHy0RawPCGl9afpyIPZMZzICq0WrFLW+TAknIvZHsH9ajdw9W/fh6vTPTYgU/er4YLeiNenh7K
WDmspFY4o7A/kOU6x+ote7KYQXbn9s0vS50+kk2/JNoPI5SwfwcF/cqMrkzFpRGCNz/3mtVP0Tx5
hE6d0OVZi0cGyVLnrd29IYCDAaDGBFsabWei3AdvrVsASV33RENwQpTV8gfBRshQ5xmNQpA+a/nd
1WODOQdKwTvRhEBCwvZtyAitW2k2WOasLaI/qV5qo73nB8ojXxixniUzTMlYTdJYHpD1l6arbJvx
5pZAW5sOIV6cXs/qxXyNJUuKDU4UZda3XAvHQ3T/RBoHK0sfY2szTU/+dP9Qj9LWtzV49T7du75F
iolHEL6fD1cIxpeEk6qN1CUv7n7rDpoYZ8o6YbiS7t2/Vh+1JPm5vPucVyPsna9oXR2VH/ZloZZC
0DK6zlAdOZAvqjqAjGW77ISCmiTbQNJK5N1NvZUcLYcRkTcB441k6QJDBIv0E8691imyDG2H8LlM
KK2DFS8c/vPmDEQ+S1P+O4sSx5ubM7lnDFFx2FqsjUabm3ZuGYfaljzG/uTo1ih73OQfn2xv0FjU
2DUmkPMqn0jT3NWnp+tfOz769RYwn9h4d38lMb3uXGadNEriOWQUiIdrg9ZfNGqKs125uu8tlaSw
rYY4VJ9iRu1RLwsCI1YATVtYwW/rzY1EI54LjQIHTTYqXo0H89EugTNvWoIeCYzDbdc8NOHG8589
tlJv48hRDGm+nEuW1aViLPlqdAXHE4S0I/EJvcckzNEphbmyZ7j712I9kB+Dk+QMcH+Wsnm7Edpl
7J/dLMi7Am5C3SDkUQPB0mkLucHb1/v9mnQFn3rWvRU77JohbxJTuqW2QmXGyfYa6oRzMlEybcRH
uFymA3PVGOgCJKkOjR66dxgPiYjvfqI5TB+REBhknKbWWhzV1I4clkPlDCHj18RCmGP2rx18EPfX
HGJl3vkt1socOp35942H5fCTLkvZwELHm4p3wthhtpLdLpP5zFkQbi2rMHNZSCLDbixXq/FcEd7Y
dxAxQ5hsiViQD1fhCjLh2VEhEeToLlJSubQHGJs78w6srSQI9eSpTIo1s5s3wwlbRWq5GgYKWTtv
Pbx2u29f8v0FjwTjItYw5dyCUrD0LzQWVa7wiwK3QqrZPa1XdbMGGzTZdoGgUTvBqYDtnk/kR/w0
9ZH6bIgPsVWtatswn+WmcEjCezdSUaZrZ8fUFZyiFRnIL8t/eNPDCgUxtLoLJvzfpNvH00wXiKE1
L+UQyDFhuESQ2fdU5VNROPbcivmAOslf88FbgiscSLK/1RLu9M+6XQMW9+KV54ql6YqUxUSEG3n0
3Dsjf6b9bLHqoQbN3kfZNUnzo+cYPRvlJo/O0cOg+6axdmrLvOa/AiMHG8BxAz5GQwzQPkNTlZCs
CroalzxK/9Ut6cb1jmWoSaQwwD3vWbJe1QyZyncqmk6b4+gB80IxN/RKjQrt0BaiqVHHAKUCLXfH
Leb2WJ0SZuaeMeJ34dNlOxdznqIdBsWqU+3v0GNwtGDzy1oxEUMq0jgOfgmG0sLQD25bnghc91s2
Q2bDW3SDXFmaU7m+qPzyb5DtAUz9jk3mGoMgDTrBI8QK2NoyuK35uJE//VBDXBRIQFXTUy0RsDAX
0mG5vYnVPyVbtUZV1uz5mfEtfd+SLjrh4XSIPJgXncfJSKOAsuJG14eKduT/58uTtocmxXEVXvqA
0AxPjxGRu0u5AxUNSFwdu0Vl/EJgN4rTwq7uwSUyHfP6gGbuTd2wn/au4aQ4YscLPga9jZNLw/tm
pAeZUa5HY7ib925Ci+hFhJlDcEbIxU/zQvz+M4zqRE2oiI45xhV4QCdxUdSa93w7hcFC3KJIvciH
P7fu9OutuF++Sfy0x6eZ4EK64er5KCt7G7EmY1V7fu9g8wPfeBcLThDMeBuMXbizQGWZ94hcFUPH
FsrQozMpd5BsYnBwMFnFM30y4aFQAljkYDMOCM7llztUSjrGy/KHeOAqVmyxzAM0zOCQVavLtn20
6UIwmdiuBdhQdaaDHy+lA/N409zqVg8RSwKhEaameYBTlaJWIvNxGV6AMBPMqtIGAsSUG1lTBrJS
Yts8JXjioaBoekVAkQwAI2eTVm//mAolk5TAQAqBKTlDuu8JI6EZlR8O/lV7Pt6aFXJv/idZEP1x
1OJfnWs6I6QzUuXkdemdduqRW4D2UMkW0CJnW5XYFJTpfGVI+iWX68XOAIPILVXW9cjI4XibPh23
53s2AVMRhJ1ldN/HmZUOIlc4kCvzjHmvGSnuOEENrAL0zDrnYeHUi7kF8T6FUD461OLGsj1DRmHc
pWvWaMQs6extS3wKVZelpfNpyGH9EIgL/ifKB/iQSxgpAs6AbQPK99IPZsOcwZ8osapJrZmeM7V/
H4Y1XjLQ635Dejk3DXH2fySVxx5zSGwc9mjhMbi1htZQvZP8lc0KcVy7JbAbI8SNuSulB4W0YOgP
hoEAsasDB8runbbLEXMfiVRUlRxhSP18C9AydXTBYjB4svk1e+akOrkabevkk5+bbog8AjQLXDWN
A5jzaqG0tPdWcbKfu/79YEl+dpchGzOrNK9gID0eT5NQ/8rybN4N5vM7/d5lREQRbBEe+2c/mvtF
1DYeyfMQ6SMI/773ewcrawB8x6cJpYtKeUJb/5ffVzeb8Vdm+jjOkuGp+4zvy4KZH/YMgRMdlW0Q
HVL4lAs/DqzXWWqdyI3cOafES9Bu+uIZ7bWgbUoXEfR5Xe10qAEqy53hzTXxyWKcr27CmqjGc9yz
HuMkUW1gZSd+gTCw2fvPVFJPWGbZHq1woINM4XwcHfnX3I6CZI9P54mK
%%% protect end_protected
