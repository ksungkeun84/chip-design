%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
NJ/H0nzvFsvYOxnmjbh6Yf28UlUk8UrfVn8Vrx3G6SEkMIFcAPTrf5Xum7tJD4GdP3Hss1I6pH9/
GALrZ7kspIZ6uu/8JZkqI30AQYjZHJZsOgJZZEzZNtTjxpERrSlJcJz/Fo8aBvb8K/CAS6rFkE+U
k9MgVb2KMA/suLQY0NO9taZGeYF+iw1vuDGLU6iV15Xl8Cjm6Pq0+/esiOEGosgepDlreMypfamY
fZxK7R5Zi8ajgjaOxdskJtsSXSABeAxIJ4mc2pTmU+a+MROoEDj73ImrOG/okN3f1MphGHeIwQz9
9nlMQWwUXTeZoRCVvGtKjwXMpb0hff867oQsXA==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
RqFgAV1dGlcSwRJKM0HHoZmAyBf58JNAi2Klv4AwodOzbRORr504HBZ7FUqJNRdbjp3VBo4H1NtO
qSA6YXs3NWo0BDG8c7CS95iIZgiphVDSlkXGGZIAj4ufsPy1moVATAaUyfCTFTglbGJorA/6GFSV
WPx+RFRGzS5+JZpgoCy5w4cYHARKJrpSWJSNTKM25tdKefGB5iaemhsSOikWIlMXCOFMrRMy65Xh
E4FD2COi9fb/VDawZkV+3g8CbKpUbDmAebOQJgu/ax4gLvOc/vDGM2LGbQZmC/HLSyMNphMuSLSA
clQh1VCXla5zTe80orrOyC7+lvtgRkvzyMH6Lpqi6wCqPeDcQVqotiZcusvb0avWsZrnxfP95PLS
KefCzwn8iR1/cQGK9lYMakAKqfFx6Yx6PpmHPfemN6lU8oUhlfvQNeDKiSEPm3SXK/AyOr6GOxSN
bn5lskvLmUel5bkzpL4t8strjde+v+oswiFGRJjL9ReQQigHAvVGcGG19uvZXvLdlCAVpsoa47JM
PahWCoXpAuvFeLNeR+mHLnvVI47ma/UDgvUkP0sHcY2eX+F7v2d1WWNNdGnrfal7wqnFSrpInkzo
C3L6yPq5jv8e8e1WCEi3bzoAusZ9zPDd74uQw8BYfcK+uxxB828o7UQ29Tfjj8HAKMJiWBvPRLxw
AuQ0BsrgjseXMCXlUisYeWCfvX6U1eKSwsyW9BNYSeVqx14ymVCEYXG8Mm+R/Do33wF5trtMTFEi
ykBMMq4S+1szJBqFV5h9Rq4VC5BMgqCcsa2+JK0uXlMmcXJATz0dLpvE7EqxWKJU+fOMwjtQAlcP
HfGqkJ8UjwrB0Vke2iCDCeAIZp5ztlT7urevyESf4Cpzwh02G37xuF8j49/nlq0GJ7g3WhromVv7
pMmH3S06eNkWfsw5l5eFbRFZut3use78tECZO9TBbIsgA98W85N5FvzbTfRHImNA148Xfbier3lA
sDnheZ/8RFEfMQL3nD6gB0Ta6JZ6F0eGoiOoyBTPnsKB11m5ylGRDvnDs5/Ej6gHEMjsxrXauh9W
OCGjViZWfbLOnFxwISDuhh/E9MWybmQFzWSAR1rt6WMBe4PDI0BgfOTPa6ra8BzNifcGuBNGcQxW
LvTiRtCgpN+uIS5NJT8Lk3Q7ThKEX4URSQyTZa96i+XddDNbXJMJrJZkwYKB7MsRwk9HmSuxasmT
Nb17XbHsL1k/BQAMugrqxrpEIItXQi7GORSidFhYh0IPFr5yBmvJLk54tJZ7OIdvp2YKSr61YXpH
R/xEWuIw6KltQ+GZ1kqavCHG8gvNXHLr0cKJPNUMpDKlbJwi4TnyjSJJ+q9Wdy82NhW75P0dq8Sk
G/GZhpcOxyO83AHgZ5boKk56Szt4bErhoFecY/dyjGNwsZb/wwIMX/8bopF7mIcqV8AqSnsWBIh6
XCN3N1P7A8YYzeX/e6pg+jQ4rN6wW+d4czfioVzY5SZ0rY+qvIiaYDRkz5FErCa7UPGvHzh5vqgI
ElQF3peovy95TMDxJ7fP4AALWCozgVFNktzabaLoOdG6r6qRGslA8I8LSFJzeKT7CbAbelpynqRV
Ew0teHwzeEoLV85DAGjcLfs3tWJ663eUi+L2d6FDtwQqVcO2CEQIdzBjn3xNZ8DoPUFjIJzFWM5W
gLqK/XMzvx1NCgIstv/Z7wqnz4QMiEylpGfKZEUbegIgCf5Jyv3kFnFAS2/cuylfEw9/ZH8Jq43A
TFdKN8RKEmbU+ZpZXM1NScJmWVPFNrqlOl+NZ55JL5gas6VG/CCLiIAf90ttKIfnwa5VmmmqMD5h
t+NJPlQsOhQop5kw0reJmUECfIWpYsoquVkTbRO/czgVzBzvB5EvHj1sHqRH3Bno1v6/iqyf5i1u
xnKfNo6pvic1vM3Kog3cNm1iUFyM8kwq8h++6XuyQaq9H9Gy7tgKQ7ainoInGmdUhDlEk2Xgw+SA
fPPrvNIVRXvEzDTobG2YvE6A5gSJhN+Voyv9lOAMQjR6KdjJu45pCL6iXdo9OfQTI3vVsriz+qpA
EY+P68wGY0vCTBsmEB8Ux/5HlFE4dDw7bzrjDnW9yH/nnuFvNm9NUJsBrchZ5kG0nBsRARq01l6Z
IR1LMeAM5ykPbB5GNgJetV+ec9O+UblcEnf9jbBjLEsAVYtXazna9kCd4A/SyGSiNo6UILwE4Afr
WBMYJGoOzznlDXifT5FcOO09WX9RW/3a5wSLRSwCA3zHu6ZTquYhKeOntcYQkwCYpDopjEY6LGTU
jTEJxyKL+8sFCcTqa9OA48DObvXdgSx2n7f4Z5g2D1tDRobxbsFfVCKJ8NDKHzFf0Dzv5o3+lSDi
oGcodWkQooKX8AEazunXyOBJddZayM/6jkQVBaXtklH1KwucSl5MqtbEBbx+2N00TR7uzsxspAAG
k9MgEAsNO2pN/ekW1+gFp7QUS+6n8KpHGa4fVsI5ZosxL/dzyamxX3CaMg0Ue+dW4I5/3jf7e0ka
DHI4lFXb5gf+rbEsBdU6O5EU6uDQQAMNyeDSGzTHL6FlwgjcH6KYOjTU5KXXkLZqaNgqtdNX74P7
plK/6/AhMSK9X9DzUY65TqcIvETN5E6s+ToJfuDwhja8xxxKZzjsIjq+aizwWAqvGMVqUuM3EElf
saniDsfdO0NBYAgKVy31uA2rXUOPPOgK0lhpgl19VNavtOykmvIUgOeXGDKeX+XUjWn/uwXNW91g
xYZ0guqFq4CVPhij+7/KJYfrKRUvoION4JiTuNgl2Zx73RiEY54bP79LdeI9iZKRorrcz0shZupR
PFf6CckjC/L3reBKkIKB7iTyA7uVf0UxZMDPoandGRYKzI86YIBRzbaovZhJ3fc7SQ1sg0xbtjir
8TJ1zW82XSzdpfJecuy6eriLIJP1/TOSQrpWaig2GYckTgpIlstHu7asYzJlOIdS7p5aVEmFT4p1
hLlJ1z2EY+i6VrWuCXU6Tzx3nNPZKagButnaIe8KtsmUNCM0moO9baBYyIcaeVafmQzhaOXmRFLv
QsDafQNaeM4MUVp8Kv9BdZXWVBoORuHinyjzByMjUrFozKWTYuAAAo4jYC39bU4QuC4YicWzcpIy
0/taUG8o0cPBlo6as9AGhxImuATCZmGzbyiM1uNxi81cwZNaVKfhKMyeRgoTmClHY6GFFR2Mb5ev
aCTTe8/lxSawAFb4Kqn0tTk0DC6P5IsYJ7BRFUcTG2Un5dQIiNUyk0pL13C13Xc1/AJvnYpGVILR
jHyagm5Se39fRrJMRQ2+6qiFufTVZ7Oi+/WwvVjIVxBqro6zm4OmU1gfNTStP3kaNdPmp8TlbR1W
Yx8wqT5VtvD5baDL35c8L/+DeZIc7nFE3PVwx8YSEpnr46BxJY+IZ0boLcpQ6N4A/HpXAO9qv25o
UGdoXdT1xeANDgDsMa4JJMXDLs5UnZMJ04NBBvTQwheRtXCv+n5/rPddaWjdW7l7dZLYRapnlafm
vdN/KZkS1HWclx08YlBUPjMjpfx0zDiXQRhFFB+JGNEEgNasZMuvNjbZbQdvnXV3P56NLIB/824g
3IvvNSr0b0YY7TTLfqvC95yeUP7zbt4AZYd9qwUdXHL2VGVvqfjjf2ggFr1T5ofVl5ohl2zdJzQA
rSaqv5Uynrp95wLHdtaQg1Fv1JQrtleUD1BnQ2VlSfMBzX20f0d/U6BaoN1Ci/nfnE45uKM3Feyi
0II2GixE3sralJsT3mjcp0W7vCOAzBvqW9YTB/9QpnV4Z0sUuAMmSBYp824FOVzx7DRkJZ1RMT0L
Sj6V0mLtIvivb03eFcDwFU0NI7THKVFo2jDecPfBxF6SiFjvBWgPAJ7mt7BXo6uS0RC3uGoeufUw
VM4fLffRUyV9lCOrhMtKsFszW6fUgIGU0tLr1ICyuJdquLOTKlUZknn0r/NS/33vfz77yvlhtIr4
vS3SIG4tmgL3UnAZxIxpel+AMEl8o9+PtvPzugip68zOsyFVr3fyYI38IDF0lenW3G6qKsnAveKz
k8PGxIA83TnAptwx8Xz2Yw5zbE7x0CRl1yDhtF+BKUk3onPfjHodQNZSjtim2cV+n5Z6/5tRiZIZ
9dDF7vTtZkKlMMzkWeVfBdDzLoAybB9IDdNI5n34/sCbgU/njywD70P5WFy/jWgwXRusmJGcvC9s
V6SBL2k5moSNgVO31wTyguqwkRsc6pTuRKpJI7A+upmGoK4Ov6ryI1KGmECNfr3YUr5CKZiK6Ujb
0Bi5VxXiOzuBIyEbRjc9WXCbTSOKTZaZ/LqKXAKXAmBGEtd86+Nkrm5lPZ8tXzWdB8mXqKMSyPjH
e6HtOTiKn04X9SD82ylBhd5Cg+Kqt9reEIsX83+wRd5iV2Z7v6E2wzgD064IACg5NQgn0PUTpuYk
PnTNjgipscvumsQOqGHEE4NwsX1YNyvncH5FLsYl+bwqgTF4YPKaArr2edjAfo1aTJR1cVXH0BT5
mYQnT2zzuoFvkaSwxtYcMgjFO4dW5LiTzejhza9jScgIeJ9usu7U0ICFp7j/u5LmTU0Pu2kOWZLp
mtvm3k1Uis35sUhQvjkLH+Nf8W2OXlh+zmDF1fA4OG81zJbzItzgimWuCSwPIiumgtu0Dk+np0wm
YdIpvd7dVxW23qdGsH4d6tkxtdxa66HDce7lu6kp0q4NTXma7H59+IAIMynTpduZZ2UEWeLCBGY+
HHRoOJJSKnppvQt6jzGDw2LXxpHSx/VSfH9uh3TLyySYI6gZ9eBNvppGmA1N+XLnAJQP/MbcCi48
bzEip/rk6qCGp/shRQQM5WnGTpOH3P7zoNhbKqe8lgCPQrAEoUBdem2Ef45umzoX5ovzSriprF9/
ns8S0RHLgsAQ/ltqVAYIdjPhaCs9zew5A4CIfEmRQeunEdDr8ekxV9/EVf81Yyz6PCDm70+IJwCj
DJ13ksmDJSfeX/6bmvUlyaD5n6/lJn17YYt6HnIfyywdtYC68GSDUhoclDmTG669wHx62ISRLnlo
W4idQZsxId5odP05JN67/ma4582iAOYxR3XbnYIt/+pVK7ANqrPN+P9iG8LTHWu3ss1MzWFyhQyL
xbHKD+9V2rLN5oQhdC7+YwwsDVAaMFWcD40F9NRDiEdSDvatvAYdxFH5nsf0BISLRjTgM+2K/tbT
gGi+z/sIupexnVKYBliSfy5XMzXNdPAu8UQ9daPTKdaDI9K7qb2X8xAyVBjOmvdH55twD06g2WHf
C4+fUG0VctmfRIB8EsDY0cp2zkFW77omRPASOAYN8+XX3VHDMnHDJsWrcdJue7Z/JRfBjVo1rw4r
Pa5hCDnV3/fXVQAp/DLUqZfnyG/eaQcWv+5KmvJBoTq74bfQs4JLf5OE7//+ZQQHMsAJXIMJ6Nr0
Pq6IV3td2A/C/L8RH+HxhUt5+6ZllsmaQ2ox7AEZr/1Tb97o9jZF9bAxkPO0pIO1mlUS30A8RSvo
16+kTq/++Marrt4VIA1pseT7UhjF5CgpCfM6jfHMUnbYuVGHaXdux3+oRghTWArFE83gXxq8iEXs
TPbne6tn9QHLjvO7YI1aeICZ7xVoIf3W3AgsDmDQC5fdLMiw/CKeuwbnFRTGPqTJru7ozTn1kN6v
z/RwZJhnX2hosJY924VB+jjEK7peaCzGJf1x7l78lCCKnRMfN4UweWViz/f3rQsdKALamL7mpk69
JJ/Q9aSCUnft1KUpJTy4DV5IxoQE4QIeZalbf+ze4P5rVV+OSEMamdN7WqQQuAIEqPVunEUTmNFl
x9fkDYC98+L0+v2PCn/oHnaQQUEcsfirnDt6z+oW6VsXp5ZiNLs78iXimf8fMm3qb2OSJxrBd7PL
XxtNge+VImPv/AWZMufdgTe9pXjrKlIYlPra2+bDCX8X7zzhK8ZNrvh8NhdK6dywBZ5ey7gWa0mc
V6YIZuuaTLtQvqi/UVnKb6A/NY9Phd7po3lZBxZsj4mTG+AjmeEaj60WQB5K0cTHHC3chA1/Y4+q
m5DaOsdDyn6+H048neM+CZzAIx1rByUS6aICrJ8nSnajHoMWSUmcS4IPTBdwOkOG4NNe0HXXzJAJ
BtmWa+Px7cFpS/xGg5RWcyz/dmU0JdeA4yJy8uLuM1CfdwdD2/k5ZPCnvh8ZyRIBwddXdi6rcwM/
RpoqQrehRw5sBKqERezX1fcx6rjV6DspAu/UZhfc+o2hmkXibNv0lAaoR47FcacmRNBiXvBkFWJa
th1AFeXgKIUMk1PhHoNh53guotShDuROkjsyV4Qc9fycFbsTIeFzOUkHq7lkwVGULOCbpEb2Ympm
i2I21cV8e+Or7FeiTtfkyekYCZJxSCqzTURBGTQJ6p4lDDn90N0OzaZAhSeNMMRq5dYcLqWURPu+
6HnNYfXVTf8Z5xwx6UYf0cczrNcNoTqU23Xpy0jZ3qTDcQ6tViqL51s0PgFRpzCgafpH6XcPHNMs
+yuo8NgtNcKu89xL3riPh7Sh4SoRsvm7ZQR4h95UQJS2IyUhfm5j8E51IBNjCwHfjdL8dm0G2G8E
9WsU377tiS7M4/dzmITvWj16LxJGouixeSFvjhUgLRsZl3fCX0FaFXZqW3KsVnhBv6xGtKGLXDJd
X+xNRVQ/DQJ87kctBq58vUE9i5+koW50VacTSsN+4USaZs2TecP944eFx9/EUo0PiNXlGnr78shP
lkm97rQyQ/wtdpNEvFaOkPUhwY8o7iY07L0u4trl0hU84sKL4pfcZHtUEo8J+hsMKH5hLpObTCDn
rnwqqno26FgA3dPVoMiR9gTyBpufDUTGeMq++NjPy4jC0+hqb7jrHUSKYWeSO9SVNdATOAAlJHtJ
bVI70Gqsa5R8bsW4H66+2MNeIjdhQJCp/GF0ihQbuYmXpZzSckZuwGGFgCMILv4wJcmlboparXGb
wtEfqMgtI/2ITIgAdtP3N8LZJKHAW3bm5RGdrrg0xzNm+7xQhODI+367S0MRqWROKFZJmCGZ8Tev
yuwEwzf9+I0tVVxpEyej0E3prVjk8aYFP6lMKchPzWJNmbqIxen/w2AWHP/IF0uir6oTC7RyoN1E
YOBRMTr/M3dtD+UJKKjthDGfxS17VerLn2p1f476FdjIl/GsL7XIm4pcapTYUhHLewt5GYwE7SW8
qTNLoZVZqzP/tiZlSrUA6z9b/IC/qnUWD+rxRKCPung70Y2uZ04RTDWFNNRjYxFx5W8zy3BNNc+7
mP01zs/qd9rvY/qon6129hL0x6zArqSGpuR9N5yoNXn0oQkQLGQYURDgHEFNFgrF9s6vu2trq8sD
FwqNWGkkZfaI+5rvUR8qcQBXDyf3wPOum/Y3UzA05Y/ScoL/b4JzQXHeI5JaKVkW6TIkfwnsEK8i
8Nw7IqHWJ0QrvSnqYoiTJ3M4Dlzgkt++L3hZ630ChEe0XrSOd764VJrAbjUx8ot+G+FRQ1htT31I
jBKw741s//0WE2MxpQ2neuei49VzkGHFsFBWTNN52j1JZuNSVXe0z8M0lJXQIg+QIvTW0UFZf8KY
ChsNzYn/Xn2OjoYicIpQFpURyoKIdLTNt9pbKvMlVVg7Y275uomJmLRPjBchw8rDrKGdhxprYI0H
KGnvmXZih2MZnxbIXkDZ9Qc7m1rKODW8cXfxZ22vMoXakyyB9VSxg5SS8oWXHIuONeGBifx3yIwx
KGVCSY2cx5pF+LUMz6jPFNyJBdqZWVKlxlCkbAGN3q9xbgv1pOCQq75pz0OVG6u4jN3T8Lx2SZrX
G7FUhp0HuO8+ZMNzhmjS2UMjmwrbhWYe7KSClEsfALQi0mPcWiVqkoz+RNkzNsAe5zFLTsBwKJV9
0zhFbw0c0+8yDJNpTdOChJk4RgbZgpK66zQJtleWRTpQCy0rg0RaVxCBuE2qO3+pFWZqyEPWqa5U
JTLGB24mDSRxJ1T9dYeDwHICRVSByuLtVF6kGVg+kq7GQhYwzaR6zrwh8PJdLjbHkA1Kl4YrxBOu
FuvK899aIfEXoqgEk+Xqq8sfdVrF7AxP4Kh0ad7UIBS9mcirGp9xbbmXArmIvAXrl9Ryv+Xp6zDs
R6eywnQ83DWf09AXHp2mwESFVknyT55leKSBu0tODsJ4ptLQYIVj+kvKNSiFRTMlLTYb9wnP9dFP
zkIDau+vY2EwLCk5wdbTuTagnjM3EMOXjcNGyYf+Q7M+V7FRsGqW2vNXg/V5dZjMxZs9ei//yw5A
p+P7Rh9MHNUMrMmmaPPt6S/hUyNb13B6TOLHzEFuzCww7/MJbKDZa45ZH2TMghx1HnlNaANuDeX6
3V1W4gVGQhYk2jhw3GkS1b/gRrLrPhUQ2xTTIXE2OfVhl4KQh+bR5YxrCw9EpRny0JGSP9EO7ytY
y8Q15Obdg/HJpJ0Nz3eFtqs2paZ1TpQUjaygyj8CgL316Mq44TJh4jcironi2B9eaFSeG7iL1Y9f
R7l9O/7k4sVR4VLsN8FViamiJw59z13zSDuwdBKqI9oVf6415TOrInWkjqir/528NsEEH4frhsDE
7zzc6JJcDG5W5WoJrkir34kOlN7FDGe0RsX8GF0AHaWbPCLJbZOsJoDZczgvYbrKoYRfWfeATUyv
uqRauGNfmKo0spIbgQVAqz0+4yUxWdurbUFZGHuLcZy1tdjEI/TVcH4K6s6LIDc8gCjPXdgBLGyT
fIRrHHLC/X91NGe0cu1fbcJegbAariDN/GvpqIkHvQFxrb5chhWYT6AF5ZMOPMUCto3TVGMOIyOu
FoUW8whfgUym55lwon7/6gycr3xkxgCGIqhHde0ZZHyXzPFLnJIGHgqYCveSzbexB1zHbXsY0B/V
tLirlj0Hn0hKMoKNC/+eteBV91lqZjltuCeO+KhvrYxfdGk/JE/EcnTZkT9Nfc1kD4v5RC+OLKy1
FxWQWUlq/UtRgguH+Zf2FqLQxCe8UpcYX+r4+621sMcZnaZ2ru+y8yF3JsbTkDG0DioCQr49lNYX
HYdDqP++qPKtta4rCEk1AJOKptrhAzDw6LrQLfzwXZkdv6jganGOH1o64DREmLNug1JZa1cc1ouE
V4MAF92uLcBB578l0qZxWAd8bzyu3c1wv7jd2qNh9tawKRjrbzWiUV/fFQ4DLyJ27/HGBj3aGP0i
ODOdLI9cpzEuKkBvnuVU4pOWwv1bW3ecTAenv7myWmY/StRmmgmJj823n6mXYoxfF9DJkrp6qD9T
3hyeIp54h9HZmL9MuKzi/gm5XHx8gdqMPxeiuI/PpqHEXT7BSMGPYTdRowL97Ucs7Lr/o85wHQxr
nwCrZr7r+bwcWP2nd7h/xneF9uvutJjnuNfzHCkBkMg/9Hfv5ZsHlSX+Dybe7m2iYM2N9Ot3v8HV
pLk0AsZwaNj63wZ3YnaQuyLqSBdqEn0pC1zyj4HhjvetQLWg9IqsioGjieQQw52RWzqDdptYxRw/
pFOM2FsoeNoxMhk80QyTco26UEVnUa0dINs/ZVjO8GbRjtUCe/TMACNFJRRa7GHjKCIZFMYESm8B
A9pqJ6VQkWlYg51pxs4ivKj7pFgUQQBpMY0AXH1dlSCuDrzshthJHbh+N+nVqQqGs5T1s0bc4pG0
GIOTEs+bNErW+F9NYxzBvhX5u8/0jM0b3kUx/4QwU3pcb9iPIE5sWRdpbiHeM4Yoiwd0SMysIYLQ
Yywk9YczcfL/737gjtthuKd+54OyOsAdyNu3RSiluI4pNK33BgrK51cfebk64zoVPqXEf3jFxoVS
zz+1XkCaJJGiilxTr8IrXWU6ERZXFl/BLbcGZw/OL8VL5KDgJuIsTYLRk4da24bXW6cCumoOBPJL
D3dVSo6ktwu7PhskPsXOy57YHrTdUXOdhIngDrtAV7fdAgUYniQgCsZaFkTAFvuzd3+bJ7/OdFB6
xSWWb7c6cybolirmK6DvArrQkYDO1uTLFMMWhCTidcQ/9LH4AHJl4TwFENRwLQ6HOkNYmrGnnh3Y
6FMIO6/9ThCWgpe7mbBLuDWXgu8eVgwqxzMdl3/5seHBWjI273eNZtmftjKQA8FgNpuHQCzRwn+o
HpJ7GWfKbPdQHX0yQ+TxS9+FVF3roNNnsAfzQskmw4E7vufYRCqSquPtE1Q+70XQ80kbJgiK1F70
fgzLiHoegfT2HIAK4UZzZbA4CbA1kL9ctg1/pLtlg6yDVnB9hHJJCrrarO8Lk5IDyXYtEFvBV/55
yJIUESFl2GeR4KqIktsPXYxYQh66QE6+Vrxywk1DFxcqSD3DBpVjVQ+wzGA+aeTJLxZWijreg/4f
XK6b9zOQCFwYYIimhXuLj0Ni44krkX3n5Rd26iXQw3ztb/Mzw+7t1/H+4y/m99LFkhOuTEB7B41z
oKfe1SuoZ6ibPKCekeeQIfdFWatQeXlcv2ifl15xT3wgfg7xLiX21Rm/g06IkAt+NZUKTkmBU3J/
y6vHtjtEKkVb4f3TNRACy7P6G577QU0unYVfP1UELoteApqNehblWDKYSO0+UmZMw121+aXtnAyB
0zoGshmvCc1PIX8Io3zr4XLrk3BsPoTvqy1Nms6DmMf84AhLKenZBaUidXeUTf2RkUm0NusXIWjB
f5az+FiBwl5T2eHDhRqN+GMcKH2UWID5lsiVfnIyJ/71TsWxGmnumg3Sp96ug3n3D4XySMBAzp18
tjHmoaHnQ3PZSm0EZW3InHr1xQaLjVThtVbmsQHsD9MEAqULWhjv2xRxcGLkhl6GpVwKFNUZUCuY
BjSul/5Dtgop9WXaKI24P93+vXYtyLZ8t2Z8VlMk0IRup3FJB0NE1zI0t3DukWSZWEevzDs0FbMY
XAy60p9H672r5QAyAm9D4DM0eVhTX+zYeQo+LOu/T/cJgwGsCjz1slDrlm/M+d4NyrZmksCQ3Fde
RGVXKM4Sc/vmVEbyB/E7Y8XTZ7A+p/Q9VaRs3/LtfnHZIexsPnDS+Lh5WgBRNwY+swe7O8/WeIN2
ryc88ES8+uxWaBsCR7h2nD/6pM+OQao2WOU16VJbbUHIiT778nKB5nxEO5VISb/HSfc9bifcFH7C
WqWTrK/oYzcmV/e2jnGavoUFsqom2/ormuEyPz6OE7dEIdtZN79Mtc8LpDk0ophUYRk7+o9JIyp3
Li8JeikSW5K0STkztQdr2Btxa06PZTJKWTlmAcZFPLRnKZVokmv+/khsqsb4jOsbydIlsr7Sgxqm
WiMDE+gxFv2QmT8qXdv4ANUCWCN/HaoHD0IYcPzvzb2Moo9jI2W6Fw4uuKpBLMiMExeBax1bSqLO
9CnS4dWgmhnawZZwkcJ4WdRda2OuHcGLppRK2+bUvqFJIQiVa9NHaHmtEbSWBCkW87/g9Hsjdd1+
5YIUeMaDGWmRsujKJ9nJlBmh+eXxV3xF6O72wOAUFQKyRX8wgjDEeSgWWQ6fz2Z5h+cak2TAqI4g
jjm+7Ft86XxFTDTVTj0zZz0wb9cK8HJ4oItIIjj5LcVGadUetI+W7j0E1cbgwAtMG23xcAUWqbUH
CQm5v241u0kYfFE0QMVsU30zlsZfn0+sipL6dP/m/CzbD7RygdoFTY0mhm+YbDJHIt5hzOtnFbBi
48md3IkhnkVuPWD39aFlOL4fAIHA8ftu/w3Po/AQfcFx7abk0HIEiCm0fbCS1QYjJNwRr/fvu6MQ
mOfVHQZGp4nTH13JKI2G0OooIo5y0jgJi+DlPUMaSjsQ9OO37+nTK8Y6lnG/VSCwRScDyNZpt3z+
oywindnZeNwgEptXyKMR2farDleYqQy6tosayDt+osdyzl8MCQf+x9SRlBk3g3mFiNd3Fq9rWKOh
DwZAUdLsLvUg3qF4r4zbaZ4acsWH2nwmOuMH6qUIboCs4watBTuwMcyb4gBZq4pvr6GejFIYGr/m
cLBFuxjGQaI1PTkYwXAIGUg4pIvvh28wnkxrDb5Kmq0uqgniCenu0feNdMfs2YkBG7fCkcshD3DB
SkP5kUkQS525XcLzJByNlxicaRkYEkI9R7opsXCPslTp2IkQ9fkoY50jZGoxVMrm7aUV5lj2H/29
i7GaEh7CLioviA2yEHdUv8srnufAOXPwdJNSkPahXSWkmn+RnQXniuneAToHsaPvZ6YNazgvyRIe
xqNAUDTTYoKKWmldzvtwMPh0vRxY2Icxnmt/ul6YMdRfoq6BBnvzmpRH3xuRVEmucIo7m6S9RdO2
hOyH6629Byu0mpAZhX5UjeejeLe5H1ToApjgaHQ13ZpoRSNAFs2VTjMeUXWOzlCwqure0Kf8o/Ev
wOl4vwzAOQIy6b0+O97LT2blHucDL85p74NZh2fAc1uEagmr58ZE0JzNCzLNiThF6DRu5AsJumEL
VGdNSDyITaH422LXdBesntLW+Tb0uvDKLiMIK3MoJwPn/B86i7J1QYN2ysM7UaY9YFxe7nFCwNQ7
C61GeLGDkAS0k4Be2boOA0LNwMk9zWn0s2A4N77UmAptJlFwjXXHnJj67fBJWhFqKVkUgzTHGJr1
+RAXipY9QAo8qn6NeeDoJrE3gdumHXN+Q49JVXUfOsRHSwjTS5fMNm6wuT3j2HlNYaIHxsPDJ1Iq
QKXSMNIdUu46EpluLhJoh2m8gPe0ornA9511YbpR5MYWVnrX6XuE3/PbLZBIkJNtE3cvCxE2g1YW
bCgqSpeOJKRVJWUuwwyu2451MuDdYvoZ3qWresfidRB01L0b1VI+DgQL/cNRW5vGrm7sc0AujERL
rfM5+z7ONGvzRqOphczLLBF26ZHBJ5zoyz8XSl80zG2d9VpuE+dInqSqpj4dDAuC+mxyf6IY/uF0
ItDxVOWtmmHZox/jeloLbMq1NziwwbVNrj54nI+CMJWaar9SqfME8V8mfPeDF4x/bK0LDeQ1UXP9
IV+cECpv/s8tMp0B+j7jjELqawdLJCW1EJ2X6guB7Zt/ngX5WD6da+7IdxHuRBrLlEpyoMPUa9dy
T4BU3yS0tDu+uSj7eWAdRKwkkybwNnCaCSkWxzL9zeDOgkdAwdfzVIfZx6MhUIXA++Laje7qjdxM
NGuQK5eNTE89QT5p8unwJ+yTxZukp3C2YEGTINiJ2KIae5c5wNqso3Oc0OS2znW40bUS8iBr+/bh
DZLEIDhhtJ4UeXMUEs59jfQGcIo8s8wFRaUbjcqvJ+NInB+wY7YxUfmzcIFo8vunAVlDhmLKNS5b
Gc1KXxCmO81Bd8IdLG3GsjdjHFwOWYwaXQNu0ZFxQbSjcdfPuUGnynD6kwHmvu65R9YlsSJvk4yN
wnT6zjpKL0SPkTRqFzBWho6STY/yIeewn3lpFbreV/cY4yCPoZfUySGwqGgkYFhaRc+nEfyrYD1o
rkO7RhDKV7cwcoFiTlI3d7XRDPmInFf52o/7EDf/6u98UcVk//iBGn8EIlU6Db7NiUbCMikkFaZW
n6e8rN1Rb17LRmRH80569Drzaudj+KoOQJ6hQ8DxGLReeObM0blHIys3bDJpsxG+IUXo3GVMtvCB
nNNeEllwSJdNaaKELNw9o6dfxZKeg6Ac/SY58s6hf+KrRFmT1LptKENNCIJpYttWLTh3lPCU4Eh6
J9elu6Z5pM6S7NG0DCq+0wLy6hHyByxlbtG7NvDpWZmSeqBhFE+yOS5zyeqagzZfl/5yHuFyWB6f
xbHqinhD+bXFajeYCkDMWzGZqNU2sciORF6qz8oh9E/vL1dGLCJUlns5rtAI55WCbagcclzXWJeK
b/aeoZe8YiZlvDtM86O5741KRtsq+GSvggGBp4xJ7JLbdv0jIYKOnrUrCadAsSJJ4ceIH9/7iKoi
tN49YaQO4P+rZdfUA0zQYADPezWJ/yNfhUigQ+5vr9Jod2uGhCS2dxnRTLRInUwgXviXIx0m3mPv
AA2bvxBXRfn/bEVSwFtgWWsNR3Lmuc2BvjWOUuFZZEmHI6eZg9BARg3q+rYjcwI0qhXZcRWfpcHd
q6kj233BMXA4MGsOAIuDfwBDf1RtoJO9yspajv6qe3VX0FHW+VwcGuEBpUC9abSQMNCSHGY/eeUn
ZbKrzfsSUbUz4KBQOUDAbOnJkCr33AX+JdG5zjrEQqRaQxHVF0Q/VoaHxKp7s7lncDcCsN3aLuTu
JJkBR7MxgVPTiCA/+Y6LiBTgW/q6nEDdgXT4ymOkkhMCQUzAjq3s4aq/tdE1c3CRLiWdWJ1Zvpjr
oHYOZamYv0Ecq0qzkdU9haWmYFpRL0DiY8WiIyL7ZVLzSAwxmJAQvZCP3GXtyrejAZV5plyO74xc
F1uclna9jauZUPUfJiF8T/IENgAZowXdbOS2NOQKgjHN8UG5jDzXSAo/DgsJCac0DaMVa2Hw++Pl
PZLlSh7z8LVvo3xxR6jjGoDUeF79wA+xw/bMRZOgsWi/gRjuJMnx7se2VS4jygRUBLRO6vI+W0tS
dNnCYZKX8aGWmhxU6Yb0c1i0RFzJf2Q0AtUVfrFfO+BTZZprMDBC4E6f/9TTISp6jCQgst/WI/lJ
bXO5TPf6YUkc/r8NuNql0ktr5tf0cJqgEVr8hAN+lYaMfqqiK90e6IFzBVETN7LAOlzVOD8lYPDF
W5dLdBLGFxlRp4ZLiColwcQFU5uXNWatQUBG1bM49oLzNQbfXmiTzHoU3Di2O34ttWKcGrPjtz+i
aH7+mmJib29IObjhG3Q1K86z4zVH9AzCI0Kfu+V5ku7QCcD49u8GbtgmF8g4lVZgNxoGMMPpXCvL
iIkofD3+m9OGBAkg6nHfmuOYgpxu6yKfjCOAo4iy/pSjA7QDlft/GJV0jbLr0UithzWCEWAseH4w
YY0EO6i+z14eHlHRKmUr+0yocH1AROvfa0kT/33wKdXKalLmS+QYJemTUAKhWcK47/TVQwr2wTDp
0yJVUZ+1XLCO2Sr9cy05SJWmkFYi49S3GWdFdKiiC7GHFzEHL9WAcyLBR4Qn77+Gt4hCIem57DAc
bwpdSHtiMfcEKp9fDuarjlQyWiJvxmBGbw8WRtPwcwEgaZmiL+XpLou5uAXs3e7CmhRUW2YPG+sw
28n4cADelFTu2QDpHigB6tI2cZdMx9GeuhGy6+ykY1XM2KHfLG5rFA9xwQX/fGA+hYg1SfdVOgv+
svvBXcDrOP3OzHBjzModJfF6v+gkKG9mcWzQg8aKH1Tt+UtLcyBJ7594ZeGR/VQcvx4pdWWkBbyF
plbsJ8YAd1bQX7WCkmEabeUkVHPBiOAbcaQghVAtSZ+qnuy+BcCeO1BVB1z5Ytkih/sn5E8MvFMa
0Z7BRjS762RmOWDoaLRv7etYNRuajFEb98IMiKPQo73bW5pg8VKo8A9gwAmp92UTi+/zSUszot3D
1ICsswKHsKYV/5x6Y0HEY8HK3B437SDF9nxk0V+vMqXBH3oAvepau9FedsfYIzP/pxeORgk1JlHP
YQf7ZsJ7YrvdnMjA8rnv48YSChWPUefsYOQhkcdu5fTsXyiVXtmS3CYgwzqsJB+7o8rqS5t1qsRx
d6lQSyRaLFMNlfwq4VF/1uQysYeSBYxAH80Ofaa0Plm+Y9SDsHpUytzybJWjuU9BN29TwHcs/hqu
6eYNzYLFvA47ojnoVp4ERziawOdSmite+CnctlkWb5tqCsRlSV1uyAgEMZ4u5+HQGHHJh3UD+Y7d
L2BjTVkkqg7ojCXRYXeHc0Qr9/rnTrXS3uFjhHJf0T43GCgNKqvv/W6FuR6HyCDjUtPUPP6iyERG
Kax9RUr824R/SH4NW64csXQBL/uEkCrdgcAhnb+SX49yC6WbAoiVr5bz0rpIvXqwma7lDFG3awqh
l8T1tGfjH4YKAPOidzmlbk0iifKjB2xgMDPt5gAOajXehEsqw9SPa3aP3yolZ/oGetKCNT0WTAVp
MvIOWHwJxtxS5l0Dx9BdsqIUxTMrnyf9BW5owzq6wYNGtKtQqFpAFwcGYLMHvG+aaoa3O7Ma+r/Y
1OPq/KYQMRzbKMCOu+TyA2vlGBwRXI4KUVvCIGJ5eMZb0rFpU3AujHhwgKmnuKnmRbDe1n2d+2pr
He1cK2UU4xqHce3pjNxtNNmsLJj4AC6/pienGUc8CRcZDfkiRWvlWDV2aa6VZwX8v7BM2XQBxP8L
Bc9zVcm/knUeZkrunGX+cfjPY3AaDjjWk+vH8KUHGXn+5OeuoikmYFDINP02+vvcVJ9vMVVWVeaj
RycOGTlffLZLQMab4ilbFpEjBInAxsg0XnrqlV+a5VSbB3xMCCXVrr7CQX/tIndy4QFeuHjj4ggG
oMs/jG8ApJQIPzMuAfzrjQIVNEdPei5bkIVDvZYpfdRQkCClw8VGTFRnQ46cTUGspWhUtUk6pjdN
vap+Et1iNWa9Vt+D4sixgu39w9jk2dqq3ID5OnUjg2CvSgR1XB7XCKA/WWQ8G7BD8fxyRzFjyRef
5QozDaqGWrrJ+4Ojmuu+U2JmUGzKv2ouReJCTQ+dHb57j7itQ0Tcj+7WCPD+IzmYa0MumK9Hot3o
eCGF5Vm1gZ1DP+NS2JuQwzNXsosalZP7BEAH5OBrEaPQiblVIQ4OHxER37buV8nJl3ZkVyaZmmsb
I/Dxk2HJ4pNSAP6B20KGs5IoN2F9HWE3jnQsVusa4qXarIjhLK9Optk0luIgGqmFvO/lxUVYL4NZ
+Jn8MV410j4E7Eq6LFp7YvbIkPIZwJoMwAnAcnqsqaURYnh2w29Gs5ehHlGwFVap6MTUrue8sLjz
3i+tamupWr5Gl+nY0Wo0Uuizs10HS6i41D/9fztCjIhrOuzRKB3duC9Pwnam3SvZaO4q7Jn2gv5n
IU+1jqV4296GFigNPmpyzv2QYIiZw18g6EP2Sxb/fNZIyCZE9tH4wSBbdZtRLYjuRKYHcjgs6nlO
E8My7NCcPVvreTBFs9dbyaekLRZ5BlfDITRu4KLsKtaKJXm3lXoYLWFY350vyu1NXFAsq833PbXy
8QrMT5kkQu9Qoymt/WtDlzsjq754RAVieQTvKWZThLg4APLT3w2xZc06jNiujCp+TifgVldlw92x
c6rFRHBQBiOprb1csZRJyHNdr0PT8YWBwpKnmZeOiztKstk5MyzcXRtPuoFI4TXr94QG1RFHrANG
5I0qMn+lUihbC7H2yRyT4BOLwcupB1dgVByXahMdo0K0ylUYva+tvxrtEvavdIvAZO3r72BMvpV3
mD7Miw6e3sTsHTPwS+NAtgTGCAt1InFwKtO7uA7KkeltlrLV2RVNiTpWUzVqfcECrKEJWl+bPU44
+9lNW9zf7asGwtIsvkR7IEqQv3AfwXnUNgs3ZhHS4NwCHyaUbuIQAjuxk80tez6WPuJKbrNpFad1
IX20sCBPrduC/TP7Zm9WYdW6M2EWTYHreIMf5rP00owoM+D2lC42FHkuk1hgw/Bi+h4tZ1DDKL9G
V+BZVvYvS1jmY7QYQVKpkI4oPXR3HuMWke7FYveq+qE8w0kP8LELdgASs2Lbyie4Fim3WiM7xG+N
yZeqPNf03SQ5ACea1QtknSXN4LuMeadVKHmIFALul69uoFWxYlasEnoxpmVPQbl46fyclXF/0eFs
jTVk8az3m9tP3Ndc4777jUBnUfquc6ZiRvfhi5rsnTQfA/A8EmE1WnnZYr1EFC0723sebt6EmOED
V++AptlCha9O3b5QkJa4GoVjZyRcrX84Ktn2DW/x90d3e4bNOpcoULbIxnqIMobyJeHf5bxTUWAJ
GwKo6UP4FNR+0eYNRgPOgvsrjzem1P9TFp6dT7aMoZlYUjRrkQjCNEoZNfCZmTYaahj+JlrDfJPj
TP39wUE+1TN1mxUM9mVttSVB9RP1bEpztRa+6d3UmGZGYYcWo9jtym4XE2w6eLOE8J7twcWnVxVQ
nRn/1lpmpEk8mTd2+WNY+u68GpmCKFDp27/7rcXR2S+UQMX30ws4D3lG7bTR/H0s/Q6dlMDpUhPD
mBIPjZO+8dAXBVXLfzB2sbbxL2NkcvX2++jf/pUP1bdJv4LTUKw5OUb5aEI9sx/qMJZPF7JB58DD
WonW9z2XSPRXhyj6FSi1Ydhlk9NS86UR0FnfRiRuxQFvL8ul+o3vIkzGCCJMNf7ZNbIbupxxgMMt
KMXa4o8WwQwfGy1uloBTyGdld1OCpbc+ZBSgFv7C3yPIZiSUT1oMn/THP9zfPIAY2KPwHfHd6Kp6
F0Wnzal5aMyFRR0SOCy5Sadm92bXZoO8O7m/nqot6eWQv1wLb5X0VozBD5afWAhVlBqs6W+2+FhS
hPcI3KMpwGKAiFE+j0/vvHTx1ao8aZyXIdcCoBdwewtz7kTQKSCjrOGA2KNLeFT+cZOd3h9l9IjA
pzAxyszu2h8bX6oieUXNELndsqj2YK79XPcy9UN8lageZtPJrYfmG6hQGYR/lbfRK9ceJwJHyI/J
ZrFiZcx0RBgam2b9iPRdZm7pSRZRHVvidemDkXlksiXRoC6haEhTwYap4nNwZhMqsa3oRm1BtVah
MIkYGafDl+uUWKuCyG47nVVUxbRg89oF/Js75SRkfelLbzS4VRFSVbLji/2QEnMWrfRelpXr1jXa
VAQxO/jAaKzYPy9X84SdC+rWQf0bx/9+dO9P1Xt0JrIkN347apU+rGQrfnDGvRmDqbpfs2ihjxIe
movH/JSKrNIJOqwi10xWwqsavhdmJNi1RhLio8zaxJ8VyosZC/ubxKNtxv3Wr1p8mVtfBk21N+RT
CDSnHwaNTXvfweRFIaofgPFIhD3eT1m45GWu2xS35comAJT+jCszdCvYjqcyQ+S6UxtPXkGiEzW1
VOBNr2KYv4bfStQAtqnTZ3fKJkin9zgk9zIyOG9fxaH8o81V+M/cwn4HOeY1XjjIjJJ9mtgTaSqS
XSMfDmfZnWEd09kIt29JEB0mzGIN8wAlt6iw6jBbkCaiPCh0UVohxO9qhzexejFYc4FrlzZ5zdm2
X9oKd2iy9vzLp2qHgCIMIvUJfoZTFLaKJCvDUBt801LXqirCjvxUxusR9Bswf0036D5IptjEq5jj
I6ArNgS4sm13bBf8HrSj3WO+NVU2lvMYuvdWD2TUtbNSyP2HQWFFplfW5xqZCLcjD6v+I4eT0Gj9
ZuP1ye3GTppTv/yvUAYhwzxJNqA7k5KX6aJLf/f82f9alVfht6kdtpVDo+4gMykjEEJVz5gJHxxg
+o9NGN/DK/XjGqnmaRCXSHt+q+B3GR2KiQCR1v5dpefa1yIxx3ZshA53R1zP2StCBBaGzmGlCNAx
RFMJjmc8gorcu2dH0kVBM5shJo1f3zSpr4aYBdMvprmn9g0cNC4ba7+Yvulr7y2zQLXh+CZBoDU7
nPsUTbtrki90oTZ1kc6RLdwzblVSjm+088LSPEIDRi/xf+mXEC2thaHqZbSQqCuEqVHyPd5jjTQ1
JLO54tcMp4YXhnTHVQVUGDm60XyGTJPyr7BCi2JFF2kMo+iFTb7dxIWi0qkBWGOxIH8rd9OjQYSD
8qlMR1Ns/I5nux5OqRsPgoWAG/w6MaagRQODf2t6MUC17/CLkW/a7JFnFsshvDLCiGrNPxRKjc+j
X/h3ZJz64xR7iIfoi1HdoLoKsHp7c48EPNZ2Ax9LnZqKuKhHBl7SaM/ILh4+6f9Mks0CrKn1M//6
vol7QWYwivzD85foE6g6Kd4Luu0rSW5DT4ok6OCuvc4JwFklqSZawkUEX4oXr3sHyHAun+wdO1bv
mwlg6a5QBHpcUWYRSH+5qNwwfG+88Oj2m6K8zNn2/4HqM1JEqUliX8ud9+sD1lPCfaPlTrfvP2Tq
yt8tNg6KrpMoRNKyH1Qz9i5IGxlBsZZzpkJ3PgX7DUz1TDSgpCgynGP3stl+VzIDZ6kw5xwN1y+N
u4PApdPcQCDFWWiRDpviQKh7FWepAEDnlCOhcciNCmPk+JSn5eRDF0bQ2xFluU8Hskco4+KIyqMP
2urdhZZV83ysFmvDiQt3hmuZ81OrgEEhy3ICJSblWs+ZciRv8od/B55XNVskcW8EIRj36mukCJVE
GzIVUC0L3kKvn8r2tsPEF5B03qNLXLtvDiuFq0Fl4/FfP1mTvciLsGxhkdnGUCiey6HMODQBDtD+
4fZ1Tj/JGFAedwzFvDqjsrE8FYwGE2qgn+eqN1i7lDZ+py5XGV3qetl8Htx2ophz44Fn4sYaLcDd
a6t9YOQNBcTMn0GljBNmiKEp1H0O/oL2/VjolZDP9cozp8ypHRAH77F4PbHtlb9PqUii75FOrOOs
2ZVzqc732JcS/9fXgsSPprCR7e5658IcQGCnR4zRkruCB94sMgdIvB3QncVYFGmhc2+Jc8hJ0Fma
a3E8HEeU8LfFd6fIIz/Awx57Py726txy2bYlw3/ptncTbLqYWOuxhTIllXxiB/dRN6uDhqTs3ouW
M677aXg99IogKuR5k0vP7zpLPNrdbhCYYLGVMLS6qZLGh9eV5Jc+eJjvK4UzOxmIkyiNP38pGCZ6
RMnqlRXU7HlE+8rR0sWdK0JaMC0ZPox5/3WZe6EqISBED4Vv7KYRO0V6LxJWF+2NRKMKXAuOmJvb
8kuX4V/+pXGYNZIIKd/qjjkOHMMo+3rCOVcl8CFCM9Tngsy6m3ZFVrWDPRvN/38CCeHO4xi41eZu
yG9bTIX6vrZDGpoxIaBgWVpsW7YhHsYQMsuMIPSLmNWNEAVDlHP3YiQCukLmyFfg7WjAK7QE3B34
T/X0VwLl4T/DW4+E1AimDJI7dKbMz/GBOgT/MYDgRN37+FFoee4NUtrVsYkx11bDxobCvZ61ZmYj
e2+GycDp64EWRTE8XEUP+9ymvE9nJ/SQz7pPxi0w5w8qdpgcA8vjy+HGIqmGix6ky625/EsRGLy7
em24WtMFgCwPZ+p3f21NMIAws0/AUgVdXw6lsz+UdkKzCusiBMoMnwWOKwWYDg07+ts4Wo6tqh9s
XvzEox8anRJZPBW3rFNutYBVe/gmJOFqRvZnhXl54gQwvYBQRyw0T8eBySkZPwb89Hxo/IQzbawu
48HG/FTqA50GYYRr26VpzLphjgKlDzWZifmVGlg8zctCVS4NRtEysDRgdoAhwDOqNSSvZszI8/T1
F5U+66Jd9Fs5EeN5pM0zYKXmzPGEPPVBSOoUn0oXas99QUuQM7U44NUhf+ru0qjy3tjBaBQP4SnH
tbBIXRXSKtwtJcqNuxDCEOyGWGXMtYAQVHzohkmFRiBeucJf/5OTC1HbYMUkdAxozK4Zg5CFZPBO
vP/Fe51jyXJ3t+UA5y40ZHhhcQUTCwqYKX95DM07YUxEGg3OK8m4V2y1aSHcb5SiybFTlmwgqUll
cuSClZteB0fYYfoWDm2Te5zDWaQvGx4l4IQJioK4g2OGyvsYkp2pAFgenSlRwJHHkDSHAiAwQhet
SpkwDZGqXhlfR3xD6wHjpnOzFclIyZeBJD0J75ofIEm7aMzO/lf/LWGZ0Qyczo9QdOF5CVPOIb6l
oAbqCZ02BTJVlP8l1ii4UrcD1OKGTiD39/jt5oGErvNqDdveNIPJXqA32g+OUojcR9LRq3okAK4Q
x+wo2JmVMRSJLzr1JEabtKwUoCGh86eOz/vQnpsyS4KOUuf7OrI65imRCTGrBQ5ZE7DebDbQT+YU
WT7VUTBZRutAGUrF6VTmO26iNUWd4fxS3U5eZtyV9aE1fkB1SMtU/M9n8qr954fOMCtcUd806iBA
ylOS5PWTS2Lqg7GkToTxip46+0m0TQgpp4IRNIRs6rXHIe1k0XV/YvQ5TTFf5Lvuu7mISOae5+2O
f1DXBRk/Fa8Gwfgf0+5YaV2KF5e9NH/Y1HznPI6W/N+yWEqsPQnvZWZ81fbBLFdTEhLbRNZsj9fA
MCtHeklDWUNhjeHyMIZDv6OMy9QelWK6PbsSxyEcnZe/Wc60qvL5toitvAPugZ2CLlNFyL5VFxn0
GOy6RCLwWOBIiH62y0Yi4W6523kZGauiJ3AIwNl8OnZt/itPkGF2HJ14zr/kRqi9ndJJ5KZce98K
AL85ib9Ck3+BqrhpgBamOiEleMivgMgoyrHSp6LnAk6zNNWUkFU5XVwotQ5EBeTZSXYdQiOpt4uX
BQa65TBG7M4PxFS5Vq5bIoeIbcWLbUsyufFgJ4z9a0g5yyI/9xdF8ygxg5UF9WI9zqADmZLUOPhq
FeuEHhHZM4+hXmioY3okXu4vNlS3P934PTmluqTvKjL5shUE1bi4ukspl+4pLg9YBMXyDJeNtMB2
qJj0YoXFsFo7qXQ7T/4MnhMfyrtenWBJkaJcYTghvaFUNFspc45gXjjUA5dr5uO55vT26BNwb04z
dNyMh50THE8zwwpO4E26/Wi6k+9n3F79QU+mUf0DwdntJ9pbKlNbqV6vbe4S8S92+hl/61WVIN0X
gqNnBdC9/qxSNtapRrkxcEe6qeGj51FJ0VGuAnch6z+O4L5RmzjdAmO/3xOyRodUfpJ4IwIaE4Ez
azR09hn/CoNplZ2eKj1WBufbMkR96sO47xkylcsS0GCeHrzaQvJZGPeURiBiQhXmMdC8jYTDyHkT
ozGehJ6VTzcZ62Z772j7H1GzfCUJJrANesGUnrkhJ1Ol4mkKbK7ygzG/ftQqYiiPi08Dqxd/RhUI
vZh3vmhAGclhYIs3my5z7Zzlewqj7DWYHQhmwU4oFTtuy3Tx0To6x+nmyWLueqa9CcGq4gGkr5Vc
ZyrXbpNDMqZgVpsD0T5tBlDqYLgaZad6b8xt6xUAORHuBtqi5GrXEuxF4x2wZ6cRcUU9PKijAYWe
3I6uAChs3tjOoi1NHqrW5eADZq55Xo/CRFaWZ8XpgkwvNZRfvDYO8LyKKeezX7bIQpwtMIvzewBk
8IJXG3pXc9p3yb1MPMkRW4O6suTEWzRlQNJrORuwIcxzxcQr0AB8Oes6m5p6tlRX34dEFwLJEj+V
3hK8Mj0TmY9tU3/cG+hLOUT2Pw00S+vJed+0DEyR2pd8V2dUidgQ38w8V+Wqdp9LNKzjlU3st6zI
VbfaCDsOSE19jzUbA23zmSWoBN6sK9bLY1SeDsLmTkiuvMxKErn++zYeD0C2m1YKzs4TcPBMMFIy
Vg6V4QmcsarRLSHEukecxOBVuNK+Dsfcp5KTtAdTUCwdZ6PdmxDiBiubtBHlXCUUZGW7aYuPbUSk
RcBg9CEH6vAEWFWK3yPW1m4LNIr6fHGHVl1UmO1wErbPJ6ovy8u92MzKIe9bnuOTY4Ulet3VVUQg
TzpIu8U42ql8O6Tifc2p3TvVZHaZFE6ZgKtcd05Mix3uMyVSIfAz0N+m1g+XXUXvPcqw4IwuZB53
fULNB3qCb4+4wY74l1rAKYeRgatAes1wHFyFRcGqM+ndhVpuRnp6k6akDQ7ikTw8GuGECOcWA6JK
OjE/xFcfMAJrPh8b6M2qPqdH1yRM1ZZ/Q5LU6qLVD53zaw/Awpj6N56ZrVwvqOZD6A54pL4aUMhw
5uYz6H6Zslgh0HtLkKvVVYtPvZr7/wF7Prk3TQWNQLp2J6K7m7cdCROHVQFiJZlx/KRiQVWfitUX
vXRufh66Sky7D7swUXVMqtMcJe9A8tAlf5+YjH8ALQRR+eiqUy+DRx0suqgl5Ezlq8aGiDhCmDEP
9T9WqnRD7sLVbNU9L4DH6V67R6/0fludgH6aFjE9zQAiEo0vpmbHugNbdAdiYApwR6EiI3ohH4Yd
9cwitUVVyTAAq7HUzJSRECn7eB54iVcM2g946juc5qUvCy1kFA1NCBpACXCoo9XizvNxb5Gs3uAE
WqSEE35MsHDummiH9KcL7VLstN7o1kX9AnbRXoxoVdN0cWJrqGcEwe+6xGhevGOhUM1X9a9oW6Jx
XvoDk92cgN3jn17DOPeQ2A7HIiMwTB9edgdW2Cj44PexERV166mc+YKEUAUDzW+VjxLGEjzU02lY
xVsRi/US+z9UIBL1rANIRN9oZicITw/8NRv39DucFMbVykRAs5xwLFpqoqaMNpWCg0Ky5eybLIS8
Htzd3b62LRFX2jEKPewv5oJ3HkRDz2AWtcvExCTiMzsklwMQxmCt6LprtO66HcGOmP5w87pSPSfC
J2ORStQHfcH/IA40Dq3ryZep2H/Mcem/nhTVEYnphVTmeD2FZmxL6JNX658kdU0TPaEQNkQh7FVB
AsmVaHhgLflDLdQ2FBGhgLed3ceLVwYFVQbXjjJY+VnHmrRLy90MEipUU9w0udfQMuGw2k+UxZYq
aHZEL/h1d6gcMZeXlp/1+q19KXg1kNGL19GLQA5jvms9Wg4O9U+rPJxikEPi4UKnWDsVL7DWDSSC
4uXQ/G8BIVGg+LKZ2AFEn+aBfpPzDY4/aw9fNF0mhyu3O9INGCdYLJqUqTj/8FFVEY2ODj+Pl7wY
VZuWhaS7F4Xp9plGddpPMP2dDdH62natDkrRSrDF714NnRW/IH/xeZSv6w7Ock/D/dVYaxFUNGmr
RhO01veAdsfHnEqSR7WiqkMnGLJNy2B/kJoudEV46vx0/sf0P+2x0jYvHoG6AYot83GKRVh2v7nX
322MMXqBHp+i95Qgz8uXdoUe/Jt9LsFEh95y7kstaGAWOGG7d+7egPNqq4U6mv4ec5+ZkGZkIspo
oCF2NOZ+A4YEV3J9BiT6MbS1Pdlw8z/8LO7tHTflOtv70/8WW72kx1g9bQZxClyyOayqeesB+J7J
vSp6tOv2e2q8hL93q24VueNhVtnpv3a44RMAbyWehkwLEV4CvOWeQxeKRyQvCoohEDsWZ7EEJ53k
mi4Zh1y+F+KpMwVokRYZpEQFDrAtJ7TEbuD1f52nYnjGg+n8484U4Th7r553inSV+FMHuylsojw4
lI6GGHVBRaxUufr6WiglPxwSVmkLHsSlAqM4xKpDwVV3ErM9SH116ZrD3BwvUvbJ5uLFXFJv3zn+
8VjKNWBuEB233bqCKDKUsEkJGm1tOhvV4duPxsVw2f8fRzou4TZuV6IRC5Dq7wPKOm2CtiPDqZRf
PKQG+DJ8HTAgHzfXFMmGgLdY8xYV7VgDK9DLX+sJgcqUFkcMWZhKvWhsT9F74QcRrjS5kPLGHJlF
xiQvilM7wrVTRHpUn2LjWxMPadsGzQQQbmVkyVsHTMlSifWaohXDt1CFw2R6ObnbrcU5DXQP1/Yi
DbEsSeDqjS4DSLSMdNQUpoMs7VUWiodNXqEjCJEpgUVhWvtupOxW1WR2pia50HLJnu4yjHHY3uOw
7KFA4Yf3CZZsYtZ9or79q7Zc6is4X01jdole1MYf8Zd06AYS191AL0Z6bULJZuQzSXk8TzwliR07
kE8Yusx+SMhVETLkQx2t7MS8w/N2oGiXkvJ22SFxnUwluOyIyjBXO+5ulf8XiAgyRKumfTfxJCny
Y5NaIPRNRWNB4L95ecJzmVRGYZIJyeCQkJhjXZGWoSCNmO5AV2fhtllZDmqIZgvqL/ac1UgvMhK1
r+TFEh1krbrw9J7NXuSdJIbc+ukl5VIlbVM1wLf7ppYdTAUdeGyG8mhscX46SPI0wwR1U6HXmNM+
ZpWf12lSfjEvwhI/S2fMALZjEGT3RyRAsc9sA+UAN0T+dCUs/41lIGO+UGd+kFbFekaXNAd84mNx
iDZLhaw74OWiiKlN4I68Jt1B2s8sqQHBcVfYUnvXpLyWzyTodLom3/app6IcTUHWdju3Mg3qWRl/
xMxC9QeYVd8Jlysb26Mtw0hP7fP1rNGWATg1T6xe5gO4uvQhnw8Uj1ATtUOl4p9E5WoqSUK0EceJ
cyLVBrmWRwVevc4RvzmOEWMaQZPJWAtYfaI0nlCpGCitVkWP8P33P9rtHHioz3s3OID6/3y4f9os
f0eZ9HylzSeSAukVMFpo1o5NuaWbHm7D6hsofeaEK8wnD789HTUshMQVjXIzy1zj701RkWjoK/W+
MUn0ZdQe/bP78Y08yKqxokfmUduk2pVeXD5bz963gKntjlWdJcjkzGKZ0FM53Dui29I6JmZSk9zv
dpWjNaWN7j+pW50pxqPb/5IqGqQ4pOTPeSHlJh58TQcQLDWaoJwHSFw1UOJdMrENbKnOtWL/Ckko
F1EmJLsUJpZsnaswDqOb/fylxnTp9BgHcXPdPYmAVciIEx5W6WlzXLebi70HienbPqubeU25CYa2
Ae3wY0rR7SqFv7vJdt+3YRgMIeJqYODZzAOvBLlKrZfcsnpAglHkWk+MjgKkaFPkWOJqjdsa26aN
7o/PxLcIFK/ikg9qm+gFdrEFkIB2CmPYsLHamUyj+JbvbAB6xFNsRMy/xhkRXbZewAUTPF++9dI/
ypOwcnULQ0ZlNuGUv26zmJZM8n3GBYiiHCwt8tvDtjCpHCkECf82n0woaSe+54R57PkZ9OkO7azM
v97FbGI1dJ59r+tOSzn55nR9cmarv7PTRSi8W8PaxOdcfocECsgAF2i4QZ/4kemM4F94gA1Sh+Ro
c5rDSDqS+89WfVmuPFnY6hNuJJ+GyrZrNA0+PT+yYvcszIYJh3q8lT0KrOzviOkBrPynK9lUSdnX
+xMs5mMivFySMi8LYRFzj5unau24h2+uJBeK7sOQdn2/6XH5JJ8iyJz6r1KxSSZPsOjzGAeasiIO
ISTNjSY8Led3+zuWBiMQx69uycPV44Vfl0XMB5sC7icRIYstAmgXZ5ZeXNvJnAWkKMWsjXKRV9jo
YXJrOxaKo47zmgp2ch7Pkl4ZjpJooff5QztrYSSGg0z2ibAWljSEhAQ7tSJFMGqtXH3ugVwyi84+
ntyyHE/wBeMoYyLyjzSIh81fDnwUpD7WSCWHARluOaumW/L4DrUmUkwXaIMhOJL2cWDaY9K1e953
LgLQ5qq8GbLBrWL3bErxO6sHPWNS/CvghB6AwFidgBQ3rHu4mOc4bf71LcJ17DyxwJ9kfR1bKFTm
T0Mflyq/4i7wyxeFgMhjE9/WiQ4fEL/UgE5J32GQqUDcfK9d2pw2bG4HeTzVJwZFkeeVDdt0OBXV
OzporodmONf6FfeRcwHnHszEUPtwt0dvx7eTv4NG6KONk058F6rwyb7T5OM1aAVoZUm5rPK0/2td
yEp40Qy2+vHPAfi7O53lnbV+EFulLa7n3vWqg4z89o/1gxQx9HSXPecaVXMWE9SZHIUZVbq1xOqq
HeYeYIhVjxC23orZwvb6HuAC1I1ATt64y2htt3CdlM8+C7KYviJ75XDcpBDpd7mAZcwboDimLTZ9
LRlj0tlJhBwwTZFwZY+e+F4fk2vwb0NKkY7YmruRjT64/YIlBTFGkHSObXFyfdrjHXQuGcWiJa0v
512UDF8pBfnFNNaJyGiErtaZV5iVXuo7xZvhj1rPDhXta3xn/WNpuTDRrZzShwcR+ptxF1hjVvCi
s80G5fJuy0AKAQ8JUls81Az7/AuJV8LhoD3b9If2TpMZ0NwWO6W5OndxPtnAKEaNr+tKugATghAT
Ytw2phONjySi3aGlaJHRKmBlJoz6RvCS4QDof04BLewz2jofzT9K4EgSJEUI7r/+cS6px5FhAr2M
BOC8ghEVuiqoFXKrdybIb4W4Js6CSNr2w/J8v4GoFR+RsFy6Dd6gKe7vxVFFzv0Dng9BNoC6xyad
kaF3ajnDKEd2Djgo1PTDPTSd8Yr76NPc88Z2gE+VlbsC/ZbmkN1Y6/ZpPPvP8g0tcHLgpAWQINvB
lq/A9xnFdk1HvoEpXLIiemF4+GVDN1YghhQcjZb/pbcyR4g0fXwY+wM1M7tdTpX6+WoAsz39gCKH
FNVZ3g9egPP3NY32lIRDzOH658dcZD7s5wWFx53NuDnSWJI3G7LjV0EIggZMbQ2XrnNcxJUKazqj
DNZoNc0RYWc0StaWBt5+I6diBhnN7CO36hj9BIIl1Hvfp/CKc9hUyfD/7gb1Imv4JnYgmU5Tcxz2
iYNPcoH7VhLfnXOwkyiSGCGrQ41fJ1oKLm1fSdQ3LEOFaI5Mlh8GlFcTdH5Rcj0Zzmt2pFSRmHV5
ub9mkeolIWxBn+sC/ra6Xa5CR8MH/8h7UYOgKRZyy+s5nj2O2mytS4iFhTBIO5JVN2hAE5aX4WoW
WtaJ68gTZDOlQQFE8CMBmGXebHbxGorx7Fdn52B09K9wkz5uENaPeUoRUodX4zMlExZlnJWmHF2C
QD8pmoXk5yYMWASKGoAtVNkjKFTCOBHHENSAYKX3drUelmahaGupnXexyDoM5I1g+flO68GaTX94
DugSukPdaGLKCBURUXdZaXhEimsu1tZlzCswSCSsgOYNrKI3SwYZg1n4rIQJlNkef6/yDIMIcYLQ
MNP8QIlHoSMLyc62WK8XCabmBJbkijWph486Wqz/0RAX/CMHoXTLCT3ykPoSz9gF15GoQmH9eiGu
hWbHMSHtmRYZo58QgRO5/OAR7fFP9+YBwid4hT72U4IWLd2rBCiaBJfPrAjKrr0bTfImTHgnEBJ3
qDAF5sI/p17NKwFyJWwUXEPQQWIhdw0OuXeUiSiWKyy4UJinhzopa2CDciNejh/a1ZABMXxslh2e
lE+EzLYM2rOKSu8DjH7WVshNiPF3H/JQG5JgzX9jrGYFud+nqJsUlJ0vVuRLgs3eL4V8kwoy3r7B
kv7/NdVJOkvo20gXi3gGei8EDkBugIFCzfX5FdeVl40OnxD+SbgAD8qociMQjCkkiNhRAc/08aQ2
c5WAS7b+YGO7hmqaEQH7PRbyTB5yLi3UNyKwt9GdbxzS66gypjXKmxaNq/fOoPBsAbbg44M3nA1l
yqmwWk88WV7gBCetn4VXo9jQV6egVaePqMfOtQwNX3cguhsTk83v8OIS+3NK8yUlbyTI+2yypxSy
5s6Gm2f0Z/3rifoddD64PUrsLx8fZ1qnS8ifhioYGytGNVLhORBnVFO/bjuQTADblRmt2rmQk4QX
w8ChKqzOTXiDcaKEg84ybtrbMkLccuyeKJiqmHwDX56wp34VvzetvYRbVaxrtfaiYQamXc5GiATT
rHgborHVfAT/x4t86bbQd8Dj2czk3r2Baukuna1dGGRRz/j3HpjTeDSOu7T3W1aeFO9YoVKhi/8K
co98rwsSt0r4j7R/RlKwSddwyF5c6X8Txu91LzANOY3baayd/E5i5VIBJM3ICwokKyzNloZkGnyB
jWDci6QUGSjLEy6ENoznv4Jm2b9KqCw8iQcNHcQSV8Y2CjYM4b59RgI5VH9l6w1jicEV9NRLryxj
qq/ZOlwQyrLVDNDb2ttaaLT7S0uOQ5X2aYsVwFPzlv2taUT+7P9bEvqnKasSn6+Q6iC3LGMIzEgm
jKSQnZ2W8hR5iVUMDXKqlNI60dBn5Eascr67XkL/Nfd8BggPTX7qfFdLUUb/o2ihMFu/DWEHQzvs
ce7UzdT0D9OnlYAFcCIF9R5yZUgE5VDyHYHZsIRRI8963U5XHwmCSMnRkgnDr49ZbKUFQkZ4+guE
/yr53wddWArGHrstZziARZJMn6f/Cwly6jmmBP6UXve2TyyCb+G8+uNOPGy+OzWW6WN+Ir++4J46
SuB8ZEf3cnEXk7ykYp30Fs2aw/WV6FL+MvUVF9TMVKWPcAO2y8diT/DSiynJwlznuxvRHdiUtrn/
VwCilWT3t7nHQUwzzR8vs1KQEf8vJ43vXtwhDHDD75QOCNUMCWX+tTRxFEk9I8ZZS9Z5C6XaoHjL
p7CBA5NoiV8jYno0BbVzCshFzvU37p/REkMz55SMY8E3ijLd/as+QYQUBC+MkVfm4t9DFj37iwt3
A950nr0szWBl0Y22Q9KvSiP2lwuHR0b7EZiBuj62+A6OdJAF/H07rCgRJx8Mpq/1PXKO6ydB6P6X
sDYzbCZju/e0aBgsXeJrx3rbD8TSa6ASx/UrNioYhCCoU7BAQ9D+n8ohkLJ2wek1TyTDDfrSGlrK
KPJA+5Lyr2skmOl+ccyY7VkGjeYkq1z5I9gFmAeGRVvyG3DhuEU2QUyOwMLgbznXKQPmmG++Za3p
W51SYuT7ZxattTpG6GOvX7pAsN2SUH20hxwwe0ajOkpshCiRIMXNoOiZrMsSHAdeup6yYUxfxIfi
/3zyeMnyPx1vSfjPmCUpiEgXGGwhLqpjNwIELsYJSlSWxGt6RngNcln1m2jFnv9nbe30sjT4ss93
1WHMQ28fSlXXsqzB+H9jEyryTz0vjpX49TOBdVJSkOSslqpZhsYwNolCpYC2IrDiXgVkaywYShvF
KNXrQlYV2hVTDFsrjQ0NSsmYQH4Sz+kQl9vmCWXOCvEe1H9NQUqjWshk11NKHVLjw3RUoo2YYia0
hw97czps1ZmCI7RRc/WaSQEFQmYjN8+Tv/337MCK0uaemI0q42MmorE5SHLYRwh5HfmXMreNMiuH
wSnQHKLkMBX38nBAhDYgMbWgZLhxezHhZIGk7x0K1DpXn1WkjmDL2aQdd/tGGP+UGi5DG3PFzqfL
Fj+Bnoj2AN/iAoumSOGHTSFHOrKlWiPBkXrjrpICDhH7YCvGu70p54YXXitRmgFePhFx5w50oHdj
ChI6Sc5d4IpmENFOdlprba1WyiYh/UQWxcZq6jjYuiOA2tf6+IEbE7NyDPLEZ8osQMAwcb9W7+x8
DOG9dQ3ijp0Bznr3NwdpbfkuRXrLohVmdxvHVk+0hPC6U1as32j1z3CFlxbEGEXwu6aMLjzO8hIy
SaCeViInKFvz+ZyT96+EgtXObNp/w/G9Ey6hz5dGa7Ae1bgKCUnZ0g2gUXmfxuhmrFtiUa6rtQs5
PabQyLueDYy2jqnmcDXsCuDkGY0Q/oSS+hNdbwCMusQaf5m+MIiTfnm+tplrTEbMVunFAR/kRL7N
kQq6zjk3CaSkefinltyVMrHRfbVcn1aXBSHlNAN6KPGDet0pKAIknfl+35yeq/VltYMbv2XFAnCm
L4nozgwj+E+i1O4zbBFLW/pVHRVbAi0d0P0FMskOjTIPxbgiZtAV0/RrX4I5sP5kzyHDbPJeyXlk
FuyY60rKfysYEZoYqHIOVpRriLLXTQRZG+oVe5Og2piatGtQEyxU0PR8BxuirrNoZZIwXIUeQrZi
LQjQRpk4TElNbUeVWNwBBBrlmM4/B2/A0MhJ8yQ7z+VwBiTKtSTE9un4O3Vn+Qi6v1hSetUVXZqI
Hu30d4Mpe4X3HT/FN161aVUjCLaHMrj6Em7YkrsMYr+SXjVNzZvNxfGvjRkYlsvXKEN0sij2DquI
B4nN5bPs/f5NANvmfzUcIyzDVoafhh2qKW6ej2cr9C9uvbWaQX0fQFJ5v2rcXJChLpUjaopT9XDJ
Vju8jaLjkojKRVB2ak2E7OBXMxNX10MT0zKgye2gSiCzXIv6tTKJwmXOCKo0isYmFgLVX/mz2aSN
obju3P6SULrCSOANqSzGntolDz7tXFtQe2tMrMeK+xooATiCwbGkiJ6d3YjfIEg9Q37r2/sYAAfd
6ZvjqG6rI0rZVWL290u04Pj+ZFeH8hgQLoqUZBWf6P1paMPyg0Ialg+P1p6f5s3QNEtqEUdGchri
RxdQN+vtmhncXU5cWLZa1pQIJRXgiJhVyD/ft5xEek2rZKBoJbeeM5tlKsxCr7koxLapMIXQEPQr
ShdouMrkXTpO+w8+RN+1vfaKVNLy2SAhaTrEEZidqJhYVyAHK1QPK6hA15rUuqGXpMDdR+ahtBhE
4/DZ1CZLrVrzNsV6j2hUgFa8Hdb+e7f7dF+EMqIuVT/1PPX7jbbG1rWA7SSHYIYH5PqpEJYDl9ky
eDj7gdWA4KzalpVKfZQ5jp0GfpA85D38W0gFrr8tkn1ji7GtAN+gHz2eDcs8/YgFSHFh/seSTvHS
iMsU3jkveVR7YZ6jyB2CkjT8qR3rj4qurkaDEuLw9rHaMWejmQFBp0ik1T3XhHk7yZJYMTW209S7
A/eWBV/P/OADfRDGQLQlexyFfpYvr2/95w7+pg52rZWyhxz+xWI7jzd7eNweN45AF0BTBRY/W6kx
UBcKAwhbRA15hOlWtzEEwC1huXdIuWmaybb38G5L5XSa+2x7uYpSqc+03fZ1abDx6y1UDHg9oDry
DaixozFkCKQFdoMVO/r3+7szUITS1PRqLxEF0hBRUQJB86hSmfouIZtbTnAV9ut2zjIqA8yOqhtY
GgmmVbSGJm3NaiWFqlreUBzc3/JcPbS34OWGlCSh8av9T2fGIT+xmBo/l5rdezN+F7SKzsPMIAls
SvfDqcobDH5oOCCAwuWwjH/5R5ueOlTV4YkpumB64GAE1wN6/HQegD/U0sX93jp2Fi/JdTC3EvPr
mjE4Vl+1nTi/MZfK9R3F93SIBLdcMUJ6bvBjaNx0+GBLnnGdo99BEdHVSitHlVsMu7GLrCf11HKG
/2Z8vaRFlhhZmnS2Pfb6o3SQkTpG5NHv2a7ZAWbd6MO80bwGYq6tW09xXrheDu8PxeWsGtVRqp2n
k1XgcpEku0l7Nq/mmg9kBRDyj9yqXjckCSAEJjbVkI/1BuiOvx+B0AsAW9Y4IgJRt7QjVQKt87sW
ywvkz8eU0frWauYUtGHEuNPpRZLb0Ii0Ta55Jtx64EcJOqvn0N/7Et6Fu0q7+fLdY393zzDZPaEd
C36iFIRX03lThsB0laZUxuJkcixIfuq1a1H9qYvGQoI0gyG8BNx8BRv7SIlog1IjM7ETVu1TaDqS
UQK1kr/gQT+EQIABd6bs26rmuBVKQcmSGqGl0ETm1lVRuoD0nuSZ3BBEgZAZ4u7yDW34ylEhWHu3
uUaFXTQnkzGQOYAur7ryYLYxHtag9iWTzgkFHbSrfkMwqtS1L3ezbRE05BCJZeNgqaye4URsQ6CE
bofrk87VmDdwqeu8QV9ahHOgajg9tK4nkSGAnLXmL5NMG6uns7F51R9t8RsJYy6CAxmb54Zh3C7B
J2e16wn6o3uBSushbDdqnDdAF8H7AlkGsD6gxYqugEhbMTFNgI8TQy77B4RYUxm3B7HBObe34gjE
NU5BVI3aurhiIrlXHrC/MK6SK5bytOcOHpCnKw5F7IFqciXwit3yDzPJ0dyO4tjwbM1CaIxmiA4J
mmlYgfc0BvFmT3bQY8TTiy+jxWhg0UYPf6hIyQaWcb2xHMEz5TJGvX8Pua5tT2yEiUMDpeLcDljB
jFJgVE9hTtV3CondixDTLsri3PDsIZy+XVHHSAoiCCx8PqFDBCTfYO/r4mnhsIZ0PNcEuZebIKEa
Rk+LiCfKfhPav7xeH8aGMuK+ieDUCFdpy2kEI+Ek/A0KZBHuW2Q+TzAORdJ1nNv0h9+0a6sIY9rX
+qk2nRSFMf5e/8iXpYQZ1PSFtnG939eKC6+Jqm8jyjKMgVkgyO6C2um3lIiY6Aud4LDG0cSxY71I
xVTVg/ZFoqBoMHi4GIv+ZiW9VbXfb8aU4VU/lA8kRzot9LSFGFSLyNaHQJPKPp1LxI2Qm689JvPZ
Pm3ikyln645FDqbPtk/tl+Dtt9EVLXZdQqH2lcBsGpQlw0r6HRmPfQdbqnt0pp+BVz09MNzgjpyD
3jscyme44AbGL7xszTEwYlIGI8zWsbKux81MvhSIltz7sfaK++8ZK14SHVb3T+4LrSoN+XUrlXOT
GFeHWXXfBrJ4Ik4fGy/p6iRBPJ8LYgW9cVUIEyV7mnaqm/kp3+MaFP6TSdaMUrcR84oTSXzM/B2I
e7EEU5YpM5gqXWfiAaofYG3aqM72NFb2LtxRZ31ps46MBKdu/bCG40j/qR5AVKo5uo/mwhQY5t8r
JIM9W076DUippgdoc6xnZLQkRmiQijXAPe9qi2bZS3q2ZZYrznUwZKHevH71/qO0ofsrChqHGeYI
7ahRAsITvew0d1J/QARi9+if3D91kv15IRtASiBUHQE3WcVpPKfYIFN8TItLejmQdl5tRMNTGB8J
r/hVFvCBsm3fZKQQgdFGv2krKWidocq/qxNUR0D28dN78/43B4g5qdQMryyM+9ZiZ+RAqNuyhGST
7ogi7N6xNuex2AzJuuYx55XnHTgTz5ngCT31JndMOKb6QiGEgMc+DKdXOpFooiz/J+7fl4tOQIKF
uffeh2IUP0k2F/EXpfrzJ71ftx0cpM/vuF15iV/5+gTNbcOu7TKJxb3j75/b8TGQlqAYrBTo2cer
HXQSM2RKX6PZaxXiDAw4Ok4cjT87qVJW65PNqZEn5AvLzFrrgu5PyvImERy6Qw0KI13QCZ45NCmK
4gEFFbAVh1ND53M1d4tIM/M/33EtTLAHbcxy8gjX4bY42Hb9LNqkou3SIcJHSRs5sdfEaP8KFFRw
NWEHwQsf6Sk+xup6I17z/EQMbMLS2d7ny71+4ceB6SVqYMjHDKM59HIyVKvZeqEtRnM10j3/qHS/
J4oeYwtQ7Rj67ZYHHPeVxfDAEJ7YCvqaTQpjuChmPXd0SiuE6P83XSM0shphF+5X9QP0TuAT7z1y
GTOdukBE5aBjMUhRdg0J7Zm3H7EYruTbiL6kqsTzX8RDeKKFzk7p/Uz0nR9FNHRQ7yKnQVKqseFk
W3nLESDQ9BhPvoCEp1uKBiINEYwo2MiAoRI1PDWBtlbUweaCrDj1IYOB0N4p3/8D2UFkDmrHRgDm
brX/g3VsQ5y2qntzXo8f3gSdifyd5vXSMfMQx+qsfsPJYCT+y+Hk000FndoC/UECz4/V0hsJ3gmt
XGnV1WGN7e/nX2vysYYdlx4alQ7NGqv/IfYYv/G7dgsWr67cyKnw/gg14OSF0+ludwVCx/a1o9rG
FZraZq9SmdmEHkkEZwQyZ41nqJmSsJZFS3M0/kjTGRWaGcmH5pxx749Wl1lhdNIMysFzzoU5w7UE
balvEtYqyzFoU/wQuP8T13JiIR4CIE8owuXWPHPYxmO5gZ5kf9vtGiYlhG/FtvLxy1y060gjn4Kj
v+qttzFgwRI8B+5DEzVSMcFKBD8s+KDFQ7/9Nl0wb/hxG7mLX0DswfScI4xd+zZTcFcV8ftC1U79
TMmGP76yBQ2D4bHTVIjZD87/s3RAZUG8YvA5VRHGy9p3BUhLZJSB3y16R70Hin13q0W5RVCj51A1
VXkk3O9pidT7/TJ9XyIe4JE0ESC08Z7g7qCdkwwA1iyXje7O9zfti/7nK4I+N4Vbzh2YQb9eUutF
WtB7zs4VsdesnvjGzW+WuJiTPfywFrWPg5kXdr6jP0RjrCUvnSMoZ+u+7syye5Q5et9IWwWitCQl
86tlKZMVBNgF5LlGwSOPMZ2EY0pPJEeqk2uzQwx8pOBLYFu5cIe/G68HjjNIAJokJIQ52zmpQdtI
ByebKs2gs1Ebsr0lqmRAcCZzRdeM7aw9Ta4BdsFaYqFIOhSfUsMrbtOJoz05ISXD0Gyrdufu7Kya
TxbIA2ok8K5namvS7nOLlRxpBK/ZKq05Rwy/jqbhW6xsFmNeY7+sUvo9vuk3d/AKDyFfJnjeERyt
Ph0QBQ2ERO7WMFfzplejKXYmQ0RykL2hRKIqHbAvbI8DLRq+qquxf0lwMCA5rXCQW8A1eNVEnCf5
CFE4tkeHQzQ5SLJl9gnmjXycsL4mUhN2WVR44Lvvua1YSM6C9Ce2wT8C9onmSRqVIDRiomUmYDDf
40qebKufsLAvAHGFYYBoiQG7cuAxqlCwlcCw2Nj2hI/+FBMRtkSd5+Yf+Eph8WxIqWypsapgG+ZM
6u6z0VaxSkaA5yja+AVvCr0//HaaHXTfxDwcwLUI2UYoaj1P/9gfupn7GJBlOR5y/XfnfTCfiBDU
5LD/AmMgO4AP1uqZHsnd8aNUzb5mZdAcDzdmo5rls2cG7zUGNAC9Kz5Yqnzl8IqzmtRa4p/IT+Zi
M8zfSHNuA+E8NwpeNf0CV36h07/Sm8+HMs2Ko5UA+IinQ1/Q6I54aD2hhY6DTsMBDaJqbx5+sZFq
ohwUliYOqaU+qL0LSM2DVvi8gT/VFnBC8zQuWlLb8QuO+m9Kg5tfC5wlSRi7uKxRiSqhSHil8vee
ftQX3HMT+nfnMpYX/BPAZtdYgc23ssehy5REY4NsTo8GhFhqLSqn2Kvr3WKnnIFCqJAvKYqcWbUt
iRlG530kqHEVJC9aPbHd8cGVQwVTTF78oSKt0nrGj54XCFTIM5HFO5JAJ4dLp2pLNbB+3HGQCfeA
UsGY5YZ/Q8ElULB2DdZhD+f3j/zJc1qzkj+QRuYDwsTrYfsS/52TAXeUkJxFmCr8z6KwjuyLhG0t
r7evAFqaqgWaV3vSL1g0f+4oRWSOGiYqkFMOgSVisnTtJB3tic0yicvPCxYU2hbglCndCTWxIUlN
9CxKYM2g8XISaY2h+TWDtEOoCNL3nPYhtANaUib91Mb4fE7aSgZk8grHy+dH799P0+bpB5EBZays
SMkKAc2E9IEItWTLzP/y3UtPV5XQrbnGbenjmHc+c4WFFLnad5WPB0ZEACvSHrqzEMhAeKHi0/WI
dFXWscPIHOt2nlZgDaeviRK0ofee+0Hf/d7gGaKfMgBq3PHN45SXlEkGHWqSj0hc5rzEUhhSqK2Y
8L3UbhTIE+CS18chdxMdgIgSPWGeS4ATpr6odfTFeIVyqHyHSzHKE0vxgN91QCevjU9X4pwKJ0KL
42m1nqxzZ6h17Mbhb5M4MVMWkyy5kHG3lkM0mocSLrsMf88ybEgIw4ecRVouYZFEYL7gWl/hDrIm
u5s8JE4gQGknDRTGRF8GgSXX0apXV+j6Ygm00r3sgk+BmjcZw5RsaQ/L2/oYd+tGk7CQjDN/31VB
EJ6/YPIZrzQ6wB8D2pk8D7LY+VQb/DmT+vX2Utv6VzrH34ZPMTL/4WxUNS78ZrQ9PENCrqeaFD4n
CIYR+/EDfhHFL7zIzskxl6PjSzcKvO5tm+Vo21d0VyQLGpIoBzVw93wcf9m2t22Pb7dPDJrzf7vA
TcF1LHXdEmK7eneFccM9ocAhg5sKRo+mgKdqGVMY20vhSyIgHirBIo6UR6ThdHDzSC6xE4K/7GDv
USo8+FDjaT3Dziv+MmmCVzUS0RG2dxEqYJZsmB8vMpDGRW0a0tPAu7hY4egZ0Se+YPjGnrVKAGdJ
msEdo7CHzKFXoHKqdQWD8sHL4J3DlXV6qwjFbirhfYQZoQUeaIe87jDdDffd3e2xQzp6zXhLkaWx
GtOjnKjRS3YtGVEDivl/XEJ/H0IhA24+adb5uVsaZwkY8Ftk5bHIFRkAjiZaDDTl+pyTF3Dgsmuw
e9vvsUC8lr07sNhHrfSrAjeQhXuV8zfwPHjYXBe2EWKjpLEUoPDJMgC43dUj6pirrKUTOAdMS2p5
k5ZxZM4i0uymA5o5lCDsSxb43F8Whu0fY2BLSzghW12063k8HTSMT3g0P7t8WAQkPN8QesJ3/ABT
WL8B26dRYD9EaHLLQ42yvkTSCsnvmyq9xj/t6TQ5zKLEP3wMko2DK+A+gGNE5Yf2qvyvZn/JU3FX
R4SyvZG8pCJT3RjDG5dhHeFKngShPylk7y2D9JrzxSernX9ROSdPB5A16drnKylmHDGzgdRv2uE7
k5ayqCtFhbsw5KcdWUJxllQZ3sk7Do6/F7v1FSx3s6rppUxu5DLO7y4baF5/nHuk57HxqNhJXkNX
grep5h37GHcCdjIwi08J1IHrfHtpFyCiW+6xONWRG+YyfZoBjwdT+1vY3OuarkTIBhMBo5EmLzq1
IhsalB6ZED43GG8mAPiJ+UMd/+GYk0/gREDTeJLzXlG0ygxnpNjjSHYi7jX9C+6Cshufp8zNf/Md
wBvXnfjuzYkNYCoSQzKPY35XfJgsccIaoCQmEtvNAzGISwx0AQqMCrsqto/X8jrUAkuyUKVJpbJY
VM1HOoa3s+zGjXusxrbhz6o6dsm2dYwebSYxmDbwE7Y48NUfxlDcZ6FPP2/sXkn+awZnzx954smr
e7t5ET/buIz8Vm45f/ukAKDegiPySiSaUiq4A/Yv2wpyB7osdPmqBTIz4TT7Rt5VTrraUIdSqcpu
cv4vrk0Tlxw+yWActC6/GzSuMkynPFUG23Sr8dQkLEQEfKHugj5LthDFYoacxA1ndARSa2FEDxcW
/L0n5DP0w03+k03rtszztXOWToc97il8U+r7r4lIuTzPUBhvGhQKuO3UaDe3vhuhq2WGTHayDmPG
K3zbanu5QUZcE6k9GQsG6augVmucDIlYqdRkmeX39pPsvpmQSsbkuWjZQjka1/9kZ2OfX18cF8cf
T2hBxmKwMI0uYCL5Dwm+qmLk8vqJpRa/mbvnE6antj79l4wkOFAAwLiXO3fQZQy5szw/bkrv5sP3
i1ulbaYNECxuq6zZpMfL3ovt6H+ZlrJSp38ihONAZUywK67iT76TIihWXO0a8yObeQ4SN7+Kxg/v
Fo8QUAIy0iDmXT0WivkQ5Q6zV9/nvsfN5jhSrltzSmlJxlZfRlF1pgrvOi9IqcChWsj57Rop/jsW
UGjxZeqiGCRko+GYosrBmvF7XLHZOeE07zljYbCs9RTqmBZwuJFGKj03l45P0l//J9qo0a4LyxXX
qD08kRE9LQfZS6LUBSR/M3S48TkM2dovTZansKlODDO49SR6zfD5tb53CbOl+faFP78PSbNsBlFf
HrlrUWN5TZiSb/k9/SeeibSx2O7Gftv4+1BthrEvYfXFqeRfS3qGRU332dtXzb7aAzI3D1j1rmMa
eLwquoUCwSO2yTl1a6CYHAXTCjqaWb/5+4VQJofS/FOOoji1J5lxHop3AN+bYREi7lPfGDz2bNlW
jv8L5rzbNlNACr4bvVUQrYgnRZ4LmNnw16JuXzWYYfcwwqnopv7zgz6SDf1Kp0KBF8i5e04Duaih
J9tyznPkyGhrulosqnuIR9wRvahLsel/IWhPT2n4n/fjbnn4FICq+9MnEG5xdCZOCELbYYXSdI5B
MBuxlfWOfIY+nGg/Fq9sb2ETXOiEIdzaYiFfIo/5+H+fcKTg0hO/4RCH8sO7ya0u4OJIY40wsDxU
cYWeFe+mMO6OgUP4rh5PPm0QvMvC5fNOfFrNHhO2kfOsEuU9WJear1+XtHIVStyRV/2G7kNAZMuv
A7K9xxsZ6OgG0ucHsBDu5PlZCZJMRrfLL3exUqowNa950LAPmWRrMQgmgNFOgL5wAaBlBKe5J9Zv
Y4AFci3LvciHCMrjTClNknzDPFqZ7MnxqzS0umf28TGYzncgX7l5Yhwf8hyHzjrZvf7hAxDWVGnV
zNhUpRXNtqiz5V0pQAqx823t6j6llpg8Nsq3LpukmrQ+plHAAPR5c91gWNTk3sOhhJ4HNwaS3vNm
CppNeKitKUhuLGglYptBGcRWZq/lUftzd/KKx7jxdOEgFMkamIWxNRhllq/LHB1HLxFmYJQ/p1xL
k2U6rRmedNAJOKWtk+tnqZhZD5HjmByBCz4RZwZC/5SlyMs49laDfcoTK6vVM96bR5gAuHrK8OLa
RtYg238ql2ol1HD+yvg5x8E1TeF46j+C9PlQMjFL0DR8rb/KXB2tu6eV02ksBg+sy1CSPf6YpR8k
MfSM03iEc+oxlJVJ3nCsV4TxdcJoxdyD5E0z12VDuCGdi5I7QLD9ga/T03Hy83ASfZC0wMvSZsNS
KzGMOgyXf2SeK/JNvjTeNywpXja8U5Qp1uej/rUmvyUz/TWkN9GerOqGY+X2AKm4Lm4yFh+Eu2Bj
uRNVqvScQxaZWuL1lK3oUQhLPoeF80jcporB/ncprOr1Uhz2aYdGNvI0tAXk92Isr7ESt2Gtx+Vu
w2+w6YRaPELNy2nlOiTJ2GxNuhTmhQaWL41qGANM3uHnXpe17Dua5kUMcYTgP+W5fRAFeYxbXwsw
x3O7tC9rq/C9+QlbsbUDT4mWz2X26eZ4sFZ52+uSUwu+Hi2G8/OKISOWjjexIoBLjwr2P9RsyFPV
iKJKWvILpmPoKCYgY4lEZdj4XZzsh6CT2kpCb3GG3Eswqx7DimGBif3Zziat3O4GftBVT3xq3t87
cDzJdg7gJBs9R5azcDk+NjxnQWTekVV0TYnaPflgXTt7QXrbpeTiuLQfis0CPxdNW7Y3OWgFKVqS
q4BtARKAoL1Hxaxty0S3qOvL1cgO4dFIkxRKC2pJM0UEMjMZ7rMvX7U4rAVs6RfcOi4NzAwUlj1Y
Urao3XuowUKkr05/7mH4of/g3BnKTg4KFBAR/zHyG731+HDQsyVrgYcHvq/Ne5Jw837eSbBR4KrD
Tz4QLPaMgqLpvgBSGWkt7SISncyvROQtFAJrZJx0tjsYzWZ2CXj7xGDQB9j+vIdfGD4O4mM8JwHz
cg8N6BOzH0qFf41mYEnpNuDGYNs0uHZkHBpxgq8300bn03rEKsMx3nlks0i3L7+xGJ60s8u+KjRg
dkVJpH4Fm9fu/euiIJzV9YGMNSko56ByEg3X8LkibzCQeIi6uKPO7reJgWZWmNdwO6ZOppsV+ko7
/uSWV7+csoZMvDWq+sU9BOIcSBQLAinTkDDAkz+kxmTvtqHrh3orii1JILRqrt0l1Bm6I+24eZOu
KLRrj2tEZcGjlCC5KylmHJNViUVCESv7BdHjTSYPaV0ZatFSv9iJH3vvQadXp59kTeLgNHuBzIjV
Y6x+K2uD5IpofX8Hs1Ee1Vcj0PYRcWmj6wC4oOin4TGUbOmatecThIAJbnIgyt+gBIigOBhv7zpX
7wNg3ebrjMjVGhHv/gzvGOkl7+0mMCB2W4txp1Fn8CfIQLMX+Vly4PWgNqV6fhEjd8aWWr5qcW4J
0UL58na4nGB3/8ZTasg/0o0jpQSpNy/OG3D4o9rdcJlsl7OWNBBnnbpZsHk/7sY1v+QqPOfFYAAg
xB0h3n9WWLowLpdvlM/lHCqukmIqGhm7gc0bpq/VHqYmNZPOhL+KFH7wo6gQ/yxdcHd/bgtIpk1A
laEoVCeQMnhneOQ3SK48qfl3MNXOJG4MHbWWfNaITFZKFQDXV4i/P4MG0iugRxrcXvWoGZjyAfvl
JVTkt5W5WboazT/lKeOGZ1q51Xrxk/3fBHHkvsjYYhd4MVPE1LpOiRZCd1YtCfeyvl0LKALA1HoD
XB0P2wYFW2EMrtmAX/+Zcce+/nCx7iZL5Uikd18igXMjJ6oQ26PvK3HpUjzUskUmUg189rP92b2/
ob+D6Hi41Bkj3qQW9DwF7WyKTGZ9Ch1KBUkKNDE6t+qJccC+RgtFdUAWAQ38P1gjMFXY8/aIw3zA
BAI7Yu+N8eEJA5NFHEB/cfncfU/5YEiADnEsCrp3Py828RH91gy2x2Rj4v7oYr205FQYQCQ6bdK0
dPZDsnfdobXkvip1H3y+W0J8E/zrj/+MMaxXHjdPPlUpMCWWLsuz3Dk/d+SdEFHwJUOMaZsrgSa1
s6Ey/XZGEHQPN1xNVYe5zqssUc0wClqEmtX+OxCpKwApw4lP8RV4BSOJcl0zVbu7s9frGekrrYFj
dWKAIgGp2Fnm+S/1HKeiXqUZHXwg+VrOYLsMtvyFSorV0+vNZTjdEHcJq1jHQFJzo52F1+SPwrI7
mxf5eo4/3lIj0QPjOCv+SVz/OfgT8Wi4bF3fAbCWBBnW80fZVsbr6zAn8E/p8plEtIqftZVuVlLU
AdWZGqM81GWAgA/wdP/MG8uGZ1m4Z/LylL0s3PXlLmbZWNf3HB7heYsJwakyPQ/+hmZg4narRSzA
2/NynpHFrP38N74mDUhP6gz8PUUfmklKASzlYp/ZyD2xJnKTjTmDZfe3LPZDK+UGWqPhqV4o9AMM
3s0Zth1janG3OvfTooSVOwsFwxsFZS7lc/h70VR4sTp8bey8vSybp3U4a6LIgnoDI6HqTKJvx9S6
M1Q9ACfNqRsrbAozC377U1LI3NV/tyk5F8jgFAPo2o/ZjdKwyj1FEBl6+sdcT+cyIlK9wbWR0Kfv
YnceyuydOk+NQz8tJuhewcr7ysLSIhVdaYdijgzqMe8Vdse5aOHmbG1cDIZu2TjdUQxU9VlTTOYJ
ZO0QOrkDqnoRdQBdGsGiD/GVOt1hNNoCDPhCQl3U639Ec/0PxYznwVBCyZcOu2NMkyDuN371yxYb
/MrdAVh8B8bB+KvxcG/LjejvlqPALpBm1dvwlQGs3mTXOOnUhadg76LzxhcVrZVUvNZQ2ww4LwpK
EcvwR04g7WBgD6pBsUQM5bQZ0kgsuvzH/5B9pgp1w+YCmxywfe7tVkuhtdbIBYEodgrLznAJ8n3/
puUfToz7guBd/dW5v3+tT0w1ubY4n32RxMFeIMF2gMKSwhig9XibkTBy9DpnIlOkUXU7n1io00xh
9YcBH3B25PVf6WPLj3SebvPXHuca7A3XacIKv0g8ccGG1Qxb771jVeJtTu1aVKgAhdvKnvonTnoU
icDECpJZopPqt8+ZgnV6nbkQ5+9qSYEOtsXnlsMVDssaINDUP22hNsm9vGi4QXJ0jyA+m58V4nS6
9x6h/gmtMUJKS4FYC84LCgV5L4whnnB2bD84SZAD6+0E/b5BGYAeuUjJf9VlKtHOYl/4j2mcHfOF
KO/6X1KkPWDhO8dG08N8tRPonEBZbEWlNcXLr1NhU1cLIy3vV+nWdRPYwOpjEziwlgZc7V6T6vhS
mt1XXYfoQ3cuW9vsFpO06sD4LdhSBfJbg+iKjJyGXKgyCqzUWECLjfnxQcQbZFt1JxzAeLbdWjPL
J8SaKRbtqbsYjCl3rvKKi7discIcg5bDVN3WCNrQPde66GwfGxEJHE/qvdY8d/HfknLxWz+CNuLm
sNmENXbAPe0J+VNoM56ihanYrWU28db7eC/uglJqhcr8lqxeqHv2vvrI/62xOD6UYiZHshi/zCrp
4t5LphcxBccWCgxDzwd8pDKrGwqGbMjGpdKGlYkIThU52iDxCnrmvcRtDujy1iigBq6c8wZYv94g
vZX8Z1ZBf5DxkzOn9lH/FxUykhoZTjSUbuJDXbAAyjnoESkBrZExk07afOqH8AT/L/z1IJ7cjKp3
lF121NP+wX0sY4YjluSAD73fLaQYjd+njPszBJUuZny4VxJzIPMDGNJCMiZ0to8fUnDTVREg6IWY
9h3yiJHP3sFTt7Y8UVe3lWfV2g1+/ausG+315Ml5kGEMMclXigKCO4Ssf+jbfy3byym7wSSrtQNC
vQFj1FXQuD7f0UcbuNzNq/n2+qjC5U/vT6gQIMIcyVnsPjIypn2UGHsE15/mJFm95eNxcU/hzgvg
/gXAMsJEldG5Cu+mJ4UIV3vlsKKpJsxwavUPW9joDiZrX0G8D5ys6BmE8eS76yJUZam8ez4UliV7
9h/FtDB086yYynM1+QNdI9o53I+dDmfPA02y6cSX+V6EImT4Jqcfg70op1xlVSZHfR9f0oBleqpL
xl6anObo9i3iYKYIAiol6enKjiMqJYJGHV1+hpqOfmNGupJLD/Vt5h08l0iRzWZuh0/vRoPsvuEQ
uePwXBpk9FLCIvBWgzk52C8H73bNsG/qk7m8v/crRUPIClNKXGxNRHL0shrhrjdm+5iGAKqiYFPK
eN1dM/CwBKUt/4IdqWCFAltxo0DomkGLHVma7M9g+weGoc8qiOvL75NONNkxtD9drzTmJWnEsweW
nTTZRlvo42C0Z8kDefZyP/0wdRhYmRftxH7KzM2R/MV529uxS6a9M2iuqgNJm8kSf+PvKgHfnLqD
UJrFnS5Prg7HEoqqChcTevkMdM+uTrT8+Gua3C6OVtnqbUsPYdihHoDQpGxSNnAKMYmsdoe+DiPL
sXTZhRXIIJ5qPpVTsCLhvNnktgoeWJNMJosrjrnoghs9C/W5Xs5kUfoueNMKm1RrhWFj+I2p8AG1
s+ja+icQ7/3jsMJG8O4ulQWaFXPI7PiduOId+Z8vMj1em6DSxUijFDUEq5dVhMTqRomQMkzUPhpW
l9SZX3YCoKhfbVPWjC6+S+lu7Cx7+EPGCTwYP9KKKBDnQK4XcCoklkkxOsHtQFjeYlL/3baJ6Npb
xZPEjsr5jofEODKQmPd97MDKpdtCwQL3gcdD1QcG+q13uBMijZu93TrPw9zf7Ce/TeEai9RQCsiX
G5aARhI9TpE3MA3RTe0GJRByNKmkhHwmTWvvtQMZQE1rPztkXW6/xUl8VLko9TuLzIUpOsq6mpt6
rbxBUzk/ukiROcbN+IA4/eugYRSAjC4yWoUIP+eExTALfDlT6x/J1x5nQR8ub+7DEe284GGZ1o9q
o65s4vYB2oQUSDaMX9pgE2qzJEn+sZfInzoYtL7KU3cSVbveJI0ASvVZ5ffURmIu38kK/qGNtVkF
1qNJLuxXGQ9IzTbdHXnY+K4rJigL2afkzJXKwNnu3EXsSbyqs5rq1QJZQ7qf5rS8eMxo1m+BbjcA
woNudliTXFp/7moVWBhI2MUV2sKaOeHUQeK6FH4W4eiBVkmRZnt5PODw6LxVSAsvmkHQXWJlX7tO
iPSAuRUUSU+Uj52bSIJhSfmj2pcN44NgVrfwqQIXlWApLdpXuKMbnMoQoRIWcNZ8AXp/zp4ptKYH
DJ2uONfI+gYFzvm71zhUoWaSE7v4dlkJqb5/UGok9w8NEiSYjj773v63wvAjwOvEdJzj8ZtBsyke
UmINoALKY/VCUqHfLFyIFwIMvZIE+d5yPpuuUprwmwMM5ZhN6/XLoHNlrxbGRwmx8GtfOHNm6w1X
/sWpjKzBg/OJSfZkzfi/5+/Goap/bZj/ILOLfLH40cACPD0mqVRhX45ZXRqF1zLfO9wrtYakGjoI
7t1ewzC9yrR56G3hFNF2XX+b7gFoMhDMwdoBAIE+cocstX6bxKlVRII9PZiUnRsdhNM3o8HUVm2L
yvCQ2JA16qCJlHej+X5BL/lT2xqD0plKCyI4zPU+6i/fxOg/4GhttYEkRcVfEENvL9arrK+EBZwz
loMCKHwWi1zjvQj35/zsVCgdvuLhQ/i9o28Bu6ulvMGefhOhvt7rnteCQfTZZJYP7TpNCudwuJYA
Iw3mvqItWBhhu/Ve/V2vCWk4B2nJEb1UDsgShHk3PBC+CyMt83d+4NaF/hXa5v4EPPFt/kGXfTS6
ihKZj2cQ0cqr0miRVvdAjlhYdJ/RDXTte93r14fxpv+rBLzOLIkc3cl1KpcdLOvEdM/N3sYXrzjK
WW54bqhPgzT7lGdcjUR4sqHCQTNkknOks3/T2GK/ShtAHmZ5aZ2za0Zs05oJfwMKg7btC7Txz/HB
hFIb3OeJjLVuHnF13j8h5uaIPv6J3MpxnySjIIpCsBuR0OiLpVqhJjQ2QPeNUdD8PwvZB8uVDaEp
3VRuUcmyM6i1G9TtQdkleNoNlQijKfMY3cd7mylXN0p6qC0c0Ncdhr4oFsoCwPNelPu60rcA2Sbd
LTag+i1tm6UcZDYXVwJ7/ClR6sLjZXAqYfa3Qa6EVSXKVAuNiI8rP+nZJZteCi8MLvjLh/fFHeSg
F3g93ruiw2EacpDECeRnreD5oNS0MdmZ4WPiRAlpCp5KGoJ7CO+2csaSvrC+hPUyspZNi4alfjP0
ZcO9ASOSn2GPvemVNbsSoEDVseyjUBwXDcnVgPftW6c6oKB1EMth92dxfrVu0kGTLWuzqnfltrb/
owTPwWd8u0VZfl0j3gv9ix4IgBgxI/4BrbyW17hgGdnVePs1benZSFnKb1iPmqs4s2UcSmswsI7B
AhRcaJdLrErHWHF6RLdq5m7dN9D+4DcS6wkL45K7GEMoWt2BxkmvYY44xr0tk35UXpo5VoDLlef9
CxD/OEmhgp9AHCXxXWeZmQgiTxYqFdV/xJg8sOw9bcFnjGEeIJsHlLrA9WN50GPmC4/LVuU6kaXM
R0SwPQMIzt5Uu7ED2sN5vg8G56cWLREYJpj9Rd4kD1YzSM/WLPSNiSVH3nrfzTw30FGrdYARPuU8
w4dK+NlnM/bv+nUZYrLqpQYcS5BGeiHr4CXo0RpxNsTSeGhqP9OTL4oRaY6X05sfwRuR4aqVRT51
1IKGNTHoUhvdxU8pvi9jla2d/TsvZTVxuxPrL8Vv1kS/O4/qcY0rrvb77irZxWEYsVLQdYXdlzt8
8aPW+RDHXnRsEOx2YSzOS7XQzEs5Ce5WGWSZuxfpH9L3vMtueTGKOidIPWj6e7mc8mTvrgcx8h+T
yt7tjtspGWpehN/VKNNl27a4l5NWvOZHY9Ay8sEqawxnHpEOUpjbgfxT2r1QVUz2Qklbvo4E2hbQ
+6NwOOW4TllB5aXC/RHuM8DR8z5EXfw6wSNzsBJYTsrwA4qcKo3sVnfUkhHct5hnJ+1H06lT+Rmh
JCyX+69emujvPhtjF78lLP5CL+qqo/8I8k7Hdvg5kfaQoL+jfKXUb6k2uwcPMkcl/29nnOWsrOrQ
NJyyffNoxE+jdaPh46UTWqvDBjchvTnvIOcI7cfZJgZMmkpy9juh/2MZ6073zWFeyTxg6z+9LTXR
xadANg6tGiYA5uyENYx4BPtpVGWAhKQ7o90+gQZzwIpZ3Mw3s7yvcueiFZvzP7pFanlRjdZjjBZN
47MAzK0vgmqzrVi4pihcPns7zOcAUObXwF2V68Nrg3Z2TZhtW4Hocg8Ku09ZVx+jZ3mwkdXE8Bwz
WV2+g4DUoq/TaqZOigxypmU9pygDcO4n27bIHWROC6Ad+yLOIM2qIuRX/Q81EO3RdlcaUrjtEQXD
1gsBtCjY0Wi6ksBUy/RUNGybxCPGw+VmEBRkZ0E+G/kQhIo3WYwk3yNYHAoKFk01K2/6RHrJJeWF
2RsibC8pFitE3afixJrNlyE0V3RPrTjUidb2DmPBD1X3OMTtpFjTu6kwoiEQ3TtcBKsYodURyE1c
xfnUsZo+/4sesgdbyV6mn62yKpGCEFxXwbvf+55JquU8lJUbCzGH1d5eLqObSJywNGWnx7Y6q6X2
NO77ATwZ9BIX/eHC82772l6NgrXiqodJ6xKlMWluIw87i51u1gYYI36vrVVgAbK/02a+yb0GhXEi
v5PKaZFqG2cv97FmkAMg0c+o/yTYv344NVGDTqf5YPh0g0sHyGmYlz05tAn6cFTbD0SCSqZj8ax0
x/1jbJf8CuT4RF7VEayszG6fILwO4NSYn35DlS5pbvMicVXMPSu8awnRvbWkHyI7sdrVnHP9n1sS
IMxQzMKYS0BIH8Upsq81fnColK4DXzMsTtx4zerPIgqCasLXSe+eaDLxnBm58C8WRF4rDWUF3HwA
wKZhNbGey2G3MDG+xadu+k+Chp5EAA3ubojiTifBGcpyfyoqy6QJDwpQP5q001Frk6xJRdzdobZV
O9pK+i5qbF4zcm4vWhNeRwk82FvV7kUwTwoUWLXfRE59kso3NTEtdtlLpJ+FmRAD5QvHLDOgdHj0
NgCMyyRLY4IrNpJqWtGeBKqVGKN1oyYiObNlcZFZaTiyxQxD1YVZSAbc4/VzltCKSDwjIxoOMdwJ
bOiKqe89w+PICTJ/wBf+HPTIdtakzTJh/o8ZkJZVfGwB10Nf7bYGTIUqzIYLCc86AfKogPGeJSS8
fCvmYXGqVr5A4vcuZcRn5QauirA8Pq8e9VLA4b3vP5ogncIttsIM4CbQEK2+LRn14EAGn0zIxByb
V8SPlqMz9wrd61SN3DCFbDfPKj/aHF3GTbpn7NkISlAw1gIW9UP7ZpSI6VywrD8gJFfzs8laL0FY
hNsyuyg4Ad6VL6XiIMYNEiPQ509swDdaYTInUbmeB6eWEbyU3cg+9btNZW4jSmClJtxhN+PsL94S
YTzxfKQ90rPihu7rFAYQ74sOkA+eujLJoqr7Z8GRBeYIcuhXl06NWvneM1ClGRqiXJuO4qaVSEIP
7rv8CJQmy1ZFdtjPpPpQMcVlaFG7JOzR+5VWMzn/4IDeWiB/3vAR++E0q4PK/2/HWD8R8folSpKi
N6hhM0kjB0hIZqoVhT2TGArITdoVesRqx2D0bXfAOQ9LJnYk7edG1hx0GRjbXr8hxF3tmmlqlzjJ
QRYS5RhVc75tTz1LthtIoaHpKR1G39SuaStclYfERvo7Y6pd36jFzAcoSlw9rn+n0eVBXw5yxEnh
Jyx3I8TO2xN9EKX3q83n8c5UW0Jlfop3+aYwQS+v418TuUmhVbq20v7lnmxB4XTHIearM73XuXF0
ycaLxkJDgxJr0/rKUP4oHY51vtCBgYEBeloDGlEYZlGDGZKg0LHzNkojhRTnYhznAsowdJITtoae
1mv3d+oaF3LGbnp/cDYsSwkS1INdMEdfunahT+iYSFMtcRi/cH+AkITVrN+OFvz92bIt+kTGEg6a
FiJ5XrTRXDi6jQDvxPF/xnUTc4YIpLUeuLI6GUj/qwCVbb1Sq2zz1sWzVCZ6/DrOX2pUMwuCr09B
PCEiE8gF/kFqwvbaP3HPA1vO7Y0EsVR0+mLZy+XhjyfTcwO/6Y+jFTqAu/LOJmkiaqdhTpJjyOqP
ff7C+/m7B06CB1+OZqgUUdlyN/E5D3lDSvPHAbxe7j3Rhqql1aesWI5Xyo+ISE2Td2FK32HTrKDM
j6iHZIRe7AcU0u0oazm/wzVD3ecS70rPA901yIX6tVtIr10a3LblOVkuNR4FXvwyt+WzY6VSe7lM
nZe/7Fb8eSX2ZHL/gh5JIqzD483h4Tq3rblnpHn1GSQaENwzjCWlD7QOfrk97dYw4rIjMEfZ5/zs
8jbNQI4JmyFjPShZu1/ZXnFK04zYr2OcJtMto5UP91bnOyIjJPE5inqWe0jzJ/SFFU6q778vqYdc
aXcu6SYng8vju3iB8uZtFXoEo4M/uTqd780UHmlzYY48WrErBbNVYmUfr3cEEmhs0yIwjwdlz6so
sQRy/UpJU8Lo9hzQOdKJG4VdrNo2xlt70+rse0PA3Oo8Og1jRr1/8yZdb1tv9T6QEIb+9M6TyUcr
e7BLw1ZER/ZV8SpBJq6OMJzRuV4Id2Roe9igjKKIGjKSPbaxs5zJxR7yQZW7ptjxtDUqmbpWUy88
jg34iwoO2GSZvUywuwOeGqOye5PjuVKMzmOVfx+GdO/s+1hWCdR6PilPDVrB6eFCGBapCvKnV4P0
nst/YNy7Mbptk8ZsDPW9AZRg+HiCeLaTXJTCA8SOK6ooHMEmlxUW0luaQlBAWZF6FWTjjIDN7UGG
8LVN2Y9lfFBT3pZanak+87OoiHcfOFX069EOY2wNIgivbXY+z83/W26qNFI932u778AZir8mSsuf
cQcXtBlp0zBXzpL6YHAYnuI40anrS1Txz6O1uMgdVKcPNc6shbDRmb9oZHnBZPYObIfeUMaizRcs
KHZuCCFUbh6cTXEX26tIuWzc+UICqUEKJ4jD5PRx0MFumf+d56mHMjGPztdhStVWIrkUuL20gNF8
u0OycL2EoTqFptk6UljHrz3YLaQAmVPxauCSvr4gUdCdxwlXbFk4A6e5S/60PCaJYTmySA+M+bU6
uw1LcJ4wPftM1iB83pMt50dqT6xgzXGUvynMXctnjUfukIvlZB7465CfDP9v5FejuL3Tz8nP9/UJ
X/gTEIm/6CcQlLFlrTm3dXree+zqzIixL2WUa6y6/2N2y3yPMoOxUIUWUFr/a3jtxQzUCDTGd36t
/qGe9f0ij9+sIYvGVhptAIAtlLy7GVDCU23Yhg/ruRNKPGWukOcOtBprd1lXmbc4z/WzD6SjmP/4
YASzghxsGRQ7+WcZkBuC9Wqa+WVkTMupuCThRpiabmqFe/jSv/RzcSU/MIXoKXX778ePbl9a06KA
OiP9mv9//qom2QZKM/50a0RqXHaYGr/WaDo7y6cyhXsskf7riDvkBZFiaJQqpoJ4fPnKwMGP829U
SVHEyxK0WIiM4hylU+J/ReE+UCO1CmY+nHv1KtWI5t/OqejL109zJgWosDOKCG1D5rAIQJgCYQEq
hX7ROidX/Egf0t4HDMJtOfi6cZVNMWaXdbK6eRD1xSZN+Cbfbm+CBMEAhTJT6i+wRfeu1JC72vYd
IvL2PRkWkrOAygW26ZyQn1BqILqbtnJ0VM1BX7V9uU2k/qEVvAXNjhpkyLpg8eW9It8n+/UtEtMy
kMo89BtObrBKcJUyutRCWuLr1k3kuvCa5sKtMt9CZjwT2tKiyoKqUfSvL/EuWz62MZwBkJFlEgFm
5IeZiAcvx+PLq0PT5ZM+I5oObMmWT8gCOMySRFOkW/7gD8cYjEooFUbfPQ2nOj2+s3X7HR3yqRZ7
LQBcjB41vHDk0xsjOAv954LgQL115wcqGLQJUe/oPF/nsNlxecdu0RGydVberUnLkkr7CIUG9HAu
DbxIkIOBmYHjg4jVTVMD0EAk1o9lNO1kEHM4iL4vOzF1hHNJvd2U9yyoAIJCPhcfa51xxIqU0/mQ
KKRSTt0Mc1nqTYBHs2Ws2ljSs/QEorHTjxTpYtnmSpWR42vsprUvxpvS7aAseVFtgLXRmd18y3qP
dIiNC0RQSccvumuBZEWpYr+LSN6pduwMJiLLsC+IPwPpfhfc3lArU29tvESnvDJpP8ky826Zbedl
PM+yAlWR5SdQS7mm0+kbBhk2KBJGZIjep+PQ11G/RaXltCwmhCJpxYLD1BJThJtNX0Hhd2VzlH7a
UlwhDzUQJKIdILwi3AmZ7FeotJlsr7GzpwE422y7oab0GvFvG65zVoUAN9iGErxoKbXA/T5h8ou2
8sjJtN3YDptAuT134gGDngdDSTIjYImwNrHKwVbhPYtkHiEYALaAo2zKgwO85EgcmDiYe9nYP/SF
9NN9RKEVL0PJyBYBEX80cy7YtEHzH0IiqPFnBUukeHLOlDKpTTbCB7UwjUipJ+Mhc0y/fKTYlweA
6Ziz+GfloQfbEyj02dezCvCbT0zxLOi8blErCkSzfdD8Rilscn7R5YsOaQQaPSPWKfPQXcIVNyE4
NxU+bUGeLGoWkHG1EtdnU4EwiMtd8MUa6zibZfAgaHfKv0yNZrQpER0Bc79MeQtxzteUfoMMTyUI
r/TpureRGGbKoH9d9FpTUipF+lhQHd2UWHA3sAtEsBAmo+ORNzC0Fz1rsQCjXndoiSXAnxvKmCLK
KQIUQS3bfwnaRO+f38qv2HCCdAhWh8pSSNi1q7613ekRfDwyfeU+4s8SoSynPWoBTKJdaKHWFsRR
+XiLVUPI3C1kxzzbE17AdLx8SE2uWmSuRSAWwcUB3kilfjkYknIAkEGhBaBHRq8CQ7KFjoniQw5s
3I6m8d1zNudg3Q7Y2l1q7Y6FpUUaUUx3YrIhmhiPFqGhL2uROy5aJWv9hWv7JxXT0i71m8udvU7c
gvoWA8Pb0e/leS3vi856UbubI2k9Cm/VHmeNcA2/VtViH+6yDfsZM1R03P3dLqKZDEVXy7f5PGvf
s6K6J0Umzyn8EJcFCp9fd3k9LJX8fLQfLWiCX9FRlZnwo5SiBdxYbta6FpLdaRfHGPsX0kWV8SC4
4Qu482oX7InUM9SzpKvw4FeYswuKz8m9//Bu7rgvYtUxwkwWrnRuvVONP967+p1F62TEqdwawIs6
hyUtdkj3PFIQtdvdz2SFGbpJNd4gk+QUlo7Bv1HSIps59R6d479Y+JW5H+u4PjmALHY0axC5xanZ
1uBLhRQ3s8FNx9gbWQx6dWILDnnsiGfXb1mT6pIihHPlL/tymaxeX1U0Y7Ax/2vDugK5WaXkzHOO
yHEZH+lm419xnl2GC2DFpU9DbvN3KpREzU+K0oDsjhTYcHizFsD//cSX5IcDWasPcQGwnovBgB6S
0IKVRtGnKK29Y0bQFYks8kxEa2A/EqY26+cFHQQh2qv20jXjqggU6cTzc47u1zY6OiIMjJ4sneVv
a8IAYBwiuQ3KnyJC7vPUk1trroMvNf5UJhJpnlxCn6B+dfdKB7k0rZZQCfnH/32kPAUBY6HW2mOY
s/rqBTC5+9nilv2Ln9fZvJ/Xow9OlHZJTvdGc3TEc1C9lIurpL/lXiJlCsy8qGMe/ugkErw8kgnc
OdcpVXtP4kFMZfaMt/Db5t83TzJ7Xx3sO86+xpNsZAYHp3NSzVLMxcflMFZowu0hCRrs/0mwjvIV
Je1lDIWbD2Y9b/4fxPXZnck1INGwKknGPg4mhjvBlnzXhQVlCqj351cfwE9/PGdW8uaqH23mJ/72
WkdEK2+S1yZwfBbR/9fhm8o50ZA02YoUnO87vnqMOPjubAcQnACU2ivx6YMANhpEvjWPgaMFzItF
GDXJViNtHOFq+Gj/2KAf7BmPpkuC0UAqul9i301ZTgifms/4lheAfXnpsPAhlvYStj1qz8DJsb8s
IU4vQUe2CnZ0KVYv/brrOySwGSax5/4+KwEu+ranP+eoVlg8DN6LGhO2YVLzSX3ckeMJU/bl342u
eWjbCpROYrkvz1KAb2ylxCZwNhHp6YX9vh6PdadWLXNX1Oy9kBaRmdIvoJVxlqjiYoDoYLERTYXu
bsSg2+IlBvcYWblOkZyn9HvFf9ZuIolgEgcAtEj8gUSQ24wQAntIGs7gbskdM3TmfyQhr0Eag1sc
6XP1EijCdQeUo5GPgDm4rGDDgT9RBosvgiH09AamUqF+LglQ2KUUm7neVUh0E+tO/G1ujYmmqB1Z
nHM1Y+9w3cspMfF9AbR0q+eSc4WITFfmvKjcmc+vnvDsme/MKEyoNzRkoE+LtwhklJoEzjMO7GV1
fLtbMLLOhKz6AseLB2IrJZi6VMfMDLWil2hhkWL9ICLNY0+ZmO3bFPUMaQ3O26Jd15by1YgEjNuX
y7ZtTGTSKenoI7wgNAPpF86ro03xRvjNm3UJlH7yGeGeXVe033IDSRGO1Mr+4knSAOcVZvikL2H/
shNX3NKo/L5VzPTZATIQ89cIZyVvOhPW+JmupZc9cMKRzPKfkMqYhYXlXzljaYRjvm4FKAJyaOFF
OQuBgi2m6LMipsv6E8z6P8n8oUJCrUprkjEUMxogr/ca+qKeF+0emcdJd19iWOZt64qC+EBysYvg
M3BF5s9n9kYVVnAquOCX6GfQ9pogNzFDIsKo/1Eo0FBXA62ZuoQjTMMGnOBiY729vuM2DGucmsfq
HoYNkypg68xkeg8YTHdq9ru14Hzldq3dK+Se+wnMGpIAdwaR/Xg7YGTsf9fgcv+eUBezcqjVm5yU
6JZ9+GricPCnvBMWum1xxyBi/Ck8THx3Lm3e5QEewdsCeaDLAft5kv76YpfTEJTsjfahXVQlfJuX
8GJheIDchLMGLWewfsrobFnYoQ/0v+et8n2p36WhSnOqDQ7uCSHxnvwOAN1I1Jd8buNQEn40M1js
YDPAzz9LL+2V5EDVo1yfpx45ncyx6AHmNg9GEpPtepQ0VvsDZO0wscFtblZxrrvmVufU5w1y7Jxf
SYlQL/1jEDQsdfg/5550eMWZbX7tiRA7t3dxq23axF2TY4Tv8Km8vdjECOSmmTqq9FiL/F2L3Qcx
8gIApskZCnMRShCtsD7dwkETBYGHBSrL/j1hVvdhkoIlOuA5GdVqxRZViOrCScuOQm5cBvYP8Dz7
/tu7R+nWf2U8reZTCUI9bvbaTyku+nmXNiakbM5QxiLToAxAgsW1vsVxcMoxyMQWZpFVyRyjVN26
JgEDoirqBCrw6GbuQBZCVoJA8HCce1xtpPLnmBFP+MVqm1p+DwQfwKqRiVen5dRxS57g68GU5NjS
Uc1yAEtUTh9tR0OnzBgx6HNaEiW7gE0OKZmbmsojPnzyKh7BBXO/zOEyrkognfF+4PfCDLCCVXut
JwHFgnT8drOHHmZ4TXWn3EhhNsCVlHSF0ks+M+qvm6Hz2Qq3lZxBe4xSfBPGR+qBizEYuJl75CQW
vrJTuQMIpsvxFOyPfidPrEjvTY8iagVPNVZR6fMU4YMCTKzPdnVfApyTvuhrvscY42xAIB2f4662
rko/uyL6Cqte+QLhyUxQ6nsCu4THqCF7GTUA8QlmmWfEZ3QEEc45/1gzU5uQiBrCHjbUPgJRskuv
X8ISXppqLoOKjk6jFKsHmRj1SffoHk9qpSf225ho1pNa6S8O8MhbXnPIuydmJS3U+NnzHSATwIX/
NopnFn8wuvGT78OCvjnef79dabzH5zrFnlWG4Pp3b3cew++hVFNN+GZ4E8ogU8nLMmwogMV0FUUr
ozflpkekpevCoob/r+AFtaU/qlpgVApvhNfrTzvin6iFnoVlDQlctDdNguYBynPjFOjw4iOPEOz4
BGNhneSVwzEOS77RSmTq5cGTDAJNAn02O32nxjXH/lkHzJRQy5ZETWFONIvdfdJxox15R/t7eswo
bEWS1WQ1NWBQClQdh+pTHHw+J26yVokaZG1dwnc6scWsnmCzH43Af1KUCwsIASirv+i5claXNbuk
FcVXUI5osL6J7VpKUfBycBvK4BOf6oeHhcm5S/N2kt31NNHg3gHjdfm6BUQXfqQxiCccVMYECQ6C
/TTVHM62ZL5FqXO/6Paf6qHEH/JzRwJTCDwadu7Nzl1PS9wC4CyxiH7y9PYiOfe/uD5NDwEcl8/u
u3ciTCpUTvmxjJsnKufdiivn4qE2C25EPmYaHROcs0xNuwfpr5wwEIgIiKyYVbouRqxJXkfP+pnn
4Q1KlXcd8LccUtQjrcCnwT6wnT/hXP7BJ28TcQ3V3F8sR9/+Rdp4yd2E0dr/SzKeQQEBGgpDqbWx
v/KwP2a8/kMH3sloTUvLaYPqq0r1p8CS8XuLEpxB6kXoX49Iz2Fb0ff/ANYVG0MIwo27atqwOalR
cHZOFkDMLxjFXgnv7Ik22CcjZ/7nHucJreJGzBYAKS12jMjFTE3uJi5tznYd3M5FH7cKivMX/5mx
7XL+3RNLgK6OeOiolNRMs5x+SLCf9CS2V8ikMSy1OolzwYnGi85ii3VwjJwcKO5Z4du2S+JQTYYk
TbnuuU8IAavQdEdxHIfS7lb8Ac3wL5bchMdpBE/DYJ7on1LZ0j50wk0LvuzeyfxByiaEYU1lgz5y
KbDvXMVv5ccrmsMKuPJq+gK9zP6qwKKSOQ9nwr1N0yISNSOkCkQ7oqepWcAFiGHohx3D1EmMwcO9
HyuQjyxhjnpBNto3/hj4vUkAruZKdaIw9VzwY0OwyYOGY6fp4A3+pIdjzAH/osvIFZizh5K43D5h
UBH/80cSlPZs7M0B66C9nmLpt5jBNM49OmwgwYONY9HSMJsJ8MXnX4Q7EOYidHT+OoDL4WyRPecQ
4m5CfbuZWnmtA/EGos9bRGxLO9sLxyXXe56/QTeeHB42KvItXYvtgKxyo4cZ1Og5+BwsIB+6g+6H
SRGjsDOrY88/ZLfruef/BbHdXM3OEd02EmwUO16CqbqRS5xf17KkIecMzJY9Bmm7wMnm96O0VLDp
dHGT+UpgQnJIpSGyR5npRC9x00Kkfl+yUgkWXZMcSFB7/vBp3n/XRUMg9y/e618i10hrbFSU4nBN
Vs6tmZjKKLbSniRJML4zCR57q5fglrQRKBmUrIbz5fFkwmDMcJrMQ4IarTEHsI8WBFtY1YXWI9Si
fBzCGk+LLgOm8/b6UWtMxXURnTf1lwYxbpKCuqzj5quPWTafxGqOqqZKgsDBm6Ww4WpXJiW5KpjX
+RztMCejCdH6l5HivsGrw+N7szrC0UmFmYXtYzbQb4HEM+BYAJjLAUFOwupo9TDuV21hF0kS1BGg
ivml2h9fCdWTfRi4GZMS95Evw8Z4laQRS/7MXNSLP22qMf7hYol6g4XDNTg6Vd/fdcZ33+wNqt7F
CXjFl7vaDsyv8piDsWbvZR/bf8VCWZ/9MiM7TAAY1/dh03SwWhNwYdlhtPNkDO/Vr+hFYu2S3LTL
8l1oWMCqovY261s+9WoAJP2vm87HLbphadaUI/Vtf4lc7hM3eOO0Tba0+DqiDupBtho1GRCRTD2I
25Q6hJvIUW2H1lKnjckQByGSrTfSSb1Z3xx6gdQxOC61ZFANHBY6ILAExesaoztbHGFWTZUHBd8K
rwDayxaoM8eAECoKITnKkXlaKtDwFZdaa2sJwqew30AJDtw6f+frQRNBvlXhLYMF/9NzTccPT9UW
0XwvfVLXnhgGcmcjdhArj5ijIToSnC5s58UDuC+olMDhgo3s0hoSH0wCdEgxAAqUYWuh+Gblryso
V1enSrpDnPoBHmMbTWyniyMl6TVQWy/K8z3Nxufi4mtRdRveMVk6Q+TPwf29rTlLtVErDdx+ft0N
IPq7u2b9fq6BGEvEKocZtZ/BhAb4urONBSy2SG+JJUAm++TxnB12n9ypio1aK0+EUjP9PsykThNw
mdGogn2qSB8gkDXlFSuUadXK1aAyOOaniUdaYF2gi0XMV/tCOSHsZoy5VaDZKF7IsiGFCMEziiAQ
wKuYEaorqbuxziMkTePCteXgYhcgmvzDbIZ6E4uorgZciD8PUwEs2D1gVPG2/D1pR4vqCpk4+vkW
0SsibMvD3nKDyV8+6gLkB3eqadyVjkZoUeh589d0if7y0ExqE+6zKSICDGyvAI8tnncMUN+iJzof
w5ctYAelwDInTMZNVVQXYNHKATW7ik+9ciwRrDFse+u54If/mtw0MLB58c8RIMP3L2fm5wcRGJ8r
XNQ9R9iYXUlN2qVcyPOu0WvcUP01Ugxs3WMkZLENC1cr3yPO4svBzeURnrGKXZDetKBk4ALVLRCw
HIK3e+FKOtYBiGn5QZCZahzGQe2o55qguOnab2ye8v4nFFx16gNwjvs61eQIadEjTgOk8gpkiemQ
gTzHD4ZeyGVPP1iOKY//GO8At4NK5dR64kn2naqYng0v2aXJSGlzLJA/LtbFWo2XWwBrQw/5HPzh
GkXEWTvCRb5DWPymOzCKv7kzWOmIoI3d6L3oZPbNl+klwmWWh4dPdMUZQ4gIzpsEg1ygWkg7Xq61
0s5oOJIHswIJYMlYtXqIDTXwIqvwn4mg3doxaURWkzNWZFSbGVpUSfVsuwff3xz3u3OCuRS8KsDV
5JpoYnE0kWv+PxUJsfn/12PAXSGdXCkkQQIAB7Uk2yrK0KGmdGU7TlyMB/XXbfj/pf3IkuMmBT8b
khnn9qLxWMlRwvnwR8U31gvPAdVFgSoHwPHHACMO/Z4SsjWDtGDnx6Jx0CHtYmpkb7mrt8JVXUi6
EgYoOURyNj8zFfK5dijJKN8izaliCuVnDNd7C3kUT3/2dbEtu7e9SLQjy2RPR38KWHPyQUkJCo+Q
vAPV8gwKJPec9lAfSvjeEq0dKaZl59wDE+7NzAhnNaVcfqWNadW5j7yVO6y7tmjGTezzHicGqIur
Kg1ADYO7P8fGHHkTz9dQj3587KvQ8a85TMje4F1LOQnljEfku7IJMdOnyCWRFH00z6Kv/Z/3YW/e
ultjGNb5/yKYdOslONpaWIwfzjwDpsCS4MDGUO3CDb+97NIdUmZrUucIuqPw8BNWqokjEDSG7atj
ic5osvGuuxL6Mf+RKiojZ/BnOzLr8BTzdwySiECeiM4EfZ3COIMWyEEG2rEdE6iCCjJdkDwgMdqZ
bFnvlUSgCx9SKAZAMRTyGvw2Z9OosL6qQcDweJfNJQIygfGEkyRBJo4IvTarA3Me+uSTRrwy+UiN
FEx785CH0oAKdVnq/H/6XYpBxt9wer7EBLaWra/1NcHp4tjIg4d4pdUZNBf8e6Lfg6k4xe/yF4zm
3h+2JvBh7vldJIylSFmao4GthF/PdbrpAECTHl8xpBQopkFlgZIE6cbRxjcy80tG6sO+E5mFMr2h
RWgkhAcPS2P4y+XYjob8lHcVxoLPY7LIjmlT4JrWVKhbm0ACzs+QKiAz8C0doCDVEsJgNx2nLjYZ
lCj21JI+gup9pqzrmYnHmJsb4JIyMGN3BGo74izsWLF905Rbw61rDtu6cVD9uULn0EhEknICCXVm
kqkxlsed26OT/bHA7FlahS+TmdfwdiYKIOL1sYJXpVnJeTzFfoPQCuTH397aV0FkGaK8WPJZiB89
qZwWVPUk+RBiraLsRW8FePCgpgJlahmk1xMABRJpglMdF2Ug21oczFKVncwlrUkfzX9UV4O9SawS
HuBfVRSFQToS769BwanIKX27fbHruYy7G1Toc1+Dl/hTh6OaYQ6iLA/tX0FS1TCevDY/sg5cmiN+
4LRReAiD2MIpYcq9fRGUd2/KHrOklwC1v96vTT/h4V5sz4Z8VjwdWC4vpmk1geCIE1HFH0Jx7U+s
Bb8NOyvNxQOVK787bbEA2Ol4kwjank0FKQg8ruGCfJbuZ93ITwjJFKAEH0iVhSpgdLW/uygvqFfl
6rAkfUmacw3+6DE3B4l9ChO+/t4v5QcdVNPMPIrgJ4pJ4zIkjsFrqYKGis2Ez7DrB76idZgTjeIc
Y/WrpvKkXXli87x+vVxjkpmezPpU25nkk/XzWJsnE4NrlthmRphs/qa1POnEr8lM9XufJIrYBBfI
5Hntr6+b/P0d+iLseTTb1TYGOjnd9F2pVpdaF9xuyoXTtMfG30T0MQsxDPthEdKocM5GX7Gxm1iR
z5IyUu2SPiuhtrmnXpdpaOjAdfQs/2omSKK7Cq+fzCOg6y21W4HCqjb0Qx+NoK5Ttm93rJjDWsM0
+CHtgKVXu1B2aUIdwdG9garw3Sf610vVusZ8AamAY2ppPT/9EH0Ctl9kxMm11B4xhU/9dhX2i0WR
M1cl316NzWPEZQF0ZdONL8MAWYfxWY9jFhNAx7leU0ALi+APZG1uc99/zXqvisu97nPeagOJZoet
nh7Qjzlqoh1u78J8hivG3noH6hHWXY9DVaixbOBlX/7GHh3MJ9mqkdBJgqvSIlE5wjORsTLPXGU6
QRM9gjQVwT+156fh9Xh1QP9JD3ZzLvvAEzD0w++vWSaIm8eOnJ55b/PSf02sMjtAFFW/4oYBzJo6
T4bJTO6pqS7cwsYZIs8JG4VP4OctEm16GD+a37+VSlfvsh1D0F1WQbBW9HFsN1sQDdFz/FdowW5Y
JBE1URGBUlgF1y8QWX0debVESUwQWEeeqsa0f9AsEsmNqM4hoNu+QH+eDPClUYnFG/b7kHSJ8IxS
ifj46VEXbfxiDImjE3EQ27FKQU6sufpjhRSPW8Gm/aEVDMcZ6ailCMMXDm3vm1291x+UYT1OAyVH
qjsnLTzUzisHKQJLIQHp96066dXlFdanv4eQZnzPj58mRx8XUevnzZclETuAKIY9f27aplKbnZkY
uyDCcBXQnO/1EoGa8a0pzgprwE6DYap2JANpeGLI/ncNddkmEkK7bVhbkKOsDqhrr1bWj5kgi5HO
YE9M2yFhil8CKjYGPCtH2rkP0NWK/iAB1vQEP3tdP/i6ZGyCgIvmeVxXJKo4BBt6IJtj30IB9jw9
YNLVm3+SCYWCatwrF+//A5gtLPerNJhCoDNkew+ebR8gaCbgpAHpoa340+vjTnuOGVQfwq8guHlg
41emdJjEUO2N0YvdpWX6nYLUwOsjpBkm+yLx/fIOwHW6qSHyxlvXMQV61bqQFzPzGvAFrdsH8d3k
W1DsPLqBNooZrgFrY7KWgt72X8XYOtLnCanrut/weX9GGck46mjMz0D0Nz1SC49c7u3uhM0SxSXs
Xrw0qcyTwbnaUI/JvdiP5AdFWMeE2ZqP9CpMhMIcrLLtCRRUfR9rYFRpXPF4YAQ+uHLaBdvJmhm3
4v/npCkWz3O8RIXqInAz0onqF7l2rt8EQyidXgQNU9DcV0glJvcLI/2XJdHlW8YjXj9yF2UsqRFH
0F2UEtfvJqUDLXB8V7OZk40+5gyWQVvJInpUcIuuO+4oCIoDiykwMHoRhbFRexVrcePKFF558Lr/
fnl/KMQfXFMncJ/pJCkLeXc04gQm7JBu+yiCcw+mZkoZr8AMbt8TuvL6QdyqzOfPiimgvCYcSqz7
7k9AtBIkh9+/FEVORL4g6NfhedyTAgLn0lc/Hf2GobktMO+yxI5yuYPm502Uqt320/fd0yzbte19
abOvNF1Pec8NSPnLzOEaz7rM5hzsVYfQUOStyXNdB4hBKFPRlujvpZNPfRMRaHveaTLybW5jPFSd
zftQvM2kk0k9loBamz1hI2ZWUc36aJRXD6OSqg2zPIQfxRrUiawoD565M04+KnCbXl+iWJEaSecr
KveQ6vQ4cadlEZH+iZTDKyK6VBmHwgH7od8/wvs/Y7L57kAW9wkRinjQVFGrso2SKG31FnDYm+Mh
7kx8FNEmkQCkjMibFwCWfoZd7DMuYivOF+cabgEYoBk5qLEqUAwVGEL4ipqBKj7R5j/UiO3V+UR/
+BOg6yJTteEUh/qu5WS/EEGb5i9hSmwtTCWJ943peKBVuHGm4ZwRZDZOD5E2rOFdna48YQz0Udje
JHAQWXsXjchXF7grOWLjkVdQoEeR/Tpvj2wEYYNDsvqnReW02qo/03JxLui0az1USisCymtxX3T6
uCP7s9UteM6BfX3TfJ3SWcq3LfUok5KGgDj0K3iQL89iVR1CsqTpJ2/8fni3bmQjnCJWPVNYz1/F
6Bbre7FzE35koFZ44LuHFMVVz7Tf9hfrE0QeC7cTQvrzMsaGG4xt0ojG0cL8WdBuIupIXCJWYFAs
+lzkJGtQep/dU5orPxn/qcX7bJ+814AMGU5Czv2Z6xK1EhmMJuqkyHgq40yvs9nPZxrTQTVSC7e6
tW7MryVi2uBKCPMKU4K0uln3bjfbXWexnrPk847fKxxInbT3aDpkS4Ztv1oA1Fjaq/vVGzeT/xPI
ZUSjw2mq3JQGqTfoJaq12s1jOENlD6M0O54rMSSF1JXgjTC78iI10Vtf3ehMkuf2i/VQ9Q3Frje/
UDf6TVOifCDYmsAbXw+SAK476oXa9YK5Kz8bWqqU7gQzL/8UIBMbeoMNCCkX3vX3CsCCuOMB91nY
5deJvk1Gb/xkDO8J8+0B1cQkTncN2uYV6rSuk8U7ro0h9UceX38RxTJGG8t2WrJWJRBSJd+yxruY
zwTxNd3bK8Z7S/IX9VcR+dEoUja8Ln/nKyWZFpBEasdkgojUI/Pht56wXMvcp4S/pmDI3MH2wGc3
HxgvOtetagGIbRhip6gW7ftT0I/Bb6d104WX5vRiH64B13JywX8LELZaiS+Q2g0BYtT4rJ2NGmYc
v9hFzvv5qnIr7u1yK2rTr3gtjTjsgmzYGsQqqrVZbmf0zfliNLUPgNHdE1pNE5ykUMmc3N6WX3Wy
H20TNNpTzqjumuCxjWr6RS4HRDBlbPCZ6uZk8KG+XilozV8kwMtONAitDAkNfQYpenudQMX6WMux
Ia1Yakz33zm6UqZyUBmci1eGdRUI5LvcrkG0IdCcDQNq0ncLoQQubpnBjypjzIXh5SBj8N3AAUXt
G7iSEZ4z4ilqPjZPq3PE0ywwQGXKXxb5cefaei8sb9zdtccVJ6jYSfscnUYt2RuKVqmZRAq/J+Fd
G/aLRz9OQhguCG3SopO5nV0dC5pKE39qKfWvig8VSr/mzstqCyaHpvVHxEr4jupVg6/tONCd3NPg
ma/kP9ExhNkfhLjqu2HPd5s0Ou4FAGzPfmLXMaaqxE3xUtN5lmJH/uYMvelZNTwkO6y5Yai4UY3K
pRCvdWOj7z88zVfUrN9TK78zohWcG/s+zZiioH1fk0l92TTKtp7FQVujgBru2GUnraE41Wz5GjxX
inbWmc7BSzV4IQkr2cUfIXIXNxmYrvw429QDjM4EsbntjIqM7IpzLdTQWJ+OAEamgG+5PuPncDrf
uHqvM/W6USxajzu1BqBJmXRnvEHdMOcpcTjQcTPoKpObq9lN1//QPojvmVGHyMTIZRSifcyeT+jh
JHWNMY9ds8SKUMxxNCfPPp3TMGCI+NMb5F7i8wppXZgYs+HscLusLph3bnhTg1RE0Zb+Y3KJ0e5o
H81YPaCg/3qyzrgFiiypLgM70eaCoBBb9hsgyt7sJ4XaelfPrp0BG2/Wzl10aqFUl1vmAohmqQMM
a3QeNeX2kgkFHWq7sbWfs4n3805qTcWAmVcEA7H/ybu1jnWM/OtUNqGLjEr/vLpRw54IMyW22BHe
fbicuJsBerUvI7OI11BbnYtj9XAP1bPLkbXPuaIjWjokE4rc0d3BbDav43suo+MZ8CuvdaGICpmu
iC6Xs7dm0ey9CaPPIUHD9hJj+rgsybpEJOkZVJY93EPnKYoHp1VX4DboN7S4Gygc5d4NCOCquPOS
ELVPCCk2yYWD2zw6+eHr0FBs73Oqjh+o+0RvdkLiyYCzg5l1eAEcKNRUevj91cxdDcoXwxhb0BAZ
JhbiS+95jZF6hyU0SzjcZ6Uwv6lzB1bpRMWINkpJ2pPy5U/VvuGFTQEgtYTPC2PAaqKy2Tmt3lO1
dwOAT5xWWw3foTKk2j4CcTx2A4u/XZzgoW3zFJ0rmgzTWqzXNumftLvUW8M+Uu9n6AcoZFl1gQtu
S5V2doy1v+mnKga2Tnmy4tVFsX2GQw/XjxnC2uiiSltP7MMkXbpq3WcRr0UjRVQv+TqZRgMBAZ2t
U9yuewqpQ18AV6/kQXPb4co4iNZ0BUPzQtXWX+bnkGJvnlZaeUx0vxzCsYEG5+cBQFWIdKB+c1A2
8+axos7Hbg7KkivHKP7aoJskXsJQQ/jQLaiUUpLGgD/52TE9SwJr6a/dITSqHPb0aoXcJ8ELeKY2
P8qWw1wi/vn8aVNDQ8nsirvOxhMvFASxgOdeZQ0LIBbMRe/hyIt+kHWSZfVGVVlOP+hGecjJHHX6
8eFcy40N28/Xu42ZLLju+LzlMr5/OClWW9p8fEZAohYZd9xC6+An8E7tJS6539QGLijpSx4/cQtf
2QFarqgpEBugxaOClC9UHr/3mq000h7q/sgPfF/CRKYTolar9FNSm4Ji4mnyathK48BFx+7Dvvm4
d6NaKCPPBjinS/OoOEVeLBPH2fLh3inUhwrf7Pze9L7aCpT8OjF3eM8pVmK/fbmsrPawSdL2v64C
2pCpnesPyWVHwSYhk5jNAoDYS0Ty+GwwSR/NrkUx4kiXmikjKMO4CA4EatifcI5SZSiW+IiBGKCl
CO3KEPvXnV10UiTCCWB2ruJYgtGIsDAC9A9r04UEnT1gpLrfo0QvueE5Wli/hmqZh7BBXNlPIqbV
3rzrXejgdCK3q0HOnxMZWXVRYcPXUUPgRRHENJlUy3s85yGN9Xb/DoPgjnT0LtB/5NxcEX4DzX0j
vXp/iDg5cXIiPxOCkCUJUVvoCcUrFSPoY/VjqasLeCSDjLtnX+ARFgrfJCikX/aKj3qRZXASAUlq
EF4pYaDYUqVYUTwZ/IqjpJmgh0diloUpzns9oPOkRDR1f2izxLbHtSb6IpTyqfvU+M0AuFdnpP0c
g4R5xIF0WZ3OfezdkVXO8FY5fBXbI6dpuAPaJZ4K0qq8VitAXnqZ4q30QynJTNVk0zjaAlKLUDm9
OFbMj9H4HZY4um+OktdtGsoqVwLA5rxfyxS8yJquOfqc+cmCBgE5d/vHONwk1OpOUPZhAzXVwGbj
fofQcjUmA3G2UI1D0Fin34AVWCqMtezcEVkDutX63NyIKk1VvgQcJ4o+T2UC9fNVU1ngt/5KUcZS
76PCZJ3qoULaXAZWWHp8ODUuCbdy6APCsjjykB+9yd/1bognZ4RAzhb55MveQMFpkGa2vLQdQQSg
Vs0OOe3MKS/uVAsUPSqhFymYEWVO2H1/ER8UwvneQTigCpwiPOeOBAOLP/gbax8E7s5HNJWxQjx+
RTstYriVyIxQhKI8s1sOy4hLk6AdLXpoj98sb8PCtwPF1VBOkrfxW6JeHZ7dIx9NDcwRycYJARe/
bHQJWPB13Hh8lh2WJ9QgOhu74krmcm6Q/QlNxmntPASosl0jOyiv1nlqdyDaVrTZwUzksvOLptlF
h+XJrFhiypXFY105yXCaSBo2FAA9np64MioxO4f+Eu042dC3dWol3KyMGIq5uaEPAvC5jmyBEaAr
iYgGvtyAJFICXirEDI4x603CovCHvN+NyHrCkmpdNBQXw+fy/UIaEvv06ivyR2WWsLjmgK9+fBEA
fRtIejxcPgxxJ14EmnpGoiE1DB3Q5Nlbc3IXKkqW9qCEm8EkrzlUX3WmePh44DT1AsePzf/c5P5i
i2y6+gCm5D0HNXuZuPH4ZqOl7d4b0749Ml5SQCCRTi7bD/mpRrqyL1uhqc/aiWyf+xSIJkVRFIS7
hfO4inRBD/Jm03r+I8+cvOdVqdCGcMt2MFxfudMWw5NG4szv0S/Lx1dzHzOxszlsvy5oHKIn3pRY
kQ8HwtcaKkte0X1fJxTonX7bkrPOEUg7tyrp9yLaennWKev9hg6gyuJ9uHBdFlRFYCAE7tciZiBC
yOa1bCB1wl7lL6Tmy0NvBYEjL5NLKYc1IMyIQzbjk6bZtethn/BS1j77CYi3ux0L33WGe/wDclWD
podXjC+lp0Ag/65LmLonioxCADvh+CanGnmFR5cty8QBFrFI17BZ5jJJzwdj+HgEX+NHE4V0XHjA
JWkhzARM+RZrQYYWDdrkUXrrCLJooNvNlr35lMlhCfnhXqu/qxjyIYSuhT92aoaxkObJkBGyTWiy
b7W9AR2wFs0DiiIgRJOJVHQIjzRN60sh18fVyPD2r2yJPrVRtdWj2fmdo4FjU7NeE8RYJsImgyX1
jJdn8M8pkc2uupbk/UAAanDjvFTVFVRjQaq8K2cVfdoW7J4ntUM01cx+ool1/WsPJby1hiexTrgz
pod/xlLix6BgA/JshWLXlZxGT8tFsSXYt46Jse28gu6LAjWHbhdF4duVsD3jC5BNu3AR3lsOOK7D
TeuFF+X6dqdqJV0tyxp208MFqK+aNKtejO4MxdaYXyc5Ej3PBfgN6A3PQuzUd7V9wrYiMmGzalJq
RMA9rbM3Bov7nODcBEYGMUcwvqv3Aug90NlRGrPKECNfmlUN6gOGw/5NQwWRfg+KCjRN96DUgqI1
suN5vjS0dZ1YuQw7ceye3VjKwZ62y0BUQ4zqNL5B738B1UnAS6hi0EwQalnuKFJAPCps+t10E4tB
snyNwrBsppWjQCK7axJUbBR7v2VP2DdNuP2J5RGorGYbXWJEr/At1xNW8FsLP9Ov62q5zHEVOfq1
0j3YpxqdFZnuu/ywNFvxuq+2YhXdP38Hm6MX4+KPeXKFfCZkaT9ZwFXbALGh9BpWI5hf+uZ0vCbL
7oU0VY7TJWZidGUe1BpATRgnBrQBxi+jP2p8VRK7fWT6+JdBU1C1panhSIIBRE7mVgx/AtJeIg37
r8fA9j1eGaP8LHi5uKKKIBQCbkd4WAqYolmaF6AVxpThHBOfpZk7POcHwAgApjDfDbC0+A+aZ1Di
wPXSUmQyj4qJrMQjGnj5AJ/onWvEmRRFs+DeIzT7GAKmW1qaJjq7j1qABn+QbXyJXUXpc6z9QSXM
CfrGXVY1ylcjl4jd0ZqgJFLaR67qLVy2WAyjVvrRZQiisXbZ3wceFTL2LBuFrjRFztgUmoQnoBuS
t1M+8934zDPki/3G6hwGeGlZ2devcGgruTw9lDkuZzAfZtGcJsvhBhyPRgx2gIgIdQcexAq1k0I0
0wv+Y0Nyzgu0lqbHPInA0k8aSzB66r3pOOLFR2K8nCKInF4UY3jKvUY2HS7W8bhUSwEG+rORU9GE
Nr2Y9UFKFBzcc9f6PGG+/b847o2Q8gpzpYkNGAwKW2opChic6q0I85mQWwGlJtcQ4Y3VUJQtsGVD
k+laTZXB95fCxILLPfI5UYAYMIvhoCmQC91Dg71MOBDS6bvgxp2jzq0HCLWLesz1itxDHjbLjSN2
VsagBIQjHie0bhQpGEzkhW4yZKVdoIVpaliNEd6sAdG6dKIgjGUV2aqyx0uWSFzePSqO3+b1RXJV
ixPq+xxv6gPgItBHxgw9W1mb6oHrC+86eQIg02vXzKtvjrlWSbTlKFFPwTExsZQmPDDQJ6TYiDLF
p/OmODUjNaNTs2aHHjhkbR0r2R75QArRbvKfNA3YBIx5uk+dMaWrAInGC3K42Qplo5A5FUVGlUBN
Xwq1OH/pkS2OahT0Uz4FCbtTOEUieCX2Mrd+UZQmqYM4dV/kjR9bh3/zuF0OXw3o11BvxNfrNR/o
0N5G09jzJ/bNDvr3XB9D4BQ1pikkT/TA8Nz5N3hDour7J9H7L2O1cr+ETqOzaIxZlTwjqElZ2YZN
nHmrAXSSf2vL780bT9081v/nXrGGXC18ApalpBPpp4FH38kRAzqD7gtWKK1dIQj4u1/+45OJs159
AjLoeVqPH82DhGXMnlOoo1UQrAewM98TB8MRo6Xf6KtEabQ3w+TsNz73v6U0m+QPV7+v7yEM7nD3
+FndMZ37S9cyl/dztbqquli98Dra2ESmqFe0RYcpwnp9KR8hL7p716GzamooKBwRa5ugq3TDDEMK
plpKDK30F43Bfs+JplWriLRL/GNGXh9UON6sRe8s0LlFmX7T8KzkTMZ4GbRAYT1nCUVPm4QQ6ZZ2
yLoOLqKtdrmCojbboxw667jf2+xSBcb53ZLBmCJ9gRNwVwU8glkvowUivbtABfv/CFz3WB7boaQt
ztJ/YZKslQCfHtcdJ8gJHg6bvtZ7pwf6A5LLwq/rHJDwFzSEEL1hg13mnjqgt8sh38zN1szKVRsL
3M0fhM+XQNTpgAQ1BA4UAucQaIFCZlAsR3o/kVOyF2Ij4NZ0XetRkoB1ehNBxXbQ0CGcw7ca3tUP
mcFETOeVDeHue52F8aBcf+tAVTEhhi105AYTaeFRfI3H7lfWvFx07JhxBkWe2HNXFN1ISSwDPXVC
+jvFJk5PA/LhXUnnH500+XdRCJiRltKw3L6fbZs5P3Q7Kpn2sCGfGA4IarNI4UAVFWYDsxf90oh+
w2tuUifYqBB4nXBVQyRdnrKxIuY06NsUqVvnyemS2iQ6eAzaYck6ND5OSQuCzp/l1g7R93RCmVDd
/E6TFXgcI3TWpsuMqyST0TPl+xNvl7wTUCntTJbUpykeQhHh0BajY+YSFxhfrYYhKC24AD3iRVT1
yImASH6QXE7tcJ1uqBbdRz5beytgskJT3NmXonOF86eaDDiFnVtFcmwR1+Bh0fPvKS/jr4qojct7
dqu7iDrBLSbIsb02SNzUrSohiInvOZxZ1DnsINHbi6roiKn35lKu9/uL4ePbAwEAbsNfW1YLDqol
z3lSJIPYm2jqh+sq5TuQyQRxgjRPey3rY+MYkD620ZB7Ib56+sVXlvWHTLb+yvgCPbO65JXDjx+g
saRj/2Hjn/2cWr9R3Rag46GGXWaOQcCe+5OV3j0GIntdcjooOY+QW2KOofkU5FtL149KkAWggdjB
Ya6fWTqeYu2HyI00Un6qe3pZ8xEXRsIoowsGdUVZIGJAQ3dzNPFz1H7X+bu4H5ENkFlSbvLAm0qc
dDQhN3JximWFCHZfwogFkvNSDjjWpd5XVWb3MU/n0wdy72FbLUt61IYZhPoPZ41QSuS1XcqTRH7X
A6j4Rm9eqmHz2Luvkt1UqCrrbzO//xn4XWq6fH2GQ3VfO4y2WrP8WAFdJzWjFFF6jJOLRfFKRVJx
BVWW/rCTuYHJtwvXC/i2HmYeS2rAkUptkOiVFEFBsFOpUnehMmHjILyZgHE09OxuuUi/P2n93bEt
5LEEtrZutMOztMNrEEYLjkGBeiY6F/uhw9vrGu0bfOd64cvseYf1FImQUtwSFneOa51n1JMx80rD
rLfIABGv9SN27rKx3f6PqXMNeDBKI7AyHGf+IJrcpdNHuUcXTuGJNKJ/Uk8OfWRRMWqDrr4438Dn
TGcHcSTZbp1U+aQPln/g4qmK/zIJAPbOKOhClrdFueyjCEx9wEzq58i0w0J+wfBNmqJPbAik6NjN
sETu7gLJ5k3CV+763PRHsReNR7SUCwlWceWbSyw6LtqgFWpffuINhSnsLgHORYJWU+GWvAveXhV6
H0h0nAVa6hM44aFh1DxL6kPFokFtZAbJuUsH6v7k5IiiTeiJfg+585ebYSVQpGs9hUs6neE6swwD
JOf2grW83K2/U/9rmMN73p2yf+F85RjtdgrbgP3xIz+pJHBBP9BDj5OvWH/l+rZAHLQhexjGAxos
rGzoZAU28CjP7kVLQ1g1TS+RUz00MJB4KawfjNvlon4U2u2cO5dOUvkCJDSpVFbr8Ta6TwMHt1QW
9fprl2oAAjK7ddl/QNhylxg1X5+MoaxxplKaSW6+mdJJBbgMv2OY8o7K2Okdn39GgptfFmTezegy
81hlgcWOLBPdWYdwdUGPyB6oewnIUh4nNgni0VRxcx0pNAfITisKjTF0r7HzPWeq3F5EMcEu8G91
Oz7SweiLXmghagjyn1Ts5wkrVK2JLAQdJ1G/6y9N/3ZC/ydkfM5ZwKWWFEK84506GylItvD4pP91
j2VGW4zMrj+lElrZ4t98SIuhakJkU7GWWntBRYryG8a3Q6/ttZFguQLQ/XONKtTs/zUCVY9n1q/G
odKd1/CmdpXc/sdGqb3LVfo0xVAAf0JlvYwtEmbQu7bJIwhZB/90oBUJZs5y72awWCpL4NcuMthL
7EmACqRvbxe8F0B/2sIX+OXkPeREp995sZ18R65IQnxQAdS89x08xsz2wvJwm0hfKGIy7OmIBZ6r
O6G9OOVUfmtudg/rWpe5tQK7V6XcNhNXibpKO8IV1EC4fWXeNwIZN/uqkcrmsAbvzqrW3oMmsdOZ
IVWNtgs5amXuseltyD/L+4HinW+gpNnYr+TXwj9Q7RLhZry5+geY8HrlBMIiVA9p5vpuczKhUm2Y
ljN19cLE4rBEUZYKD1upV36KuvMOh/7SCslyPfiFsZmXGi2UaUB7R3jlPirJ2kleN8KuzvDgDMTy
zTIfa1nJoDoA9iJwshQClJy7eF0/GEwJZxfXemaYmW/xIcwZt+FZdtffnOqdguSfNOdpgZXQq6ni
83pm7fY3inLYs5iSCpcrcvgNIPiU4mLoxpWqWbhDNRJrS+hmUXprD2RTWIqkfvWOakcl0miKgB2S
YaAAYxcr4vSKXGgsVh9qC5G3r5HFJjRXNXSupCeW5jaR45YFJA+ytRZcO3gH6Rv/PeorSDdFegGU
CcMAaGT2OvQkQ/lukjewm+SDPOzgoTYLmUPHphiIVMR9HlM4TkpTICKdvQozpcYSkSoUEGSZ27p9
+WBr4ixIRrUgUAkds9G6/mah1No6oiJOnR270qnZPAhAtqQA5GFNcmowmKzwSzgxWibuV+RJgbUF
kouWPG3mb8rcbSq8X9GsrpgbaBAqsGQwFdeIm7K8rnFMEmOj1LaLZtmnjwnHotZ3AXsD6+v6bCV8
q9bi20wo/X86bboQE4h5e4rshdF70CSeQoNwyH5AjSNdXB9XbDGLT1tp7j0oQbHqgS/T5eFJ6/bd
O1AF2zT8y9H9wFAjyHLfP4wAtUUeM4FbB4iYEeWITWPJVMtrAz7fpNIIfeVNxQqLKAFS+MT6B1Lf
YUH55KPcBC1LWd2/hrwEejWILrllL8n9YM7CoFwJCCsOIVDNEuJsltIrcDdO29hZ5hsH79OTxZeu
7z5bWqKpkyCdQTfClMoa0ThT2gV/baUwPzfdDt/e03MY6ZDKJaXezWRzmGLCkJr9B4ppudH4vbYA
5rdsMpadV0DSHSvGHy1NKG7fDPQUrJ1Tzi7al/43168laeUtfDgKFusxNooksyfu3NiLVBSHhyvg
igONA2BbW0CPYa7rV0l1hsbXqFp4ZgDwlziQBwhD5HzZtdcSLGZM0FGKpbR7MtMl7GaLKQ9MtfOJ
iQjBd26QAJpRGDz5Rp18PMJ9VuYcvvSQMuuebSz/Mz7C2Yn/op0ucm8qhj35VnJWLwQuFLTf6Qdv
7CH0GMMmkF5KoJocdCdTdz7dXRHQ+1SAdpWocJdarKbfqDmI2PsFBNrwh1O77Ij9q3tozOx3X90C
qSPu/ZBlU4GFno883AfKGtzj5gVBDwgkfv57bPfc10xSjtu6qzqJNKLLoEiJ5tFDNdDQdYP9V1dc
/1/uocRA+SJf9Ey/Q+5Y7NGN3r4Fe4WZn81rOEtbTzOjEm2Fmv+jsaFt+YqvS+sh4tkPmdIofItO
A03+q+mcAGt+tP1fk3b4HPFnnkw9NveIvLfVkaZkUL60MFxb/hcI1jopGy8aGTd6BbST07E+OY4G
KIlc09OdO5UF9O20AaY9C6jyLnXMMNQrIbdpf/Td13ADCBa6169xDCu9lmSUUKtlDHv3ZbWjTqmA
Q2RHCm+KVd9dsJ/wuufM6hwD7COadj8d+cvsOsPY+8YO3dEnBjLySVfzgyYLRmqS/kwmIbYvhJ67
rq35NXJx9y/0mstYbRAACgEQKD3OT3HAAx1lH7OdWmfP25O6IYoMHuQt+0wpxhwEx6Fgc4qkxCqu
Sj51815ntjuGIfjMSpyo4OCwb8qc14SpOOL26n6lHhsqoF2tlQNh1ZRcxXT2qXDmzlOvmlN9jrDz
rwLHDdPuczLEIvwOr222LCsHFLm6IXUwdkK+DBwluHmzmJhDLa/ousdcib/xyMY/lCiwyIBgnlGp
atuTgHbkJaH6UFP07wt6mPA2EjXLx9rDbbzovgLB1zYeo42W7c0SU5KzVFAzJVZPQMXt1Nn0kV6q
7qBA31TcirtRSDHjVNZ/kv8F6W44r4zgkwqznwM7fZ4KTQ8hjJabd16E18zLaDkSVrLi0CC3ApWe
ZFWZwmm5pLlHSolAsRmqF5DuzGknjIkfVTpviE0scdO6HdJmfTQCHjfWhrjAc50ha/AUhIflBa6j
8KfFTQkK7Z0X69GSNSF9nJ7yQlJ6SFZXW44K2KZmsPIc2GEI0XDRZtyShG2zWVMFzq5jYsxAT1kY
uCQP+VOJSk5UOMsYhEc3zsiutcf+29GzwC7e65zGv09TLtO03RcUCEQ2a8NElNnJL1JLqSjzdkzs
vvegzVno7sB6nNSo1fn5gskQuxJp0Cey9wvm/+gPbS5I336nxMJgrB7m1/T2qml7y75WqP9KEP/e
6xp7ZUvM6QrhPaJrrAcyk5K9MPIdKP4/qOlvFSsyesAx1GcHN2RuiBKZZJcuFASs7LEjvFK+TMfs
F9R4Ppt3sA/vubmwKJ0/7FSLiRP/Mt7V8mExH9OXOLoEwzvnFYWNS+OSOrNOyI9sExS0VNYB5YXN
09h/2dhLL+TkuBkLkrT75sM0QI7pmYiaA5A1l/YSEAUHjHqLcpJHl+9oeHT7wDUMX1DcLP7+2xOW
UjXB2gtTfdotSAf/Shfo8vebKPmtcaI70bmcaZzDPBBAs53NxU4iRBMTRFN3fSAMxhrSUtYLTq0Y
7ktqA1OZ7LTMl6YV7F5mmtDYaDPWgBoFnKmuzs99ireH0CdAgHLQ+f624DcMnKpFeVNeVqQX+/a9
qNMC/E0jIQ8Oeb9QYjlEGNgWaL3sD4NmXmGil8vf6iFFX3hPVY4t+G1Jvh7hwqnyFlwzBGiFY0z1
32TCZdZjnKMBTqZgEeM+cMrALZG4Y2stYWNZptPk0/nE63Dlft4ZpMgrKOnUitn+TkgahGv5XBW2
xLZl9Mgs7r6n9gUxuhb9mIIGENg+n2IdCzpnSenh9fCl4ipQQsb0NX58iYosqIaH8j2WPeIwHXAA
MAOfKi4M1q39i3wQaWNfOyfC20hGDYhtekgTVzFsAC70svNlO3D/HWOVM7b011ii06UFWSxCUD/Z
/9EN6qQjt919dX5j9NI5nUcW36EbMPA2jcMEdPTAuXA6NzvnRGcWLDd5AvSgzbgHkbkNAIkhkS5+
zdTlA/ALvD5ilYJOnpml8tGsqZ1pepvmh+u/Szb9jkmeoA+A7aJ6Iw6u42QS2yOM+g6QT1gJhL50
dz8/3WSgqL7g91wpAzmaNgx9pVztqojcubPYmorDFnGfufXc1H2rKWVMqe35t8IWTNFPMOFR85aO
jcTr5tdNyR5qEAYozngwn8ASC75+fakV10LkPeDMP9SBfBtbohhLMeP0cWeWEtR0ZO6WRnW0Sqar
mfqhBGUJnklqzcQrmAQOrHgBu+G/EA1SRqJOT60RkAhQukcez6ymxtwY1dIOVRGc6YVkSmOI6+EQ
LRaRhX2tjxDQ/qzwszEc6eA4iBchjN9JLsLYKOXbFhS5d7rPoWxANGTcFfCzjqp7KIrBbY5XjHR6
Q7Jh9WSNAhjtOxNcP6ACt6kK7GYqnB9BUJkt/XnTBETpK5uSwOUeH/fpEEswY75jDSZmt3dld7sW
Pc1dR6thSkCNt8brzvS5tYYf86eCUWet2svFFMLLtgs5ODYAGIho3wUPdI/GYofunySF8JrxoPTV
XlVGt95BW+YsY5mmL0X2jK74j6PEnGV3Yyx6VsOLVGSW7YDHXsxVcfFJQ8IC47N6GjCE0hsS8Jr4
ZyTcokw+cOYsU9NUAr01UcZtpZccz6b1rNW3WZu496FJIorPaiTJh49PyEl2X25RJTCECnADA+5J
cU/XrNG3vkHpa1FiEMCLf751/X0NQA+56a1aL3YuWjTj5BUbUXvPVmQ9LPCAqDqO9/X2VYBOOW8o
JkO79Jo5cSEEIt6Od5meQxVOeL/TzEgRi+5Ot/GERf1kHBIMZ11OrswLogMpXAB/mXCKqqJbH9kl
5TkABxjfMjXK2s2B1W8UWXhDcSptedcYhMOHfI+DzCvVw2J0YBB1btMpkufHeenoSsOOcDHUhNJE
AINSWy71Dc6CBUQvkHnWYRWsloFyt2B9pUUFsOC/EcEKyboAHKKqdtJQUjivwTBQlyDVYE4OcJ2P
ISAuqVi2oMAPHyGwi8CVquSlC/gwoIH1LxlwHuYmGykyAW4sNNy8DdA2dMJTWcVDGPDnHQZwBoUb
aFBzIY17sa8XHrZLhbKQ9EWlwEeSPRvTnN3rIKOwbvcHdjqpkkFlhD7EMfkO8L0qQDNdLI81EUgC
XzD1HLIhcxo9mhOdZaGZHxfQ1E5E1OlX/v2e34kOZFyNnd7aHbRLX8UsCYvd+pB/ZZIbqZrYxaLV
+XykLnDNWic5HfQ9lu8ToCI5iAF4tBgCn38xIleNQy6p1sKDavgjcBPG2cBgP4cwppdMtSeBDbs/
3gR4J5UV02QvtAkxNHTsz5C8i2rUqsSBxZ09xWPbVvNHuNdVNn7/UXHtDGXBaSJgbOFISjvg3IIg
r0qdbKhizZby7D8K131dx/5gxJI9yErtU2i8RGwx65cwX7kqgOM8fFx5ZJhxOwYTUHbWHWwtzlKX
vmoI/UTrwYRVb4BP1yRGr06gBslEQhaxB9+bAr6NyXc7LFOl4ZlLS6uZ3KHBEJdgU5hrEwj9bUU8
oXoB4Rp8LMTcp3LKA/sHzRzZWWPY90Az6bA8Gx6Ahgn4q7f9M2mPf0jbIVQv0hTvTp43VTCYY8kI
sCBWGe0SZPI7xd3/9a56/K79ge5ztBWmn+3MIqmxqaUVqceCzgXNOOrXKJtDSfSZzYIMY4El8rEw
WRrNOCYpW09BreTUDqq51/Sq46WSMx0XZxGpOkwg2yklTKbiR0C6rukwrAh9NcZvMWJ1kF0eEROj
WOlYVjP0mZT85IOxZ2IlAZTpp+kp8OwgOGYZExY8tuyq4cM3W5ZizYAPM50C9bAzcDzIeklqGr2L
15/+CXL0lJ5yU87P7KEwccDh1sdRu6Tq2DL+rkLz8Ld9CQUOetosRb7DYM15w2qhEm8IWy2gqJnI
2CSzR3z7GH355IB2TBAjnrCcWhbVATQkgsfTWoJlhzB6VDUru5JVeIowSYTQumeQ9UXuVNwyLHE3
6nl/bE6aAZHJa9NrrLEzAfFiCyiphCDifc4ljs+416TFghJ84LChfHFpLHnZOy8VWChGpGKPrYyJ
DXQGA+9mhTAxhhLpurjy8MnpsZhcdFNNXWaUl7/IJO5NfqPj0lhsHRQttFu49DvOaHZQgcGov3kI
J9Q8kr0XSgVt28GzqszUN+NJ0AWg5dlpfgkDfjjFVBBJg9w8bsf8k3iviq/cSnrYrXHI4tUN5JJf
FMIale80dSLVjgutZxNtq8omcKwbcqoaNzYK8Fn4XJZJFKccyI6QUdGlUIFOqenxKR9lEWFOSyXq
6BtEhgoGri3B6whP8SYVZ2K6/jKO3F7pS4OXGUcKiX0/HNwx4ddV8pq07rAZVj12s6H9mK+6rj6b
MNLbKQcy2JrrnPS6w90PNg2GAMjVcH6HZr05EhzfvIpi/HxISZ6kYb3XsX7BB0EMav0IAK5T37Xs
O/J53j4APt9nVJ4RJpbp1c6EpAFn2D0o2uq3rcbyvtdBRo7UAsNWWSy8qZowxFwk8UbAhGkv3r6a
RNfSSNHNDuDV6UTg4dqwegXVOBWUdAkseNrS1Mgw+jH4FbmWuxA90k1T0a0MmtydpeL1TLl9YWU+
/yzbw6m2Y7XwxbqeI2Xneyc/jx/3tCwkq4az3l9oMCpzidBLp72dT3ItwDKynfxNWNa2WKlbHTLz
+sd7skpR6oHr/Opruks1BZC1yZgeNa8yCBWCLMweyU8YGeq2tbmxgim5zrvPBLIaTu6yCoYWkG8k
2H3yZD7Qr/Zdt1pKY3wS7ZQtBWefsMghp6IYBP5faPP1QopoBA9p4JuaX8FIdMLyr27+uUn+yosm
y7U4WhPTOHuKOAWzuUnRzkHItzAPSuIThwwyulh2K7zA14CRbBNp9nOu8giJUgrFsuOJygdmTVsY
FUyDL6K3jWvOelr4o6Yb06BukSX8839YVM9f2VO+ITg6BuUyShbAN4bKt5IMlIMeRj4KLgW/xhNJ
NWAqOi0vLlcN/P6Jepg9NqgN8Tml/mdQmGeBmI7b5ytt0i00EJbsm8dHLR9mdiR0blaPNk6mxLRw
VJ9t2cF5hSsCFY6CpGiuw9716va68GPL4u0BrgNGRflpMFHMFf6fFtC0OVLIpRiNEyQRmQdIXPWn
h9qpVtmo+4tqrZF9GJN7n2P5xrEI7fW2mtoEYokkh9t2Id93gjNEH2y+RcZZlN4ktjsmC3OCYrbH
irv1SZqKnEzw647EaH+SYKSM+epdP4pgQz54TX9MbCDMyFTUyqnLZ4S2FtwU/gxmA6RqPj6GTJn5
ui+Otn4E8CwWpvKnxibf331bB3Xt3ZlbTL3RfCnbvVqVeYr/oKdk0dcjgIQX/GEbCYK5okgOQUcD
G4IlC2iMMe5wpzpmtAw6M1Jayh81tH+k8c5HclK5uIS6EYpYIpaub44/BYWimwSMarVzZa4JD8kQ
zIW5l6aw/KzZ+iNmk2dgLX1tIjrFdYDVIvlvLMQYNAnwSLSUo6eLmt9aPk9wQ1fnLsLqiQdqhzCn
KXfOw6ZbswlUfm6rv4NSBB1pEnbqZLVK4f6RoM46Bii7O4rAaHDzUJoR+JnZf3Q+Rn4NIJJI5qv1
2q0FBW1Iey/sISD5H6i3dxnL/0Bzq55ozdmL+QZdgkIjiYORZWCYYZwFg9QMW+ZNIy1eM8wBAKTV
xCH64pcvpoSCMn9onSV6YVO2mr9n7uvQXEZ1FgwfUMt5QlMkIhiYlT0gGF0/EzxWJXu9EmHgblHS
uJAIDl8wAgakzjz63zy4KLNAAabc3Q8bPc8la2vf3GjdgBjU1WX3Jrm2XFRdwNUPFJTzKiyNJZSw
OQ0JTr0Zn/Zi0/95qWxa81hgMheF2IzzB42hMpgG/Op9YahjAGmUxRc3lwDXhbVLd5kHyvWZLAti
N/RIztKDMEMzQ53iKCMnIOCYCJFyPOPO5lkOHNPb38n6zS8TV555MUrmtawKZc1snhqt6pc5kUaV
r2Hy6+zmBSI8Y+I6UEVP++9B6WMb8cb2rIdivDrP6mFyo58+/Bo29I4ZiR1UuDgsLHawClKiVa+b
Dgg+chbaPFPVITo71dHNrXb0p5gtF4FrsHfleCPBj7BFw7PGxvgcZBHE4Cj5m/VaxOP//JL0zsrY
v8ppUxaVPeljLfZXesqg5iNlNPUdRbNiAcLp1eyzCLZswg3mS+y8xicqB5ohCpZ28Pa93g+KwKIo
Kbw0mOa2PWW9vvgq/x6Mo/V+K5Up3Y94nltUesqmu99KIQgNpTF3T1OC0yXikLgQYUIHKWSMORm2
XxP26vTR/V57UZXtgpsiBDVAaiJ2esAmXrwZUdJkAT9lpo/QJYetoIyLBBwsYPkx+hhQ3I01iKrz
cqivHQSo4O3F8sLSypVfdVY1a0tBshP/MKqn4rdVFGlySBGJn/rnGaOxYwhH9tMvUsrQFBLCduo1
eurSgYy5klwbXN1+9Ub9YrgtE2xdOos9pK3fK6A/kzNyJf9PqZj3MXwWnTDT6RxJh8NpMYYoXZa0
C/KRgB4An5wnEhC6DNPgr1rZbuIaZ94vwp6Z20mIrTI9I/RObybqRpthy9m7YhWu1cSioP5G6tfQ
1m3sGMtt93paP91AhWCT6yDarzBOLvV90QkJTlF6NVKOoCJlz8b0b0P0diEUaJ1dbLxjYd7qMhBX
sy2+ak9B/28V0AyguQyfY99QBKhYCjaKWu5mUNQ5bWIFmi8dzRliPOChFwoxuFdcyr/yRr02HscC
VhKntWGWglcL0ZAHLwfU9r5B+8RIK7cxtnwbuYoT2dMGz+Nveb+w8wtyjmhjHfVDogsKARAcXWEX
kirImDJtFo/hzFODAVtaVDa85sh7vh5l5PvlaMq5FBx81vsHFwJyBLmlziqLTGd/zLatcAMKzlJh
86+dYeXT3unmea7ocmmTJpJQOLRR8pmZYCWLUV8tdpCb3BvIF8VYIr29QcsFnLbYa4hjCzpm74eF
GjbIvX3V1oigb83mYS35POBCWUVA7IdwpoOEOyM0bM1p5wBlc7yVTQJ1U1mE70CQnsTmou89ObfV
ZAHg6GBRwmbfNLmyOcoSmzZFSSqdtY8xcBF+/do0oPfH1Flyc4t5nv4jGtuRz5m/swBfvHIKGP3U
8/vYTlmO+LAvt/1Yl26xpJHc4jWaimMN62Vd/kTHBUhjiy3DNKnBIrtMcq2gVKBJ2CxWCkuHrMmP
Vk4BdvOmuk8sNm8Wg20Kybfy3q4O+6jnclZ6cP2BtW+dBtBhFcsLvRIKuw/g+xrAyohsmAq/0YH5
H/CJ+NCsMi0t3fgNxxU6A8lSiTXqrjZfEvMyOdB6qBH5qy39NRh7iy8RR6WYrsEs9KkbXFTStm9a
DcCDniljbZG6pE8Y14vnLLv3aghb2QTW+BNnnj79OzRyZcc2oeKmw0acriel+Fneye24LveJTCAG
+xCNBw2JGZn5LWuTvTXfNOcRV50EYb1xU5bmd+1Z/OiFtoLG2IY/d2ACAeG1lDv/06kmvGX0W8jJ
UluTjtJLGxukba4Fiv/OJwn8uyEg/RDE3BGrZiMs4RYOq6LsbYhXneSwX5GuviIqtYjYFBqM+d9T
47tui/2bniIJcEwPQE2QR7d5M9pp9+0UDSos3L8S2RFpZY0QAttDwmD+3KVNFPt6MWBMP+EkxLZY
879fNjVDHMbuD3lB4aaEcHgw/yIQSjPQVbG0VRAjm9GEo8D8yeV/FRcJqV0wxqAYxAC5ebz9uOr3
TgMKXbCRvRN6Olz8ykAJVSK62Cj4dfKJeKQNGOyB3i02kHpHMF/10F3EOqGlBgtfFwVhq7v2u9LT
6hWYL47BwSY0hLKf8W0AtEIw+9FOE1weYSL9m+Jbiy83um5D6gT3dPChA6cz2PuoLNUj/BEcck6A
IQvKRjPSa/DC6NE/IssaznH6oJuhO1G7sKVmtVBcz6oNpHSa1KBzXorOQjVyWbSDyjvEIyzUw2/y
C6vTshO1HEDO2OIbA5gPaVZvFLZ1SIsGE8MpUNq0LRL255rAC14Ac12tuMCmmS60btFXFBvBOuHH
o5ySSsrrklnyuZ5nrnWhkL93TKwZ5HeEHGzlUCz3XPFbE3mpqcj1zw8lJDO5qzR/vwAGG/IZgPju
gVIv+CvTE8A7U8p4RIg6zbLrlOuM70slmTqkw1DTS5if6p+Ws1OBrKf49ZovYoCnbOEgUhcHx6C3
Ig/JC7zG2D8FXvb2F2hXaIANNS5nHlUdQiSzygGpiIFbGTaVSY+PDo1mrzXq1YM3Ke7yBJLgQ5G0
LSgeHWBT8pPM33uxbBjYOhbzcMngpxtaTY47kw3UJwDb6NoRSBTZk8b7RefjPuq6d9wMSiqh3RCa
+s3u7YBlO8jjmrt0slEzixGQ0PXKJi6DjyAILISFpLHG61it0xRw2A/ms36u1+6Qjz4iT0xodMeq
/dWi5uagc0I3yp99z9l5IXMJUApVSj8TQIoyL8eoGbu8pKnTmODH+ziBFvL8mSNVjdwJBqMELhix
YkMYIBefd1+EnvMVzl++ZsY6sP97/wXR1hoaTXZdFRhW+d65vpgJaKmJN/b/2uDF+nWyU/6qdm9Y
+CbNT1JWkfhbxuWP/taZg0q7JKpY/MwVg6BZKW5lfZJtb0LFI46I4hcepZziAS6ftRDJbdpWAAaV
dlGPc0QJVeiLnmHocCY4ST2KCLIpUsEcwTaqQS0bli6MI9oJI3UeT9SIB8HaK32qm+rEoZz2IFLT
81scUosV+qL27I32ksQGKPuG/QzbFCNLqtUG8VnVoc+0V0WB2+nRuSfQb37ey+K1lS948EdDtDHK
DHfrcI1M458t8inOemA4Bn7PzlImAcfEpCVMwrAOwHlEOwVHOLD8Rs4MbcdWq5WWin1cXZQgYfZC
fJ2j2phGiOVyVsMLqEm0DJKtjRHv7aYsFCrSpqKJpXd/9woydfMAIJ566g/FILMLyROwrtIBdCyQ
WBb6qigMZtjTC18dZpyB1KEqHsL8TIJB2WWHaMiaQvafHuSI3kz86kfvrRHBSAAqKv1JRayGoztQ
VVvd4Fl5G/I1bKpRocJZ92RzPgnr0wc4d8JFDoNibkLa3vKlp6O0/MPUG9YKlXUeu2doe29mckcf
67h71IE2d+c39vIR1qY/6qBPRlRZmWUbDtHeBfQ/+u5omDJ1/ZgsIsrSgT4l/fBBwSlKMmFdUyCR
VEz6whqgsWne+KNhY8qVM6yZan5UOUjJd3/ayiEG95dOlGAxOxs0CCzri7xpvWOLOXvxa10cO5D1
4UItHfLihJ9oJVBl1zB+8Zi9vcPe71DRAkUd0p9Zr7ZTDS7SiYRL/qpywKdn3mjPWsrJ5MvANXgH
+8YAJvqNa715KjD4KScreM2FNz5f0BGaQLpIbzfRcj8GJaS3Xy5vdD7tForm/swLaUsbsYIlZlD8
wEzB+/jCfEhUlEKAMQjchm9quiyrLpzw9buFQ8O8t7N1To9YWbNhHOJjXmoQWVWj6PBPMY5aB8YZ
FKpK8fQ7ZaLZ0G28kJEjl5HoW6r4Ydrwe83+aOBLBULeV6HO73yETqFVXCN6EILtiztgGBxi64h6
csSXmBJFczic1umMDkTEJXj11Ci7WUbZR/ZJDEMybAr8MpMjz/0XVkQaivfun8bZCdJyNTfBVcI1
I1RyoFHz719Tqm+v3nswq1uMITEHfkFXchlpfjZARNI/vy34ZjCiimD49/j2AfIVGGG3mnJhCFoM
ozIfYbPjeDS7Iibxmr9NemojWbEs3X6wRzeUbv2AIsDp7m9jYDFKMRhKZZ6X7Z+Emf2qxVSrzuSK
GIB41SDVcYovUBYtpGRTM7FQ/p3KRi1QiS8sVsFKZwFeTP0/BiGQ2a4+2y35hbTBOR6RhBgqx3/8
/xO/cV+SWeAt7o0AGHE7dEdNy1LPZ6kKyU3zzOx394QXwM0jpcYf9u3evmlFVwGTmnkxsuUBOnww
O9hp5wjZkvWt023mYP3bptt2oihv5AUOf3eICjj0eS0HmVrt/hkK6ziW6T5on1clWY+N6ztOah88
8iljh8NgXEuJtXc6vAWY2u/Fx60k2KBZxBtatopXDbNoNsehYyATi/jCx2PMNf77lJvhZwCl8FOM
gjkOjVDsbSBNyb4MKL7O+n2VM1QCTbHYcPPysksXTOuN1Noi8LBM4d9fJFRb1r6Wd0FNOENC1aTb
c6oQWFguWrYfG4qzoRG5rsMwH2GKIwwvQe0mgcWYcH7dVqn4op18Ub/gz9Xm5YvSxZlpGeP63Qh/
SF3W/vrbUBPqRS9sytCWRjDpv/9R9RmqJhTupO6kFY5yXAD+3+Fvv0wQWNALBomcJ5e5AVDc1FgE
xj79i01XNmRPYiGwHhhPX1xC7yLWbY/C/lTeInwpotQ03XHfEeOZJWbKjLa3yE8A0N4xpT4hozN+
/zKiUwPzR4i41uaVLSKYQwb0+ByXZzkxG0tudYXvC3GRgjNh9r4bfwQDIZ/FYS0g/5jzy+vM46Vd
g9mbEzQ8UBiWul8ndd1ztFyy6e4au4LmnYv7NNu+iRkjfjxKrR38WdgcJ0sqjgLE4Iao4U8+ksbX
cVpHfUwZEu7DqSWTG4HsDkoU6xsv8K7JkM+DTAg0kA2fgyTmZSkAbrNq+AfggG3m9C2z2OATokTM
FsTEYt3MpS9mwexRoe8AS+bMITVwC9gM3t6/PMi3y5v0nNCtn21exf+b4YvzFc47bhzDi2cvN6EX
z9UdYypJkIoLURrDX2+9QFay4Gk+GVRtbkAbQ8+ARThIIeGkkG+FINn95RiLPWpK/WdPZs3lgtQz
j1oYIx+0pItorUi3VHmWP77rewcrAa4L6M/wi+YAx64kPfbZrIrjVHYB/hNiGgcMVnXDug0nCBXU
n/4HtwQpMtO1ovqUBdBs/iztDX9dmXw4bH5Ar28n/yJ6tQEJvsxyJj02VbB0ZMZDeDZ3gAAD3knD
VckiUVkPcs3Asff8fdDFkow+EAlr0NN4l4wyCzd7nWhbja3xGc4fRCu7FnF0Z5LoyYoJPgm9SL57
SroHZPLTTPbAILrIDvHFJJQmAc2RwcUAKDC+nWb6M616lenT8QjQc5dICVV+u7yOn0shBs0ReoDo
Q+Upwi+uRf38CKa8Nqqp3bVoOSgplf3rQhN7WaOpSNqIMEEfK4MFbBHzG+cXzq0pYjR7lgVkKQ5J
qOgLbmHlS+/j/HBNwK3nPQCgW0lNi3oo7BPPR7+IBHLaNg8Mq/OKZIyYaxlRKafvxq2PKu7dTq5K
Y50p429xjJfQ7E8VUnuTQbmMsLGWPtB3+LmH20iSFDzj2Lr2YzOacBV4F2A61hLncbwCtgt0WG16
8IvrsOg7McGpMjQJi3JE0zthwebwgv/gS7Y8nT8z4vzuUOPV/+6Z/LhoQ1j1a8YZmexmhuarcBKm
sTLt5T2dgGegFoNzHiPOPfX+xrAdcxNgxqkAKQIP1wZIpciAVWTKmuW0ht+9265zYQwF3HlVnYmZ
PhnZA0pxsuipwP3f+0lSeECEitBAjmGXkomKHa++92SPQ3VV6BmVPQXrL4gGERQn3RuxhhYP5CY3
0FjX7lezCkZG/upy/YH3neWeWgzTOd3JTXAfUKB61mXMZCl6de4QvJ8vCvPegMn1oWLL+VAiEqLt
WvjXbAr8txFM6wYMNc3tGn33Ho8OOsn+zRpw9CHRB0xZox4BBWb/o13vXA2enQf24boTjrfrEKJR
/rtC0ZqSAEZIC19FkdbU8ZA7NDvJZBXOjmWDWVEceOyu1y9vr1do4erIJxUsEAdf50pDUfniUoOR
txcbvmCezI7gchjkeorBfhsON50o3yc9InQfsuIStHgHsE7c527AwAPABEdbvlINVwZAf1ovG1mc
43UXV7mRCLMBLMXxstBZHR/wfIxGNztHCwXF2iPrl/Fgd5PiWGyskgikqnAWn/xmaFU21p6YLygv
wUq+v01CwjAxY+pjKLiUdVEeslF16Uru9srTKU+UFlD1WxmG1Qcr9QW6REwv4cwWq9g1iEoBIr6e
2TqurO/9jn734g34IrCIU2YI+zCG5q5nUkVo4/h/9MYE0BOHtMb7pFI9wWJ/7U+icF7PnbSXzXjB
2RtgpQmuI72V9zd4+lkyJobdXrhovR27avdjOxiYw6tabSPImv14ms+CurhyBoOJW40pqqmRwxEg
wlIrGCsMDnz41KxJX+jrTbSrd/0gha8AY497rPheuR/b7mh7n1WHTOlIWErfsSPTwo6mDa0tdaLS
4xaKM2+PECsOCYm9JvwjZmgcXOdUZ22T5xUVHADJai+JvMIKp6y9TAXrc+oy0z1qP3xIMKodylSg
M9dPfM0j+6tY6YxaWRZxrhD8d8jyLATe98M8O0QW+MqCH6uA3ZvbiMYcOUFdr7beuKd89W4Ltz2g
iVLwcozQAkhyz0lhx16CGyaAaECjheBbI0Kd1Z5FOMdhew8dxbhY1qY07Zg/h9r5yzuC2Jx6y9DF
smCwowQ0gTAWmTalFL5RVJbgOGlTFcZvFpVKHr+yeeRrZXS7NRvDCwgkadfY610VH7HoQMv/YXT1
bROyRVI8o8QpEgrNlqAkA0HM6L/rpn7y0LfqO8nEIu0VZ/1spHIn9iAXGD95WeU2zy30d+0iR6H/
5id0dgnuzH22SSmOYF9iUh/Roj2i3ocXtlhTpRPdSFxVc/s6ghz6UxkGTr2yYRiWSuj+iho9xF6x
/8j2WvgCp8831gHlI6/iI+b241th7CNSh2rOs24GcQNcDGXRPEwZIw3zXXCXQ58t5MK0c0PvtkQd
VKei1qwd4+GtZSNrNSweAT4Sd9HTQj1huQYUXTp61wgPCS8hnGPvS5EOEzVJVM/b7Ln6gf7Tj41v
EB6FmeGqvr8/nqwS9dYMB0fpprk8ACo0dVjjgwTO/pn3qxM+G/QcuHAq03YraZaLZuwZZyqyPQlU
7Z6bVBtqLWJS8B4OpCwsJajWjP+7hRKHEyPOfHxOK9Xo9ZGZG5iG8W1UHsvMFCprSDErEmjhfdYX
uq1cZWXgm36alJEYVkFCTRVIxpWMohojmi8iGyuBnbXDdY/i1H9j4zCGjhfDSnWsAwMk6Zc4/3qH
NNed75VaHj7yw9MbPZzVBUwwR/esVzFydEYKHfMSKYEnhtRdu2GcWCGzBW4votO0rJslCi7P3Uq3
esIjzGGXUjwWpRh+Xj515aLTAqcMDWgT4IovgUG4OpmQVEKQh+26trgon++it+yngzyPEP5cjfMQ
GEK19BX0of0hpTFsc3KDP253nO7rrf7ybCzUqckwlsQltd5zRzO4Ut117+u/IIk575MrxFkb1QMD
a4wr1sy2aY/OsfkEtojkhFKhB/sBG66rr/6r550GYLPqpvIKNd+/oxtizoLFEw1uxqQM96+6ffWu
UEajXfCq0b9kWq8f4qkIyOS7FGq6TNNAFWG5fH0sNCr/7Zs+jl2D1W1noAT4gwCC+uOBzgXFGJ4+
ejGJRoYtVw4vcHlpxl2jS0G1hUUXmBWVEOib3OfwbagWgjuAPOO1TEmXTD/I5oDRxvhfWEMRc/gY
WCAPyxpb7K97NswuPRB0e8bUT7/TxWPdWwN3uYsNl1r0ZfF/t6uc+8c1gMHagbFacTrLBxnXNzN+
2y4Vqp+BPX6k3UzhEFuDQ0uKX12+L/ZNRC9AII5oGIanwN3v9H5e5+BiMnO7jWy8CwUpvAjkYMBO
7ueatEjBZO3IKYXSZmuWeojFQgTKLYKxu9lQEFgVN0L4SZCxH/IMvrMDnA+jeLi4zy4higRzj3AD
YsLPrV1U+YM1R3mMxNhM5QM+dJIldrZgsVIopaJqspVSQLXU4G6mpEbGZNDqNO1O4PWlw+cWqqcY
etFEXdYjk9DeNTnShfBb3zR3MYkihXA+18sWXSVIWGFYwdTCT752Cj/jWxGlxitQ8DX6KBd+SWs1
DevEVV1NpFJ78GTNFWu427fuUVoXzpA3+rlQsAldtaiPRgSPlAdVXVYjfT1SiwLrHed2cdgx5lrW
KlIJsNfp4+S7pjGU0Wo/9YA2eRr8ZmP601tel1jwzHjX2seOjqO4SyFsztcEnDzpBW9II1KH02hV
uDBBwOZN0JdnYkbBKSQRVAoqoy/joqxMENgjaVKUspiaJoQjl3p/5DV3mYfRF0F9l94d+qk2jxF9
APZVbDXhbK5bvlL6kfAAawHo9paLjz+zWEDzjmV/C2XWSRc8zRMG05lWt/ixklJzwDZfr6+aeb3t
yorEJa7Lg2urbTJ7eutmlw5Qv3caJsbaZZbvcKScKIPfccjeKjx9o0TwiGTbf0EV658da7qoYGlb
EZ88XR8+HOYfO3ozYD3FA75j4bqw+897qIZCZ+AIxiB7ZnG9w8d0mkqpX3gWHouUQiRECdr9SXOC
b6DPAZGeGiNgrEUFTorRZnA5mdKhsMn+BaZl847I8ND0dpq4hCvbmgzi/uloEjurL6pamJigewp6
RSmPye4EdjA6NB3JSk34ymPwkIttAb++Y7Df6gmigzEUQvuR0dAWTcgXBLmTiU28TuTBEfgD47ev
AjspMN6xjso7dp5Pkpoq5bUwN47sOU+e3FioGv3fct7bmDF3j3F0VAhrDYJB+M1xG8RFXdfJoawv
yQnutYxaPOXABiR6/okzIHkr4vZj2lEc4DqCe7KfCsaO2cVqg70pPs8lPIbhfSpg7K7gz50A2ljg
q723WzlZDZlI+/6BKsxFcPa29PF/pAeAt5AWd/+q3hJl19b8yQzIYn5h+VeoVxOYxHIUOaNqP2i7
gbhdGcnUVQASOtnS2aqPZkuYVpOfOYk7qTz3Nr4RSi2ysqB2al5qHBFp1Av5E/BQ0QzbEC3S7kad
T7iJa6IQD6Kal2uJYZrtFKteTBOfhVnxVXCNML/8aHrFdCYgtrErxG7O2eSfEP/zCrsmejuCcUsH
X3ZWym/ooBN4uTstMrZjcIvq9r6DRvYzoUAo4NQxuMsTUVkGRXyidgL4N9hJuDod7aBClVXmCK+k
NsDN3e2TTwBmcvM88ExuGyJG0RpWfKV+7yMg6gtIskLO1He+9lP/C4ApG7oqQHGjmTyTD1v2C8UC
PXWQ2hXb0FYx2SPsXQzjEZdRUvzCPsSDXtLl40e1GKoj9w+CwWGNhZEdpAoWR4tfU01v/HZHxBz0
IFiUKcbwddIgtayNhiyWlRvzv6+p+jFuge4L9omO8Lr/QRV7MKZppufXDM7UF1IAWMGAfyqJKX7q
hlVF64lYwz1I/ZKkuJe+k11mXIdJXoOZfamcjaLgP7UvSZlH5i/laaNVa2PDjgNleHqB/naxfRAs
RmpaCNtWiz/IccoovyDz6OkCNTpyMjC0huJPcNNbA+C7atZ3ZtZ1qwLkGD0P9/i4bR7dnmSiuR0u
NF6r700CSFI9uEUmJml2LlKShBNSx8eyN+PYVBMJQwYbvZ8FrN9l9utJSVHWKhBUydC6npAGuHA5
IDnnh8CjuTRp1ugCExROZiGpkK8s7BKnNYQYPvu22cV1NigdofmaiXkOq4FkD6bSN/QvW4kYJ10V
gKDXgBlCrQ/dPWjXVkLG51HKKcNrbpKnscUfH38XkoAM55f8xUJ3v+7o4LQ3EFuO4ZAZK3WUWJlQ
B3rsdxVbeUqrNtQqjHjd+vTGh8IDQPZ2ROh1LPvOu/zWaJ0uDUE85mq6S4t3Zuw3XEf+OkrTFzJi
b70jBye2PckhzZmLu+P/MZKMi673JgJ6+NE4mtV+e/BF6pWyHwWKMZTGDaeDNS0Gq+iGtVtKZ48G
nmgHybrEl8jgquOTo7GiaJ1X8m48F5C4ualyXhFACADQyX292HxMIT52G2l9WuNMFbU3GAwxXYXN
YtuERGk8jbtIf1eyJFX7p7T1vO/Y3uoEoIqqTugdmPT1QhE8HO5KPbu6cTOZEf1kFZnEbm+gZKGp
H9oziwVwsDM+MkmX6nJCZV4CASEWzZvXLCkXqc5ZW8f3N5h2zcUk4xqq+z1eCOHct5STpmam5HZS
uCn0VQkpoQOVfkIGGaH0M7Xb6iX6x+pGjC9X88e6H6WfJRFZ9OOLbV7VCOBLIsr8eXuXpaMx4XF7
naMpCpbXHzOMyuiE2ACjuosMRy0oN3u0wNZF+yBjnaI/lh7QsHHqFhMKR8iaOKWJ/9cHXpJRi1Qr
M2ZQb/u+JFgmI/Q1wUfS0qMh9OYB7yMS0pKYYhXKyyxLYRUazjxr1JBGFyZDEVNlRfp7OugUja8N
j2KhSFoXd4pcPbRvHZf18wRAXPirE8FWPQUuabk/Y79z9Oc9c93mYxMqMPoXFKGcq5DHaXmAXSYu
wK97O7xNE/7E4czz4coVkWNiCTxCfXTp1jdiRIX8ZFZlBkayKOcAcaihflqV+TMcmEyOROTq4TXm
5sPj3mi2NBSAQ6IcMIE0Y8G6Bm8Yxh91Kpt28GUtI4F66oeo1gHdLDcgU9eiujLUYVi7TIrnv8A+
mJ/zHLvTAvQCNOAgRkjt4Ril6EVzeYfioM3KkwkgSqYF67b63MqE/GYQv14IGFzP+H+wdVIXCIVI
WV+5fT6kmydtCN1BD6PYHU1MRVGSOzrW/E3TvsTHy0fHfkiktXmsJkN02qhouSwRviSrXSHqrqWH
/K5qGzy6cFpQnDsrfkuk5VFfXSk0C0OaGJowMZrgIHUd/yUDxZgrFTcm9z/7WWBiOabfo6E0MraS
7W6OuMVfgjiRFESsTTnqr50kRDMPcrxDYweSpNBeSmhX1z4gJouc+O/Tf/SKMggGe9Ozb50wR0ng
1tqKvTnMPwezcYo1cQeI3h3B2nNt1098sKveuqBl5RmRVMv4qf8cFyBlmV4VxxkqN+FTfkdpbcWS
R4vGTJgKfiT06R788FgXU65eBZozHdi1x4mVdBTQRfqHkjN5q3tjAN0MERIQyWndKaxavSSS8rkC
cG9OcrnNoF5ciOo9EfSivgx+hswdF97CM65GX/qg+c01ao/mNo/JCtwSD3jzlF6/Zb9idRWcLNNj
VOsR/xaQmgfEJVnle8Nm/zgaadBU4RKTg+Lxwcug3zsEKgDr4FBnTgMKZu3WmGenaqM2DtjDfHOo
LZ8CLo6PLk7r8QybGIrUOJuqYG5a3AQ70R9Ys7OWyCa98jUSoQ6yaV/7t5k6QOXxL/mgSBduA8+d
tLZb9kcYIp0lZ1OWrKL0qPvcvn9Y4pc6ys11ImX6f42TC8Y6PBFNJ8ntmZRHBoO9KnBPrOrz9iqf
NJfcimqBUxM9KuQ0UKeLwhSOrEckL2QhTwGpmocM5TP2kpjLfTPZJusDCphUjRt6ria0tLzFqLDO
9XFktTi+P4y44LGuCLZul5db37qNEGZ/sSUr8KQRhPhzOt3+oYyqFkoSh1Aj67LGtave//sOcwAE
HUBr1tBifQG6I62AP/cJxtXSEtpO1ojAsW/VCgjb8tLGvjvwelh/YahBQXXm6/hz9jM+vOpAKAzA
xfXd3eJpD2lrdHznzCH7Oms6Fgo8GUq2OMW5JdZcpWNUl5CTpIjzqK5Xr56fKsTMoUb7Rkrq425T
l8ZNBfp3TJRs9VboYbOD+UexcmRgq6bhXRCnRmHBn3/hwCgl3s6jlFNAeekvZfhhoLs9vUz4DlEw
kjIfF+/n8P/pQkxmORuCaImVv71Xq5fLCjWtLNyvG91G3qetkYenNRM/WTGS42/lHzDFSdv5PZkX
vpV0oN+mc2OnjnSGtErI4ofDd9zbvAD2G8cIXDczWch7JGycAeICPQiWdV3Ggi1Zq/0e8zB6h+lx
EHzOznfb01KN7KMjpCzWPA68Ki35nTb2XWUByDIrAGACwrae7SkWjQgtZ8XOjQsIfy0HQTgzPqsp
K0cJPF1/TBDkROyWtDp32lJrH2wF9eM2HDRIMCh0xYMEGwYr0f8AdGdJP2P5HhG1uygzeIwn0Sps
W8EvVI10ZRL8yG1cHLUrOyhS5fxP5RdClgy0wblpOTQvLIbY83pcoJ3p4xFPHw5sQetRa0Ct9P+t
lHRAMMrqH2FjxBgDWTdrZ/eXBjNeWIjZMTGVoAF9Mw3N9IfEXbdcp+d47tDlTxggHD9zcAU9rJrv
UdgGJdQNC3U3E05xLMElRrxZuUpw542tAG+4Gcsrf43/erotnUxTfMxhbFBOqFFhkd+p9cRIMCAy
/u4GJgxNdOfq09aTq4C4kvp6wqmp2ayMpLRbBNWMj7vyACTHN3GiTkmuFhVz0T4YJB2C0K+Tmz7r
HbyICwD/En+kbjrrjdetb0uEQotQ7qBmRYj0c9kXgmuvH/Lsv8Cvzb49pSGmRvh/a0QGBkqBdya+
/zbkN17tmM/HXIFZbrsgeRaq1iX1LaJLqg7ujX1ZED5xxccT+6xbisQNTqjQ2qozefsaRuuyunYl
hh4M3Bc0713ZgRkljQ0nYzmSZGADuOlwuneCwrBcNXMd0Mtmdjy1eWbLM/LX0FBhelKp+L9PfxMM
WYWlIt6NXy68D+tJDZNFRqmozua4kbnmHo5QRCnZeqllR7aLGi6o2ano+xAy2z+gjAF02E+jFQra
TzBEZ71oJbs1G5gWMgcSZ3ZCivKJ2mhSCpyIy6DfP8R1gl5Z2+cx4sCHspyZfOJMMPBMGhlGHvct
DBQGaIN2DR/YmUCGlYFgHhGqJ+4bSNfGXgwgVBE5OuMi5BEHcjBhb3k9RFGswtZ5TtA1uz6KrqxU
ZhBJBkD5mldX/yxBAFqV2lueZsxDCP4NpIS0N7in0i7FZFvUT/1b9RZGI5CLj+PP0CVkvZSJmrU1
Dw29Nf3H5OI3U3mD5s4vyZcJQtexsqSw2c0gHY2HKX7VdVtMvnMZ/gT+3+xQ0GsF8/M/fNuA4omL
Yt0xgxtUb4kZTeH1xzVDjTySbjJ40rHCyoDVCAHbwKw0DvSyupOGuYndWq6KXcBvmkeXu+iQ5bNe
kn3cofLhwrfk5crDxQdEqD3OG7q7SgmEW2Ew8zyWOdVLIzDCIkjwfI9R4/0Cn3sCpMIR6J3I1lnN
PmFHvJLDraLs/KBcnshR2CS25kVfsh7WY/OuGGmJwwFnfAt7KOpQNiXe9tsJGhfLPTIOUPlLxo53
UjMGQ6fGwD2ByC4rQbHCsoAVDWf1URbwQyoWyihxs6hPyTZMsnJscMTCBOjenVtwQv2rfrapQlFV
cgIpmy6ylqHsHZlTxnl0uyq6vIj/5IayfriTXZ+9d3dGXTX8L1nrO0guTT77L7pM5YtFB5HJrfb3
A3TSkAZsfHzaLJB3ja8ZsZqxKpzPOpneOr+6BZFcVEUabi0YCOfc/CNHVMeAXtIQPOXT+qMagpYl
NJloLXYLAmxZVm7F8EXAb2C/kInsepX8QG4p5dv6nOwXB7ZxQvHnAszpSYedAwqSawRFLiY9DtO6
v2xDi8kkZEnwbXE50JcOyQgicr1A7U2ASx7BoYpdJqM/0GAfD5MqpdzlP/xFbC0EZwjn6lOovyqD
bhv4Pa3X9dq0Oc5B5NV0R6zTc7vJb2pZN1xHLD/GjoKjoSX606WvbnVi5rP1aPx+4pG6ukmPa5bC
DNdFv1aFPzLjCLsAtKoSYI6/PSQCn/isEIOOh/tZ6HrdqXEvlF9q0V2538RDKwfNhsR1jGB2mgci
negZyvPvfgtaaGvQSNb9JvVrDWZInGRO4MPpthFMDbwIko9z7qfigGiBkNcRDH0tRMBtder0xm6z
7m3z4Qa084WV5KBx3Hwvc+inpUNkOFmTOCs6DJ4FwwI31M0in2/BBONajlKfmDfHDubwCIbd8bm5
8Auk1Y8APqyuaoJKlR6fYn4CypliknkE+V0EQACn+uCtNpa4SKiHr2Sevzba48K5o8A+f7uBJl2H
mKNDQ9Y5sXaHJLRD57jMo1CRXmlDiiGirli6TY8tP7eYFv3RoNhsYaqSck7R6ta/X6cwVZNSnxbA
LMnMp6Wz51el/usKYLID1B9QYIrhe4PBOqdOnz700xJlX9cT9yZVmY8kXz1j0hWsVcV6OWgDx9SI
HZq5eLptKZgNTiANqS1iYkir9y/eISdjaS2qwS7QO01Xa3d7GrJOdzAFIEiMoa5WDVXEKlR1Tr9u
b20MCO6GjtfAPPWEHFj6hlsXO87qBeKwPbvmx3gEzPC62dzFayBGhBsFz6R4WqvvatXMQRAEHdld
1ecdW4HJFhXyh28aJ7egRTyi56MghL5yBdfs5VU8KRMixMt0nu7p9o72x0RK1yj6tGlPZDGp2ynn
C9JVMOYffXxt4E31I9rssyVEyt7R2rD7AA4a0PKKzLaZ1k/pqd+PWQJHf/c1nKi0Co1m4EehjJaw
GzBwcriSRQSPjBeh0D+omBA2jVyYzgqrzw/jGA0KKd/sLULz57rHn5GA5z1fboq+Iw4+VQjhugdK
V9X2WfD2T8duL3yxNiHFx2HIHc0EKCzQ02AylQzRKbinbjdNnn9hEH8mxwGeAvC97DOx2XNV4TOm
/2d3517zC299Bhr08LDl4yIQBSnJ5sKTVyZIwRc3pafV8hmocbP7vzywAc9B3/RUAKiU+Revleg3
9WJH4vXO4n2EI29wx/D16nVf2xmgb28cWxOUCDbJA+VXUeCK+GZ/YtqK2zwAJWs7BbAF/54Tclq7
0VKCtQYKBq9xrvxidN72hTn196gKgoQhDHE9Fx6Rd+52I/CGsrZpkZWrKxMnJbEO84pR1KP1FQ3f
nHcaB0xCZ0FYwf21NQRtOBSchNYJbxDNsJWgXjMm8kFuhXYbHn2iFQvk8Y8hqZNbBYqOz8M/GkBm
jkhvlJBisLUVauuXZ8DCkrh/CDV5Bpf/ZQkBP5JDWAboBhm5URtp+Hai8ge+xz/tiuqn+INH3u49
4l4AKgTqvQS+FwLVQnrfhXPhOKPdx9UwpHVuUhhZ3F5258BWVCioe/pbJCrgYoH6vxn1xCTlH1fJ
Uuq4HGIYTA79GYcuYk6NBrKtg1xyGyFuYv1YkFt9o9xZCi5HeVLz6VQYqj8zOegyxOPI4mgmveny
9bo0H358i9qpCYycrmMKcYn1DuqDbEzskldwRQADV0mKVIdD+qjzN6qx9u279I1COyX/o8yXYDUA
73t31xlZDS6ZPPktb7yk2GmCZgkNCeYX6I9FE1BrUAQ6Y4taY7jfZcyKjsF6vP3h3qz8HmpKNZl1
4P7d+5lVDGW9csq0LsHZnpaoGRdPg8Wb+nYwyU1Jb4pR0NowaJTi2B85FGh5ABys0IAhO5ZXCr+p
+ZaCa9lqBIuIPb+9WMjJd9ko9onnFsVDlJ8pYtS/vfWyg3bnuOhFNb5YYAH2GensofkUkI7M3gI2
+RFzXj88gDnihdBQNOq7bWuR5m86QOyxJaVM62IQIyoznKYJvPuNOjISDpwsC+w3Ze4ybOhpuZxW
r0ENzRlypMi9+dCxlG50sjt1EXhrhjExnvYWE5RbotAwRuVMDe/q0ZOf8rOY+YA9yxc3QvKapl7z
lH5Ql0NLTycB1gkz34hKWbzUEjMAtoeYByODPCYRoG4FBPb/su94WmTDwsVlhWOAWgms1KZjXlyl
Sh48hSfjGmg+1+xT5LFqqXaqbklm8QSbELp/MgVrSsypGbiR8Xz6TSKDWYyMCHxVVoidEDGJT4ir
OoCgjKAmKP1qJSBv0xcuhGgTAYSFfTqXKjZF6cMJGy7gBHgnM1R4yvQ4+bHlowBKaZDopfySmIy5
4TiUWWhSVzUDH4Dw49hXLYhJ5zRe7VXYX9T7k3kQ7XN+8+wUydsR9uTCDJOePwoF5oy8+BSZe6Gt
Nxpf3pIIe8mGMtYYX4vFygO/fWN/LK8sk/gsd2znE83Yb+EC19Tkz53pYO1wW/NCawc9tmTytwEH
NVk9JyFIL3UAg0FwlbyNrEcgjSAQg027csvSWS4lVO/IXp8TjwqJ4FhuQakz/TM+4gGXsYIOgp7F
SWGXPSmcxrwBgPKpksctTxMkt5DZeX9fusnGQBkuJ/qEFhw+n0dwB4WoP7d1caFpzfWy786qDA9N
5BdcDPc7/T/MtOACiIyZ78qjzVprA40HeNxiinZVGFqxpmcD6OQ2OvGtmfC/GdvYJ/Fs9fJNC18X
sCHSabfEMV/8ppAeRdByab/82rohWoBf4eFEqh4ZKl9pVMP56TPL7wnWEMGR6kEnxOsnzENcisV1
7Wm3PPQzPpgE5AiugRgtZh7Td27X3AIrQcD1kY8UA1QP4emOH+sMA5VY0JYkb+uAfkh5ft55CWHV
zlEiDRNj48y9cEu7rhvZsukCof9TeqEDJodMe5v0EYeLT+dzhXbXNo5jElHjAc0p9M0MJnmDOlcG
ibs+O4p9uTTJnpas0SU4jIwox8MlEkQ5UoNSTUZrEzr7/gtIuMH+IpZrmYg1Fw3WYTe22UGSVOFP
kU0/HQgqNMk1z9qD1qdFwDjUtvEvNmxLcw3VZMaABZd+0p5IazbJQWcPla9uq+aLymn7c3T3rZyQ
RUnkoqKaKR+wgxMC1ILmisbervsOtJmKSyHhsuvHK/9oYINpzaWl0zOfneAE6o1IgZtI4oFWGjxT
l5FCSgEnnTHtIESe5aKM9/fp4OJ2DvRcOiZvibnY9ALs8Q7UDdWxIXOp/Den6Z5q1KKWF72+fn5c
rqFKqOlojtWlGj2yEff4Vvg2UbKr43IFF8UoDuCimIfUyKxB9ktMrD1zW5UHnSIPU8lwMtxzI5Qi
YyrF3ObikI3dzb/VPG+asFb6kw+aMUqmaJxJN3/qnttLe5QxNlHiSDL1Kkg9Zq9XcExPhf/PVkNp
o3JhygRqc8t+g6X50KRHkxBd6wbyiOFwn18rdv+XFzxXOJHlJiDUuuFoKMCZ6riiihsrH2hJFngT
Aq9PLU+tpyz8wwWxvNsiH+x2GRiguQpJoxDWu5k9qKX19Muhj3DTboDc/FcDYbJG7eqKAFU4zosK
dfqsERv9m5xnt/pwQTgeeTfpkSLdMWogPSxLoyZerDghaqB0+Vn6mYoplWCbi/ZXBF7G9nGwX7iG
UeT1Im62D/lfzKlYyoI3lp23VqASiEYZbHw5SSwxWnsTBiADvMw72SQHf+sDWUYnMNQFf6YofU+j
cmdSpwZDLiigwvcjV2EB/c//TCPFaaynHzXUKzcOJ+XJOwVlQoUWSWjozULM52Beskbm4RsUTvzy
/8xJJZ1qgiBu15gWnks3xhlBLKYoehWn1M5trQtgiZzBZDIbNkA8nkbf8DyruIu+g73410iI8tf5
FaP7bE7yMKxG3pFqZMyqMnhRPSP1OAPnN6OVuTfoviK9OgDSBDBdhRCljpjQUo8RqBDhkfFWfatI
49pxXyP7UzJbpkyUKweBK1UEFfuznxiuBhfNFr5fy+S8L4gebVvSf7xPV+ihiFKb+tGKadO/aR3Q
yLAtSYhNIbOrfVIc3DNl3Gin8NbTWRt5L9FYGhJkS2Qwyk4sttNc2m2dvIQNVlheIMIjX0VIUbKI
iVU82tfb7tL6LxzQuSdxRQq6pfHjU7KlEscz1ApEciwqEMnsqd/Cvz3z06Qap+pzXrt6VsXZvn6p
9i6QdSQXWL9xKQsc/1Na0tBwdTOJn11Y1m8Aca13Y9C3EXfB4Yz4nYOsaKou6+8uqMLeDE5ssvWM
iVjMlB+DEo3i1oDcuDt7flioGgp9Hg3PNk353O1r3aoxUcRHCi/46CHt6hv7iDe8TWkFImdI1wjA
VRjhJwIcvqCSW8spXEfgiTAGLz/6mrokOfLLBdXXUUuyfUk2fJkJuDHz5+FIGKoo8lKyzBUi/mLa
CHNUqPZxixoOmMkAuRhFyGKJpwpaOVCj+xP0NCbeMN8IjB/bAKL2WMniIZhmwHWaSaYmNxeWRNNy
KQ/HNjywvbSBr6x4XjoU+QX0tOQsR0bAq0sRtunZ2fOPDZcnc1hcl4QeoKPeArKtEu6LdqeWDEBz
eDqjJEfId1dGo76jL/gi3lqPZnEm/s1TIq3cx4T0QkTB6tfoTCqlom8Xw0i2m4PmRIy+GxjrRi3f
6mbnJT+1ssjcFEqmC74LrWfTsSDoFKw5Z0NsU2m67pqUbaQXPW7wHRS3aDYOK4yKK3uUxLAK5pcM
75jUY/2LrLUOUrp2hBYF1heo2mtWeA7hNfdknHKVI/JPtswn7uRgUogqLbqm4acDDx+jaC7r9k4z
W7fOG4aK7P2jwTafHjmclkaAP3lIbYw8kTC1DQQcqWeOyNx3RpZYx4ARw3BBWMqtbpa9vInzMrZ4
Oro4W6kYXpIx56HaaUrjisumcvd8WNzsxQIoXW1frT8wwnUxCUcyPHltm5ybb4NFZVmaBwAlAlLX
dYnmvr053Pm3tGH4idn6I3ep9NZdfZoATNm4lkBCybTEegmQL0THwsKSkPN/kaiJF17obrtMODCg
HQt2WvhDldMJRTTumYrueITsLf1aX7N/Ea3+c6LouQ50H1kIvnAF8YzTeUdnhfDJn3DACrNcqqu9
Ati3wMQOPamBfuMyvh3lMvngZgDcthjK5NOv0tBKXNDR2Jlzmm2zfdJzmE3pA/n01Pn1hcuvI31A
PXjeUX/Mw7rqNSWBilleJhUCvQY7TzDBo/71fNKv995wdB95240NV4pnY8eZJoWi/45MKCO1S2yA
TW65/29ouZeo4aRrP/koSQSKYpLt9Qxo9k1YJMfrBMnZNIVL30tJexHBRiump/4sEPmhwZ/c5AjV
Vsko5lFu91QTkRLUwIVfFE57d5juNUZx+47H+HqILRDx0/KnHSfjUuPm31ZQQ7MD4ooT2IbYCUSB
pNZgCsDpJWshOo8eXIN/DCAwDPO0pr52U/P2ZJEm6rmjio6tJNxpuI7/DhzAuoq6B8IRsyMG5tiY
C/KIudphpukjPvOaHJND+OSsyqdxC+a2sBBeBspg8YZb4UPRzLyV4tPYmP+EMZEmo5pXk4oPur3z
7jZhE0qexbbm6JuloEAQ2bSx3tFEUIV/Z2+pIR6Ca27aNGBr1vlNISmnOZtHqI9T71CVkpyQsCqL
pvKjt30MhRbO10+saHR0eR1ExhhYbXOyD8+1+WAFT3wBrfAnftV3km1b1NKkeVyfxwHTNdwqM1Ld
zWL5/+C3cGRWFrFEzAF4VtzZPAzvvNfrmZ27K1Iy2Yd1zeMSkTqivzjlMzkhgd6g1CYbzuN33H3C
y9S9Kj+SgmZPm4D3kY9x/Q9isWQeecQzCfP3GOt7Wn6cJWzpx7Xyybx5PNETIBlxQXtOMiIgHPs8
JX5/G3VCjEsIyz7nv4k5DdZz2S/MPWTOYTAmc2LUoCL9/73A+L1PT99CNyygzPZ32Kp7yDlCaPoC
03wycCmb3bo269MtrvCscduJTyRwrVcSQ7+oZejV3gUrXon7bh1D/+tKBnlqVq0kFjFtQOpXXJX2
kDXunz0aITwHopsD+cZ1wM4IvdPOiJeL0PUUh2YT+W2DtXcpycMq7uZ2UvSDKe41/gEPlEQmO5NF
zzegKDRMYnGW7mo5nXMfvkjYwlj8Wj6SV0qk79qPPSVjMCifGCHgvOTj584T3tljNyRV8no4rHCe
VaHMnZS+Ob//1T2dDmHSec1Yy69s2lq6MT8LlMUbLqWxrvo1tARkwFMYHWe94AFUnuYho6owMiVH
L4x8xebTSIOixquE5fzwILyvblFB8aJ2fPxjTMtMVgQO5ejtUagUHvlsjloqKvWnftWa8VKKC5VV
V2cGvGN7HpAIoquzeS9vT7IX4pklWixZkE5I5ktSwtcOYFl9RINMT3J1HJbNYp16f0ZMXz/Xy8bR
QAT/HihjQoDjyfDgntGPw3Yr8ilPwDUnh8cXrUUcBffI06rcmfmAnCjY7USUZobE1V6qDvEMyGQF
4FU8r3RxEzLpofguVNr+3DyP019CSQWQQI64jXxuVtwAcdHg3HjBCtYZXtrWaxr0Mx87rIUf2O/a
GWcEtp+JZ7r8/xH/FsHVBnmuxCtysLP9j2qX78FM96BVSS9oe/DixUAntbV6hrdvbTJJTEVGd8my
2dZ6GfY9uyu7mm9ycKjKGgJY1mRzoAeSWvImqXapQOCpi+o2+B+adsxQpKxfHacSaLpgbdlxXsC2
JW3d53J6YALEbdp8HPXSpbQVGV7jUB/m55bV9DbQT2dAboWqUKKrUGTyNFr8TYQftPZnP6TDn0ZD
Omdzlh1AqLn8XKz/8SQRDftmeOOic5F06zRiw/1QXilc4RlnFkrWPo+kHh6qUPQYjh+CQSLEZOVt
l6pIPUJgSn+QcMVlo9U2VFky3a1jxyENXycS57Xi9fm2S17DPLMXBdw1Y2hGvgtZvn1vnKuwdJJo
0fWVvqJEG0YkNdVeYomkvKkSR0IdoaRVVNLjaXPSdkK0XhB+aptk3EoyDA7XA3/bhqE586ZiNxrJ
WZwge+yM8IYSRahnR98UskvTmh6gXqoOoEttQoVKOtEYlPI19RcSi0Lv43lkM5xonjI4TLBopFf+
24uBvSk7zB2huue+nrZoxlWjJQPAUknP/cZoe9ty9wMpyyF3Eqmj6wtBrFRkm+029a/MD2HsCd3b
XxFcF2imoU+V7K7dxzBz9xnWz76ubv+ARc/63Mta9MEC2pa8U9HdzewuV+EzNXd+hK8gVL8pnGQc
K54rmZ7v96eLk8kT2JHjxVkdSsAn1Yz2GeRFJGQiSlJjDzM+0/fCz6BZkXUGgsR2dej7IWVSO3TB
gyBxJSz4LIXy8kJAyful+vEQFzFXwPWFwBjvb9hd1uVR/kCv2Zl8yTL0VNYNlzqpCW/jgSq97/8c
Nkh2olHNLcbSqXBXUUWcSL90/fUqUsW0QlgmOUIGKBL7xnHaADeV09s9FpFW9BzYxhrboPnYzveK
j7s61IQxCfZqO88yFPlaDinqWJ5U1VfkxiRZkn/8fQP5GcbTlBdOzgckscQ2FodJe7Md8kum9bZC
85iQ6bjzoBmlbwv2UqWlbTek7tbu0YDILtrj2desTFze2rRCvqp5dVXNHoDXYKdF+2FSYNxIaTyi
//WL29X3i6mbA6G1srM60KkDvco8p2VIF8LHAJ4MhL/MxyVN2k9V15Le3SNnRnFUa9Owo9WaC6JR
3orUruR47x8krcPxM0Lk0tVxt01g+fDVznaW76vo2Z1WN24lzEt5XHzm9RyEoQ131fPJTCqVdqgZ
8qyUY+nDWUqCKwF+hMoE5ez68KhcrxOyq5VRjl3od1c6meRWYWVZIICOIuPB+m17EuzDp3rhvNnU
qjtvzZ+rMXKP6zI2I0oboUG3uStdbYAJVEn2KJdVAOVSFpszZ17+6Emq9XMVcGKP4oDp2/zQYyO/
q8GUHtC0BUEXVMLgE2GkqyBdzDUkUnakWImzMsKL4YEryEwvKout92FVZ+4/CbW7SMy7FCRlDF8H
sRu40zJ5oiMaga71sxSr4ZlrSMrnECL3qyUfqbXrsnxBQyxRX1XTyiV3IU32pbpuq7V3D3v0YomT
rXG4AnczcnRrBz4Npous+vYrnpHvRsMJ/A0EYftXNU67aOkbejAwZlBaPkPg3+wRtYhyZwL+Gmfx
mALCetGEYCiPxcsGJ2odFNqgIIoOjkOWKssV1TFTs6GpGU2Ch8OSlayTfr8yEzzfN8Kwz/dGATy9
ukuesvzOmpu2P0zqE7GITELZaPL3+SWIUjiIp37UVpC3E4uRk3WZjerNxMlA/awcFc11L4u949dj
2iNjuxtx9a7YMtMPsv9s/vGnrzrSiwStFM+8AEaKitmQphqqz43GWELLz/eVGF+HVdvCW7yZQ3T7
Li01tS9SEHZme3OY+IdLtkuqMdsdsml3cw2KIMt0tlSclFqo4vVWoErq1D6kzSc50BtQAkw16rSd
c9AcArWAn3E14MBaMtJ2YG2ALWy9Fx+/eXv+5qU8U7VTJweqNSxSS2S1l2F/KrlwonbZxOQH2fiR
djYHDMiGMfWGmvgQWxM2YRWVTegaKckgEYFOwl5ejPdBSGiD19EZNr0U6EedPxQuqoXtTwPoiG/d
bE1R1pUW23XpJhmI5HjSr/3TJDvaCg+q1B/vYC76dqs3gSUX1SMhsQRiPTYvTnWbPoRUJCJbXPhX
WhmH7A2VxXrhInokuwqB6+sJDqiyxAoQ5FwmfbCV4dFXpUgZYncNGh/m9nlXT1GU3m+rgPLAt7Nn
iEwAOcuK95xKv0vev7Zb0lHpXA90Na3IbC51vHkrV+FkbdpaW9FjJLxWqtv4mm8r184S3BrHeTNU
lzJ1Lb+y2iAg/x09I9EQItQ5yhffCzTiiviYJbDknLRijpTGRGcTXEK7fZlUUMTlezvmAtC+/seS
VfoPX82xzcmAEVT/c1bY32mIyz0Ok4s/r5bbBZtEOvRIwxaDcJRldvOkGhyNRMxb136t7SPF2joP
ukXUsnjT/XUtqh53eBkuyIN+Gs8/XQwyBWHEIGXv5WExeIcJ8bsIOnUXoyLJe4hfptfBQKmGtxCw
Qz3eHCikV3GdyMxnWOT9szPFcHryig08Makk2+48GZCh2acT66zgVqEFMbiFoB4zDqkm3Jc4OVk4
rLKf0tmXcelIzdhLahI7JGjdPlc0n2p3nI+X1l1VmiQ7TnX2DVxBb3Xw7TQEYLkA1cQrY2MWpOoR
rCH1tDzSVCg/v9rO2zUV0OOTRtwqw8tqQZGsWQczM/wd+sGoWoZkn0h3UYbh2q2/ucTwzL0aBhgS
wgNkQ/sX/bEDrpvRnEAq69Lj3QSrjg9Pgx/IPHKXTGHXRYbanQiMb1x9pcM3C/opIhriIcYf+Iz+
tfnE/QovHY+B3XUEwF3GoQL44o1DdyNN2+Pxt/lXaeEVrBNfrmVrCokdIJ+xvregzfMJNvZaAYsw
cEAOq6XMRyZqHwfU2umEEM1JaEJt0mwi+N9jzOUW3h8K0+o67I1FDhtxZqA6XdlV/0dQlv1hp/GZ
NGXU4OzP2nEOa2yxyaar6t2Mtrh5+Nk5dEnV2IeaFZmfIW6UlFy5JHdgs0ytupJZkYVr0LWeecKS
rtLPBtc8yyf1kT8o19NyCNMMGrX/FePv1tVxgDpdNUtGIvEtHqJm5RhYip2N7WogljQcEr3m1RAI
qqpPtSj+4KBbUw6d3D0FOhX3LB48lzGmYVGJTrY+VJhFV64YuknUNCWNr7Uqi/6tIC7vgR7zUfcX
LarIWZ2mRfxfxyQRNoWSsjuK7nLDALAMT8AcOab5gmZu/kUjJ4qOi9GdVweTStExTHR0p6jXLU4Z
/zN2GzNfIRBGOhCdPDUsF56sG7u67W/yPvPmfLHkPFmZB70X6Ue02W484od+L64RplNl7BdH6PV6
ujtVYVxy4N1dJHFwrQJ2C3JilSw8uSUHa2SQJOk5N6WTZQKgmzKnsh1/suv9FU9YFaKjHHUj7mv0
ZMAS+7xNLrFlN8qjchQ8Xyo2xbiC/aJWBfSlpZcrpm3urg3n0vehLZREIflNcfrIZv9XvhqkKzby
0d5qu5Nm+i4AkqmqAnnGEf9OhdV5IIk7IiZsq1L/HFpeQpTw/YU1R9H1wJUMPRwSEbp7YI6iU25z
uo2HQGdANnQwsE1Njm9XUbD5cKLrS90RIAE5/7VNQxux/Xl0Wu2+3TTXE92gYy3pyeuIy7QG4JDN
RSwy4oaNapSlhoUcKLX4kXh9XySaYORQDo2v0Eh95rFFrwIwLnYfmlMJ/oUCp5eVGXER2x96VIJn
gkj+7R0ydKny9z9IEcMoznCd4842xlThtY6huZgXQDIaXvkwDvcVGIn3BGzx+qtM+OMP+BHz6dry
ZnDBAIHtI3Xeithf3VuCF3mkeTmmqAXX/lYmJ8HN9gT3daZWNEuaeZbVVeGQwuNjSG5pd6xab9Ca
y80JDwj9r7cfxf1c/GzpACt3cfKD+1lLe4Ck1TMQ+LCvff0id9svrwH9RDqo8TyBUh3/zUnzHEQr
S+6qlyGyXfFM894Yc9YykPFVEufsmd3zlYYX+ZJlMP04YXX2Rv8uXlk9mTNiGlI+uCsdxVsixxWa
nzdRafV4Dya6Tw3Lk0kK/caA4cFv5dCK8XF7CV1vghRuYyEyFK5W4jeF7gyfXQzrFtgdEW8Gog3B
2BpzlPID0ssMeW86eqFUi5Ogaz76cLkBpKw6w2uB1BMoojr/w0WHxenLZAHpt902gwEpznPAlpra
B9QxOCTn2qm4vkEhpHCCUok9nYgp9LEc3ZAVKNpnX3xa0gBZ4wxU8ZxGEbc1MCyHXpj2xmOFkDcD
S6fbytY1CM8E+/dkpccPkbklK9ernJiPO2NHwIOSewnHroENiuCH3O3gdZaGzKdyztZyf4h1GUBn
BIDLYK9BY4X2E/owbc/8vB9wqjGFTor6t8EoT0P/NNYNEHHvb/asTb0/VnDszbPVUepb06a6090f
HfHkl07fID7zh9eQ48cXaUnJZhCUA3JqY9x5egdu90TsId799MosfGuWZ7HgFsvMdNAeAIdcHDKP
msQTcQJvmMVdAlzxRVdXQhxuxBCGjccQhVjjZOdbusT+qotvVYOzdJ3kdZhCDzHjwOMsiMj2XO3o
IIklkiSasoCqMKptKy/alt7d+M5vQzcDOct9fF1Ppa9i3tFSyaSritNE4Z41E5FPtDif4qxxjA8r
ZVedsfKR5anCiq9+jOjICLJ2TkCBqfa44fXpZwbPXVXhr6LACv/ixMlFalMEDAhbjEljxfQMn1Z7
tkTv9Y/pYepXGOxxAkob7WXXxPrUTtXxjR4uq1vjA8dGplXZzi3PPMOrma9vHEQH+iHM7nvqlxnE
A8OEoGyaJV26PnN1XbAWAPDQYgyISQvY186ZE6MrsVsxBr91knBUeGHWjV6RANBROzcuR/LSXgDW
TSRk/wyTcQgMToVYQOS9k279CXFcFT6z2+hZHvXABnmK/9whKQMowHfK2u4f7cLdaNeidyxwqstr
gwE4NVOz3BYQok/cLWq3PvJS6IwnMQPuHoYgPj+GEdZxMk5KFge1//JLEcz0AtURM1Rp9OZFeQYo
8uqVQsbumFjORRSsw296WdXTiMeMnGpATB7h/Yzwh27EndDBzA2XsrjxfixunF5zlv5vJNFKiYdx
/NUFb5iQROGqLzexeR4REy6f5ZTBrbQ3nbQiq+xltQYPad26+HlKCF02/kkzkxsViTekPdFNEbB7
ED/bXmpyjTOSPA4/i3G89B/8NVkSxKvPhy2jy6Qf9aiOQWwgDDzoBXqQcVn2kAtod40FRQRDZ2ON
Y5GCwY5NqqXz+cSb/wjuGRdKhYpR5nc94Ik/AiObm2lMY7YrTAoMvNh88KWZnzKmUBBKWlz30u3M
a+X1A56bkv6wT9DpkRtzm0IVpWVfvGl0U7EyTmpS71Imd7XyJlwGZ3Ir232pDOZCkjyfQXgZaRBK
ItXOxGr2goprpJyBmum60N1lps+XAxNLViZlJaqbkDr2yBUNxAGP5NqJ3kmC37Aur0VLDsRDpJuZ
iiXAXvPNDC2cWFtUFVZXHNlvHmvns1E47BUbMxtZp1whMMz7ulY/RN6PCvtBCWKFBoGuEXmGBAx/
6sj6JjJyefS+hbe6XjIDP++mEIJVOZsGnTgQpk0qh2lm+JOyiMIpVJ59FRVBf8B7UrdEu2pzHXa3
tYCBXtPRtjGzJs6YKgXy1mAoGBBjK4wpW+Prkc9K71BTVlhRSVEoMrAwRtFuM+G/TOES8B+uIYUO
sAav6PKccsKqy2FJ1LECH1PZe7vslGhXmyMuX6jt/l/GjazPqXBk4y60TDK9bFR6UoxDooDsv94v
p0/AWWJ6B1FQHzH2CVV3NRXh/vVBADHjapXzlwHZAiMJhBsv/pU2nDsMnco8gXRoxfC6u06ucYBc
VFp0WYAxzsViJ2LMxtkcMxSdxzBCUpVsHAizh33LMaTu4ESbyQ6P1oXMEOOppHPvDvhATvtcguSd
VPn5rWoWzXWfjsoE0ETVi6bLIKcS8VyoBfzEvem9fIAaT6PI/wuvAVDwQ6D7yMf4cglApgXOweO1
/jm40UHmeV7Ea09IHCBgcs5WPbmWtQIB06VKH1nNgrQ2dY1wYa8xISLZtNYnh0S2zNVlsEWYaOgd
ixo0fsOtMIX0VpnvNIDkno1kegiqKi12GO8bTVHVA88p1b9CTGZFdRThJIUxwMdCX0S+p6UIXqs/
lQqpqMnPjj25JOs0NetiY1h/nwEPtQ7BRL7twMU1U+WIYoV3fVO3jwuALiQ2PnxR2KL83fTFAxER
6VLvLALrDKCVDxvNiHF8xRUGSuyO8N3EMVJIEfz75gmDRzSykYAHAF1d0WVNHS2c09zzQlwvooIK
kRFefcQ5YO+WPvpKrxjBEGQi1Ry8FGyIxrTB1iRMkMno8fUkadQZ9cFUTW/f509PGCACqEpYMTo+
vW3f4fsmuLWYWaD67+0jPZDTqq0a3z3B1cC0TSflDxBGb0J2ikF5uNMZyiFQ1d4kfiAdqiK/cw6X
3jee6znzCXGRUs6DTl7Jl9K6jtAMlkD++b0V2uypwoekkka5u0aALXbg+69FpWIK9JioDhRiS/Ke
Dk7K70tjash/Qh5RfgI6UPr3ZD5XnbwWaR6Tn2ZcRfluzSuH9xWyD5iz+FAOv92ARZ6X/EyTDZ69
o14AWIRy4hnJtsGFHFMF0QCA4D9Ooieox5ld2cP6IzSz8fcSfT6PsNm+IUfHQ6qBOj/LJYwNdEZ3
2MXDTr/pWN0iI8VPuxHDcz16YQGjDYu87y/68jYthiDxBRN8HdGzguUTxEQpek9KYCuPIT1M36Pn
nP9wz11bv9EXkBXtqObGHsg4YRGYIOuCWRQgvagkA8N872MYVstyQJtK5EaYRXg6eHZYJPDmDI/u
RckE9Gd6SPgRkXYtFQYeTebCJTf2dsOgLvLUjnqjChEYQ7aX6frZsG2SYIxX9KFh6kFIhTq9vUFQ
kkqrKtyPZoz5b6o6XTOgird9o/EtFm779JuZfcQAuPqy9N/mQbjsmvih48eWK3GN1an6m+axJw9a
eJDnk4JNS0DuWrZbSAOkDXFM7OIdaqHjSR25vIXvcfvorWGD2tGREx9g7d1CtwvJ+vQOz57ysrj1
iKhI3KxEepDN4HBs/2XuvjVV3VjDdG1SbNF3DzrTL5oLx1KPt1CCDL24MMB+NLhgnVDwhbR8Luih
Ayj//MFhuck9E845+3gxxc2CKBf12VY9Y/fdYinMEe9XiyX9+0Gt1TNK1uanpndooWGv1kXvM3Ct
U0I8iSAHvQCSVUliU0wkHcPFeRr1wnw2ssg+JR45/3v2qe8wxy+iNlEM0VufPPw9lC1IBtL74WmI
RpYARTH8mQGs8Mo0NggpVkgWQgOHTYuC4bmzEM6mq0UTPBiyxutTdbkBT2EX8SvE0KBBC4kDeSo2
j8Ghuk4qzAqO/0hSn5xHn12ASMFFFn6cuRJowxsNwKWf7ZmOeecTlKz2FJyqkIIOtu1hL5OtGh8t
v3sfwl7Y7P66bIuk1l0WZhBzBI9RhMVTN+mD6JasG9eZaIo/vlno1oQ6qGPUtPQVpUCVLBnR/+hr
Yny6SeQ1N1EzeoARtpagnPMtPPDsom139hL5MXMI9d/6WauKRF/BbFlWZ+ElDs/a0zuIhSZTk8GF
w8i0L2DsXga2tSvggPz1qtM9ots9uOp/RvMtNimDdnME5l7H+ZoeploD3+QeSC7FnGNUvRAAtw/W
Z993LWOPoCSXSgCJTdAaqp6PPIFjkVjoRWNoWNv7hEHCPe8rS5/eDaYxrNvFjzi+5jvxBFLhaleG
JIbGVRF60qbdkacwHKO/YRU7h9vGZ9XHTn28Yp3+IzeXOwdTXkQ3NDVr+PSru+3vaKb+DE8fo/du
76XSEPjCK/j4oohhwBCnYZDKxay9KBv8vD1dJLXJ5CF7oWqeikNutBAGCpN3G72EcO07q2xJ0Uud
sZaGTkPCiMeunpkQg/5ES7vg7rKKdYrI6JLbVIoJbhz5nfNLENbgUqieQj1Alx1hRn9+gi1mtyT6
mmSfk0XeYOofwT9y7XdOM9Zl/2hzq4668GHM9bdM52UokWwtcjDs1iXl8ibWC4h++qPOdjgNhTXR
ENrO1SXpFhgNgFbN0CwSJqvXTsYoGZNAJjEJqGpytyX3wbpq9rknQNUCUUuOMkecPl8XGRnjp5dO
rDtu1JX5qvLeECCNm4r8k3I0lVH76iJ5IWetXmI4qNetjBQSevLMI8W2HchKY534Lh3eigGs3z1v
R9vtX7PVZWwYHGn0Zzh/04T3aENb5IpnPrdgYpuWFzaEF3HcL63Yu4OFjaS3aWQR0iBENxaG0xJw
v7XwXPaKu+vU3yiWCt/JEsFJP1GOzGEyyUd5jTEpW1p2M1qyygB7JEYAKn/21AeYLBRBdygcDFJb
RvX54TgOtVm9H1miE02G0AbuxXLnA1Plt2sVddmHCgChLfw7+i0Lr4tpfOz/Ae6z5L0FiixpfOQL
mSdjdVS2d6WH+9lZ6vpmby1V8rzzTP+WtePcXS7YdUxMdK6yrJzAYVYN8lecltEy98031iH9mbtk
ph14TlfR7uplPgzQiuoSqoFLQVPxruoP9gcnE8M4NUg0X6tKCRanEmH/n27YJyFagDsyee8idyga
EYe2eZ4U8NK33KxkqiMSDBGf621WIW/L5Fgfimt7Ka5mz0kGonaStLpurFP3dj88SULLvSeghV9O
ZOmCEJYSqW8LX98Zfw4EYe/Su83X9fLdninIOY3DzBxgMkIAJr2ErmGL9wNXIaGim4IR83MymE02
dqQY6qJq2GX83dz/PD/69LwUczvsTECuoFWVsY4dXD4SK+pX9Axk2cw2F2wO/jAxn/O+DrVDaG3w
8i6AOwiEsQa8EWoHNEY5FGmTXinvKvFg+Cb+70CDjrk+XT6DnzSAXlP/9S0JEXv2CIMQjiosyhc9
yN1gmCXx0K8tZneA+dN1kF4pPG7wVbkw6a/jH1ud4I82mn7dOF4YYDI41LU+A5MQrJTpMS2lwFVh
i8awHZt6yiMp5PjGSYd4UY2xrcEsLTg3VL2x3xSr+1+PsSJ3xFcvozyeTcWYJk7WprCXBRdkO/x6
h4VO6xt0koABabR3STqskghqIMg2qJ9kpRSEu0zB1RXvq3KVegv3wH2THVxGwWNLpUCqEKkO8+LG
vhhiwdPBoESKiHroejolR+Fd/NCMLH9y5XXpPnfLyN3+p1YC4VaFvHXBR1/7zZttyuH4XkaMBiNN
3vJ6I3Jjqejsn0x+Io37QZ2nPrSgYntxljnMdEja2Wyiw/sbDrxg0Pc4PpryKdYr5fYLIJwO1XHJ
Kh9YEJTovRPCgo9b9b0dilT3VWerHGvQKJM4uNbkuj0rptDBz9q2M/EnCy8v7NhoVUSUSxTjGBSS
NXNazoqkUuKQeQvNJPCQY9CCUVV9vTypFyunJ7hck3ys2lPoZnuSQWCi7+4DMvwmvs3KEeSSv+Jx
LWTCxLnTniGPTxlN3t4mt5WqOuDTBc5V+y/i6JD+GF3idWdN1fmQtH0G/wsbt0PGEW5YA+rpYfpG
eQ/eapr/Rv7TMzOw4sOzbMhLhkfcsKWfRPD85wMsDx3i8IX/WfnlOsPPe3KsDaivAON9V3byUVOl
RCHwJatXWivNvRzzSIICUQFOWJR8glOi2MPy1B8a6HHtIn/Vfo5mLzr/9j33A3uBI1rWqoh/UBp/
6xiYGhAqrWkvk0rdroBHaBQaeAhUFcjuAu0oj5wySasIcK34MBHf5Zz7aIyTKiL0jveAz1XNPbvm
D9VzpPLKev3C47rCNJYsm9GPNnvySr+XMkkiAmyG46ujJbDu/6Vtgkf6rjO24Szn19udlGOq43sn
0TwVyDXFRE5whPC0Zr1BmqjnMcPVBy8tjfLdur1yemHqoi8n4YhqgNjT2l0s+gVTdCoY/p9Gy/TG
GVHZLwgJc20gAnV7DTbS25MMN8Kuw5Y3dCBp4H4KCHQZJlI9hp0uB6xHEBmVsoJmwlhBoU72oz7c
RTpOCaXWHX/lVs4ZKcrk5cKvV+ZCGXUh2kqbYDitwv4v7HphQ7OiQLYn1VKk9UwnjWkE4viZvlBM
dF2ouGrSviturTFw/my4UfNc80G/y9ny4pZeN7WPpWNq8UY2GeqlhG/Pd2azRWYFFznCTjzX41+T
Y30V3YXFRYme639NwIcAMsEk6FwNZ/DtlFXs4OaQQeixOLxan88pZNEOEAs3NozCjeruevpZA6Nz
j8PEaMYqEpTKMBMfHHAIaK/mGprTJr6Ow6PDx3a6rm+Q3DCW9rfOFHOcLhn7wdtlyXTi0jKx9m9G
R0UcxrJp8TWa3VQ+l1F9hxkNr8WNUmdqZbatn/mMZysvuZyC+2Ojo5BbyoQBO8//hAeNHqeHfydv
ORJV87vtZsu+TimxbF1bwkZT9zg/oiENXvZ+f356j9ZokMybQECciD7cav+k39/L+3MCBNq6BZWw
tX1Q0a3JkEnwYZVWHTS50zYHGBAVkshV3IJlsEXbAJqY6mohWvZGbzqDwdatOtWVwvrG5g/3GfsC
OaUY47LabyiWnRuO2KXy7yb5WePGu+jFTwLQ5M7qXjVOn+/6AphUulpSmx00zKSuUUERFcrZTrBD
8VOnx7TeqT80GVgVJKza5mYMvwor+bzWvPY17E2suowGw7J8nRoN3re/WjE/ertxlii512/Cs33W
sc0XFzuKlLvQZMlJ5Xk3XR/fhJFZN0iqvwXwgeAIZr7AqKbm2ziyow99dviHLWgAEB/0rfBzx8+W
d3jV+VwmR8t9K1zA72FAYLW9blyDLiUeH5rWapSqXi3T5Zqosk1QFNacAmGxCYrBViQzyQZcsIDa
KcCesxZZFjSwg6G5R8PRa87qdLsy3dJ1MO/ZLKgqqZdcxyIbsUaEl68PhpYHg2AJrGTmBge/hVWM
hyQ0cp6ev+cAWyu88v5zjjpe9GDAGXMqIcYNqnw6k61+ETVlXTWw7Nm4aq2SD+pp0qktE44mwYE4
5hMqg68VvUdmZ5I2SSosxSvcEtpimCmYuR2vYfrC/tO6qP08zyS6tkXRLTbXGqEoFsQtW8SQDecR
TVSLzqIW6Hl5UD8At4znzxqkQf6cgHiPWvyWYnBL4lSw4pvwX6w7j16hdqbI/j1c6wtKtM7zC7eL
8fU9X3EKwcAhygcSK5Ze0wsMs9CRj6nDlZmvUV96Ag1UOHnoPBTWxqqR1YtrmJNrLXhMrgoi2KJV
3aTRuOyUzkpZubVby2z8kw0W3M6KQ8hoPY70NoF6HTWMqdone8xEezVq3IZXTr7vivTA1d60qKCW
nyomtEAQryrTO50Dr323xlTz4VeV04tlN3hJ9GQJrxAcAl3PRnMUAaGRbcofbsFOGmJ07T9q4+KB
uHGG3ngy83B/AYEHn23v/aXpAxAt+KeooJHul779QxkV1UTWpxqZKReTsle5Dg95MP2pRqhepec4
H/1yz+VO0wYfZAUFx9moBw9rVhzFW9ydjtjy3uRAumUJrlaykahjMyPeJdAHlz7qg+VBc7zp6PaV
ChmZ206XCR4PLiWKPly6bFljg3hmaWV1S4XfCcmzCCqxoikbq+AjYhV3U+NT3ULZrnNABnwrwnAf
mTCptmrjz+qCBPXAxTy3h7iaI0oNuYRR7KMRg0y3D7MmXo9wXmFeqc7FA3WgApNlEv99XO8oKN8C
ETTXC9Bgn0Rc7I7wqpMlKce9NKQ2ZdxJssR3ntiACKS5P84BVEmb2iexr4kNFbWY6x27/nChzLcE
jsh8Wf06YlDSKt+iMhEq8qGYmTJVA1CkpYa2O8O85xCIEVyG2Buhg+PtrsCRBJow5C7aPARVLho8
IG5gJrHEtEwYBZZyaErmL14FmyBkK9kxraG3aGuxmTgp0AIQmgLyYpirxgMcCWCLfwAYM2vg6Nx0
XkUvQEs6QoJ037QZ1x9Z/NSLSTNDNbl2UkHHLCxrKXJ9LZ+Jwow4i7b4tpV7HjuT60UHf26oVurM
RNreIQm8qRUKcZ2nJR4AyznbxzYe+fyjrw46fYiMrboMQNuz6faIebiex7L1VMOG97sCRWS8UogG
6kNGATBmYgkby12SaS0EoV7dc+N9RI1dQbjZCeklFGSE6ktiecfcGMpFRe8dlGZAA2PX8emdF8gz
DCuIqJywhbfS+/+lXHIPzilEVhZ6Rbhua+OXJOblK4K8copXQPNb9pSnnaaBisVBqKo3nC9LT+YJ
YyvAaTP4z9NQ17BUvNfOQd+V8ybdwgTltzPB3DoxHfkEOpvGHLqObcIh47oK//StzgPPC65aUEmG
q6pVD0deWoKDIREGV8f7ctAHf1u1+49HCLAUEq4bK+6Rf5OpBwaldAJ6LEsdvAC3337PxdmJw1aQ
oXa3sD4xh70Htz9JYiHylyChxMeHj5bU27resGSMC8HEN4G3/kZjZd8+iTf/oiffa9EefKfWmFyK
80L3cPx5AXi42Xhz8ji6thb4WEXp2Ig1ziiwEm3wbPyKjX1Hrl9hJRG4UAbC2dXOlf4dg5JLt4O4
1rZs0nQ9RWMYgMQcaVWcF5BhNqcsTwJRqyFvrsRLG3JN/qhb36Rs+Nf/qudffA+LD9sN67EbMMzL
Hxd1y6GBXGcMwAr3YRysDYYWPD3C0Ji439/W2n+0vQzKag0k4vmlvEeAZ7zYmF52RbzF+6PFHEoG
F1Ocl+8q2olh0OjhuVj0t/y9VIzkB5Kc4sL9pXbxST/osKvcNYW/d4X5U1gOxX1lGw0GUBtukYXP
jB4uyEsLM6zGqJePB5gOCF0s5S7YWTlkN7m2+fXaBhjkmMiArA2hxrb+PUM2ywKKd31rE6cG9+1o
PKQzGmDkxpuBhlUOqx5hzVE5M/TUCsF40JZzP3sZt1p/9zxz4t9W/IjxE5IR5dVo2Mti438iJzBi
J+mnkCp9O+R1L8PZrNFY7CHRSG+CAKivg5Fo5sfVbgi9EDXmo54mIP7z4jW6Z3qXHdYvnjfvqmtW
ZB9gfB6QcNTQctCYmguDnEPXKQ10uV5ORjrSoNeh1mnl1TQDkJQm31sZdOE0Iq9BBT2gfUrfNGxj
rVr1D+YBR6qQQMDbggV6JLLLDLbdskeSC9lzsrIq+lrl09oEIMdLDV8kQ99QJ4NLBGvce/WGxXJA
y9vPRTCv4u3r00txq4I98lJuCRvL5Hc3Ar91Bn+UryuU9NsoLYRJu1YsnyeapMLRlm6etRYH+9pj
ci5G36xn6QjB6DzD8ZoDH7j400Zl3fnds6Fw26mSYjt6ah+zqFKxppR1C2L9dUu+eE02m71I+7US
Frmpq8nW1rQloZvcHXYW2dwXlyg8S6VnUMTRVssLyRPFQhObGSb+FT+IArfiO1ib3W4SDwGexmtH
PGoNHV5JxwSKxvgrQlUvX2VGD6DO42KnZiVQLjSBa9SunI83BcdJTv5YtoCOw33EM/P0YTpDgKRQ
3iXS1S0kE28iqP43i6fJZQOZvCuN3C0eHf5T8I8bjOVJzMRwKmKHtnLePZftRGKfIt/huJa2Qf/o
OhD+oW0Ixr9YnyjpHtnPybm2Kr92SCpzdHFf70SpVDS3icLjC/aOAoaDb2fRvTRFcBNP9zkNbsQ5
pZpdagjtzsc/G48hKdfV6hiC4Ib/1gkFhD/RSSbEiWGk3kjb/Id7ma7Dk2rmzlGAn1MtpEpuW4kw
wl+gwYRwreH41829jnkBQo0wyoWwDN6ei3jDSUQjpmnj3tSvEENXyZDYuAkN5+IlecF6kudVaY30
sx5CO42aDS42mDqwiNhUJSKVBAgBCrREQ5DhLqV6lk+q8Klu2T1yTPrJNrEFLDOkG2UaIvb7Ls7W
XYU9L9StPU6u81M0hNeeJkjuB4jAsOMrtl/DqaUXK4G6QYyFHPxoC5yTgCYg9bUV7anPDhVAy9VK
al2ObIR4Ibi+20zYC+ge6cIc5R9ZiQBa9aOnFb1BLlufY5ZKfU3xQ8XjrR+33z92lchtOOGXY8zY
MDJsf92ZNjmqDhdgFnWcCo6DWVGkQ58w7X5ZyOx8k3izZAmLzq8l5vaG6pHdMoYYOFSuprdqpJPF
2N84vEkKoWZ0UKAx4LJVVQWnf2GVUe60px/OdtP9F3CbQFHvp71Hmk8Py9sgIZeFf5juE9ZOCdaD
G/hbKy5vlTDOY8zw/t6xsNzmA+JGtWoVzaXmOigXY8Jt5lx2UZYAZxWFnArLlYAdxHDa56Ib/1ZQ
largJN0HWO5ABSOwsF3gssnY9/7tPUmbuD6Jax4Htpqu3NUd64ks+ZuoBQXZWqTbAWnRfCLQVrji
HNFnEmLucMyE3V2uO8Mf9GvDsoBAkqn2raVRnDI+wz1Pyf3usiwpBTdz0FzTwExuXbksNnbnAiT1
j76uFsD6U2r5qJt3Q73o5dhEE2qPFjNT+xe03BdUaM42r89UTYG3FoaPc2b45eGfNzkgCKjxYomQ
vdSoMwUXeJk74cjo/xSKVnBCrgowrmH8kRNqiwEhhzVhOIPYi96Rp3b6CGugDothCEWVqssECfuO
BpbTZLusMWJZHlHhhtUPRnvICd3SWGkUzM0MSvR+kGjsOjQdYFzPnr0347PZKxS07QOPeomuiFVi
RaV6EqGneLQ3krw5XJxMXkiT7X8L4dKefXDWfDX+eIOWv2+SmZNJRNhkANLlCG1+2TOBq9INf8a7
u1fTI1WKMKghoFA1RSejgUCMIM444MiCIwba0/THTIEngIEZNn2oPULjR6PgmnZlQeuddi2fuRsL
L/H2BMzPGcBRcOuW5hhcyzKnaNCsx49Ucu1DycMuqbz/zonLaUcoUMTlHGXcD/GbTIoYI5y5uMax
1U2o4m6BXPP7dMDSMRIMtMBV9z3BuyS8hsRNyJwVMM8dV99at5qQEyWG4pbx4be6f9pc/1zzAE+S
4zN0YWE5qoU9CB1QXu2MI+1FbEC1TSKOS1RnRxj10B4jR89ulH5FOZUYCWonqFKbNgCRSsxKiGlo
mDi9cG8Pwo2qq8Cu5DGFPH2JoAU/5L5XtY5DUQqM0WReNMNyRZExKbKXIcRF59UsozxguFPA6T0m
AaFKeHwPbcSsqTU7ZHI5Umlhb1dKFPNF5n5yWTS+8pTxsCO/+lpLiWMcb0Gpc2dgoam1d1yXkSRj
dpG+IIC/3/eq7zaMnH4EtGEUBjVyhi4/HWRyrkxC+/MgvUz8DHQvr+UbkLJc5i74XZu5hWUzMXvU
fRNzfTA4nltwAXnwz/H/SdUwMHK0q90PtzNkdMry5c2XcWkYZrd0TvCfK2KZ+l99dRfUf8QEJWDr
sukjKHoNreFMV1wJgHwohJ5MSCMEl1KYvUwQkQJRVBz928R6Ea14oFdy4VDhDRUMAAKLvqfFvm9v
O00Ay35tbIGRNRfTlDiW1DVk8mnZXFMLF8f3YvJD5y88zuNAmHA4ivIuXQKNeDPH5LnFByDLt24Y
u4V5JeMpZk6ToBWIrwKiiTJFEJkDzgVF9MFyJfgpMYjD+TOuxBg2mpYyygSHDi6zjn71N5irTIAh
NWw1rR8gYc9GxIlJ+rWR62OtD/fzsptk7y7TQKG6xS9CAaYaDnAp1/42egwgSrQoR7AUEgJgfJOz
XYkDsDx4aD5477vQtmx8/72ZeTUdJqfVuhi6F2IvqLV6U15cv6pce3c2gLm5mKoD3DNadSUiQfP6
eqiLqpcdyh6fYLnpj8WXv0LkXurbz5GA7kW8p/Fn1jsHctJj7rk69V1vJmsGRGGmd7+MnX5humKE
GUegb/YMQtkOuO9T803VSz+AsQRG1MqrprzQPiLvrl3TYkaPoQS+dcjjdUvpCELk98GwXCvlpmPl
uiQ44cKddqBpX3wLGhxbTT1W6tcGqiY1OSdgT9vrSOniNWTISUMkte3UkJeZnjs1oqwXH6qumPS+
hOPeCRc6IV9saBklmAc/Qyv/3x5GVXKEYxibAGb14Ssmylm3iG3t6ZCL6fZEs4lWVD4eEpzw91+A
37TaaseYSinpfyh0yoH4JMXtlp12UPgEW18ph2Hiwpedlld5r1dBE8gQShkom2R0rdW1APeCLTMo
fij3kbWwRTYZ1WGOtHJPvoI8K9xRVvXx3czXyeSt/g6nSqX0E4EHhA0sQ7e2Axw/l7/xZrMAE/Sa
QoJApdC8F4+VhHHeTffc7P4xJR/00y9XDWyuJWD51b/b7aFMKKcvwFpbS2tRYB4JOnsF7TbBFsuk
kC2Zg64be7XTsgbGg8h7rWgTEoh2VUE7I1HFf4GHbNTgENiwC3ci4RzRALS6eAVpUYBkpdMVXfyn
+kPGi5FNPJimJcC8ZAEDZDRhj2XvkHnbuF0Z2AVmDea4RNi0fQHuwMkhNCA58xzqCHgzA1ZkraYe
AVn+TqP5bFRYv5krTQ6TkoLPKP33UnfJiWX9FBvUcUugBj84rQspM6963qKVfYoqbSpUQ3eFGpQf
8rw/lfKHbQICFFmRxLzEvv5NdVorrYT2m1remqWdeQjcCtQaYyJa0fg713/er2rTmnIn+ma7NHyC
AwP7Gg36DWIt5pv64egYIUolrH4RNZw5vln3LcMyccePIY0tmJAJhfuIsZYHwtqaU1bmYfvZNnNh
G9uFDzT6sWLtRSRnTMUrr7afA2MLblJ5SMGLgTGhXQOVV04FuGWZUE32tl3YYUsEYAEaeaf2KsLQ
2dVZkq/VSLT0p9ZiWjSgrYD8QkTnGp3HNGef4Q3kDu6A18znl2dvhw8D1dcsKnEcUzxy1njXdHGC
bdss7drOPGiHKcNF99TXniMgraNSEWz+TuUkUjTktoM9pdgdH8rIQyZAH3per2j3NxzFAhHh4Sag
S8MLkXGXrxC5WZygXDclGjmjK3iw/9MtDp9K4Fmv5e9kWP5+GEdkx7Lq3WUtxwOZU4X6vILjDWOX
T2Pq3JesRWr7ECF/KFtXlxTRsDt/bnKvGoNMmDQadYuqFWKvz6riwinLdpu+X8jSM05y1klQrdRx
baAmhzygJa/2f/8BcssAWH+27pzFZdn3SrRDZnS5xl5rZqoNRnQGIk9TYHjkCR4zHsaTnMsYM/xf
YKLnriAfLgH0F6CAnEvWWgCXgClIgw9paPvx7HPlcxq+uiplG4jq80JxU4b3/xKy9PRqolU8zW1I
XqBGi3leEruT8TfI00WbS3+YI9j9dZGV+1y9ivjg6rxWU+b87hYWia0PMh8mf/0qoHaBRzMK3jR5
Z2oN9Rkz8jDMFf8Lbz7xc3anpROGpEsr4j4ZtN4mRlyTbMalSC/VxkSb4tvf2FyRNycnA4bGlOuH
oFpVc58bJiW6BYFESDfOoN8D/5/9eUreOF5DSBTO0tVAau/MaslyEcLs2M+RTAsyAFN7EUDC4m+J
ilJn9+vQAhrB7JU6SJHUkixmj65vinhDmfa1YEcYktaSb6RANrOFV6ivh1EuquVDf1HBw4YXeKSZ
+cCdI5h72XelegWZMNsgm36VQ7ienl2AKTtU6ANiGod3kSrZiTexe9DxdFYKeyCNmE8LPRySNN2F
JYlUzXjSmAOvbYDFTOsQW1om/SwhtynxWUxOuPQZCvudg+t9yJC3qFQ/Rkzp6zd0/Z+ae1264T5+
A9YOYK/gFvcCs9KMGtLbGIf0MPwLrqFwZ1wK+W4yUuSxLNmtlTzyqe5RSlQTPV/3O2BEXGZKPBYk
QaucRVr+rJ89X39NyKmf1Cephj5XKbl9xbNBwn4Am/xdaeLDOEjjW6+v221g2wsIaD5HeffRoyxl
B6G49Kno3vdyNXCs7p9tfUVK43FYbvgkFb+Hd66hkh8c37ShJOWQpTE3oovFnwupiOvkkoumgiDV
wj+geO3ACgDvDCKCEac5EdkXBxXCw4xQsSDDs9Z+/zUrE3TstdPEauu6FdqfomqNj7C4GMlCVt9t
mX3KO/nCYPHTlQKnD57YjLf9gxF+kfr3+m2/+a6bbbkcGs/7UH7W3+6O/xpGxsbi3lkca4iqhdCO
rbRXDi9JCM9i6FZ+AbQyRO7A7cjPYo177CO8UvvsfrNrU4/D3gkcBC+utWRfgApd6O+iBPvfadTI
Yk3JYzzfmImEUWbqXUeZd7uP7VwWZUAmE//xoe1/4Hui2wNzvw2+Jb1fXQbqQAqY4Fmkx1XUNDPN
4z3uL7fNcdcrrAcs74GsAsDXzFgXdBH7Jm4lIDF9lom2992CUjvuksv3NMjU4sC8eElaZ+RA9P2I
Nh7TiMp3XZ/LWmNyFjbTbzUQTdP/nXWRPmrOaD09uboumfbk8qCnmCljMEy2iRD9nSDwb8X2vObX
ikIsgNvsRoq42GL41MSH3pw0dyHs7d0LC0TIGGFcVSwTLfSzIyr2S16AsSOSwzLZSZ2QFGimk3mY
sikFk4n8Qg1/3zfwf9V7+BcNggIgQGMh5Ri6fQagRE/RiOqFlh6viwJ8Mj6fTH4u8D0jLBY3B75R
wSajp3jdPsc1Fh12ITg9m4hAu3zpQt6mgF3Q0q1lvhgsZt9aOHXCRzgqUfwAbIrzdQZwdSu8Pa7G
YPebzZslleQ1zU7/6a6MJd8bP5HwV0xGWKZcKB8/VG9sFReOsBcI9rMzZpQ0Wp9lj14s+yu4/n74
kOG2f3RWFRcOMu6v0caavvSn61VAgVAUHrdARnbktUDy925G9Mmy2zriKUxlqGzSYTKw8h8U17DH
sy5+P2ETP2z0XGMuCkPg0zyUeKRfAz3pvrMdn64X//2jWaUSK9X9IK5jt7hO6FrXt9o3z5JFcobk
QF1dcG8XZEQws4OY9UyOUlh5vqPmuS6zQ61Fs5EWD423DB+C1GM4GXd6Mcmf8bFfXQcyoVHBXtg7
5YRu6d5O++Enul2XPgZueOLAiV1EtKcj9rgFE8VkJT2htH8WyFjd60o69tAjb3hiBIwUFLXJXpps
R0t6UsrDpAZYi5GkCTb0K9EMnTQKkZhOb6fywEO2sw+easeTChAJoK5hmigx0AmiPeU7NuLyvBVI
VdDNV1RHtr+Zn8ZJa3Hv8j2PSa/Hh9ES7UxvvzUCqb7ynmhNyY7w/ZewAnEBuOSX2H4K20LaJvbI
lPceCM/Uu+/wlSRqj6vwBDjcjFmZ8lrPA4j054O3BjcPhL7I6FxpcdgDTNpbXMly3Jm9HSNVmAoe
g3wF7nmYkOKMygCThMaU8e0wLEjgUo7xOPMUKNRPafxEICEJiLb2nlMj/7cJjuok/LfUlrVL4QZC
ESFK9V8g5Hj1lqBestozxwV+rC7BqkcMRzxAbVZ55gZqATiODvN1zXmaes8fRfkFMGUELr1WpOzT
lvBHikMybb1+9wl9/uhgLx8yCUrz9rWUU2fJZcEupsMCfA8W0jQKTJGRoZgOJnJ15uWLwul6RVuo
NR78zCsa0STt6JQ1pFce8AuijLSxXbUfjbXe1pNrUrN5T3mhK2zlscnpbelvW+jp64aG89YCpJdZ
Jc58j+GA8/944zUCp2dcWTdxGdC9TbLP1g0ZeRZQfrEEijrMLY1/AAdQMjmrZddxbwOvAy3G7EXD
BIfjCbavwYQ7w28WElmpt7mEPZZS0Ac3xDVJA7z09WnQLzTRdCXcT6yxXQEM2417IY7+y51lhYd8
fvZJlrZOHZmMuScuuAOse2Tqt4fhyy0npmrKGmnofc1lEsnzBA8YFVCFHpWlxMq5JKLOxYdmLPIK
v4UCWuDAoStzI7UJgALwFI1sNZxyjPpM40MrAIUDupS2DTKPJmdfKYFSR5dlgLV74d56iLM0mkIw
/ak0Zv09QowU7XkZaGxPraikifQxGegtfyi/ZvFcpp+aHiAX1ebN5vpKqZtDibIPPdqm9FTCtNk7
IYyRwhXSfJVXTkOU9E7qOzfeyXNQQbsB1ia5BJmBs8rNOmmdJnYkmX5JXgXxBUDzuWwv2thWStY+
zP7fM6nUX5LDvGLOxt+9aajjWeJx52TeFcKHg1GSXC+EXQbanGdpPKacQRE6ZvGKhI0mN2auhDbF
M8xBJ+O7KklJdDNm+uCjOweH3Ipdy8LUVowM40UlZlz4zreZP97cQRLzrQBXfWEgrTBEIX1eZlI4
HPllc/2eSXljFtYhddBRImmmJs1Rt37u4kiChILxalBN9VDfUNQ3VbWVXC1qjFmsqbuD9vSvriAq
IuNuVOKi4EFh3fhUWTMKcUK0k/UFS079MZExVHOsSWVv5SVA6ouqibviMvSKUjLXe1AJ8jLpSAeV
J/L34Nngq9l9XY1pWLjy7F5MSz40oF6d8fBLa2Gh0y+dQYvPVjGf60QpgTbyq4F+FF57If+0pKC8
cHnhRNAPjtFTo4SnwuYyA1lWc+0BYpGboEa9n46TfMfHDCrfU3qh/Kr4CTOeF2DqGMKTzX8yX7tc
ARF8fVFBGf6+u1hjpl4Qi8eKKtRHUC2R698rIBZc+bwrUcm1x9YHySHwLJLI9yqU49e3gcGtfO6g
I6wlddtWGZHWuwoqZ/O+hW/jxgFn2/tYjr0T4+tsuQ0fzuYUG3x+hWMXvgc48dfqbt8XQUtWYMqL
Y8C9psQfWG7fk9zbdzGzQFBVQt/xUZU4vGlw6mSLrA/rbUWL2b+ClCxokNxvpWS44GsS93KDf5mG
x7uh9HfSl6UYdNGDG3S54Up4ZXaidnj23UY6EzH5kbOy0ZsvdFqCaEug+Nlv6vodKX9nR/Rfj3P2
hXPH73CO43O4D8OR+Q4+eBRzrP1D+BVUjwTMXSlfAHmidum7l1O0jH58xRZg9OJabh2IZa8w0Ow9
bjPW8ghpDglMZal+3NJwm57wC3hYKevss7CG80U6Ghbi6Ellq0T6GwlSCW/oaz1Qlak6E1SAtbxe
2s5Dp9KhBUnvF+Jf3Xltl1+CS5MqssVyf3Hw7vlNsKcDcitrq8MI8YnxgD2RLM7u1O0NYdZq/pqS
/lKHQR2hbwvJ0fiPOd/d/3YpJFZ2yJAxSxSebMnriPFv0ioW72SS1JyJuD8Y+yE0cDNTLdv3dlU4
TgDi/AgfvOUcPyfuB1Zu/h2LcxTdsjn6RCLtWRZnLjacZ63rSgepG3v5psket0A471FJL6KSfKLt
qjPnyo81k+IPUMTWDb02hOtnvPxwTKWsBY2Dkl+i2tS3R3EtldFeMQIW/8kjb3JQEaBLTBOpBpy9
T/fi/w8mFSpbZVT4NS9ull+aY0AOxN/7uuW1mWNTFwwdX/wPw9AhCdB3blBn3y6S2Ba+EWfk84/7
yxoGzXCvTTpCC8XTH3p6ZlEzmn4R21V6vgjcNLbZLPJWn3iGNSiClW1GYcrEK2lpJvFvwmAt/arn
uNe4I9/jXx9Tx9jXXBF+wG+98e+U9AG2aLWjd1vUkgLQCbf/8+C4t9EOxvkd+X64Mi3Rlzs1UYhS
izYRVNw3oug7RVanconGmXjC2Js9ePsYur+TTCUFqT/Lt2KS1MklnsAd+jfjbJ0c/P35elUsnLIE
wFy19/PSS3ZhCTqNVDD0e/m4yRNj89PP1DgO3895yR/Pu4rv6FVTLF1F/pfo4aSnX8638iJFkmjH
mlFuki7zINjpxSAlTdsTB4XYaIgxYSd2iHYtNyyOvEGqRqvNUqm+PzDrhObtuuMKfC6219vdzSBl
ru26XQgsOSuak/lEBqFPGuLcRyztthBwIIIQ5KYwQBS1PRSkPEQsNDucYAsBh2s1Vesj9/JLcIi8
os9AJW5ldxb6eYynEEFdp96rK5tzJAOAKoXtoyyslmKNsst72aj04sSY+cniRmRhs2WsajV+VLrT
ta/zF84Li1JZdttyhesjix06Ya8KVaVnWd3cu55pgJVEAVIEoL1t8cf1AIWXiqLssGyqXXe3rW7T
q1z9jgdWEW6iiGQSOL7F8Otp046870DpuZ7iANoTfoA7Zk2TU22XcAzfXM0CG66ZtrsZHJN+tiRS
uS7v7+yTr9rtJDS5LzDuZn8Yuxkb0ztundNzkAjCkUyfdlCuBbmYfsLZN8wON52fNtZNUcY/R1ba
Y/fn/DtFMNrUnj2g4+eD7WbswkEUI13T2iYFMkDckBbBi+jx04SCMfWAwnmYsKbqSRnrAS1YTxFG
/d/raoxXzuW68L5/EiTtIh697icf4SL2vRl8DhnKet2C3idLuxivtXlmNzOxk4uCjWVpwdnuSfSZ
De5i5bWA5pGasLbFy0kwWkqksyTUkr8fyrNf7CFng62fX8lv9bT9uITSqMIq/5+ZeFAJtfeAm+rS
7ds1iWwIUXtX7n0l2Fkz3CRwL6Apn3HeomrBWlTmuTVbsaaDN/Yp4WL1NNLtXXSCVm9m5ShvVID5
j1/pS8CYPN5Ih3qHBNaMkKTUP2AipFG8FHI6o1pTzyLBr7+BOONa4JvIoNBTCgIy/NZhAB3Zcgy5
DHGhSB+nhcPfaZERoZqRskt6DRu+xjlylmSZdtyvb89RCAa1mmaGdqyErbi3vFKOUlfrX0fxBXyF
8cJh4gySqUFn/qsUegQ+0czNDDEfbmfmOK46XMkahun3oLZD8nxpkaytsmUWY7C/Y9zJCjFK0Pn0
XM9/ZHJ6LoAlAPRiLmVSmRGARXBLdGZzI/M/0gglLhmp/U3auuWw30BTbYKno1MjexyW4jkLS7VY
gytsgJp7Fylbk31Jj1BxmCOPScIzmbu4H4/NwTgFB2T73MMFtxdDltb1JXtzpbXvusygdAO5xEXm
m8X4G7fH2YNo7spuaVDjPSWhxZAmNMDZPRCT2/rYcxUpddghnJrbXz5T7d1LVEGFRgUanMk3z8Mz
PMtg/sUW0kSTND/zeHjfGjRwO42aBFbb8J1aqwaVWxhm16t5Nt8M7V+f21yRwtZKjB5VavF395hV
we+s8bSm2rrzel31x7MM+5zXkDz3wfwUtjBXGzVcGi8WvtQiRxyfY3jvPQvnDyXpKafAvHRCWB/X
ALpszxPvufKEY842cQoDBXrFKX8tfU1RQmHcoJPED6762RkERWbEW0YWlVxIoQ1Xn01jOKOImUwI
/sQVmW8fSs5tkP4vRw9mIa7sVeRsMe1JhxHYZfrCIrarDrZX7JdLYjtG6SbKZApCwU70HOB3xhrI
Mks/ZWbvb+U1IOtmoDjlqBfbPMV1UY+KlpKKl3Mthx8o/LUrsXxhRtPc/IQzGwOTSIatjUvfij9Z
geUZRuD78qfGBAY3irdgSZIG6uurBV0kVTwuNLEKh8e3o6+Ml20GD2PdkGVmI+NmwVHUW5dAKQs4
A7xl5nBK43xzn2yhtmYiCX6l/36kNQmrtboVtdtfs5lPJRZwFId+PnEr2cbdJUif2gbNEbnZTCZG
JJUEYENQWE3976Tp4RWg8Dv+NBBCxXesWaKK0neYZRLYNwXmNUjM9q5dt18Ox7j7pK6+FwcrUBEY
fmwksqWmYogVus5lXeYRFJGuNgLp9AOLKKY6/otcYQpiiRsx+u5D743fnhOM3qVQsuNKWD29ydfj
/v09qFDZS6Ds5krknkCz1HZoPXBNsaUvTt7GG1m0T27wmdtcaiE4B+3nosLBBbb+Gp0SEkAuhjyN
N89AKV6R1p/09Hpwk2mQRX1A46UXT/1HDhnMAYhs11bKDyGczBnnLta+g9ZP3c+M/l9+G/3C0SUS
GqwEKZqTFlqWoDidBJ2w5Fo5pRpEFkpriTA0KL2DFdN/PX6niIE8w9jmmfxYkENgL0Qyi/ta0rut
nanumbi3ZKoOKi6Jvy6Yvvwt+OuiNfmqPkQFbl9cDaJzH1wTe5TNpTMBZoq3yxPHC+NT5ZzdwVx6
TkxBnw/iI/5co+8b7nwJG/uMCrbyg7X4mBbyHkLt9HDkNu/K0bVAQJpjowBjWb67OmNlQ4RIWO4R
nSs16uHwQTrow5kBw+kbqvQ63buxIVDEP3zwR+uXXjHCTPXuD9OZwNedRq1v8007wd46pcV+Lxv8
yHiwIMdUYBtB3lqi7aibm7xy8A/mfRapCD9a9xWSi3NfTzDj+4b2O+7zuo397LP7z3k3/LdeTXjS
Bnevmx8SPSC6ZyutOvRW1tHN2LMpZ2q6TCgeJIwIvKETHUCzCIcEUWSji9zDrVrwrx6Fnu1mDrFm
LEcYxp5bYB/0wYtPPtyKdKzuC+Q5I9Eh8V6G+EVxtI7dUaB3XfPHQgUg+y/YAdB+FgHtj+yVWI9R
ww/Tnlr76ktiTXL6fzretF05ojtgy53hmiTYpN4rCuZpN9dfUrqD06fcRXFEFfdbOoiaZ5l18RSO
8p8U6wWv3u0maC4aCVfwq8aiZ6LeRed1er+KRoOpEaV+tTlNfkm2OVVdeTnCLMHttsz8AJNIHGKF
721YSD8IO/XdfMoZG4ZCtRTwjRa/WngisTzFh+7uOjs+HSD4aG+iws2T8bVo2o/ojR3caq4mqxyU
f1Iy9yLpz0WJmawRzt/truan0h+Pdl+Rr/D/ni7pylZRetCY2pDpOOxR8vGFRaasiHwv1CQ5+SMa
XjAOA7d/4E/v4zw98x5WGrn+R71dGaVHTiruS1piGPmWW1I3RkSVyrI9o2tHzdoIgIbq0IdJeOO/
Jwqgv9vQYR9NTRrfDIyvzi1IiVLjDN3Wj7Yxeh3NckDCe8jP9YOO7ngO+kmuz+dzhDN/TuKQ6NWT
mpDhe1KyytWR9Urpzj1lE1ZUU7u3lEzcET5f5BYtyRs9gGYf/WH3o58z27NWwXysjHBTvsMCuNkq
dDuG0359CeA9EGl8XJMNdY+/G5LM4GhwCwJDiutf/PQRjWdzSUgoV+Jo0twbUIGYyWHewTD2FsfA
5x9crM2VzRNPWNe7VcvtMdOlLWWPXgzQpF0ci+LtKHtrm0i3W/LAT0zS6QKdO9ntuo2MENfp5O/C
RgtY5UdWfetfjvlTtK+S8Wlb0/sWC4BPo6842IukVcqPpFGnQKK/n5eXJ/gHMcS8Q3PNos/dmjs3
OD51LNAkrZ7uUo6JbrNN8lL1FqFtPWbhPCAH2unGDCnvMsyDwwhtjJY12ZpgJ49PP8s0860CTVH0
8csxGnNJ2b8X8P6rZphFjCfnYW5z2RiL31GRGCimtDMyER90tN8IedskoqZ3xnGmaLUIsxIR9Iod
2C6ewIZ4FN1HijDZ+kZfU20ipSTaB2hf3ufFhg6a91ZhYcv5ZHiNotf13EpyygcAQdRCSrRkTPP9
jfF8QDPieX2/T4PGUGGXoCMpSZY2GRXc5yqS95ly9uDoH5Na1YnmQneuooY40GxxibInMxGrUJUN
wIcH2txnQ82OY6zDCc7Gnq0oLn3pbQbcyPSBsqvdlb8T8vDEKN5XWCPmUblv59lqMJRSYc4kBN20
LRqF76oT9vONudtSU8PvvT0HshVZ7Juxf5UT2EVoni5DSXg6dTlPwFyEpxk8PFv2HG4I6ueaqFb9
eF6sIeFaz4Lg4QrO5Z7mCVrqaofv/VzBD4bQr0sfi6NTD5j/5DGqtNoaUcZMvvEdqQlPy+shteph
P5uPx0HHgB5+b/q65HcVyFmcu2RPJNPGhtWqG/mpiPqMoaRUdSP6BPmKfKf7l7aScFjMKlOFI7yS
TIf39tAkM6xmYhV3udJy5+Jh51cm1Cgtn53SprSz1+wZCgl55I/mHLSI/O7AP5hlYbFVMroKNC0S
sdnx1rGVsbu81+88bEP8y6GX6tTOBSKbA9CSwClqZkMwnV54k/qxVUVdmWdUrQxwTBOML+jvwwSY
NRLdplaPcnxcZEsp6pauZh2h3LsZO2XkhtJeW6bXxMyOPnsisV8NroseGgrczUJooSZmJLveRwyl
a0dzT81LFSG5stFSurT17vLDg+KutWw+0kfi7GGwUICUiJBRyvefyWLUQIc4r6I/Pv7T5mejdxPq
8ypRlqTLUeeZDewxEn9qDyA4yG5S5fyTx64cVY4cvB9Zh9Ega2fbw/lFEtFOVCNFBRUyXiInozLF
fpyDRsZOUjd5KTxtXE1HZA2tujetoF/nU74iZJUC97HpVBcDWzzHIpWGvmmkcaSgT9ypFVTZkN38
lmzBezgSmPX35VvrtBC4Btbc+B85IW070lG3QIaicrKc8c/DDrExYFTYVMFVvFzuh0+rH8bL07ff
s4EkWFerg9ytL+v5lUEqBQfRyty9TmsxFwNTu2z/PyIM632p75MsMuHEMmMuJ7GUE5yrrnQK0+5J
XLHTZDMHUnIix9oQ9RZ+ovW4Sz7dP61A4wF3+nnG9FHo49BHIj/eNS3CJr3IRLW7xfnJ64un5m+E
JR0qcnS8LFbfTd0gU+OxN+wy3NBLKm8RjmDOSYqdEKt0n/Y/b1zgJgNPZlBxejBP39nlnLDSUwVn
UOygft59dy6YAKcDNu4TV3AYkEwdaPQixP2Te6wXEuNIgC6/v/3ZNv6ldqC7OifYthSYnEuWOcr+
BfBFpnea/iwW0dvLFqsUIsGIuYiVfRxhuRLs6lKSrteK06kPHvi0BrpSysx+ScIcREI2xOp7POIF
DLbzsuVRYhS08nfKk8XKxEUjpUMRamD7rGRXVSsv3mw6/FetehHlQPbpHzu1z2TDbOfTqU5DiAxU
WdxU8N8qd1EHQsZ7KTckk1/Q/eQIXqNZn44UuZWfBI6bilV1IrPFjLTJJ9yAn9Dz/x88q3O35SCy
99h51SMuZXwsQSx/C/qF7o40LzCDWI/0G31qannETv/aNAreWuudZbCBaaB6YQ0IRV6h1AevVwx4
vPZly251ffTe3IeuEctTzpUWpmU1F462dAkigXmqP7MDVUHokHfT+da6EgpYJlZydpb0oVIOQVYN
QfFiVRPy19juALDTH1QQvrQFFJWs8KshrHpyoYNN3DoKyaWcYBUtepNwmszJHp6jsYbuPxY/7EDP
nam6zXA7msLju4SQqOVdAWjz9N2Pxsf01jqISP0uJpwyu8+F+8+vMnLIIyn3hJUBv9olsystqbev
yFIKvh/hRfXP1M4dawE9/kGotQViwLvS2SmDvgan2cuN/56v8vKQJzWsHz5tA3JLO6dpovxVYoQj
tTo7NaWpbJACz5rfSKSh4ZB83t1t0dXWqR8b4WUGlPl2so9JIbiC0jJoo7+SNU2aPTAX8zvRuWiT
eoQMr/dCu9+vm04MDxxNxVS2MVY5IOIWtnDGp2qgi/xLRz65ZV1Bix0LjfGG0UZMUIno7w3nXDnJ
q3i9vgtgBC/wN+p5RBAeeyvGdUABtYwAT+Dhnm0HRKEmtq6sI0gtPWCnMAOULGe+U/oH/+vNp10y
XjvWk8NV8qqSFPnkk+0jk2skCNJEI0r4W9Kq/LJtvt1l06AUzKrrD8nHxhh0YrxZIxQEmjQEffzu
7w5UDQNTiAwBSZ5aeA/kkcy8Iu/x2h+2cwAkefVYmbql02Fw1eYzuHU0UQF75dhPPZGm6AjMD3Ga
1a8KRYwYmWcxBxmMnRvSJCwgEzovcaQ0YxPiDQdPPgj+G4WVerMIcVmB5pWVgind9JBgq+SH86YH
cZSXl36r8ubeg726AfzkSqYI/pG2/ztvJr+ldWQ1Ko25BQUt7uPF+Q5qP4sW8FCl1RFrW6Sd6OZJ
PDObNtMYfB0xRkQwjkk8CH6QS/vRWgJhJT43kX+R0gBzRAnNOrPSqPECFrHScZ/WjbTifytcg9w3
cF1v0S+OfQjoYf7qo4fdyuDCbr6dqIGmMr1RP88w7zG04mNaV7IDhNZWkwkvJAgZwOuNa+YqAlES
ygMFEKaRFmGml+PjGl+6iAkbNs/As0/B+1EYWxs+6C/EnvV4Y82xBzOlQrsx8RIpwpABSoIkE+Pq
NjccSfYIqXXsyaAcaQMfF+WGTV4bgGFa5a7rjk1pi0mfsxZcG24fVQ6IFhpnkGy8BFP+qFOdTXNF
5XpqD8TpVdsE5LQdJDpmANeJ0cXtv1vHwddVvRN913kR96LaaveBMdWmL468EplNXaT68/lHWQyV
dn2uuedQlfQJDv8e8Aj/3ZehLarfoFF3OTqwuow4UBqrGUjOtnStFIkpf0q1MlusSG8j9UW1rEuU
mwy5abpHNHr0Wd9fEYWSDphLTT8xU4QA/4huyrJoH13OC7dLoYByPo4hHq7lg74VcWeyYaYIrqzZ
VAzzGRcy8lUMCQ0bbIZSUk1ZktwP8bzbDA66wb9YpRhPdB76wZNZLiwzwYesB0H0WfnSVTYvYDsq
cPxyUFUWJFiBcHhLabBSWQ4WNON2/yvS6hPxD0YNNPIc7B5/pX9N2ZPaiN4WeP8A7uOypxs7q9JC
Zr660EpO+1OOXW8bR2jlrTS3LwPDrPcZkBO0lg5r9ljOK/whWLstT2sRbUAyJVL5DeBunNMl3jZl
CrCirLkYat8C9Dx2NO39PXFxYaVjt8Y+UJKxVzgRjcnfn34FG85insvjCyqeHbcepFtMAaYWuGNM
BltLVQzvlUcNKpstOmaXXvP0k4reed7klCX/WepeQXIOT7qa/dwh4buyCaH/D81u/Z5j99HCOfdx
RYHb/U7AIVcscYrY4uJfirb0Gf47nQRkOF+4MWUBycjXn3/CYMli1NVR3zf3ao/f+XEH0cH6uem4
LjccrIeUROzef+XRBpraEb7B9UkzzXBoiWNE4E94nNvO3Q+yhPBVqMjzYJlWKOwW0Xlk3n7BP2g7
gk1gsFCFMADLrpsB7Nf69YlRaLDg7kHEHXAHXI5cLuaPs+qckp1zxM1d41RmUiLpSqsgYYNNGrd3
Jlcyelc8oepCjFODRGnylXz3zQMAwdgvesy7e9jD/r7/b/XciqpnoZIlmjabupEUY/0Fk8dE8oaS
m6n9tY55x4iNBuKsMTj3zrI3VJfiuCNOH2+fKFiFa4/ZgQmekJJ3+F2x3SCUBOFEhGYOq2hL38V4
7SYhO6GWTArLFdV9/O3JDhl0BLeWN1IvUXDcJ+clYmLi2y8f2OddsHk65UmZYNfKKKIKr6v9+QDI
3n2UbXFsiI0SETogibGcy/ymzogPq40HXAwC9BSMpeXDeQBAQxLnjuF0ubl7IyzATPSCWk7oJuv0
GaXaQT0mwks/O0AAFohcIadPfEFuBDkpMZ9U7p9fl4tt7CoaRxM30tWrbTvzAV5qneoyg0vLHBHn
3R9Q6FN+vtmZprk2kTAHn1UGjqATLVvtp+ASHNDx0iaXRnrv5tqTkNZTOmJT2UuKMvS/RlI9Sm+v
AZN+64x30jt/dQ0gfcFy+rv/W6wBkUFP1eJGxPCZNz0R/FUD+8+QHi5BF9uqeA8KTvru+znErohM
u4puVrparmDSjlcU7PUFYJk+yRXkr5MqtgsPh6vAG9M6qnLjFnIjPyjSMpxmoaMQMAGoeFZgcFp3
3Fio4o7lVSng3GxI6Ou9eYa6bWTj8wz1CZrpj8qFZ0Ko1ZXH+0XoLPE5ULTbWV5ZdqI667RIpBtq
eG0ujjlLZjYp3F54xETYTb6C8HLerJBuXDSbT6gyutvHhpFWmlMV8mXOx+oViTQqyNUCdAhUEpD0
qxoxXXsn6+j7PLeq60a1QkO5mPyh+pq8WtNWuinyW9oP0KLaa50PWFNHSqzzv0wJwTpjGzUSIvoi
FlGTj/xeL/9TktXKwof04gKeeMK9PQBFa1C55sqQ6StvnPcN3DRCm3eNy4eYn5cjl9T9/fUJXeW2
A+Sx/ZLPtRuFr35TVJNjjTu+0PYFXPgsVFh/kuN0MkejuP3SwmvnBCGyChFsVCYGuPctdq7jqHFC
Yudxir8HXSPqtZQKpcPhh1kUocgSk9PuqzcLKayYjpYEUEGkF3k9+jQfsBaQ6uCUxOOerkdiQc1Z
CCZpo4eRwJmRhblHAOIznT/vs+im4lL+VaFx2SmMJUFOF9LWFATwDVtpWvspaNg8jLgY29omZLPd
EjN5fhWpErT+pkC80sjCFkalidcE+arvQeX63qEN3OU2N8+xhSKmddFlOeebFU9/rPUXwDiG4dzW
kVNvF1mxjp0A92sfE44ZwBLV58EtAuwg6kIMPWEtCPbuozo1uBnZObXaCS9u+R28LvrZg6imbT/4
zuUfFbZNmD/nruoPLU5rLUXrTuevsuRXJbI9+YMnMymOIcb06sIbmcJ9hr6dDnB7PJ+lLE7AKb+U
xGQKuh0zp8ZjyxaaeHGTn5BOndpQKJlAsp22INqUMmgAHMizSKBHfkSJWyeHhXcjqHLTd/h/i/oG
YbMV41DQ8LWzHVo4+5GA8oH/MAGEGgceqmCNvAsoKwJMV/L0FBjQA/jm1LwyJTJmHPisWzDKeSFy
/tY08wfz8htioS87cC4TdV20ceniHZRRLWgG7fXzdrvNAGj4PGoSg2Xb014R43NRWLZHbBxOqDef
2JpNjb3VzOTxt/iwv7aSqTMsiTUw67wMMZ9E7eo/1Ea9+TPX8rCD0P5oVx4kDYHr3zQBS5i0dvtF
iLJ6j812yUQT2C6USsjCky8O617qslyjr84UiCq/yTMWSpVhFdHp3ED0GZSGPO/UwcwNgxNxQoov
ChXcM2dT8kKZGLUS8g1j2m7dQ3Ow4i5AdPaKgVbFoRxahxLhNAmGG4uCss1MKV6MDoTj1vORqjyi
DNIs/8TynU4xXtQp3IInN0NFPk2fU5E6bYC9bDxgFo4e5Uodgu+ZX4v77aQRqxVvHifLAhpotoN8
Oxr+Fqif/vgAANgUCcoI0Jb/fOjdxzlPluw/WTFxgxGEsNrUvi8orcWyZvXG6j4seKwSIwXdPqfe
95UsH4pm5nvTHSflM0xZ/JokWLn/CVoDDmd33JMNqqhj5ULVU4uQ5AaD3WFHkee9hT4poEKFmguM
BcYWQ6jp4+6yYDAyCp3nPIqAXTkSF/8deG+rmpSdQ2BW4STopg0Pg8pYjsjxJbmqmBT4+jbW8SHT
6Pj0xgr6oZwmaq/CuOADd0lE2acgQaxgqBd1/8XZBz3CwxJxDWo99lYzAcVN2OXiDs2T7PiHqpWg
ncfEqSPpQes8vCiyFazTW6Lbu91g6YVYnqJQ1QPMbXNAH7daZkW+HE+s8QMucYQ+A6mii+P9zy3s
Ul8bCigypSt0Z5L/SGZv88Lx+0FbR9+UhIt2f33ANguu7xFULsU3UPPCRovOO1OVxCDW5/M2fUrC
oTLWF/IiFH8XegI3udERfBwOIO22ZXU2ozVvPCh3LDWcrvJ65X4bHIFLTJ32CedUflttdLtdKJZq
WpYGfK+Vhzc+iI2pplsbgEgzFKGNugebuw21qoT1PGXHjGSKZWGdFMiVQi7/MSKXrV72ltfFUiID
bZdKqN7Gf6DkLoDsTDKPdWukeWXBFB7e2Bd+bOZXgtcx2983yU70ywLS6sDTGWDyHDsP+DUiDrKY
QtJ4vJC5Mhq/b618K4wCZ6t6QOwezbpXGRaGEbKgT9DwXSzRuIKVCl5MJ9jxC5yOGS77G5btxt9N
e7aBYaOk1Jk+8FbbjLwPfwpTdHDwUybI+Ep88aOqVVMlttG3EIW4mxhKdunR8YeHxiIKuQAFPN74
MaII4vCzNgxVWDkYNyxeSn1vnzhPrLSiBM+hjaE2D1Q33X/2G6lozJe8RCq+xNk15V+TJ6qOLdYC
vb0z+GKkEx7YIvRAqj9ZMOcQvvjdszeDGC4hgGiSILEY8j4bqhltqKYTDp5yWszryFI+Vb3bWJmW
H8PF30QwgWj5sK/VKf243GLebgazSbZQ/v/5pAkXCy899fsou54AlUG747fQ9Acwvu9TWLWdRIyK
FX6oPeOx+ocNdXkSGDlTFdxZP8twWfIJuMDtMy38Wa1f19HllDaRV0kASfLh0WyOQ6yugu7o8vx8
0vRUm5kfmyKt+Y3012E3wRa+SastKGO3pXd2lD6QXVEOC/IDwzPaI9F+bUlZHUceWvL10RBGc5ID
lakZvnUlSR4wPlfxbmwnaI6qWsoVEMZBPEplFSWHRmSF5Q2A1NPJe1Atlx/tTTcgPmM/fk2pBUh9
O/2zIUqTr3CkDVglTDgXjq62M2TP8PIuTDQmKy+QCn4SyJ7MynpKmNCjw4PgTrUQy1mwuYtOSvmh
LEFKknag/+Oca6AYwv0KOSafw4+lyuH2Uxb6Q6BCm1QKyChEoCC8MXHrc35kxeOxmUj7cpi7yW7L
c9VMlff4iqunDW1uRYT/EAFHLWDxo8UTacwzcqVqGKV7vN3EhvO65F1UZEpq+vcru4uDlaPsyxSt
hcDiONT5C5gKtOZZ1wZo1dJkwG4ED7JmtBsYeGIuzuG6OeK+2D6O+ygAjEu4NKDFmG5pA0FyParh
8GZh5jwfUeRhD90reETkcCAkYqLl8/FSe0MmTn/OfzdsyCc92gCyH4DUNO2W8Al2GzaQqCaOd6De
tW+r5ob5DIKOgqtJDbOt9ZDgLEfyF+IC4GhYue5XpqmkG6CIz9jeZwvdm0bfln6dpG5QbplxJlCQ
sP+Iqw+BhDByf1GN6U61Pm1S+y2UPmOlmb+FUORFuppedLO7b4sA7h8eD0QxkC78GoJqpQPCaMGO
FVsegxnZ741/9YP7P1MB1mlteawI0OnnwMO57aNRBnC69O+JNlX4Uf13F2bHhAPf4tZivR+zkZ/U
EGqzTOsqvAV8h49LFhk2U4phKiwG/6s7vU419jbx2zB9q6zBAk48WFp8IIjsYS8VSU8Ut/pez46g
jnC2GKgOe12K4pQuTOHIbAc63aq+yv1H9k8ijvKLEBR0sWwSRQJx/N9Qs3cE0AFLOSKY0jL61AkY
CTlitlYNIdqeSmhF64rKvAKGRCUokOQD468xmC/hKP0s7HH2RixN7ZOq/hkJdMWqOZ1yCJgDsE+f
TrTGCuj4jlvbhR3iboPSbiD9peL19/AD4FpqgpEdh+99LwZoQITkEhDPHj3xpRyqKf8MdQkxyPS4
36BtmVuAHSvVxiC3lfXdKj0fLU3eXCetX8EDcrctlY4tR6CqyyzNp88WpZXKIrJ/GWUPvVg8MeGt
JrNE+Q8aLaDQ8jcg90qMexB9VmZKvEZJdsMj+60UtbhdTXvGvo6kxwc9gnDH275ryiOwJJhz6qmc
IqW2a0X1thfJ7yGatnPIJl/MhvQ4Ws9bysLLGDZGwqqgzmuYo0it5l/2VsBZlw+54LPS4gwcxc8w
IquGngiIrRNnztAfVSNM54n9kGVrCydKjRwAyDSle+ieXxrU89yxzBqrBsMZ3bLBgbciTUr+2crA
h6iPgvqWQ30jGFK9yM3Z7hg/awZAZ0PU/5L3K7nrIP3jiU+wGufdOACkW2fl9kxQipeFkuUEgRio
0S/8jt2Xfzen7djyO9oJ+9tWHIBWRUqlJkXGbfa4XklLJaed8HgV+rymv/vSaUQkdOmCOjP8kHFN
1hqoQZD4zZztJ5JwN0Z0bWN8IicQkNibCNPcGdilMXYebtBD4ReggUUv2kJPSU6IdAWxRetKwvdV
hvBM4GO6rXx0sZK4EWuVSRcaNd/PwQojnSF2v01WWIMxSWhDNouEBFKjqNFWb9JucMvFkxQ1l3lO
Cd+k4gqJAphHLiBwwpfyUT+7sb4IcZuaUIxHrUZGz18b3hqnVqzY/VHS8NLb8wMtpfXHSjCCs9hP
kdQVVY/WfBObbt+80p9aOwT2JOABO5KUDJXezsjXgfZafIaip+rGDAbgazatTLXjVF8YvKClUjuR
sko7KDEy8knlIkKDqCZUsn4RR8kPZnhTyUpMMdcgTcHkz7FdzqZJthhBZ3q2ew4Vsy1Io04U32z4
fG2nwCdIq5D7Q+Avh33ZroqIKWU94KgBmK9GFJBt5WECI2bQ/YeB66ur6+PeL+tk5wm0nOdzuyQg
siBRp9Syio3nkzDtuIT3aO8OHdmVFKbC5qSw5sGBOdUFnT+bl5wa8iJ9l0Zl8OB3NlLn+Vdywu7l
FiKonoK2VJS1cmIyk881Hw8igweXfKaqQD/GYY2yxMfo3/FlFbvHflaDm+6ztvtAPoIlRR/Tjak9
gA7hpBbOjPJLKtAzy2/yQwjPDlYDUnrujzaWsSLyLsTtWR4hGwAG+7uqfwuhkrjjg2+w1h+eVguj
8OQjiTD2JxnlbeAfsckl2WD2bhbF6hlyCXFNZjZ0ocOvp8OIWLaa5md+ArF/yGMwTcGsZXc9H8Vx
NJYOa6H5IxEe/bOy15TGOEnYl1D5Cw4Oh+W2uFmbnZIMU7ywYaHpN1id655MffBn1BoTf3kV0BNI
CDcyzx/wpYPwiEcNkBouGnccFTuZwD5f6nabtNa6DyPCWLea3ihrMuZcCxN4CeXPKzZzBiQJCsxe
/AbjnsDMDZuyaL1RtMPq2Hp2tSknpGqj1PHU0BfncU/tMA+F9CcCJcBB+rd6DafdH6+TTaT5qRoA
7e3tnhiOgsyW+S6pnOSPh7224XIjtujSqRgQzyXrgwDajF+setgpEzUktmfHP5A0AI6RqM/MP2XY
jEUlAJTLrsgzUR4/A/G4zDvF9tO0oUqaavj3Lne94ikL/OWEXbKD8q0y2HBEWqQ3JjJtRZxNft0A
NRZRDVKshmYvVzaRTbgn0E2LAUFZcyC0qF4dMJYzF6isiUmZglAfnJKAo0jqLUGOZ0fAzvyx2evb
3BiDPFz87ijTrJ7OjN8ABHKF/Fj5qQ3exabf7Btd2KUVcLSMf/ttAZ2VDF/LUvCGAjHN6ADTmAw2
WkzKELUKVnR1lE83ISPBuoL6v4XPhwF6bws29RtG63HPogvqAeogHsW+Fr83RLfY6ylmEgJYvOla
/pwebg8d0mqLc22/MsTbFpTRdO23v3qg+R5X5QFiXR+1mQMaYh0dYiw/11cOjYCLhsfAVo0xr00q
cMZVfHbNVfrgJDpTxP0E1EDggDGOamvZIxoVPivHq3XPI5V3efMOIEQ3dpmo5mUCj/gTKz8rlIkF
CSeQLIraoUgyZPygcaKf/S6fnczymSUHQFLcGvR7wbaxZ3chNvyvp4pbQDFylQRzt3BVvMSNHME4
JmwCuvSgDKrgeTubwJoMQUROl5sEgYaYM3CZCr+OYI00nfhF9aMoVJRyuVyhIunJ/Vy6N0/wWCQ4
dRNJdm7Cj3RMhshZpY+rpgCIJ9nZ3lNZdSZPc2+Rh8PqYPfuo4KFmdmmysnBPE1ZiY2Yfro6WYhV
crf/kJ+ca9g6jK2fSTCfZA1BU1kYL/gWmCZ/ff4eOzgwCLJzODVVYJ9j7aKYTkN2b961rjgpqR92
/c5E0ycLIegHp63sIy5DxWh4mdrM4RD6de1FCfvP6GnzvfXA+c8S84dZlvp0dUpsSqnh+ev+6sjJ
mExy+VN6XwyxuCwE+YtHnMRIKJbm40bAWSQMtXqO95JMf8b2p+B12xTu1LZzeSxs+7vv6vW4XkVk
V2l6ZRwDA02zH1iWnmNtbCicl31uj4lHcSfAQEHMlSKCv71i6vzDT0/MvpTUU9dNNzEhza76WAwF
3HvICoXqwDNh3yQBtPzeFnD8iwY1+doDx7FWWkUnpl/72VYkpW99qls77iyLIjvB1XcfA875g7g4
YOnNj75iTYTzEgrq6LRkkKFwQuNtzUHedS73+XcvlrTQENynJybWhxzQflUvT/shGe13OaBbmCHG
iW9HM0oSwwk44bidabsfv0mWSgoUZDgwGKVgwdy6HxFiGz2UK0VxULLyLgBREkDFwd6nm3maQker
c4JQCluB1yyprm/SNFAYcZEGc6BMB+pxUS2z/rYm0DdX1h5DKoT8qpYO3+EdgJHMH1UejL2kuiIs
zYdAsv55T+mHzxFm+chMiuT1AiEbm8nnqYwLQnCqB+wdki8W1UtxWv2Y7r+FVSBzJtRXI+6NSTN9
BHHIV82FL/P/1sDnh/orPPvLGYKYORjeqyCdJsPvMzDwpxlhAdOfvJQM5oo8hL52HSR8n2VnrGJq
CiXJdbm+izRUQMEW9BPMIg/Sc+j8bMb89N4iSPWl940fOVX7wQlQjN1j+Npe+qgtYxBaiplTccU+
Rk4eZHutgmbB9ahUTeRxAbQeapHkuCQR5G/nX/Ukc9ChWbG7qe9Yjv6psi5JaO5pv6rRrvkbEHCf
2QzWUAPJN2tSvArs+2K7iXrLp/jnF8WTF3G0wsjXtb+5aNTvj/e1j1VIQhNXy5QBD3/hUm6PjRlJ
8x325rkkHxZBZjXmPpV6eGNW324JnbgZLfxGf4uvpa8TP0ZQvgx/Uryz8hRoANLlaNfyJY4rf1gf
zfwDE4v/NRAggWOhd4453q5ETdmSWgCbSk4ce2Jz9j53hdKdnvv7t+VSMrBADmY8DldcgU+7kpFC
a06p3gaaeC7CdI5ZIZblQgIdqgC/5nWZhICl0zBPggk4MSRovRdHSqhmQl9h5LRE8oGXRnfQZyN+
fx1sneyJyKXZBwY7eoaHRLYDBsjQETPiE8X8yrzyx85ONsmRF9+f6EU8IEau2LngIyc8TSTjllQJ
FpgRisRoVl9sMYSZkeSHu3itV24sZGjIDnaLuAb4AjWN3ccnkeF9eS5sPgccxYSXGhsQQrmVL49S
3VTlFaXgc/fMV+CiPitgqDsKYR9/3dM7mRf8ftwzWgbqQHScJbuJXJ24mXPqTgE92VVdYFwqYd67
mHLm4KVZqO+VQmpmlRE5qn2EN+UFozogg4ukHRVAJlrbPhIw41HjBXj4fPboR3kmNgy85c3wwvyo
4Ysub8C+/9fx81CMb7cVDKnAn8/efBj4gynal3QwbPecdaQt2Vc0uWP1+KAcxqCxuXiFTWBDZaqg
IcJOBgtuWeMw+pZxZt7eX+/6/AaCUH6KDkMUdsgIdXvK6ap842u0zpJTS9pKeBXHIFYqqT3TFp+v
OwM8KxX2PQn5zhWZHvL0rQEoS4ABk+OXe6GzI7ORFEll+fLCycYOI+iS6EcwDY5jgvG7HhIO4WlA
sFtdxuZ/hs/AAcL6Jn4eEfBuEy4FbXuYafd/aQpLxyq6QzKJTw4xtJIZqv55NMFIuzczhXktOdmU
HpSSFlD2W2o+d6cUrmj/GwocZ2JSDhl6j16ocuEFRc1cXGpi92ZhcM5PcBRARJwyH3p+DBH5bTvH
6RSIgcaohGOtWXhp3qfoWSfzg8ZAE++cv/rG6DrJ9EALtke0201jdHokpaLA9QszmkjSyIErXEN7
FBBga3PA5XbMg0qW3rPaLO96i3Gsgonu32o58C8fj+LZMSTBfP3HiRsGGT6Iq3uSkKsw1fies5gq
hHX0nf5eeywO/YGass9eag3so+puSdTRnEMwJm9io88//ML58loJGvhpAwRLCiZZNZGD2oLVQH5v
gbdwzhHv5QxY08Itpl5isDxQ3T33i2X1Zxpc+cqyOru/2vAkemLPE8ZeURh2Hyc6z1Y+euRzyC2y
K+cqLheviKeldh/PZ0mBKiwUgUgrobfQUVihrm8g28Uu5huuh0LpLJVCd4Vmdp8tsclB9I5sFEIx
eT9a7Fz3Bi9mq7gJlaa2QZixNHENN6Fnrd8wQmMYSttzGY46oNBN24qzMvB9BcQNQiPFapzwCiw8
fDvk3OMwTEdpWFolEHKx623fUVEHdLvbwN546RzOhXdhllCt5xOtvVQSX5bfQCPayynedm9nr1fv
a7BmhQ1lrewX1+Wjd2bD09gxHhK+FPyQNoY1YpUAvifR4Fxx1h57yrxDfOTGY1dmEZUWbNT5YTq8
TIxBBe25w6PIoyU0h5YvXNihVbmAwzEiFWtNo5gDdZDSbqPIhVPD0j/fWxPrh64tdiikesKO7i46
TU7rWA9PTwkst1KKMGTHwKFdQsF1Bl8+ADNtBojJ4JLUe5RszMV09q+adYVKzUsj+CIAX10YxubV
rN5vcNIwoXNYGyaSRN/1S/Ps/3dXadlJ38b0ARSc9LI5vUVrfS8WYL3fBYEJeJvQZv0CR7H3F/h4
kCGQpkvvYxyXHQoNSjyXcPoJ8TKFvakut122T+XA6quglzG+MrdTXryZeeHuP0anveg4AG1SugOQ
1ACwgffHDup51bR3ZBeEYvY1Boq8dgcz7NdflrD/RlJVAKBq6yaOB2UtuCOva+CqY13MoJzHxj+z
MWPHp6yx7ndEgQN1gxzQf/ZahtJ9XDSvZNROIjuf7uFBHQ2RKqT1x5iBsHMYyqeR2qC1GnohkXTS
Iprl3nAJThumWJWVATcDvWGz8ESJsxaCY/OE3Z63iLx15KAIyS9YNWNlkEUvHatC2RycvMM5+llK
oT9dO4E9teMJtrvOWqsfMdIIbDTEH9lq41WGaHBDZ/qsTPl39AQWyQuIV1tv+I5nuvDhpcmIq6Ym
WzmvpCk6mlB2FDy3MmEbF47U9396/Pdp8hE9ymPiPV1pppkQPH7ZH+yeh5DSFvrZk9uyghDawwh0
XcKPlCZZC2KcRFP1qyJFX4wln8ggt+hJvrhYUnx2fWcAU649ypPCn2dWVYW+cZ1b5EBQSS5wqRT+
6ytohR7kSoUcBoLVY2XoaGeTUQXHGEXyoetl27IcuRbq7frVZceETxIRTT6fXNv7RVC5eU+sjh5z
2HdfHJJMOjlVhh298XYoAIF51mXY21+0DtkYP3yEbOlbmj6KIx12SBZ1LoSMcaQN6JRFFDBlAQ9a
BL78gjF3uMSGgmNndLtdT5ODDAncEysJM/t/6QTfLhDNFNIDxYo52o1JcxDxIiIIEgTCdCOwVngT
LigZlL2hVvUxCVu2/rKvWEm1XH/NGNzdU2kFqDzo1Miq+PhZJcXZaQGgHAXXGPEPquC1dl/AU6xX
BQKkyv5Tuc4cLozJLX45bxe1r3ATpMfRzmGmpUHPy23C+ZimVIBBlrF+gMPs4UT2OtjxgIBAAHFv
Ks11JtgnhwSvt64y3WPkKe8Tpjro9qq7z/q1N92dyyZEJOV9onLH7x6BedFMRknfcIz/qPug/c5t
wTPorY+nny5VXcI45FVCc4/pXheIIh39iP0ZcjRRavmkJGUUrgPdsBgx5zn5LkXzkkqtRyULZSxG
6cMTKwv3/mUxXll7I+nn0udn79+VFMwN3I8ZmWDRgL2+W6qBqve1sJq7FLSAbfZVt2nGCoq8zbkf
q12/ufzImDNo+2wwoouMpxb3btEJ41/+rHKXHQX0mTT+kgbYO4i3n/GxcOdaanc8aFugxYFcD6+7
zZeaemHJ9zq5qgau2ddCoxWafpKS88hjQMaXh0Y49qXZTvpGyepc+0fOfnYQbosJHQTE81Jl/GMi
PMg4eAcZnbeREl/PdpkJi4XB2ZCLRst3k+IHw/vtxMaSefU/d+6zVjcKl4aaKK4UyGtdFeXZuISL
ZmEwA+nh7T309jpwOK2exdCa3Sp7KC+TFCTj3aQjHqo4OOYjFC3LVzfrMwnt1stZQHVT29ua8Egd
xJadCz7+GthEvn0i+L37EqzYY/rocejfm7OiiAXkMbELSz9u4xD1d1toeeQ6Rn867B7bBFW7j7cc
lE20rJaXGXIpBIcLR+cXkprBQuS9Qpb1QL6GDHkL+Mwzja3xX0IScvUJxg50An9meiaGM965l1pf
fQqi3BrDYKjj1rbR5mm6W5SN5UQBkS50nfPaXqWca3a9+Yp0JDQct7YP8M5MlAx4D1z9JSsQQjb0
gaE8+6PTee+ousCxY0nz6gB0Qrl3k0pjH41wPluah8cd1O2BuDBSTieWz/r9paaCPZU3t3OAufVW
rQvIXQxSMy89GUk8Ft2L36PgicyjbTs/uFp6ELutkB76AJtijBavY+S4QPAqySFErNjHG2r+WLSx
3FhXCzNJ2bDMcNxGLBr+c+n0IGCuVMMIbisR9ZLmnaYaeqXKeJNyiR+DieLT9/wwhx30/PtY7QuZ
u8PSvC3wFAPIGt5E6Fr8gKKShZGipkBwb58k4R7/dQzeSOdt5ulIdnETE/XgykMv3O4hoK3GA7vf
yzq2nqz6z13pIqE/oIUjxlr3nUW9jLxhdHzmQIhPuoKWEVSAH1ZDUCPO92dO6lWLwT0tZVeNMO+W
cVFoG/XrYFXGg84wu4RmogqHOBIPwdzBAiKtXa5Ju+O1124DtvCE1+gDCRdIRVkM5FaiFnZjNVf1
KwbjoYbCZJwLpZPLH/wMlZ8goT3khpJ4TWXsipaPERBmlf70N/VbAkoSgLvaAI7cezO5018/D0KB
R7UDwCrDl3I2MGGSSmas8xZrDA3EQ50t8LY9L8K1FyGEJ19hQG9yp30DswcIZwqt8ibZzEbH1k+C
SjOlY7k0J3VdRTI//GMXXPlVg2qQuV0EA6X002vI6vD8wHlMZxl+oWmwlTohPyVISzzph42Ks1SK
Jd2iDXtUwdMZmo0V1nBI3h3DAj7Gs6qRQK/qlOFptCdAKaZN7YCz3cyLstwM0FKrjqEu+nq4Q7k1
vJhD+EsS9tsGyjgHhBgFqD0fkh8Uh62B/Rn35S2wwlLoc1XPb80HBwCzrdaMCKXsjYwt+iLSSANM
Bxmi1yCakF29qepkyh99T/N7zzv3mkSIoA+NWzv+d7oruG6cFn15myTWYC7tNRKrrQERprJESiFp
Av69EOeswXHj00ytmsxqbn2iII7kcSIEPc59by+krEdL97QZHpfAR1wD3mu+UpW0NqpaQsxyF63k
G7SzC5ayuAuNBWoed2L7+R9/5Bfj/qOKNqu9ebjgGp1ISIz2jXJIyWBtTVG445bHenFMa+HT5zcJ
iVfKqr2iBX+fuUoAXkPBC8qAcjp+Bjfxa0BkAYlUlak/Uh2X3kke8aKvdgFLgkhR24OGPxmtgci5
jsgjiNri6xbOfigUNPomRZOyJTLA7rL2DFIF48mHUG0YA2g31UOZBadKjM9rByGn4PpQHoGTUvin
u7T39H7Cc6WTODBq6rR3+WA+dKrlwhw8mK3tYkINru76n8VL6aowzHErXMnvAwH+WGJbMrgxsQcm
R9ffv/2O+JxgdL0ENi259EqhU/AlT/ur0PhGlKdssz/5Ir2V0/HhgRE8Zp9JndxdLKyTQrARv/Jp
s6CEmriN6Sup2e0S9Uc0h6zJ1t1VDNGRk+hi3R6bZgtwgnE5kffuEQxCcwiWeyG9TWGD9WfvQ1iK
eRfsIDOojuIiGB/ctDZCeAyhwihKEwi+zCZ/KzPsXAB9xl+I+l/o+1VBBK9dyWYuknDn9YmjFidy
8mhgkQQ6QPXGN3saBaidEkdJZcHpJot7JgNfNwGlspTFpl66/xE66jwoMcSetdWpywtefsRFT0LE
hrH0RdaXY9dUFeZ2Gbw+TjWiFnKN8af5iqGpyaRqBKSNRthvQD+4SvK61uOTmLGPffDZ72RjqHDG
EoIuE00wSiNyEW5atTB/sHzX/JnoFMHKKB2EpiU/rCmpl4HZJExMRLmxpJaVuxY4pTmPvCsjSGQk
Uh+hDRnzMr0Lz2NvH+w8ASCrAy5Zvs/vYLgd9oEWcc4s0rdTsOHYEEyOkTNa/ZXMwG9zJsMlM1S3
8uKRZmioTbGS8fCgxGyD5pIgFWBd2N2qVepybNMVf6rkNBHM76qAqFu4jdizQbf1Gho9Tmcye1Mz
ti1LJB0/8AxF0nh3nTocu2iCe1kg580KWOygnIvFaVm5KNtHlFkaJM3pWcpcgbH39UUi2dVhxdK7
EgFdjrwrLkLwCbs9jXhxFd5S6OH+4aK0oeEN4gX4Hw1veibcp5ns9oVkhcGnBFXDpRKJLzMwbbk1
X92VoLXEaNkIeOvHbWaRVTNdNyEgseC0QdzIv5t9oc9feoGsi/3grvnFSenL55M2fw4W/dB8zmO6
k56K7OUoNhFi8EdOGcNSk92JcI9MVszVcyovuMLIR1bFGOQu6CAnA0ncUnHOzHN66uRBn6gs88CG
TVCMrd1JVhTX3ANbU99kN6n/frTCXok87zH00IsV4NXYxfPMWPsB1dGv2TkrgA4gN3NSZFvbKnSU
GfuU9mF7R8GSqb8XXRBd3r53gvmRO0jOLoMajTMBPIfODpt7GAFOhZ50oyBbYJN6NFvHENMq4oVT
sSoqXGoqrVuyvVhgHBc3Gum4UmX+tgkt+zUOhliqUrehvK6Xb5E654hWADyDY3DCQ0CZwkQzdevT
VUkHKl9sDB5j9DEF9KuaFxZUHN6Fj/L2dSRMQGaHyAodi6IRAenwV61ZNLR/zsf2KOU4JSJpTcN/
PHrQ/jSg9/bWAekGTSOvZYTfJdKsLK1v/xi7DxyrUClgaM9euTaUd3SUyERuajcSCDeBgvpCEOE0
i4phMoPnqRjBFjRo3X2NFDo15irV78OvJ4zhT43tGeq8q9z5KXpLKQx7ZjTT6Z1AZWAeq5dbkiEw
+OouWpkjGTshHcMLmLQDahI2eGQf1Cxu0fj4UxyZBSR8LTSWGIjfXihKC43mzP/AlTjW1Rr3OUE2
P/6QteH7pKmAeY6XNxAns59S63yCFrSEXY2KUf8hFAv9l6kFRrX44yMJmIh+4zF+gubYKuONkd0s
IOTZO3E9MWmxcsYWGqfnEDdfb30omTcLbj1yr/1RDe59nAUqdT8kC74eQQAosvozY1fowX/5Gqwf
VjfOSMOVuec4NewF4mHCJKFqgrtlLo/2bqjyuqSnd24dAcDOqnP55ewQLZ0wycQfmcu68BT9oT5m
nD5N45HLDHRRQfdYaMS5GWq67CSVJXJ/P8RIU4DFoCqdIIc4n1xupcU8GmexwzD1/IPkWjD6yqg3
BQ73kVN4tNxPJdnd91d3sysY5m7+NMzUvqFJeQXpnYP8ZlOHYhCdjNDWwRMz5pXsSdmfcvvy9gys
b18X6hqQRB2Hi+pqNb7CuDmWwwteRgOLJ1VP4qfg2M8g8laOLy2vjj+Q9O1KPXCv7wWp4u2VA8V2
BDxlq1AnQVoU3y15f+QlrUmElrBOANMaseJVPdMcYaAjEZVflun7RG/fPIjMV9rFsuS8QsTB4axO
aYlnHW4e5LdiUWayEtNAaPZ9oZdBhirIhfMOdokGCTIxeLQkszVmgxMmJQZLh0izAZSNLVLblRfd
2C9b9BnboAZrw54If7wJngIvV3BTDMgaRvqv/dp6imLxAi7YRuY7aFrSTYJ2V+lD+Myo5JBlMBFX
kmEB6TLF+sNfzYyreIo5HfSXqUrlR3VlSaoleCuJ3fWdroun8rGdKg7t7VT9/P7bNr5d7K3totZ5
tLz5KdCQ5/PH8GTQI5h6yNYrBp3ahJuqRJTHDqfzLOVtZzkF4sdWrf0dXTjVTYiqE+Qu/U3Ue7+3
HpyJahO2WpTXGttk8qlxxZuw0FKrxgk4RmFRNYrLuYVBsTuOO8SzxOrT8apgOfmr1cAT6ynzD1to
yk+CFZl9rqK4Ia4ewoOaI/PtNxQNvoZFRhgAPxIORuYmvF9h6xpEiKIIZUgbigqHs9IWDhMIJx5X
fCOQXZMvkR//0pLkfkQJTv5xAwDAq96ukC04B8MF0duxV2MxJOShsZOduXIpSZARqBBazUnxTrSi
LiWs/UX9dwJfI2EOykypkHYLkamkQBdPcfxKAcP7hEfW+ENsDDnLM7gv0/EqAhXYLTIhWjhUg7ag
e0j6tjPJ3WOGj/VOHWDw+/xl+2rwKbd3KFSSH/V9nbypwiX584Ux+/qJEJIXpHcAFUwZu5FmNMcp
Ix6M4RIGJ8lLkLLzh4DHg3aBc9iB62Bnx7lOcGodNlq6IJDJPrmoZq11SAZnV6xrY4++ljM5D8t+
NPrATYirRqkSOmhENL+YpjcWtKmTAB/2DJJ2HLce/fj8ch2ubNRPQO7EmN2EHVxdA7S1k8e4LmeD
EI4zVcb5wtckPCkYyGZcyrWRgHqD3j1k1s1peNsAcFdtyWhnoS5iq+2kohNZDLEbjcW2KsEFRG6l
4KHssg/wbvXpmsybiZ1Sr/wMNbC1A5Gks/J6S0y5ahIbgP8+WqVQ3MZE08pxVB8INUdDVBHxXAik
DJcp47ToeD2gDNwPqpqrv6MO3L1Z5uT9UMhNv53FE9RwzSR5PaDNtMvQITH9igTqd81KqG/brGoW
y01yNbGWN9RhPBKJwl7kKm3/oeho4wDFLGgUP8vPuHST7RxR0ivDT7izwARNAQRocQX8dmbbhTug
fYF5AVekij8495Ejv9Mau4zYL1Xrnqbc5WKWyRgoXVLVGYyK69U3rG8lLzZdj0sdP78ZhjQ27aaI
Z/eRqu2nJfNqwL+DF83V6RnvDTqBK9/On1NVfPnI2s3eQAAWUkUwdkiMh115z5eN89hGY9bMVP18
17sMd3vdKhd/U9sRM1Pu+lg7HQgPiowj1OmYcJ0xuGKDinu0pesWGk+MaBuS4SjKYzh9+R7YA+JU
Ld/wKlIpQcoP9DO/UafE6iHRAs7ffZ5bWtyjwQHYesIA9pyHfquxUvcVAhbTykuqPsAzY9NNoIlb
JbMDIbvPaNG+dzDoHRL1mYabiLVYBn2GFh6NSXy03MUybYdajEgfpZtx5e0PZaGXkfa/JQXW/hnU
AmYRIDaf5Ed4/45FIXw4WriBeTCAVeNMEWTJFXEMIEmIwNofHFTOQEGRk8Cs9HVolf7E5PftRe3J
zppQdpZ3wEPwwm5nRd4mCv53t/cRfIOxy8xhvq/sqq6CHssaTULoBAXQ7JzK3MmqA0Yp/1HEXrqP
WS4G9xMOu/VrTzbaNPmGnWokgwYoWpQ95XAkwyewEN0yxgrwD4kQ/rhYrd2fTvCK9h8vxDOetzAd
QIsGTGX8VG+NWUXmNHPGIoBSA5Oth7j6SABUYg3N7b625hrEtv6gVv4mIpXRMURy0wSpJWZ3xVK8
C9VZ3cAC6Nf/iRRHbFLcDKBDKcjCkbz95Zvu7V552PdjKpVAPFTAJOQvlYtNijKTgYf92Vm2ro3h
otAG6IYEsONRYNCdfrQZaOTJtz2IQtKfIl2Wa44RHAoDDjgOW612Prwf3S9pA14mjtJmDIucPaqT
L8epvQi9VPujqpNkkHNhhZiv5PT06PjPlh7MhYg8K3926D+epBpNL2RZpgQ8l48gMZ66o7zWWcUR
BP2ksoXKuSMLuzQlRjxfpFiYiflUwUOQkJ37ILQGkeEVhlkov08jvt5AQK2naoWSIz6CsSfc8C5h
SlAf8gqfuhHC4nM1s740zKsmhnKM3NG2HKewiHQlrsAGp6oXcV1BEmQvKLGMj8kbEAzuegyNssZn
4FUAeO+RIFjuJg3LRYW+PHmcIne4zD/fHL2CZ3J4fLVouqPfE8LOlE3jYtcH16dPd9zA/HeQRiGD
s8sX/Y0esUjIXYFLQoAl55IOm0ZPZ0VusbalBjQIsiL6f94N6E6Ok7og4gdfSoBxULwgMrKkm54K
vAssEs+I7rE8ee3TOegSiv1YeQ5IgbQT6zB7H5Es5nyzS+1PDCEth+9IiyKuSTahSexrdpYrhYhR
iiuhjqxDvqmyaF3Wa5O43F1X3eCnMgfMOXI+On3MnucxDJXP5HWkvd2eYWCqUcMmHSLNgd2zsVCI
CchLzQzd/He5zTqjoiLboMK6K1w9Jf3mSCEXDhdmez1zy+CBgZyT/HW18Dxt9H4pwTy64ZBw9MA2
ePLYk+g7DFNaCkT8TidEzrg2ab8SECuDVb8Yxvj5fisSYVDxRucBO4Ytc5AhC92VssC5oYTgMWl0
CxQIheMD7Sy+PFtAiu6qclQ5Y6ctWNdWnXjd85SP3u4TOmB7bctPTerOtMDLf0M5qt7PLdnRKBNV
Yq5oTNxyQGevmH3+P6Qji5PuBR/wRWSYuUJfdpDJy065Ud3WU+0WK9boqgxkhVUShjhZhz/9mfNY
5iGz0Du2R9325GC6J8GjBP1YDN5LBalPJdq/zW888rizC39ZTy76O7TQ6KT8rG+WKDe/j89Re5hu
/lCV969U0bKgq76OoIiFu7S4pZfkaVvRWd6pIsGdOH6/ijZkmfBLXXN1mT4ZwvliML40yKGGWKhO
VNmLCdQqCnDNdRByloh0nWxP3zIqwUNwnvIAEBiPcw0qLTkP7Cy/o9js3PSGg70v7+LQk3dK1N51
Z0R0om0sD1tcFwr5a4ZV/Q/z7pfwTndagWiC8pAn+/Klizjq5kSLIxX7mUzOfta8DNihnzUTpCdZ
DtUvw7ICLBEkZXwGbWFqLZKf9pclNgNqXFJNuyG9KK9F01OuDDpGNPXU+JuJve3rnCUoG1Y4dT+9
C8HuyCFGuRumubA4GhAdt6HpkWYkFkDCLP5RRKoc+W4CDMpytilhE9ChfjeaMSVFDnuq4QIrkr7C
vXAgJXWqJsIJjgMQZniyqVXMGeQ41LWenkARgHOpAvAJhaJdkpYGxNPeCOgHOTDNx5TYRwdd5Duz
F7pEeSfGQFZRmJKfarfTvmnitmzzqwWmW2xeRGEPAmTULbvxXfteNzxHhZggnINjPctUJtR+kQg+
WhY5qLw07/Z7Qc6EgiYRCJr5n75XTdnWfu+9Xa1LzUlM33W8Pxfm93eObR3ycTjYSrEYUAZXF49O
9sYmdeC1x0pPI9AguAe1C4IN/PCRD1Vi5mNQ/A9lHLtEYHJRXMAqJNCvNDHJRjEiaRemp3ggqEls
MS6dUzQrB+8WXNrI8xJEi6a43955MwP9BsZzqulzw/UlUje4DX3rPkuKiGu4rfCNpHWiXNmVTbh4
AjB3BmYxY81KnMlvxcUrByGtBjZWoxcskQyAm5gAnKREMPOed/PqEmeoI3AYPY7IWFPILq8csFRA
7LmcVbIjyDvfgi/snVU3NwxSvC4utcCa34P7YCv+18WP7pNspXaseHscUrHvhJw4KzfQZV7zaj16
HTSX0ciySIwgfeUDqNuWHdSyRAuljyGg6bAkW2O/B1kuhTXhkfUU9oq9Ej9Tc1Qg+FIo9Q/2msP2
wSPN72R9UIsUMnxKe8sX2uzcuoLY8lMsyySY6xlNCizKW6rCFJhESaBJhBewMiqWPXdkiVCKq1cV
xnkyldNXBUfcd/v8J6SZIobzjP3S9g4z7tW9tMk6VzYS1aP3vxo3EhW8IY6PWM9VO6lABPspGOfF
kfIoNlJAEzvb7nH9SjoFyvvlRc4MToPxfdnBG6d7VN9n2HN3n80g2aohW05CYeoNGC/JDQKq4Mqf
sMytwJZF8ODNJroXUATIpn0USWhS9Sip9mccHJDv48b/ku4PXKUDhvzI2bBLV8hUUg2uMlAULvA6
vVa4W1AtIZvaxIzjcAUGrzixoT24UUJFpXy6wYTxB+6RqoEFMLxQEhZgzsifvzJc+rQAty/XAosK
6GwqGswnh9pDWhDYViFaewv9B/W4R2hGcB7NjDSR/adO28xnvcLoFGUylWdgt7nFv3hJVz24NXJR
I77d1pmUoMXpdYvB55JUdofwMSaavEi2VJv2wNfocsogdq/O70z8zOkBq7JxUtWzrg1TS3EWJXi1
tGUM5JEekLW9Kx0sfuqkdXfBwpNdu6s9W/zADPb2NPxe7fhVLvrEw7D/rOPnuP/4PPPf7Y8THwfB
K0DGBcL0cxae8bS5cqBE1uUU1GGlKY99aSmZiOjCukc/kj4CG94YUl/2K5l2kYYzYf/KxXNv1u7q
OiwnJQcCbAsAMkaQCaUVUesylN0+nYd2+0imNuPpSmFTiE2bzovIAfKLXkaAs5kQySWYVIoKCEwu
p6bwaCkipm+xYYIcjMiAM41dMh4CKoUcZ+K2OhG2QBWFmBp6/P3Rwf99fHlIwRfL0bYPANW/FdJP
7dmXst0ZwvT0Ktv3L+ugjvK0aZf/wFlJxmBzxClrwoB5Lr4coVBthAApi350mi9q6hGhpXRAXGZV
sX4DbjuclIMSMOU9xVQBio5fO8evwkRduwwFD6gk8l86iPJge8XnZGgTMb4wBxJNANRijBvdri9v
KO/o3sxRulrK2p0Oe5DxX9+TJ4hMxYVQ+p4Y5fqt0q/rIv93j730PG87oEkWrUkGHDLwdl6Pq+ZY
8yBe0LenA3BSONUrKvLrbzvK7t43CQG0M+lC+Y412RVW6hoMsAQwravM5QQtkpBGB2zxZ4zHrxRt
8w25Eq0rcJLzYDQE/bIPsCUDQBYmjXPNXnP4qdFCCSd4ep7AoKKDcl05xrGbV6m1GeSVRlbGEzYs
IAqEg+4PDZVl5xfVDFT1lQ1stdBcuF+ncAiMRyPRdBwu6E1FTu+gRDNdL5UIpv7uwm27IlAwwW59
Um1QKbLjF6UPfrxWOnQ8ty5WkCh9Vjwct0UPuZRHgkFKg7hQtiZE4xrOzcG6qCcSkbQgkcS2v8rm
JQfbh6F3OrINML8uxflpFISN2GJaKz4wG+bNzG1QqLxvXaU3VRi6DyDC806FcToXgA5+gd436JA+
N0zXUpiKnD+pq1Pia6vHbFdSxldHCYoeJgcYV2/UduLqo/BP9buEfooOVF76xFEPBJOEo3yq9u2v
9hJZ1UGPXH1OmZ1cGHMi2fE/qKhkLjdBkW195f6SEaSM2EF9/1MS/GeeWpMCT2SMaasJOI+5H7EJ
qIenki/Vqxt+dkdcd7xvNbFWryemzcboVpL61BjE5w39DsNdoZijtP84An/Ox6L9esHFH8aW2ysS
Oj6ggVcbZT9ElRCYpDCaR5DyMFus9T8CLnxb4vkRXrVyolC+6DsUi7WNkzwdmdepOJPEoZogpZHL
EZttLUvpOLLv9UZxZE6CXPS65E+H/59YqA97SQYU2zLMPOCF4cS3xoJyHjjKQUx667v5ZQo5YElX
e1e/CIFj90jHsHwzbXfIxnp99szR7XyY0kMx0XxkGH0JBHO6AHC66SoAHOMWWq7Asg44ZzUEs1rh
oy8XJ9YOcv4KfPDEaZFSjxKvpPnDa3iaqR0O6UIpPWd7dXVbo3kYK6eMayajQDb9+q3DKOU0hFO1
HibkhMwqvCMkjJg1A2Eyq9QmEDIFWiHmN5aFwmXpA2ca2+sQ2EZj/oVd8bnIK+XcUOhIzZeIWRCM
yrYNfsfZsR7LTPATAZ/cyVS7cac7NcWhlHDNE2eLZAAbXc1yudI307MK/+vbD2zi0GRRYHrXE3Cd
uuVA3u2b+kCQhbNo+95sQeYrZhh5ZCht55SXm/KhKlVryEewkzRyttVJmwPdifcd9ZLSkfOFsj8W
AWH0cOW642TVXsnf63xxTVMkTJGi1Zil+6DajHlK14KLObpTc302oMQNtzqfTAyfM5QSUThuADGy
J6zgHEJqwFcp1biZNiwhdqrYObV8/cQhMBuDjJcbjlz91fVg4RzizRQctSekWuLGhoOzogJhe5go
l8s1dJHzbugNvnCaEMqtlmKHO4b6rhsTvXOmeH3RcWMZB3K14VBtZ+Us7p5ofMdVDoANdZw6K7lK
4ooZNGzDrZZ/4aBawFcHhw7dzSarHuDPxIafuhYrRn0fJNlL4xcpMI/Se8rPdiVv3rD7714EbdlE
FnzEt7X+Ejii6nCmxaL98FREfYXHOK26FIxrbrxyUXwIi47X06J4uazZBcAYOEmqSyfahncb0ZvU
VClL7eqEER0m9ZmHlqSfem+OOhk+JUF1ok7SbmJX4BPtinn6Ostk1Yi61C1vrIfCO1n+894MrEuh
xFVYIaU4wcAGqmhDAv/Rned5EaODxXhLFnQgK+OHBMFPoxrUes4zloj3ZISVGZldV4g06Syf3w4/
ZK/+g6r4jf/R8w+UMMVMwUEqwyTGYUC4+lSZIZNJtNIqSsy/E5l+Rpn11Ar+E/5EX7B0Wc8S8pIS
J/6AZVbXO/oWP3Lxjwvx+0h32ftVHu5sWwVfWELxeFkhtpeNCqOEseKDvv29YSLkgjW8EZkZz8ik
UxoqXJXqAmESqMqdqv9VPOokQt2zMf29IxPsW71Q60R97PwrA9cC/XyEhQqlgNXFRIZ42MZX4Rnb
hALdqi/y5MVA664jKs8u5/ulcsVz9YQQLBJ4Tq+90em1i7Dp0CccMryvSFuVCeSxbbnpu923CVXr
HasXxfJnlXmJQwf5gRGle+LpgNYcSlxh/CvXwbaRtYyDqmV69+jaLiC9h1+mLbRWOcRguGSmxGcS
Jq5HBHlHo6pjxT9yiKZCprr75w6pB2TJWL82eex8HzbRXgFA8sIUMgIVRic7AhyX+bdMWONmbykZ
lf6MIker6Lamw9Cpb4JZjOMddAc8ohCEYD9WlAt7cbx0edmA75Lm/ptVoamxVkzayIzwGXCALmca
YaDkeQSIV9MI+GCBxZpKwNFVrSsEFhS4jXVM0B7Fhg9yuDRe+XQ1OIRYaxDH5NbGqReabIdGDXXo
7tgj68X2XxKYTgWAkOX4nxoCRG0mjNxCEbhRcP+bpChzgkO/gobwov/H+uJQ2SZ6EU+ifFd/CJWd
gjTiKy20W5q10Co19OIIuGGuV/7mWH9PGMq0On2+d39ap9D6+gU9fRgjSZgMLWQ3qAaQcetrXSCn
AOVJ28NDuDHjCDEbzT1PapgEKmQRMSY4J/zK1EMTRX08ODCAGwq1uZ2RPZ7I1R+wS/EjSxFdqYV0
eudxZq8GAA+xS1ltlnKB+VKunyIXLaYomPpf4I89Lkp6SKKcwixaeddTJSf3JfPpjoEpJ61oUyNY
yAzM9C3RNC9I1quwAljx+TQjuie7G8HXy4HWKxjuuHeTZHYkYT4LScoGTXS8sEZlCgf5TnMgK1re
hnttkWe8V5zetHLWkyvQZ8MMERXQeJNC12qv2gThXkgN85tWRUNxSdTIZFZiIitZti13WhSxpygn
iig78TE6bAOUUk98A18a1UMBYysw2z9245WkySOLxthOHmyJuWQU1H8UcUL2WeE/cLj7bS4seX7O
H1bjI7wQGF6tf31cIJfdC2jxtSdlWNKVi1IKxL9x4kFQmajbSJUgoArCDSWY/ZfW7ySAaMgmKiEZ
JvPa9jtAoUDV+BEog0NfXOjbRL1vbCW0hQ1vD5hs5yCMniLDSsgpgAJ6hAW8r9PfMQfu7HXTyqus
8JtaTZx0KWs1JIIN1q+Nb1SmDdzzd17SPOp7DI36g5AODWSVsq8xaBfDCzx3dvrZLb/MzxpCGQcg
BhFjvGOI3G5y5RuP9qP1Ct/eyD6Ogvdlx3+ydUc/dIwDh8X5JsDQdjfruMVaezjWHdUv7XbXiF3h
OJh9/LryFtmFa5j15Hjkq2ZUg6jJlHI5m11c9/hDKzeYw+hiRBS6ZHauzlrvtsM+WtBm2MKJa+0K
ReQ8c3HqYqpqyWoMVlgaBRUxF9sfpwgDV3em7Bmtrt7n+iZ2M1ulyQj3ANG3KPRzbpjwnhfFF+Ta
BnG/drkDG/EOTzyxxCyvsqHrX5djDtUCmcflxhBG2gqmYi+nwW794gWqwPqzV/u5/8hCYiChL/AJ
V4HEHV1oadGbsVuPiHb8mXXjw+ZIpitET35yD8wT8C06nAPWwf76dPk2rCm7vSayavaLU4iyKMt2
UMcq7uNueo6XfcBgzXhyPm1tWjmZZ7QGUWW6k4AOMHx8bHr7dyE7b2rgi24eJwssEq+6RbDaRqnp
DZ20j0dyU+CX3e/lVtvkbbEaFhMmqgDWQb419bahoT4Fxl0hYLp4FaiaiWtFY6iZEsjGFPUgp3OI
vbETSWNDMq78+qr+vaGcYT1ggdB1p4dk+q/LGACumhseL8maf0bmDsbDEkKgdDMkSptmzGILZ23K
PJsSA/bRGcxXV8L33hhFXTZhE/BJr9z6GpNsb+iJtbT65QxlI8MEpR8SegQhNOa9pTRQ2awE4/FD
2OzeBn4cLOHld+EgFT6MENRp9YlCSwvTsVYfYH3UVa6RTlVTxzD7jExWVaBdoeYqXClzESA7Lxck
wosm6VejrhN8OYWQt12NTZxaIz95BeQ4eiSwwHcw6/eIllKA90P93CCVrg4wgdrJbXroKREZpb89
3i8R4c0uN/JFSCEktZdg80j2SBdEb7D4MecY43NRL4WZdLXEsk+t5fXVZMmkV1IpFepgEQhZ5SYk
bLQgOqBUcOJLLHn9qWwxIiRk12RatIgGUKdWe5Vt4BgNG4BK6G6p9NFcIlg8c89Bs04wZB1GLmgS
XPIb8jcwHI5cGqVCtiTe1yy37vRtM+auUmHKi1x8NEpBpjIHp+YG+hLhc8T87BuQCLSd1OGqfuWS
vyPBBO4GpEP7vRvsS1tlNDwB/WcrAnEBJT4baAm8dk51vD+Ua8aNGYCVchT3ZMFJ8W4YoZYgFPnG
15/gg8FjZy/hyNEuSdf6tEqA2cXusmao3R4QNySPSQuwGISLop0dMj07ALiPHSx0XggMd0HiQ6x+
0YdIw5Moe/5IiwWB7jD+Dqz1qlnfTuDJyhEzDyO6t/Ms9U2PqWySqmCNJ73chqibAE7kVqhcWQf5
EIpUNr91d0mRakQTjsltDqgtpFEQnzVh9AvDDEzACZ0wcJXG0X3Hbum7mk9F8//wLJaPObUPHeGi
DQqULpdYKiBum6wsYUy0ftO479nfL3lH1W9yUxqZb9hQ2HbTQPxehu3qVgL2cPoTnn0feTR17u6m
Ka4MHS07D8Kw0oW97UGK54H3uXBQVcByuk4JLfL24fq79+/ldliq/yznCSp7kVniYRuR/8JEcbXl
OkTNVkMMgHW9vdVKjy/FteWFdFNPdq/Z4BVeSah9qEUa8zDqpB8NK/3LU2j7k0f5RUOfUdRjZDIg
15Z7BUxrOKqcRfUZy/uAcCqsTttae8W8FBHWgLud0BfSpcumFGIaeloVcMWgY5YW6z97qxRaLjZN
A4KSkwLp4jfgpYYPJwVWbjcvmYcqvCWgvInaIVpYv783eKvkhE00sDL8bhLfflZBT3FtRLklcw4G
98wP6Z5KwkdJIx0KndH85Ed2ovQ1ggbwLL7vbWQf++NVtG+h2JHnLwAWrRXyff4MhHcDZEc2SY3+
nywh6O+z3KTj+YhQBVNUasBma5XTqMaZrj0OGrNxnMTanL+BWN6wH6hGSptuscOMIPT6JdrferGG
sSGiXOVh3FH1FF9lGLoi358BnxIpwxRFur2pFmMLgMrrN1urT5uqAZ7qgEgXEHtKuCNmu4tJ70ui
y8cHV/MMLKI+b9x9nOBtyqH55nwkyv1B+pYHSqiq7rUXaFdjdzUuelqgVNufXjw3Kx7D1CwoovA5
ZdEYhxir0JGaDRC9U3ukYjXE1XyW2LskFJgDK7M++hz0IptvJAjlyLBATEEuO/c8wr3RA0zyqaAj
6yz9CDsmXcta84QRvT/r1JpX0r5Xvmk3hGsu5Roy4hyXNHmR61cJbGfhoSY3x1Q1IRz8U+ju0h6i
KPrX44pXhaNKl0KaTlQN6gkXw2BTmI1Ff2RF/VmvFPW35pmXJZSW44x4h3Awsm5jF3SXEs3LWw1Q
d66JSpwdJBgPabg8U76cstgi9vKJC/I8QlvLsO7JNFjMGAs0OaVuLHS6gx2G+Q7qz13mZi4hRqj6
eC3mZOVjEOdR2WfB3nFAYvSHLoiorVqnUyxQCkTpIbOMf8Qc6Wr3E7mOFnsD90Iy5LnC8C9Esxh/
qLm0igexsFDM1ch7yFo8NhR2RTCEbk5YFV5K76Hd+R4gsoK+4ESSMQAmEej6f6s99wcn+p56qgMZ
NJ7J+CpiuE2iNE8IErHunf7wik89Z16JdmIWGdyjnZloVxnUvNEaB7mm7dvtHKrk7RCQJCqWnMzM
9x9++IPLzF5cGgrHhor5v/F0Ii+wXaJcv/1XJfbuH0apueEEpwWrlUC+aZorpqfnqtFS6TTPUFfA
xuuuChkYwYz3DXYVVy3lMw+Vcil1hroag8Rj0awRZFU9DQYxn8CUTEHDnYiNWIbghwr9DEcsQ6bM
teJdPQmQ/10k5iUWBTaSmctVMatxxELgleCKXZDD732lbpMsBiC3wat55tVCveGY1k/mQYTYUH2Q
lU3j8aoeyQ6NFmYVXs3r+t8Upvv7AFrWw8FMOz3p4sweq+aOnKC9FMTbU8Y6vsae7I9n+/b7iegC
8OmNWoRu+SFNO5aMQXnAq2U1nxzUqYcx+NFdPKe+OoardWV3M25Kn5M+J+wiyKfMRk4CKPf5ftT8
Qio+vMKVUyTxbxvai24J1ZcYL+1x6Yiw/kjRe0M4b5aFaSUPU9mdSF2maD7njjK3lRJyN73yT+Vq
UdShtZZFfOz1P4+05mhKaBZnufggNCpWUtf4gSitQ4kYsK5B2TbeyUfDsrrKohr+ZMiotcbpWOpc
sdE5T31EQ+QpX4HlY/Ha1STZ25TA/Ts3/0+UfbgjveFo+vTj4ygDFd5CmWCbDmYjzqQnnLYsvGxE
v4xajWNubi3wY45MW8yeRcvAI+1vsnILQBQuViQq0PKtqMgi2syRVp5S6A43QmQjjEJVGQlJTcKg
CUeDPcvoCN3B1gsvYzGgJTFbdESMDo9JKoy+TQfHvk8pPATO5hFTquqyrpuivMTU0IglZCMCStw7
CxVZaez/CPYKzp399wKm+NEFlU0DrEcn/9+uMW76g2h202mZu2OHpi06a++7IJTNa8GJT8XGqdvJ
ds20Sd9lncbQru8OVMbhijVd33oIxQJdWYMxtyZqBvTW02DJIMW8G7Iwsm3U0KWmySONrBn7a7Ij
SjT+e6zcMogQyudjYjOe/nQRhjhkogYceAUhqNhV0+9nnIVTHdx6p9FSTxe/tndpXTA5/V/dLxKn
p0nRSWrAOKbUZWVsY5Ye3FpC9XwkP5/mA00zS6f36CfNs6o4XbN1E5uIK00A7KBBO14M9ON3p44b
DwR0cQjw0w5pRJ3wUlMLGtBCKGdz3dE+3N8nHu1+0NlE5/qJVU6zpRy6RoGyMSFy4t0Sj3qpuQgp
IsYLYu90R7hasxzTkrsjRaMsFZUz6Y4uDozebUmX8yqFJAKgzz3N+uesyLUGArjxc2nPoIexopfT
76irYPi6sxTcKulgMMNBx6l3gh1U0Icu6IW/RwIW0rVe4scbdS8zWyTDmSZpZIfx5bTZDxRzLyB5
ViLjSV1nHKpWpg+C8Q6TFzmHe1TevNWl3d08oYU2KGmRKeuIsix1nJ3x2MUKsxyeMqy1xP2vQBNR
3gawJT8NRkPArlfZhcz1Gx8V9s62gkus/2IWWIwZJx9WPtEHti+NTBUYDVNiLjup/odR4+Pmtsv/
6kWxAlVJ7YZ+p37DjfpwsVF62NwOrYNRhONHS2fu5bbMLC8TPhGa9Pl0q0Jw3i2foXxCHv26S4gw
dADxF4vhyRpSIeLuxivxeCBEdrTdZsaYxjBvXx0bNa+8rTUJbqfXqMXqMp6ZFgt99ZTt4QBm8578
KwvSvhiLLvHm8AJ/+6vJ9/K9rgKD1R7Q0xVoUvEt7VexlKg9awDynSar2W5GDcWLdF45wWqMEzJC
7rkQnZOThmr25Ha1cod5rBsOxcrNp1pQlTWz2SZgO1YzgABpRzUSkahjLorbi2TuRosOiDOHWZn4
97vH8YZwpWRzVP+9KtiiyprQC/E2hP7mYd1fC2aYiIInTg5O+WWLoojspgZJmnCf4394XOGdJ35I
oMP2taXr67azhVaVTdTYBeIGRjHs9kp8SFtYRQtbmZZ+MuRp7Y+cQOCsA1OPNayLUED5MQgQUy3Z
iagJaCVAaSN2WQ9kMQhzaly0ADyEBKdlNA0dq9Yh7JD0XjHtz6x9nf7LPxTfYDCHoStBg7RwNwVS
SDpPwHR91+VoOoB0f0A0K2GzSHQjiomNrnDe0okl36596aEGZiNaei0SRsfY4iYEJu5D8e2cPvAv
5dRcqOW86y0fhcRRo1GtK/MnRflsKiKOcqailF2zHrqL0osj4Pvg+wgCE32NQWRFhXU/OOwt6pEr
jjMxJ6M6ZXQu5WvZzQ+70pw8rkGTyNUtZUC76D177lRw1sRA5/aOj1s31mJH05P0OiTAPc94opIZ
z0vhkuB1rXim+COWFS3ewYduxvVRO4F6oU7/UZxpNet2Q7MVATkA5D16UZpQfsxaPp5XVhIAgcn6
n+vpjCRG81COFTNU49gQcZHS1njdoCK1VKazbreA2aI1hs9lmH0WbG9xwCoT1WiOrmh0ojEp/nqk
ShzZlLuGBHlLKFlQLHqj5tade8+7o1xYwO/eSPj5RV4WvnGtj6JhOoqXFAHEE64SNVNSiKDgvijg
kUgJrjYvFCCNkxddRDzRyLiUmiTsvqyY7rc6wo1hx8wAlFyCMOwMP/7L/WMJLe0EC2GOJG6L3Scb
HwoPBN7077OY+q/QWgk0OeMywlpe8+2J5r3xBcqmM/DXSvALE1/V9E8a6w2R+CXnMLgdZZH2bjCa
Y3uNOr8BOAXpnosvNgRWLLs5YdTsLvSAA5GfuArzUYZEl1DQ7hCMl/KwUjslyfGgqpTBr3AVrzjY
lya3cv2rSThm+SFct+H8TYTHH82C8aDHj/+1aJ1iq8XkVqMYCRl5I0sJfPpQOH6vzoHPe+UUvc4T
7SzAStHuBLVUMEB9qUW56OrdO2PJP0yvSzZ+dMqRllq3WVEiS7+5rh/cwqin8JkkKv5zQjzaAhtw
uzM5bkYiSPXWMvNKu/qaWEPyX3xdd9/rlKsiLQRWWuf12f32+MdVvJO0sdmJLqhoS1ThGljNCFNh
k7DthE+yOEZWccSsHphI0mMCNpSAGkAUXqv7WhOvZX7H0NtVlDnlYqTwcImHCdIfxtGsVcoq7TpP
rffjaebtksruGhvg8LwEiH53m7GBrOli8punjlNC3Nk8qbne4Qz/HQ8ao1FDhdEKgBDwS/TEEd4q
BZ6C52BwH0QqaY9H1wUARKuc1o8D3q0ZmsXFolgoYsB7snpNjld3iTsGZvo7Gt5ct5CqPPr0nCV6
Axf20W3yNIK0kM44Xh1iRslJu3Og6MpqQMguFQkygXj9592emhhpkmYTnzE8mSzf+fJKwVXJSJ/4
h42cv8F7UUDKWT9W61R5f2zEtqlaHDfOxYmY9u9k/SD1qViNnCuEB5NW9LBLe/Cx8tywLi+IA4Fe
S1BFbC+dK+ki671gwy7UbdFwnu0r/vmytY7WHDT2fi8+da4IvmjD50EYAWREyazhzCz5rs+uxDUy
WaJMR2grMHmUQlOkkehmysBKDm//OGwgpmJtLwg5wgpuqUCoyHKyaGQBm19+Cc48rYsIiGucpI30
Sm3Jy7+G2jO1QXGEbOclyKvaqnZtVd5iWUefSGsH6aH08cyFzPEEUhzqQ2Yqts/vYLgXal11OjRR
wSmI6CFyE2N/4iZUmDxI6YFwFVHDfH5zYHF05ujXCGk9h2NU0M0lM31uB7DA/OhC3dZYc7at22ni
XfBp21uQ+1/vIWn8AvCtL9RE8Y+IxwY4j5npsgZ5k9L3bHr/LXvQZ/3WCzmBu87JRlnPaebZx4by
hID6ZBQx7vusRALY4n2AinCHNk6FGN0/Zo1dIeTeSJArzAJyW2jWXgaunw8pwxswkynqeJmytpi0
Quen4oYWm+opT2FpzmIXiBNZiNOofXCeQ8IQ7ffXkdhI8z5Nei7oa3QjRZU679BxHjkKw3vSFMVN
ahLYPbauMSm1iIttyyCOGBDndSiw9nbXTj7e+Vq1667tRvgXTsqEIvVJYgzIFGNFJVNwAB8dduhp
9zC4AeRnkuRGe8KHz2pOXWckZ3YJWPpgI5aVeSWp3nRSPBS2cXPGinbE4qhpsOTeJGEdjvj+rDBz
auHW7L7evIfWwlU0G76UIceanhjynDFCF8XXTR57jzBIuySJrpaeHDtbtKwyjrqVUHUIwfnXXJZL
GMhcdKTxQbRFw79f+1Mv9NG2SMtY2+CPT90c9A1JQj2h+IwfZszlccKEDSZhB/hbrIS5zkAaIuRI
9U43SpU3lk4QzNjl40QxZORWraEfSCzezUcqwemwpdQpOIG115ZPWbUhdG/L3HEYwJOqvrwyuqs6
m9kQvjas2cROTMpmAWDqNYwsrZuWx67GWfUSx96J9HBoFCyKpsjkmZBTChhlPtmKYMkB8y/LDj29
OZEGOrnJLGTtRoHc3n7mfAUPxkNzn52IC7hJro2qWMFg+RAqRtPVOVHjON2+xtyqoilE4BQun3hW
PeQjAHCvIoBu21FTuWtHPV5VBfHR5XAHkWnQUONUK6UZec6PnGB339lmQXuJ1hZ54ZICf8UOumv/
0KTCWCxkHNyXCt1WgcBBFEAdVcG2+jvu6fPhutVNBAXW06114OMiL76ZduJRtzj+YTNUUbWcFH5r
dXmgET17h4LWMq9ORKBivWjTVa18XCJRzuh6e6oh6HwFnv6zTSJXd8Fp5g56Ny57QPoX8upNzt7R
TKGG1tL7Y1Fcc/cON+HT0a5OVMS6BxdKIoVH2ETY6S5pcPm1EwQj/c/k9myGAmQHVZRE6GDCHsQG
iAhOG6oaxrJQ3pDj4q4w2inBK3TaIFGjrMqXiR4nV4qRd0RrBlujSS9CXgPhGPWwMmwKyt/4si/k
0SRsQ723F5F2UCtPoqTDreTCvz6m47NddMhAf0BemcYVwoR1i1lsF8fhUcB8B/3/ihsza7946oKm
BBUoG7VtVjWsTv4yFGQn6BAWis73bGLLublKf9N/UuqmJG+Pl/rFNwggETxfBO7oeaDNc1stFg63
t3qAjVIS/O4dVRcp/0KBu1oYgWX+gfoWDh7eb0nxl4KLlqeOM50vAjI+AmjBY299NTutCUossE4g
UQp+oO47ce+94YgPKFPEmzy81AxzXYNRI2yDmAgGIHGpY87R2Ny0fzHmZu3NWCWJCZ2RK21eM+I5
h6G3CgEyyzhIGHzQLK/Wc1CSc7U3w1xkA5qN63BiOeoEheovd0VR37/GJDEKVdjovINcWz59PL0b
SwxIK/JFMH+DRi8HkXAVLDWlvuENJeH3iDOSaWFyzKDvdAf5OTSz8FVRuiJmZNJXHNs/woLEE31c
1TjUl8DjaKNy7mH9gLac/QvxHz5Ir88Lh/UlzVpwm7aH6721Wo0fgyNf3jHIbccfAceq5eAH6es2
9TOd/pWMkYiWv9KntBoVpYNhMgL4ZxPHbTDzEJ9kqRhoneHoof9RaIU2EKfSK5/Tjd4mEsU2R3bd
JjNW3EwzK23/MGsHAGpg4Se65eGSYPYey9iQmUhkjlBALLQThdUIOw5BYF0FqgtdzuJJyk8yMYa5
2GBeaB1RTtsFqCxOZHI/nnv7b6kwg+Um9EfvX7cC/REvc3tv4X8aaXc30k3/1GoKOTHc5DKAs4qY
BbbbaG/Z39ZbEWii+cmmyHQWK8orA482q7jySwDV/8QIkBiLtU/3w+ATUKuGv+iddrXDR6Ywu2S1
H3NMX3YULNfsS6Zw6O95dOVzhpaz+Y5z7zkct+9K3BwVwaQegMAxxFxyZh0iyVZju/j6Wq3PW+0H
SAsccRUO7/O7rM0Ya1kCXayYx+FuHVk7qEJWJH1UJvdnaxXaQ5QwJ70rbkAknxozhjWoDj9KVdST
ndRM0oYwiBED8B+6DjZIqME4gAPMqn2+o7XUqNdrU2l8qB0gtcZA8mesrxAP5LTi4bcyfnxd6kGW
5XbTiyoeZFzBc64SWjjCtz3Upd8BHeF4LjUN2ZQ2+Z/8GOgFznxSlnTF8MYFgc6HBnj2hpK/n3SS
f5Or65BTFx60tHcagZile+nvDzI8bVU/E8PESvNc6DFvE8jE4+UAJ1JuG5oiFHBOAZAhXK9UZU+H
W0hv6+PJkpJAK6tLsEDuK3EXDFNVyyBKfrN92udYbPBEAhwFS8i98Hut/0S1inr5+oJQWemiRNnS
F5XX1v5LGYPpHl77czC27yDWKVpmM8Gt1BNKH70bPnnd8fsYd2kBfLgqthPl9iLOIpoLrxDz2NFc
LChjOk3dYRFGzraeuAH5zcMrCkfujUYJF6FJupUQYt7lmM9hQr+GLz0dFTaf4kIdkf4p9F5tEq8I
Wbft8wzvl2MmepXgUOCwPeyt5YvB6ijrsDyn3vd6NrSA6/M6ZFa5V5pP1skpLYISvhMXYkjq2hT8
mBvKstj17WiHWFSi8r/BvxP/j6Ut800A+zmd4MpYwbNhBMmyOGgxUzFaqIVcWGZNWuE6PgljP693
h0nD6kwKSDkR/eY5I0OPlPffpeh3VWMzDj+o0hAwUqYYjjXck8mZpnG8l0jq7EwXfQoA0MMlpsmm
WodaZ2ZKNV4B6GKGRv7VN5vkrPTs5Alk0MD3ZctnmzqxgsTgv7Iwwg+PEkJ+ktzVgZ1E40crECf6
mZ9pOJSf8gFdWb5JGIgh84Fpc1Y0vzgMQaSBYMi25mjb8Fr+PVFc/8S0Rbnbm4mvEmcqF/FLuARK
WBCNXURwfT57LHkDQOYxF/kkfM0kA8gnHxFICwb+8Rup41vcVgYCrXThknoP09DWCFa7SKuO4nXo
2g4lnbxEebfzx0SOOUs32oAa2Cg9/JMr90fp+l8njHI5VBl5kE5qEZfA6fXyDlq1RJHCitdNMzTV
6JesAMO0pA/+7iRnyvyvrLniuSiqRNG7XbDxEPdtghIU+92NvEDcRDWZY1p6BJ6+KJ6RQ1sy96bW
wQ3gY3THD0JZrUGslz6kwpn+Ugwm/T50GHZQl6ArlNkX2LWgAG1cI7FB3PJiC5ub1/TY4Bsg2lMF
xRbwcomI+DgYhIM6ZlsOno84kfdr+GV32W+FN4iEN/bfKQrAP3ZR2FEhuFVi6XYVCRR/g+u/vX7M
UG4KmwAohxW9Q8+/j2z/pObmjreY968BbPQcjL8ZSQ8j8DOZwwY3aGDEVdJBXnDWK0mu7JiwmPax
T0BZXFOie9ks1pYWrBCq312C0JjUpnELHRe3hLpwHwDFuPsal3mPg4P3VVAuE/RBu2bAwOyRMEN2
vDjP2FFTzK45C0zdtNxDIQ88fm6SdffyUgIu868wJm7HlA6CHljQrkfTuE9Q1RwiGbLFHGh/dLzj
gJ+PzXx8lJO+Xcrv86YgGCZtQ0pCJ+ZroGsF1cZ12mB5FuyEsBqlpmHWq/4IOYiWugjjiSStNgv9
xIsybg9NTAQEGsZ5tE9L+mwrpRGZ/4IyQzuZvhZIMnmFGPulGr1Zg+XzNXoajpg1YMyUdGhM6H5k
iHgApkbNedNFFTrBxS/MHrIzdZ2eVlJJYqL+gToII2QuZhi2R2fJ5GBcjseOivQkzEBLFozeTxKO
pn73k0ewO7X+0EA55yhh7izXRKxW6ChFHXdHOI/8HIhjEz7q1pMj1p/SpqejYQVEJfV21tNdjQZ7
Ayu8TscsMMCaAkjI+LfeyVmBY631G8c9I2gWQHTy9dl0SjKgy9zgDw9mZa1wreVxcR8XLzFucFr9
DABw9gB24P5h1rOu4GTJiHAfyJTmGyqB/iRTGDQu58fbZpeM6FqzXu0xlGBHfuFC56iTTotW2Mu2
DUZm9Grold6AQW71N6CB2krNQ35w7KxppzlTRhTfHJgXjaTxt9tFx8d/0bHEkpSsc+PZ/zt1eDt3
Y2fbXu8ZfxPl0VFWoutGALpqkEKTtQ8cfUerSaD+vjsWmIS3hfcLJe7k15W7/nhAJ/weBPO/lmUG
PWq1o/DbwCGQD+T5QTaFB0qGLkDVMaupKbZGOMNpL9HXgm7MlyOcuVNYE3y6lHF+mbAPxe7NRXJP
UE19a+zDbbsFjI0SMrTfZUa/dHcF3rqFStg78HzB9BqdO+xsZH2l5hnL3p/h7RhNJblEz/4iNF1K
WTL/qEIQaVL9Kp8if1jXO5q65mwL0/Vo9rEmdAF1dxEOrrrauHPJeF86/B15UvpMWKwydPvmA86s
xYpIteBb6KL3oDW64rFbzVnuzs3J87mGvUUWug0YmzVbGuyTpy/LzKRIlCKA5Nhu4pmLAmFJAUzL
hdCO5fB99Dl2RTcmmEjzwkLNbhzgoiZnai+72y+tAERCjKSUCU8llFH/1bcCzZv17x7CoRZo36sd
iT42jr5x/oEldjm+KCiU/zNZZHSyjBXWyZkEem+Lh3W5GRKtNw+Pon5APDkOjWnySzb9yVnVYYev
UV6DSjBLbuWz6sKZFw/tqb+gpf9l5AS3t7iYZEEL93lFiIx3ReJNhRtspkMMWznay051SCJ+ZYd1
n+TNk/D0/WARX5kWIDmV1gF75U54Jbrb8xsKo/I+UqOf2uvaraH44cxJKqKTlzrhXlR5Yc+xZ/O+
vz2HR2fPkhcoicF/FVW8k959obULUT9ipeLGr8/Pw6FmUm9f0E7w6D6x/iifBjXv/s/ML2j7RS2q
Uut9LAR8N3vxxTecvy6YuwM3ZtelFeqjcMOLwETJObEt9Mr4aTaolEYOfY7ZybIQ0lUq5/wgXypa
D+WaFTYCcbuwwbTy1W2aI9sgR3cJbLFhq04o+2nq1TNaQGbQOevnc9EonuizAz3RKuWJLhElFu6H
ZC5DKbi1QgyOH6+32nWWusnPAhQxl3XjrPkUHNNqloLzrmXgQ0JqfeAP/MXI90y5yqSU5nojbkBk
gUGbagUH7gw6uSzUiNlFV24/lx+Do9MWfAfvgYEMk5QkrP40K/CSFsWrpqcS2MsHcXa9WTBdOsnv
XVEfZX9C/3rFaHcW9r7fSa6E37CxnijiDHpOYsAvNPaxTxn2ZJzRMhT5UQgGE3/yDHYXNp0DOwP1
ZErpJ5VJw39brNMazMJdIByq9ktrVgR0d05zAsXNK/CH4nPenwsLJH4mgHEB+5008DeQc/r49TRB
25sO8DnFt4aBKKuRAqpLJjODtJaMu6JgmcXrX4b1UmOnRqQ8pDaLlrGP3xMcdCWOgzt7J9997KEs
OEQ/kDNnuOy8XAZmXsJVc3G/7qDExMw7RbepHgDX5S3KDU8YFgSvU9kOay3xw3goz8qOpGbQg0+b
sI/Pwyb/ByVAPzcFpSR3hkfeW9Q5DVNcuib3B1X4WPCCE961gkfg9lo4Z5sfxI+6fZt/4am2rMiN
EJhkDv+4wSh8EJViJNpVyei+pDe9+qReZVT4g1cKxyZ8KizW0M3LGjPp6eoENCT4GoLmQAsQO0JT
nfEFcWV79g+QsSKJsct3cnwvJT2w48cOLP+17WUiO60gRYcf3EWe2Pczn4+38OSJfwtZw3x0hZiq
tM4KyX/En09VxLvpL4ZVK3ff4gTxTXjgOzA0Y96kIrsylfFitNbMtTIysEzwJCE9GjYTrgwMwTns
yU/zwJs2t81HzSppojSicxYJil5bfW9/bN7Z7r6OOj8i1Pkq4eP5nh0ETUXdpEbbjNZJu2hN79WR
rW9ha6jTXUVKlojoOckQKHA9laiVbXDe3CQozn+B4njnqE34OrZnd7oOVyYxsVZdk87HvKOBprrI
k28opAwwQghffd5x1Sr4JVg8q28A/7sxDTajHAg7HVQ9bq6hZAzFlQ0I6stXH4ejzo65owsig3yX
281nxW4hm+OHeqult8ikcujrFeKbQFiJJyDew7X6nYg47Jeaa4yXp3yQ0mwG2gj2aE2DH5VY1W3A
OSxYn73b1LHVG0IH8j5xahMj3Bsh1Dt2EyZNzEjMCUpx8np/nFDBVW1n4eiMZBdrtSeV+pRTXN8w
C5QfcSGF3yn/ymKrSHhUsHLBByHct0hEpfA8JT+m6eG3C5VWvHQCY4HeUhLQDL7kwy2LU/ZBhhJC
qM5N2Un2pRUJseQmjt8uw+Fvk1nCe3cNerxw44l9bWPwuWrJ23wWnJUfHGdZdPSrVIVbJhq9G54e
BZM+zJ6rSe+Zpd8xyo++EtXSOQhkphCajaO1KIAkkWr4DewqXSYcCpYxZ6CgOh4rCWDqvrWSa0/9
AkwIrQMqyOBvZDRQCBGk5W2nIf46dAosK11YvZ2Cc5BdFwzxwycbG+DLEm8+r4s0ly08eRouKAyO
fwRjKz+e0Das40Nsa7KQH8EEl3XYfdCJCPL/cDiNSM0dk4sYudH0t84U3inSGrY19lHr7HZM6QuL
NHRrY0WVZw/zTeqyFYNHv6alF1eteo2ZAOVQ94VN2f/6Ue3sUnXqJ/HMh3egF7Mj5LPzWZxi/TWH
2Af+Rx3AruMKio8x8YVaJBvImGfxUZyvoEM5FqTGzZPHvPVuu24N5xK2ztnYQzNJjsDscMG+Olfc
VSIqGEq1FPuybBNkjyl3jKIGJ1WtlLcsM6l+Xwy//4J0Uam8HAFs4GpMPDHfeg6mgURhBfEHRKb4
g0arbu+/PaYza+C7cqfVIw5SkZZ0Fk3irNzjg6XKZmLdkV029IzruaewX1YPL/U6l+ITzx5cxtvd
IW/CS1dH86tEK/8I2SlJhv7laTsRIp4jg2nGsvuyRLRoxdbLtslFF8/hqy3Rous9/5kxlwHhWwZK
2Sm8lcI3ZDiQV/nz9hnRoh1Hg7gZ6aniZS9tWEk4b7pCfQX8jp6QCcqFRHp4XlqoTFDzGTxftSjx
Io4V4Zh7sHjCCRbJWq282FoUsyFzsSH6h1Z1yl6ZCMGO3YK5rdpBsou/ihdXAPDHYZ+gKHYPmcMM
gbSQ51WlOSxJIByUbeDpSVrvoKGYwKvTxV5xpFqa9ENVq4kezz3iPxGI+eVan8IacbWUwi92u+WT
Sj/6Yksm9HU2K5vFsmS7Hgic4Aec42WEyD8pmZJReS4hIO0a/quN4qMNr97rhDTkjJcH64Sg0jgD
SygHRoEnJy7lZDgbqGt2vxlApqeVCLukbqnkjeC8VA3Is5i4SnW/2nNNKfv3svkfUy7B3WxD5U20
u7zRxPUiM2tIkKUgZ42qRwEMhfI57cfLyG8R8qdMmJD337OgrfFIK7/aB+ZjTQviu9vAwbv83O6x
Y2GDMWdO4cDbmAoTpyhrHdRCV9ZUAOk48Y3bYWZfoLGC42Oc3OaqNN56zWrf5B5CUq1jrXkHMuyj
GuS3ldcGNAlQ4aXVXubQroOacHxrU1L2X4yWFrv2p2p2ZkC4mZVTo3fLeAVm0btE9EbpO3dgNi+h
fnjJsrwTCJMqkH/jhZbfwOMQaTyiLMy+bmfL8blBIVpY7dHTBYwXYPdqIain0hlyN9OqXi9Fw/y7
5Phn705ImdOrPoK3db/8l/jq74m8nt1uky5uoQEOLF4bWHU1ziP+fPFiBHfWbpl18mx3okzxWrnY
n9KP127L1lPkvZSsQtqPon9FGJQj7xFzgVupo92Pb+OCPSzuEp1bYJU5rIHrLYnhPeJkkcdsNvbX
RzW5lUNQjdZub/AzbfHYiSra+3+HlP9Mo61FMFpSf4FFOG3VJIY9aLL4QKBqLYdiLYXifObwyaCw
rFgjltaLkogfdytil0b7WZYn30aMxVF2Jn/04fbaZAfPXl13ASsE/OsUpBGrz9MVN7n5mct0+0s+
hLqKUTadzJ41A8MmeSaER8a4R3UZwjqdzCPEpI0Zc1qxhsd2/Xcd99C4JQBga2H6XJXT5hnWyE27
MmzAdsaasPfgqeX3pC3YRqz3vN3Z3QKt4J1RP8aQkHu6nfs0BVpbISXNy2qHxZthBDLJBFi3WrNl
4g+rqS1h77uO4EMcd5tLcSqNYH2zUlYgg9hBYE3717V9voj8jlamc9KJWn4haPYguuQyVtC6jWM5
TkSKi46BiwkaUPHnU//k2aLSRv+x+ncBkICo7YJD32KjsZjkXY9iBR3DCcKApffJ0Glpdzpv36Zz
7YLe3MenmpahGMJSMQCq81Iz1mG+qLruXH8AHzDzo6gjvjClaO26CLSgsrOS0ww/mrCHYzsZWyTr
6lhlGRHJvBU7M0X1DuDGfa/CsPWvA8DxgieTw7epvuvFjH8YNagazUJsIlvpIwAiJ03id8deQUKI
U29TDgaHpCtby9jlq9PlJgxB4fYi2GChUpMWfrRC8iIzSRswPLUgk0beckRYtze4T04lB/yU9I3M
iUKsJtScwxXM9SqiMDC6gPpdIcyEqBoAIeHCc8b7cqIiSCbEsP0p8FJTOF9W+F5OukY91OOz1eEh
mjlGzr3A9nLrWvZbFE1wMzSgUIKZ4Ruf9VmxYVLP/T7UTNT1IRwfnDTI8drFiT4Q/yDNF/o3Z1xy
HLGpzyYKf0PyU3FrGKtJp/w60Atd6yjBfZMJN73Bv3olwEpyDVTNvZShgz5fQ52ow5bSaksicw2I
tl6k1LAAEw+eyGSsPQ4q+BhYaBTqgcnrQArAuC5oNIxTmufK9GTDxRjecS0fx51SHfKrCgIiz+ZX
ckW+54Ju98ObKW+U7E240S5fNuUhsUHAUo6nY3Ogfb87iBqgkfvr9gmRfco+cq1NmEFNuwBbAsdk
c5Ipkv5/Q7YDJX0Yw3HSdNwxQidSOxLJzm5oOVVy5p6TqZ6WD84n9kfr8wT8kfA7Y413yi+UcDIc
vxRTqwaTip2sccGCx2A43fic6sENB4nyYvValtNuBE+x00lxkD1nRwYHyV93WewOEirBR0beNJyu
hhysqhto4x8M0IGwYtltQF7P1REmjPFxol8ZioomQm9Ds8/MxnUueF2ppc195ofjd5T77/GICZ4O
27nmDiifx/BaSvUFmQTrK0buPlb2NXgdxq3DzRWubgd567VugGKHcsQ8ZkUFdE9gClXugZcCYVpT
7Xvm8ojXsDcI+EQXPcyK+iGLU5hEoCIC4zHFeQe7gLz1Ur0DhNaP1Js8iBjlek/IFkVjhRdWQNb9
gi5VHgNMO6aXIfLg3sk56iSfW5pZ3uzCOhsUc2IJ4BOQ8MjUOVr2ljOHrpnOObpV5BwRz6pah6ws
EFmjCVk51XeWgQemM8ATD0pbjSLJ5zsfABZncQJ5GWuDEqCfwS3dnacty7Wf5T48JH4AvnQ8DVEX
1TnTjHRRSxzSOb4nEk59Wu78EGmFeLkIvMzrvf2uZL7d/K7DHl4EEyy3dObaG6O+BRZUwpT4yxTp
xiD/sbPP4i8t35pW6WL1q9Cpro+EeD3oKwwZN0oKSOMyIU5hII5YykLh31pVlz8MqBuwXRNvKTaO
WQq93wS8rWtWQVnrQejkgcwm1pBrxfg+oiJApNaxbhYELz6DiKE+/2t6LA1DlCDPTNqo3vMXJhuZ
fi/QoL6IaiLm80Z1grrv+O56z290cIgq0LxS9MVmpEOfrXR8CJHRd3tHoOWtw+PtlJnnO8y4BcFl
jXg+VPdV/tPCNGGR18OOcPgHSbb+NANzI0/0KK5ISfYbW8keSaxieO1+yBfpH0ZzJnig7gU5Ogo3
b0fCClI7P2YcR/hu8kIu7wCuiviQguG3c5qMDhO1fiEsOgxY3be0Dbg3Y9cA5DR/uKKAhvgIjpAD
vFX/ygHci5SqSTkX+/8rvT9iCKhzGAY/JUBYv/yBigkTctOfAwfAcO39DsLojVrcyBHeMe9Uos+/
KUlZWtQW/4ygz56+XWaiYv3h+LNK8dXFlpFtoa3WHdUQAGzV3TdRR1wvPM5lFEersNyHe4JaXpto
kA9ykrxXWBf6S7t0LETJLODSN4zNo6zSJmw5vbg31SxE11iz8EKQISKlkU99smBCYyM8hqU9mH/V
ZmRjIWdC8BVl7K+gZnirMs/x/SdNkyXl4yfXpwuHY3kRWJV1YfTVLe1Ug+qFMD9VdfyOPQnAitgU
tYZ3Who5Nb5MJpIhhnEC+JwAjuWKhPGwK/uwjRUSJQ0ZaKSiBU9G+mwJcpnrhQnNvSL+22849zh8
piMShhgb9RdaENJ0mX8aet1SeIKcKapBcMAVHEH2myQnrDuRE4JVbEukQ1nNqIIvup0HtZQe2TyK
9dr4M4p7nswv08nc7saMwkU8yxkzDaCnkm921Mo84zXDu8NHlGqaF39MZiH5FmJrj5YtV/EyEVWd
j28l95IWVDlHPrA1xd871uTZPU5jlqtWZeM+NoaufIRv4Qkzq0o1dFVMdu6X7dYs0hzZBl+MKm9C
uLaB/hsz/Ro7F3B6+JJTyRPoEUNIFjU7XBs8ZAeObMCgOtPzQU9enapy+NKjnBtg50iiuRO75V61
h8/5qKetAv9nVU/iZMTE+i8lfRsSIT40OCc34D+NUpUH+tXyOxVbbhElQ6tQuQ6oWFVf+jaADe3E
0c1hSSMdZDNp8nNCC4p/lMmaKrt2W4gexXEannyMkhEZxZ3sohfqHApD7hsGd/FdO5emWdo3EWvx
NdXB7+/yD3RRXyrdSs04SK84Gyq6xBuBGizMzWV0CcpcTtb5zEWi0tstky1G0va+2axPKoyztyCn
5FwhNaYCxM7/qBK2AGDUpB68KaVoOlreF7xcv3m70k8Oi5jLPte/RYXHL0o+Bin+rqbrmxS3SpLN
42W1wItkP7eUCb/g5HHciNTvPiYBoDeIEOnDAEDP9PPc5VF2eKu/yhVzaKVnticB1O1GoeMuJkMb
yg+h3vuTSBshP6ku+e4Wf+SbPpDMkC8/DKYSN9kl1Ru86Cc1RIuLQRYnoMtw3E5URaa2JJD0Uj4F
Y1EY+QaTqHSi+MmhtbXwnGrn5gF5cfBlj0n8cLKvHCeDthWK7XAxzECCzwc4J4O0AxuuLiW5kxJt
1ChUnNBcxrXQi7ZtEIarfvgcF18ZMNfZcAdK01C4dF/mxfR11DV5CH6ZlPWq8+F7z0tyiGxcxYfP
jt9B22ZudvKf1u7xQr1u4eAU25SI2TKXgm16/vpMaU9Uy/CFRV/EKYbjRww1XZG2s9s3EveyGv7e
jk9Wbf5RF6nJt/qsaZ1ww1CU0jw/iESBZt22TYXcZSglXRUmD8J+oT5eQ/4cvSQNvFIqXcnq1sJ4
N6LyCNx4BFl/rfOFe9zvKluKZ5XCaOFXzZ8ZHZP9PWbSsGOPtXrU4GVAPotbEJTHrsoA5hqPS87e
D/5vZIr+2hwuMbJQa6+wDCuVDN9Jt9aIYK1uR+EcGdyE/BHQljEXq/0vKghRkWGCuFrdNak+rALR
WkwGzxuq+f2WvTIW5GK9XAvzHJBQUkKBGZaljkI+vE6DkXqWOK3e5x0sxlUrXfrKxATN1K+3jaRW
DmdlDKuhYta1QPiZphfZOdb+DfJZf9ah1p7TSjeS2aR49YVoCQJHobKB2RilqildHVsOKYDd0FA6
xLi/gKpcBb3uEkkjPT+NXHV0D5zO1QtL0U++rT+r5/YaeMkKcX2x2g98A6JpG4H7/EtQOeQGysX7
NtLdXmTqvd7m2eeQs6Rbq92Z3m3QrLBOgmJqDmJOUNZTa+8rbir+jfc+xo0qpPB+XHHA9YZTaW+2
5Tzc68DPSlSL5a5QDgCNHZy8vronXMLlLyYes2Umm5RSh/noJeLA9YTQLgPtvHgemUtUTWofhh97
7IEVjCR8+B4/KVGn4yfy+LhqnGebUUtHVULNlLQ5SZcot/sldQ0zNO4sdIA9mQnew05quTuhFueK
xr5pmcTou9B2umCTx8m1D4p649fjoupnGhcDgbn8xmOZSecWMHr0MVIf8t2jiMFv0ut4EAhy1QTJ
W8uxsUvQO1EwaCJKJlrgdHiMwLaEi1HrPHHu76WZcOVoN+kixaRaM3siUcPqGnCMCmTo2v32sZKh
qnnmpeEAbF1ryoHmseU1mhEUNkh2AL3JAZ1+ZN6495ngO7f/whTwrwLjV43KwnVG0qLt1C51dUnO
FZwCqBFxPSmwplfvXYIKtMxSy0Er3RtOQSZWPzyl3uSCykir4miwQtRpc/YkNDd9GtbG6FaHNPp5
D/9zrLCT2z7JnmULHQE/L3oGymKHokjY8jXCYOT0NB4//jF4St8hlsFYXB9n08nIXc0F6fu+Hs1F
TuyQV6Nghpthf3Kt9MDxkpkZV16XTDevodVE2ctoyOGHW8Je/pA5Klnh30WWqWwHgaUVycj+OW3K
AH0aYAXZEatbwnOYkxhNtp/FLhrPT/CLWzYfXTeX0Rby4psLgKcU7jSihvtBkftgL2mOAl7rFiYr
9sUiuRL0LE2H1v1JMb9hXOyvBkItwTaDOtf70t5Gx0O8eOpr86Zm5d9lKBlHoXVVPhOQ5VBWi5Yz
fR4KrF/OBQSpvfXPngVi8Zv0qZEDD6gcS40DVBTxHBBF12UWhEqXk8qqZWhp6eSXkkmGNyRnm1CH
e4UMnGvGR5IM/Pexnqr+yD/aJERJCmLzX4CZU4sBOlXWq+N5/MNQJ+d+If32UIEgCKuzSx0GCqZ6
29FmqVx2Flvgss3qqRdTjIHL+zbDhGNu8wCoQb6zhFtbFqewBg+pT2cAb5WADFaUcZN4jkKqcp2R
Q1iPj6O8AVp5hhPDNQa/ZWGnTm44GUOYcqmKt352iK+tTSBbm0h3IMnDA5Oq4e0SXI72JTP9doxn
b83IZQXtrBhztxUFwUni/DztUv1rGNB1kaB8rgN/ZnORHkU+3UmC9ovSx7+z0GcL2Mkixax6hq7n
XzhAc8jJJAvQVffhHdymIJr+oFOvMcBXGH4PNVMkQ8NK3IaWDrhCgtaGa/Qah95ZEr7Po/5Mcrc5
e+BMs7w0Bp3HsYeZXyGOBSd1elGfruW64w8YkfJuwMUp1GcnNntrHDRq/qLtlJdPCarPqp2EdgI+
/F9qH1PZqM54vzpx+r5npUSGh4LTPySLU0Z7QOZlUYqfUHwLDy5NPD6JhLX5+17paplhkG4+jzaX
Uou1brmcVQ6ij3xAuwYk59ZaqRgPvSgyJdJQ72b0i6Bkrb9+n5lCiCNRUoC4o43mN/5KYpWcL0t1
QdLPg81uYCsKHMhopZbiV5JVRiOf4SoVYLj4L3bhC4WzhUxRXwXNFwPYk4fkCkrJwjnCSkRxqkX2
mbyfpxvrdoUHvqAnTvz5o6SmnKRSUX+ynoW/DPbiZ1X671XhPh1+eDUbXsL3GF12gOI/ZhJbKZFN
X8ssbVrcNpD7WdTdUKIOAFy/IykxwJP6FJtpok0csui3m1sWxdlzSi5Nj0WP7dTHtlddCDX5jXIv
3zWHguBScLlifvB4okUYKhO5QTGyO3jfbegobIw4nTK64OnwKeU+NjqsAZ3GCGBjbNT/75vLADSC
y6owMvFp4bvJTI9WPKXzN0mzkufbGcsPVLNBOf7FeJ4JbFbgr5APAZdObYIDptA6v6DnDzDyRJQp
d34mI6sdwJ27KtCd75bl91r/vmEtQJ3Jw62dIZIp3PwuheJ9riQzKJF+LWyqGjA/Chsxs+fssV2k
O6d6umUPx6ZVRVYh65JH10V/sTbq3ZxCgeO8wIRLJFi87xa92dpzId1aPonQJTDwkRvYMT8pdrI6
X78KxrbS0zUnG/ScaVu0Y35GAOSOyr1Pd6e86vCsmkuCYWF1nmJery+qy0/rr8g477PIKfe5oRLG
oGEoYDSJlbXjl7abgrKxQu8vKZaHeaoKQuUeGN9Jq5VTZwcEPJTmae3zUzJIiiWYVwehymDcEvfz
gtupExupdiP8+vHmKx+vZhXViK75YWG4VI2X97OPotWjhoTB04KFTfM4FIFebeAARhArYHP6kDA8
3Ffyh+WbzXcdndw4gFavBF0glTA0ESoIiUljKO2BPrwVnU8SrTixDti8VUQsfhu/Z0SbVezzChBX
q9WBRkAzqsGIUTIkU+lCdudW1FaJ+BcrZjVcWFWi87HfhmbN4R9D2GeJ5vbxy3n4r6cxraOqawtW
aCKjReWTN0hfElUhTFUmB8FBMsHGj0b4V4ThYKxudyQinQu/DiOwc9BrObMPfL9OjBzMlCW/hw9s
VgRLNfotjp/SNCnqkzBvQO94wWMCoQ8NQPe9X37OMeN6D5etka7aCHO/wdA8e2m7omhccNQnXiqD
4H2DDDiIwyT31QPaHbn2fnJZ/sI1zkd+MnnI8q4RioR9NdvWaeTlISYWkBSIDgY8fwiM/53js1y7
HGmL2FJRttfkFFY9924pBRZwycBp56emcxIK9PMD5WAVsDxi/GEdfd8PQ4Uzrop5vsWaG9lRGViT
rIbubSd1Vv/bnZTutdG06Rc2pNo+GoDjviy09dl9ggGPVgIKV4WP1eA/cSvApvQtzAymNIzOWSs+
Kh7IP6T6oVSWQqPGrDuND8iwHWjc9QjWnmcBiDDXmsyWJLZST7neUX6loz9RGSBa+3AMKb64Cbin
w5kDD53a9za86mSb5S8ltII4bva2iMARlPAbzQVZuM0TpbjYeApNY2s2ueQxFRO7w8v+JbuCjSq0
WPVIaOsZn5Z+DbCc13r2/IbB0NQqeznaF9LWOMPvg6vfdotcW6nWyZFdnNNfeMHD6Z0i41jIBG25
diMPsaBdVdnbtA7s50n9yNeSdc8dPG0wTfY4joE+0tr6VkZbW0UowQGaMaw0L/1MVmB2OYfcrR5C
vSXD8FWu9fD4vku5taV3JNmq8IJMSGSWNr3wJwsAgW5o9Vyi/mQqnhJiud3wNb3YnFy+p9pFCcb6
V/pnzuP6vuDyeDWbRXErAO/HR7YYZTMxao7xnrrQa+JxGOeQ5CSoejbqtc3ApsCIl/f2qSlyPcFG
TU3vsLiLdhooEiNDVOZoT+1cG9ygtT7xw0e1J9cnKrGU6nFCSgWeKk/sP6M5n0ecSQxhbWgEeCEN
gJ2B8JmPsxJe00BmCWW+0D9J4ZtG1o4VF61ZdyIY7LrqX5j/6MlUFps0FTFUpBU/JYQz8emS/cVC
joesLhgspNY9dTXEsdoq1+y2dNjgCXe/jDrF7XHgoVSyZIe0i54ZxnU/Si9uvQu8hv+aydcg6z71
1Kymxr2bxiT54oiowre68c/pjVblrtmM1HubWeRelx4gp0Q5WG3Ds5CRMvyH2PW6jTSYeSyqQQBi
JL8SGXSnsQCTUMePFj7kRNLVFBL5CBVh0wSSf8MELIUxdsz56KiDT6jBu79QA+mZzQPKxMnF0e6P
x641qjK10HkyTTPK5d4wbRH6J14e0iYd8oRlH9o6tLZLusG2nwn3NOTrk02latXCaAxpMDW1MqS9
sGxYn0Py9jsjzrOrDA7cz7HUdzHwpq38jLGb2PHpPe/gYes7YY3ALRRnc0IQsXMp4tYzahTep8Yd
mhTLBgRoHNNqJARzEbahoeu1gt0fZqV9l5dRmiSM7+yk8d+pP2GQZjzlAeKLUHs4+bXr0fTD5MJC
syoD2JOzu9VeWOrSe97znEosEPaZ6L3DJBug86mpRJgI0T17Ld9FdPslkotKr8Uy9RS75DGugUaj
SDZbRfj9bFz+E4u3HMMDrtmXD2zk7ScXO8tqCo4+MawTUW+RTNxpy9zw7Bd3tbBinl8nRPnJNHpH
x8RS0Y2/N/qiIXEi/R1gd6BOoG9ORf5WJrplqFxkkX/qFMlddo6zZESCg82VQX+ZuBVFtzDi/omu
+/I6zHjJgnxcDfo1728SjDtsvmSgZdHQ6jaiSjC8hjZxf9RfHKz1UUBhLWWPADwwwkOFeQrhrf3f
rQqttY86b4XMAWtIrw1Ft0InNNQbif+gz+jQ7UMJ/dUQ2+GyAk32v5PXbSTH34ISairjKN5yycKQ
ezIeX8y3iFX01si5a/1gl+HT5/dwGe1IFGUJRbk3/4pobxzzFevWIw7+OO1HTF3Pw9F0WW/fTvvg
28iUGdKhWbPk0zlMlxgFPXQkQwSN1+KjRFBYXC3uizlf0COfPa6QhiOYJNWLU5Al+Z0bnzgl377h
jlhamzVC7WzGsYvtOz1OVu8TQjq9i1RKcm5Sw76pJ4WyiWj1Z0bjF1ldpp4rZXEz+nVnLyMfjy4j
n5AX1gt6CGFa5J+bHpdgz9dDtSTr8J+MQc4qoR2J6EnvG6+PBRpXJbVyn5zWoiwrkd7WTRPVmW+A
LYqO2bR5+jzOaWBgRRN1kaljsq6kN3K1RkXTjuzI3rKxZ0TfRqqzUdfg/1vIN+UJr76OVSblWYRS
Xuiq5yewVyTFIKoy6J70Iq4ctML1Lc5YPjofpb75CttzsY/jpkOojdfB6lGZ3Oa2JZEK9igvqEJe
58J07vDexgg9X2Sjs22J8uMt6AdGywOfk3ruoPp7mKEG1roRAweMN0mkFVvHiC0sREDmAY7s8pEg
n8IohCHF556CyXE7hqSrY//ruQkLLQkCpB6ZkPEw1242V3Z7MX05dUMeRXWqPl4FppVwotD9aZ8P
lwvwwH4WQRdkNwZ0PO2hNBuI4zf4wIxQ4y7Q9osPjcFUOewz+Sw7QA/F60wDD79VeK3Jv6RJHns/
UyZA7/MuAUV72Sy4b89HNGbRzaHatVuwP9wrMyRJ3WZxwXbywGBZIrVGtTVf+4/t0+90NG8yzJ/1
OOXZQUVX+88SFz0LoJkxRP+FieXLr28jHxQBBUFPhbJ5xU70IcsZ5dDXzs3yVZ1ylVe4q2tBUtz/
cB5Yugq66K8L9R8T29S79xY7r2LgD7rT5QsZ4dAEdEeKsKkfRedNbKwzIPZnzJ+g05/5boxxlmlO
vVNLFw/NB0tbzstnHks5MP72K+FWmWY5S+U2pA5tiH7QGdXLfDsbVvTd7hL/iFLMBrXFseQTmTT7
088Rx42zXyzp76Nhxhx5cVdcXzBlkwEXmJXcaQTS3ECitIBGQ+SXSSDI/o1kSSZqebq8X3rC05LQ
WF7WMueVIu82/F+AvC76DuR59KoRYFoJkleyXrBNxJYGNo9wls4peNgHNkpB66t8ZZvWl++s9t+2
IAuqCVqhFIxE6VrAynKBeN5KEhWe3t9EccEMVvsuUzQ2b+AhCx6HOoQP8K0c9qCH2my2T5uswIF3
qG5cAH6uWdr7IvB++Lgi+FpjRbAMNQsjgOmg6V/4VJmyu5He1bPvgQW9kQPCdXOQR5YWJj0ZblyV
4iIsZbMMjqTRAzaHyIIeDQGgzElSmWohboZ+LIgN/aHQlidbKRtjEa2bPfQ2PSixRnCcdLsifVae
XIdKnD92SQ8l04jQakCz+i0X9IivqeOFEJtEqNlfw+jvVbARESDkamgWYVYcV+gul988P5twoWyV
Yw3VqMS+pIh2CfWHQfQmS2pLuonk1cjtB/bG6ASdnZgUa/1BwcWxZRIoyKDJRufC7wtKCUjAUqsH
UZuX8fIPOOY67u1X2Q/I9EQksHK6vt7szDZPlu9a+ttbhJSulUmyICsWvpWkm8zCzcJbR1TtCDGz
iE7vJJpyZwr/r16d2RmapyGuRR35WGFQQI6nWRouGvDf/PhezuDWnsu5rVGHfVNC9oduFP/lVYIl
n//A/7UQ7t6qatNjKy/bH3yZ1CURVTppp4I3VjiEJADEysIlBSIOfGhT3O/kaa1Kr6r5IWZ5Hal+
iCnnPQkfOVLnC6hujDLsFAhHjRT8II+Z8Ope1SQzNpNvXFXaY/bUbCOvp/qJPQztma4pnu/O2bMk
tJrMBiBSQqJiRI142qgkf7c5LJNIph7or3fieCax6NnNjYtgr/cuoa89dDW6BtDH3b+EpzM5EtN2
zaCukWITp8c+tN3E6DE2PtVzba1EED/C+QU3giKYKSigowmx2ArUtFnrMiEyFG7eWqIoXJPNqH66
3IqoflvDVLdifuqoiSP0vARJ9e0C+DHBDii2TGAuWoajSbQto8hqdzuRETzA/GIoY49qWoQicx3x
SUHAFfm8b5V4KOXpJ9XuUvoa4ooB+Y3juf0WreJ8c8MQSIlT5qPqWLSI/DIwY/IxYX1ONSMdQfxd
FNScGOHmoMP4SHtIRTp1jfvf+gi+3aFQc+ADSdMkx1M4rFPWmyh6L2r2mSURHar1Pb5r9sPn8YhU
+kWmuhysbeyvaiWxcUzzuP0fENBCe1VIb2dkVNPoxjDijPCyKN4xBjiIBXpbzVMMQ4rvZmwkOzvq
jIMK12NBEVfYW7l9f3XVwiP7RoWmX6c4L1YBswOwNjfnaaxgCHbLXewWy5UZVjpvVQcSfFUg3nDZ
YgNvHJpIwwjKDK8gBWOjhzA26PJXlGZHh2G4fzOkRwMe4WBZbKtjxQZ01WrAH2pwS5nOpcEFwQ8A
bb2heo4NkQkU1U0HserrVO/2kIecJItstqVk38YuFoqXRRT8q8Ox3RXog1qPKQWbDraaaDeSs+UV
5gJ5Sjlx9kIYj7mEx0WH448QbO/7kQyBxBDLq5QPer6HqxTjwmtVa4bBE8rqqk4Y2VQveVBXxD3d
mis1GwbsWMeITHZa/VDHHN56tsHLtw6rnsrVyYGEz2pBkrbG8wkpp66q4sM9y3P6cZZImG1mTkdH
XWJjaM65kU1pCmVaOL7nrB65Iv8TZjag2jpo8O3RDGIt/tf+nk4n7a+K92mkPgQJ6BmHh+k1hKXg
ptOvEi0LOUWoHQX6dy4zEPWLVu/1baIbv9dspeTZZwXzfUNdLQKkNpi8I04ETXxU/xA/ORPaJIZz
YhZ/Jy+H2qlGkk0x4HpAJYGB1tEsAPuvnW2IcNpZnlpd4oWXzpFj1lzKJO+59y9CgUZCEaIlbcnH
t7Lo6SVT+FKdz2Pjsc0oFgklW65CpJUfiTFJcy3zY51gI1zpIXoayvc7y3I0cbnfhhJpbcyzYQ88
6ti+V/ps2VtONOQzSsMMYxm2fFj1CR8iST1An+03eIiCpcsjLrGc6hFEPtfAtQBMRBjsOaDdJ+i1
zKRsC89035UFPrV4fbkg1oIvUHkcs6DOCYTLqgaEyIT2tWpn1+iEJEmo0SMngzdns4EBEv5/mHdi
ZvkQlCacM/y9aMKRGfs9uoa1UXRKH8tq5oOUGLn7ID3IVgcXFBEtzrTDTB519Uljyiq3NE6z0wvU
yri7lG/crltBKTXfPVCu/YNM/0t8RAoV9ZGlO2cbR61rEIHVlcqRvnaAQS8s40pS7ibL60JZ+rgO
SxLcsOpWviaaqis82OTp0B7/IThVHr67/gZO3xDT7EYxySqQRgqDKetWGb1md0dArG0kBmwjOQkN
4oern4iJcC4hRvlZoMbkl6S/o8LbWIkI4xtByBB+C4CBzBK3JbrHFyeaOfvKSr6J+ZDF3McYeeVy
0g+hQBxbkWw93OovW1QpaoVTkqjaqKZ/ZMd3C56SlpNuaWE+d7t3/sKEDACuiZuYdJV5DtOLU+Kp
363Pk/zDe9p9P1//1ArZpk/Yh8QzB9xVLcGBDBazz37cXocCH7xEEP9588WfVDUU0O7Mb+PQmLdn
ld/qEmVOFJPUsZAiMHvwT8FzLNK5XzHgEC1L18rstcvzHugPAQJyUQaKOWwDr9wz9kf63kAWrhGt
SJN2nJyGEJSs64jyX/10ksVQ55Q5eEL1ysvQ/ZqEWvxIgFhK7EfJXCe68BK8kefgEgACf7okLxY2
7OVoFcDvJFeSviIVYOM0pxNwb4aps8zGNBQZ8MOk8OWDjn9CdDAsZ0VlFIlv0o9I/jnkYXkxnhW6
qfOtDH1Q2UYRND3ffJfTxfCAaKxAqh3/FUUR9hHhQYlpuQ2TwchKNrv4+8jjQ3maCLjYq05SLO+O
TTvujOtvlQMTWg+rx7vI/+pwZYO7Udm6gjIu9Zmnc7rsS2ihn/ABqE+hf7hwZb4QDTTXIANPhqB0
KQQn4hiE+VI34xxR/1UmOKYo+gA4Kc9jxUIoKhNC0R8Oz7iE56jvD/Yw8XrdNM2hsk3+mz+VfFgP
7BQ+dnRTB90tW3y+uuueQWxcV/HQe0FYSak3Do2oc2NAuRd28KOzIYf8GZz7KF5z2Tu/jD8NKA6K
TWWcBFQPKjOySSOAsQsZvIuEJA9i5z97sJ8TM/nWhNXTCzCEDndERVv45PvLfbBrz+kjMtnOwnIB
GMlUz85W+jNCQh68Nz+qgZTyQrmE4pDRoQBQ8zjCH9lGvqZxSr9vbib2gAMaxS8393MMLIh4HEJS
P5JC0Sl47qiP4WM7AOYvLlf/SkkH35CpEFNffmX5MpDLI6fnMCy+q6tx+vVaYzg5yZnXwh3uZ+bA
r7LB0l4W7nAbzNfP8Hs6mtWHilvdw529BFNIfCCXx+o4KAA68M01AWyyR9wXqOoD/wH0lmX39la5
sazbYZj04rYSrlgBH6FncTmL7LZF63ISukh94ikS28SaL/4lTi46PYexq2eO9CJqdMDXjID9nuwM
TDntEElRNPKNUuL2wD6RsaWnHpjhmywfqc9Qr461WxnePtPNXxDnoWK/xS0/KZwHEpxtRALyPF8/
g6VVvN1fAGsPhvONXd4Bv8xNVUCX400xUI63A2eOYHulmPmsUtBbBt6RZLgbsx6wo09/XGwZVF8E
SSoxF24n6DOcaVwc4JwtenxUnVgpDUxjDsbgZhx3H9JqAv1jl99eqLfcf1CCRe40uWfCn0hzbzOP
+zFug2E+QpIOquYD75aeoUEXTqa7iwXpIqBWxHHbEZl3ax2dI4VITBeI/bGB5letG/toSwudiOdB
/zNlNZx9Z8fx1UBAgPLwDIsKs6O7OI5G/Qphm98qXaMyFoMaf7ptmJKnC7mDdCTX3d4dVu+4n1Pr
YqDv+gPTbS++wzk3xwS8tzrTh9frqFcxde5mh8ARgD5ohFRALVM/YiKKcXFzhYhiLl2P5V2v5nRj
f8UlwjK4QSTtIulBb1FsUk0bHqjt9HjjdnjlcqC+jutPreUXuCQy+rzbYcx5Chc/h9COk+dpiZBK
ZyZ0JkRae4YKkCFdUvi6TT+yEpmFRFuLcECM/FVC3Oxm9apTwb/E5BT+Cd/Q1/htIp07/kbZNldw
X5n4hMi7h7fgDss3a4wsGivEHYiNVx4MTlVbCuw05iUJFWLFlM0cI+7qN6TCGMTcJtxMSMbOw1VI
gNQKMz3MCLoN3Ftzlw9qyF9waXiYdvlOvNv6fletZewBWuyn7fCG4RPa9Czit+tmdBa0w1UViP3c
vShthyJXcLfvdM68mL48tpO7R1Ni7P8yNKBEHHFmUIcXBXPgrFNToLTDL/q7EFWB7qr/vH/jP5A3
gCMGbwq15rj8vU/4/vpXm8IMK3PxgkHEGNESEI3EEW6nA/ldliXScenFQ1d0lfRDsEBbBZNSM7uV
21HpPdFBpkujnqeYv2HTJviP+1E6GUJVZxkzQN+FgKw9J7YAhJp86EHHZNDWwYV4KMgYVbBRUTtH
vzuLDiGIeiTiUnoaCuY5bj+kEzy9QNIZYcTLSOB6W08ftSKI2/lD4eoMeH2sHm0l/D9fyvvoZPjB
b+n+ZctDXQGlirTp62TlsMIyRj0CHo5UQyiNwjv+y3zaJQVRwqzEVmKuWuOglF4GmXjMEVkbPB8E
2IpNHk3fknhAam8NC9SwndcrkpUMqwvTsGIco9uy9jAGq0HBhISb511PJC+5uounYTSutIXg8nZB
C7/bW7cBTrEc2AbQvICBAV+OZvKoEwhNncSbvF9QHwA6j9u926Cb3kLkZ5bl6icjUPCq0NIg0eTG
3xbnlkdUzUHovdaeWydgoQzJR+nk+jW7wY6c4iimsFweHvJ/YFDSN8Hdz4BPlaASqeyLjHwztDe5
jRLRYuGcDgl+9M1SuahstmPlTrnjwRc8jVphbbBISraa39i1Jf19m947L/FFAP8TOk/FExfK8vXP
57CT3Z22YJOuq7jBOIIlvD4nNz/1Z2zLz7ZFcz6PJp4WUCCKtJaFmO18O9ZtQD5k3tmlzTPOUh8F
stbTDDbY9RV/FYzP+UlD0dCERQZ/TC/MCa0/5Hs4calQcV2IuB+jeGUJIx9hnFpbGaHcT7EQVHqg
sAdVjUYdc/OkJuDyjmISDGSyX3hLnkzMOTUFECLJI5t2bq/ae6NeUGZnPPTyWlhwlq6DjnfQkXEW
LYx3HnDSbjVcnWAHfjaO+JFRuHtu8VWsvXfE/UEcHI8vpYa/Z4+7Khl9hHzkOAbX1yPF1BNopgGk
Q/PuT0ZshIwf+d4GF7I88JgR/UJ2UISK2qgx+FXVXmC5WZYsFGio4/Ih0d3TNKEJ7sV6FqM9L5qS
1cHncpnpiUT9tZY8f8FXmJE6VUyVc1LpwX6AYyCnKHcovza96HqKGbqemG9ULn31ual6Uyx1sDWF
e5vJoQO5d2gE4DOlAewCF1BPprXAetXj8imoWbnv6IaDmSbGzTaDv8yWU6vBRTUYmIsr9Tx7TGy8
RUfLID7C4js2PkO7TEjDmHhX0jqcstz4qR5WHkpLIOz0bINJoafbPxnJT09yfvxo6OFpp/Oqymq1
pe0CHhcO0Vm9WJ0IzWFNwoX5h/6AWHmBduyzgzT65RfiggN0FKxbEpY23fOgiuf6dECQhS+qDySO
MtNEb2xjRyxVnL4h9jhSiG1AJMJB8dDIi9tyk+iQtJpSTCuOyklkiyHC+tDFEgkc7/vXY8k2nFPX
65yxeDF15lNUPdC6xY2O7EzHR/1tJS8RVOWWmYqmV9wT5TEHWYtfPj9ipAGcJ0lRvWJI6TpURva+
t5Ki5OK97MiYSa7PmcMHvZoUEtsZWBPVkv7E6Jt1Gs9d1F+egS8mMTGuMkr2qh2wgV9p2ENThvtP
AbxJmoTF8CHPt3C9Sm0YGyEjCy5NguqcldRGq+NiesSyc6c/bcz/Juci6wCytiVHyLlvqgpBFilG
zEUhhn7tqa+OoVjU9F38xB4dZqy1llG6dTAlnObPLRlTUiXg9E5xX3/gcr10kixPSWOL+4/WFFhK
rl6HyA+1vFEivy4nROyb3nNI23DJn8FKpcW7XXi/KjKwM36tMlHxiZnpDV3/8oJgEAJMnFekZAOS
xnfmlQd8rHg68NG/JtakX7Yelj5iirH4lSsgISXZSBEb21gYT6S6w6tkj+hrPi9kRY1JQL+bCJWh
8FsJFEnaslhnXf5X1Z4TsD72s5Ro7LCh/8NZxHymHaaZUBZ3lgMDVsJ7Ctkp/hTKSeFtI6AhsQKO
FMtpfI2XZ/PnImFa9p2kXEEJEIxd+nMhFMvkHAtN1tJkIk6kI0rpMBG4FQgpT7SwBwtATQEbuB/3
CWBhbJ9qSrPgHNmJbu/sGVvGBH7U3GFolwOpaCzVx0kEKgfGfO9bQCkcX35kNLj49AxefcLCpX3A
Pbc9RF8ehxyE62jzK8RX8V8rUsJPxaXXIYB80WhYIHu5QhcWS3zKmkX3q0qoc0LUj4l61lkJiC1z
B0foMX/tzBr43GBq+Vm/dzKBdm9hiVNfqqFmXmP7BaKtsbeT6pPJqdq2MWvjqiozFZfKjJjaqvCQ
wGBFH5Y9/1TnXEwNwY/BnXeRX9V2Si5uVgajv238xluCSmDZ3NY9kf7C5crL3nNc+8B+KFy34koK
rKS4HtAEv7IopBKKwxHaqX4RBdQh7NDcA36IObJDYPOsWm+H1OGPTMTbrN1EHTFrO+43rkd1sWUf
0xyQFFHEaanVCH4wfjmGeGLG2QINbyhx3VuZ68DDEfYO0AR9NYVkH1ADTEHbM8pRgeLYvnOZZnEK
sse/7+TeE1A65CrYP4YxNnKg+iZJbd28tMyR7USP5wmKezH7NaJiFnn3W9kNiXOYjSyARGq+w6S5
edLvKKWuZsUiBq11VD+zJq9o5nlV5dI376bf19UREc+sGp8CVWRz6ULVOtTHA8Xi6OrMs97l7CgG
jRIJ1QlZWnLHIOano/x//u1KU1VqFjHEv98I9smWagwY12JCcZvsI3+TDOvAnx7OzOpbFm9kw1vy
ZczeLnbhMRDMECzPawJPBUGUpLSPGSoCEHaKpz4CagcaDHHarlUl4zyapWqLe8W+ebeBcVaESQM4
as67qmQcGd9g+HLa4KpOhlKhrOgkW3AhyiPZXBRi4Zt4slK3JwRp9NH/KTKA1jcZACIL7otfHl3B
29iKInSgFCC+vMN4tBR+f8L+tbtUr12oWQkYdphxqt6CcFZH2kW9m9EhaGN9H07bD69yPvv+Oz7r
rLmRfReXhT2ajYyUqo0B5TXrXlLt8BhGrPEzq4rtJ+8mXPdxH3xl2lFZtg/eUsG9pwQ9CsEK67LW
KBdga8UooCTAK62P5g1Is3QKq6G/NazZNiycNQu91FJlZFgztFM0S8A8ESni233DG3PLCTUq7XxT
HjdOfUC0P5OfHUQbn7mPKzL9hSe3PSbj7DD8Qx/aAxhDW8W/FD5fs/gXU3CXzUxq39Kt7Pyhd5Ml
/unAI9bgfM6vTNmsGEHqB8cb3/InbZs0YR/k4l1j2tOJWEIv4Za8FbdQSwmXBZV/HTQDPX9KP9ns
u3lUV2RJassyoy6P5NM5qtutbZS+V/+Ie5oGGFz26M4+MWkjEKVRpuMXEoYWyWJPNSjYN1ALR2UC
qJkGpBzPl9++x29zvWUN6cZgwi6cH4gENXwaDc5VzNYpKqMTE76WMdPkUYcR8U1Tj27t/0Cxtxzx
zB1yozh7xQtiROqE13QPbh+Kn2AM9wZv5AkIFYXGtUOn4XtIHKkXd3CFewnY8IWGyopddVT0CSlk
CiL4oaZThislRIYJNhStOIZlYlel5ql00s19/RCFc8PrsgGIuCsZnwuAPRfh682egB7Nt8ZPnz2s
dFrWBMMZwZQ2DZnbkS4BElDTZ+e4sS8W8qMgKnvwGH8Sm14peN4nlqikfyj2hpMuaK37Wxa6E/U4
WC4h+38DmLgcBTc3Ef7SKaD0RwSsi5K54MwgHFSFF1I0TNhnmov7/GLRELNZQ2az83ovDhNb127P
yloX03iAQ9Qhha9p13dSoD+uJMXdGFLaCXx3S0+1gg360ojwyCkq0R8WQJpQcWC5c/4atSKNkzuT
eQIYoZOLW5UxiWPoFPLzuzkpQT01/nXQXwmWbJ+aE2NAj6+tUObqaGi63AF60olJyramabdWMKBL
fK9Y9J5s6gOXhKEX5GZyvpWfzhShpTr61ME8nRCi+I5TFSd6AXaxP+O06CayF2hWP949PHhpF4RY
lCfTxY1BH0BJqGMfCuG+w1jFq2vDkY64nGf2oTrrl+lQn85vCT79kyOKl85Xlmg317sD/Gxx+IDT
+qpBXiir5Y1RrDcXXWxXvWCCXKGJb8JrkpUl0eeYzeKgFxVS9aqKxIA/Gn9Ux0OkUNFmzS49NHrh
VJ6uHZtwC2sNaZq1nUdDsKYar8QS+lVF3VXTnMkxLIHy2869OyI3/d3zhwVpSAfFFfOxZjUAzqcj
8mJCzT+6kBJpKBTcMbu/6D9y1AXYK5rvw3K/hIAs1t7Fe1D9BeHeE9FQgC8yyF7F8KE2ynPeUwtk
JgdPj38ahd82j9oDJ934ceYg5WSZgp+m15LFxNm/N0BF2Ij+iU3ZXa25ZRYBFGErQtwLTB5I7BBW
FtLIiXMfHMvRODDMogu5KOxYF/l0F/yYBJ/FO24FkyjvNHL6mo6yDeO6ov12EXlF8VeKPx02XkaK
BQ3JgT/0XYIM2cYjlIVFSKybyk9X10MgwZ1R1J3agMCWvEO5F8gNWFfGcrEgj4rULiyC5OUDW4mD
8TadHKx90qTKHLO23krpRiDPtVJpL445Jaj6xtENnPRptwuWY+np/hbPoZ/hMu9KfNB1lo9QJDAL
faQRSFsHJiDYxR/wZFWWNCdpMW0SYruwCXL09GqVULqgr6eMq4NAcBRamgM+hSwEykl5D1VLSLma
nvCblVkfRojDNvHLkhgtCdwh7UxSx55tT2s/LVVzFkZhG4FALAGu0p4ulVFB+6IhRo7g3V+8MZ8a
2aDdVrrlw3Iyzy5NhMDwKiItMo65oT5zOzhyvB8gLcX6vx+eqAmn+X1W67D2efL6czBZcRQL+YXv
/WLRb3lFwCFbHMyZLaku/6GtnvWefNnJPb9SfhvKu1P6s1JOtuyYov9iqXzBlaoHnfzbsWFsBL82
RFIRQmlga9gDLhxdifb68sdzYdjWBmXyVDo320mTUXEfkg/CkYzdTaax+g/J23FMD2oBgM6j1RDK
+IcVm2DE/SrSk7xxhvHf188HsaBH48Zv0ONkD0s09N//s/oVLc9TR5eifolbHXtjYw2Nxnm+HWKG
XwHlDU2eDna5E9+RVWJKQP8UBCNqT11ggafMIPUEsDi+ES6/gEo/7FO1DoFYEZbOWHZq/R5m7Pnj
50yNmD7Qg/rEWFmACFW3x/RNoozqhX6yjV2ttTlcwyIsBhwx0EmRo7vzphb3lOM9a20F/nt1lbgX
1RnyoHYD/IFoSPDGvyd7KBRJKMtar4oHecTtNwCNrSf5K2R9HTvJzrJbTC1tMACBtXmzF2rm2HlE
KyftTEPj0f+y2V5JW3m4EepyZkm0KzA+AzSPddBUosa7wnULsz9qIhakpvezAWtNaoZALjhDXL0p
XIO8eMBWlx0cbMlUT+raozA64jVMW7iThgFBl1Puu/lrRfcK/0nSt8JeUlP5z9O0LZ/K4RFP48Cz
VG/pMpMiDB9bkhlH0I32KmT/n0OYjWlwgFBRC0avYcibIX4Evke92bAdEx5o+vQ7NcZCz0cMa+aw
HZVBHFc4II4kcEg3nPyP63Nijz2GGTAgx91fhAwQJkksokmJthEdsRvCP0X3g4mhq5S5qrsV6Ox8
26Ik7O0Xi5Et/LDNRp7XPSEpPeayy6FTLmeJWOpETfWag+PQHRMUt4APTglUMkv5yLyvkN9tQKs7
K9VGSTbaX0rXpBcVqUii9COss9gc6sCMkoiUT6WpDUz0QhgjTQlpZi87+vEK/aDmw8mCGKc4CSG0
xzGT8G6+47b7TSg+zQhb9Pi7cy+rTxQ7GfHHWilHIPlTGpLvs/bS4XnPmTySuwIVg0LOCDBiDvfc
t0sCDUfQnKazTNn62ESRHBGY3YXVFHFuzNyLbAm7Csd9JTE3g71ziDnD9mhv/mJrxlMoXNgA72JT
wxof5NCl2jQIYJrJxvjk37dhJlqjlzfQGsWkkSuGIYuGSt/zLxcyJTbgSeqP/MFYlwMcnOzg1MPp
ITwYz3zjFv/D20D3BiolwzamuIqZi8wQ4kEtVXHm4B7zM7XA4oBgdBt0U1WwPqs2ON4WTrg2Np83
4WwWcTdOnHXS0LICxYxUewlWDVQKQX7dkl35KXVWvGKQtUBcwKQQqKXys3zA1cmRS+Y+V8CT2ton
aDqdC+Mp2N7peMejgLH/gvITOgmL2bH40bKs3NMgO8Dw4uvAE2GfT4Qc40Tm3EPAcdIRXl4Yva8p
8AHhCDd6Ds1IfRnr4JltjAVStjtHSlF31/+pH/xiJC+GgC3VBZAizP54pEo6S1zA2g9jH+6BbkJB
k3xLf398ocBdGj5spxTNQUC1GEiyW9tO53BZUn7Ats/2DY5/ruFo1yjUtkswdBJ2qom1XGKkp5BX
lUg0H/Xyj6SfWaLnG4f3W5jXJluouEonJVIUTEhUsE5jem2RBqZcPwCH5GTL3iX97tlGBhoDcSu+
8vBr3Z6T9RoQgK6xgTiZhlzmKPqDtx3Z4geDVD5jBrggHiEiLuGQwXG+GFl9P4v/nPBEUAm7iMSV
pGOKr8MXZltk7WZXuh8+piGV/fEL6hb/qozgxk5ZxCxivX5WigKThLUmRNc8UhpFUh6TC39EBHP0
phNRiI47sGofnNH20MvXVcz6rpQeoumfQqAP4iN1QcbLByQWjOdBxFj35miEsAhdDAEcYSDhaapf
1xMRP93l0xh6POE2E/wuGCXYT0g96zu5E85p5LOCNfAwG5DAI5mNYu8/iorG5LJ8SSXlEvqNKxyN
rbMgRGpJ4eDOOyY8is2d2C954hvUBePEfE7enySJBeuNHglJi8sTA8W+fKji1tvuSFppmhVX+1fe
UEWCl6JT/MqXpuG87eAiJNqe/oVGKGZtubE7R40/OvhU+zn0JNHB0Uno/tBIQHhe8JCBMTqZ7eFe
qBITAms5xrFB7IYYcDKbN5wDtlb5wTuUz9Xv2bR1tI4yxT2r3goNWaa/2Oa7DQxyiZsdr52F6vpm
POdnicUfhGwobogxpywVfxLpxlm7sDKi7/C0W49ZCRHh7zgLCLUwqIowDjzlFBqKjy7IWW3scX1T
T1GjQ7NdMieIst7AFerrF6J4P+4mffiKIP6Hjn1cWCfAG98bLhWCY/LE9uEZ5RwslkDxXMUfolRy
qb1CxeePfDbAcKi49yHlpssuhAStYzEbL5NqrkV4JIaK1oD1x3npGeDhB8oH6QXnPK5iel3kCmeP
PxgVlZfjXwrWYg2KXMaSKoyVEptmIHRPezlGWG2wAvXu437R//5KToEoWjIezQsW+AQbI0esnApa
1FE4rsgcl/8SXBQdNEIwVWnEZWczUF3pxeUVjm9iuqrslfhZV5Z0qhfZIHvEkefdGLdufJAbHMnp
eEnx3OmNUJSDYhQFRTNII4OIk1DA4GUvOrmxN8KafR+vgwNpd9EFLTd901jkgzD1eO3xR/aT8LPx
OOOw+/i6rXLsswsMPLwS0q66ZTcYhAw4Msn3GMKjWrperjqaIm0pCZRsE+ze3zHxoahCqcrhQzpX
efx9bCuDf7SG8bGQGNxWFcc/FxIpPhvWnKycnGm3fjDiSdGmDXjxuNBQx2soiuh7IyXQVVuS/Jw5
rfwl7P3R/2+RH3J1f5pQ03jojcvxl+TZkE6/MI4tbpd8GPV15oSbJoPX24WU6jo0qzi3zndoZiZr
NpR+cH8kchXLwfIW4M29L+fWX8yS8ok+YOS48N63rx2ozBn9rfqaFKTfsVioqd59frG23v44HncN
qeKD3xcSgUao040WWC1nrXv5h9IuI3hlzdj65fFwvZHW4S6UhD34nfkpdpG4DVmqEFW2FarCYoLv
9YzWZH/rjwXbXzHtW9C9x8/nD1EdQBerbON6FMF3jUsPzlGesdkg8+kkDr1aEVGS44u56tdyepNc
9NS+kHe4nX/8bKIg6P/BcTGMxybfd6Or7Fj9HDd+CgyLlkuLPs0RlnLRuo1XNCNHTX2gV7Wp1Z2B
ipR3MN7f06G+rhp1iJY91EzJE1XdWqm1PECJehc21wPIzLrnu46wNNBAo3UUKTJDiI6J+0bhiTuF
VfcF3VZj/clyeupQ2ZyR2Tu8lXjm9mSIIu0U8xJ0sm0z6wGpOgMecAtXQCRoxkCMsb3z6S4xtckj
Yt6ecuRx5B2d1A3ZHZt901tv8s8k9nne2wQQdXGzB0XddsTkit4+x+rUpHAgrQhmBywBbnnmWU62
b1ZhVqvjlCkBW2Y0CRTVVC+kL2mYX3qhQGrzicwTYShcQog7Jrg0176VdrLRdIZmVsH1QN+8VetI
x44EWoMAb2L1vGCnjL3oQdVV1lQz+jou7dOGS/mbK5cKl84/WrS9/1dY7O0r+X+tPlN7TUSVGA6u
YPLXzyTGmrHbqkHODAYVC06OltcBcjb/iAET6QHGlsWaZIVueN9eCpLQS2HFfmjdiGwbC2xJ/2T9
NJKMkxoJjPaTswtrQQkno+cF+2zGafpc/2HnuA/nCOuBN40cEiM1AbwUn0TaFQTn7hA2UF4SRugL
JgJIz24RUhQB/FolR0ZjGGw8GGLb76Pu8mFrcU1tFyFTHCZiPK4taTmuz9qMiQbWXpR63C3Vs9S4
B3yTYwd0AVrrdCkPhFUvknRd604LMwTtqhNISZwoQvxBozM8MLMRCnCvbd6iWwRAGH45glq4kpPz
jpTOh2RFiLaSWyqwmNKKuECttvtZEYeLyBN4EpknUqYe3Oq0cADWzVAyNPYkxTxZDM93fZ/SdFUh
O1kPnctRYREAfaGSIadGR8NdxVUI5B+mu4prJ1JX3Y2XsPG0k1jO1bdLE28F4FNiLZB7pEWuoal1
AreS2y9Mjemo8WZkAg1ZaplTWI3Rwsr7BVsSI2VxftzRzVz5/BiUNhFW1AsvIWXH6bYjAsmHymsZ
ltU8SvmhwzrXUV0Oc5lIOHM7lRn0zw3vrIkf+3wIXqAKIFhBT5fgfeNGrIWfRENF7mVsVCFOpARK
b+4mWebeb6GCQOD5AGjMRgkCp81PFjzbtYbqpySL6MuIqmatCYPJFOmQi2fmN7HCwFbfpjDYXXms
D8DMYH7MIkwL/WlGO8i1ulacX4ojrFAcg6nlj0ccTk/KRwSIlyMJdyAArjfALbJWsNaZE/KLwIfq
3fuBZEgdlkEXwFA0olqCe1KfP+T5Ewc8KOPANg5ssOe2OMtISAKXQWWiWazXiXrQOP8XphM42TlB
nwi+MOcwIT7rIg0Kft5NSzCGFLETwuOYUORzFRAK5QmrzImjbKcEmpufYFYYNY8UBDtSRo53MBdq
J08tjElGGDRDeEcjNoFmvGwJWB5Zrznxmeblde7MM9w9UHoWd6tQ5cKH6jgE8W//fYKJYcHWTjjc
Zr1lYN7Nn+eNke1MYPTCP1+WczRV2/zQAxx7bLFV+w6XiKr31vETz3BZFK0KFwXsf0FGFJ2zso0E
zUz8OHcKlsp7eMyTzEedMKqskdrlXmv2Z7FbEevoIUkJ+bwyJLLtw/0Yowhv+a0eKOz/aDa9hs50
orKNIGQaEdm+Rb5lxeW2b88S8KyiaqaRx0HWHya5BmPOwDM0rWdn0mge5xh30qYGmorwmzVFx2BB
fnE7BH3IkPe8Bum1Dka/ZGguMjM0wdPTFG5gZTjF9rl8FunpNjSmru/jH95ZydOO8SukmSok6A0T
mnnt0cnI4qcijB0P3now6mqpJHvPwXtb2WP0Iq+kr3v/io0KRkzWa7uLp+5sXd0Ql8HQ1GS4sB8L
vL1pFaJxmrMVAXQlioZauq2DIlVYPvHOnp+xfF4Dp97PfXOa0haHsxi91whWdpT43VB3b3B3G0P4
g6SmvxR0vlZkfOF3CoPq7cK2G5TVQdafIJKbMvl2KMWpg5KaxejqGHnqdrljqRxVJAOnwSqDKpxj
EeF5wDTsXeZyZtzg4zViGgpMloYEJ7HfKNFS4pYECxfxY2eV1caQQYXYz+aqkX90V1X7Mp0d4RPD
UC+cBQ0FQvoHV137Pm4Dr031yH/TjCfkCg2QwNFQSCLbQh6mLIsjWIOqHCkId7gH/825//rb1qqm
TacmEHoD/zwkCvX/FnnqmiyDvL5qDrlWEOzoydCUco0mpYWai/nYqzKDlFDNAvDXN6hE+3NlfkL4
9KfAiQBOUPozjN+JJmFmmA6HMow5xr0QYqmalv9E5hWI7otDzwsYGCSe6aDJMY46v69zww2JhguE
t+xen1xNVY7WzHi2YSFJogJVj106MKMdQ+WB99Y9hXfWvb2auM9LI/7Posd/P+ZX2xJWMkiPGETK
Cur9yyGPGQdGWzPVFI1EtT1oXgiFJFaLNpPJWZMckd+PGCSC1iRrNiQBJXEJ9uuWEzyv93ouh3uV
7EKq5T6LvOUpfWJGzGW4Ty1LAbJLLpBBD7wjtkgbkmK9qMBPW5aZrfkw1CkOqeHvJDuR1nEIv9al
ikTkiI5YwSUXjok+CgbrxreFKCisLw//AnlakB83vzkcqno5qpT5yTeJgucoq29oz6iAWjNqg+qW
twZ29IDChzLbW7o+CSVLqK9/IQ4w9ZEbRW39PmGsMX2F4rp6NeCfQi4k006dFktfCBRLQwxi6JIw
GC4XIqesPTmPx5ADkKe+DM/HgEjo4llSSS5zwo69760BhL134O4w2Xa9bMilMURW6PKBJ8G1+x3K
h85mmV2yw5I8i9s/eh9/wuzdvG/gWbf+OXqHAXRqHdMAkFGKuhfQLISRltIxvK/1SM6DIev4pegB
GyX3/m+Oma9bOlq2cNM0zh8qXq81YUJjQjvtQVvtpEp80paDjp5UffcvXQU/hC/OT8keRLKepoxL
BfcN61H8Cpf8cFzOBvQRjSkTmHTgFuqWAcgBey1KfLKzmqtoJdJyQ2h7Nd7OWB0cLcSskNCm+Hz5
CjsYS6Ju8jBZYtZu062RzXOzxoGi+WuxZE/udo3JJaQ95V0N2CnLa7JjX1AFNFeCzQOoTAALH1kz
GOI9lvE31Z/Cg9OywEwuvY0+XcBtw82SThq5f/EhBh78CXY2uDqIseHjZHIj03ye4jIwb6rSqQRi
q/BYSZ37hbyOFsSmrOqYeWnUTqpfyNTBD72zt4rkVxYAhc9dgHTlIIXzaj6aCR4SW2sbXGYoTjYr
hk4jcqIjKHY0IFR4LMwAnLJPAG4FaHfAHFxocS/nu5MRo2ysXvfNsJm70fSGwrjnObMl/wBATErp
qwmO1Dl4o7MdxFRBppAwCZ4ZB/YombHc5ECL2SiYN6FDpVjqK+pzw8Bciv76toteyHg7cQYw8FK+
qhd2c4Y0GUfkDuth2p5Hbdlwc8G334c9AGEP/8IzBxZomQ1QsmJbRtTm2ELg1ZJ2ulrj3PIWOgqA
gpKP0u2Zc3fsh9Akew3/dsEP8YtxoYrYgl8pW6+c5x2p0JqK8EUMLrhE2LHpLn8Ht/aXhTu2lEdC
nMnjl8t1SWdv4hQQWWFwG5pji+F9si9KefPnc6pKoZc6ApSVekRbU9eWm5hPWtINuql8pKio8y2C
OboFa4YPnkYzQvOJSZel2CufV2SbN/Q/Twov/WAt4OU/2oCy/g6zI3C8l/Yf2tzGDDHETZXBIPaC
gaDkj6lFiMyNplPEhhFWOCeIHwuQ48fUd1QZAeWs4KREyKo1jQJtn8jW7PFgJA9KicWiWQY7CxNa
JichOyBb2BYr/xbzb7dDm19FcGupYxo+WaiqEj9ZZShm57gwV66HVlC31XrkJjNUBTo0ldJhZFE7
mpfpD2pVZKiCStKIQ42a3XB7bbFKyrjq+pz4B4ebVceErGOkiicIaBatdbVg/inqtxtV3UdxHn1E
EiYQW09+K3V3JtNqYicd1zKsRc0PcG1r+u3JHcGloTPayTpK8xFJvdhWXvuaS/fUuXY5jHm8NpaH
49tb3riFbWDGCMxDqTRKvyPQK9tPPxXoF09ZgUq/MMR4IS+rZID+600y4/7hGlheHM9+74Tneb84
iqPwaaZ5I4pH1uivXuYEFZHVSm9zQlb4a+FdhhvdEOlee0Kbo6LYAL2uRSQWe3hSl/hzLjiu2uwS
DQ5LNlvodBYpNCA6kBQVkT/zZXXMGII5JlD+ffYPzywww6C9Bse5BSFaFSUPAI9xUqLFB+V2XRzM
VE1578FkEf5Eomm4EcFIzh6R+/dzvLdc9ji0TB7EdXcYuJ132YijHK8RF1gc0OBWvpDp0UImowZ1
cyL5Ls79SetRNZKWAXzJDGUlPYUnW3s+PtaJBungNeXTPttDv9Ujgcm9H4aL34m2TrdKVJbcmQGe
/T7JnGO8SR/gauQ3FIl0igzp2OuTZqhU9tMyK3q6q6r51yXKqHexemQrcWESlsObo0F5dD3xScbf
MePlwViZcWxI/q2Z/RYTDQxEm8SHRXevJemfYNQvKAO2SNaxpWqs5IX+OoHRlAUD0xYrDmuTEW8A
b9yk2u/3ZmL/JYRth+AOPsORIR/KEgZSQ5MDCz5uEmdhikmRloGxKVqtznW5hZfHmeHDAvCv5egq
MKqSur1GcyYrGIjJn2/yZeWBxTHxHReeUIQugNvwOSbAaBKlIagsOYQmWfCAiC3CGuAhFM6wsK5P
yPdYgfgaxeDArWH694uSfR/hLNjGBhiaFYX8+W0YXjWhDnsnr2k2M1rkdgLS0oVx+Toc7qB2eLQb
XI5WJ399XpNuPLd0GuN59f7sgArS83t1OtSohZoKxOW7fzg/UTk/BR3L3+AEBN9223HlSVaB6Kzq
9j3STMt35ZraOQ93sSRsJ0wGZOFYye+u/ripcw1NjsIZ1ER2/dmUO8nCiwJBZ/VibMk340yD8NqD
L430ivyK6KQez8ACnCsAMDTiVF9ou2cG7vwXfJ+3YIQ+PBi4qI+PLv14K8OqW3m1uay9Bs/TY04S
79O4Klkh7d5VJmQxrZs7nA0OHdjosj5+i8EoGyKU4T+UOPmWNFgK5XigZLjXRPOZ1YXwe598CS7C
x6rV70sjv2iLhYmx5rxigOQr4LAT0Co3uvT66s7/pht2kwL3nZ/tRUrF8BQdpPwc6n1hPxkSNruw
7nyuQQk8T+jcZ2SlTF/fNCZhi2W7f658bACDWKcy0hIdxHP6z0TXlIfaV690Cj37ESPiFyyGBz3O
M45EsXtLGa5RaDfrJmNC/9bsI0vdkEMYP2Tnu51T8nymTv5DwKMAdiSnDdRc2BKyufh3Ee87H9Wo
iBCcMxmgoXymYLfzdlXcSYUXu+fXzSPSxzqaE5IaoWr1Kzix2/+nyw1pTkJe7/3ZQFkx0rSn4msL
+UiNFdKW+o/rKAFsD4wibilLVJqKDdVTTQmrmXVAmhd35nkRh4VCFDrULrtDRutHVTjcitTooldT
sopb+TSQByWTRLR90DvDa5xHp7x43VxZMIhDbn68XHaGN+VKKQ8vADmqefrT6v78gO2YO20rI5Cb
kcG4hexVyG6jtldt+tTQ/h/s0MvyxdwKhcnITceawy4FzFJU8JtCsgZKiHhPxGqFRNB85O1hCGUG
Oxr7os5lQz6ZoeR7JK75plCdynN+I2VFXu92NJvFdTMu7hyknCJK5TxURW0jgjJbCdrx3uMSsZ4p
rapEudBl6CIZbawiHjtpSGpIKtFzeJG7ltP9c8Qg7JG4/FHnc84gieuzHLWT+yAVFn3yLxR9rmJU
10HJhf66q8dYCy7400C/gNpFJYRemw80cn8ZLtnRbr//NMKQSjzEIbGnf7CGmKq4KWoGpjaWKPyB
W4PtvEYHufzAWY+c3z7hTopWtlqnkwVjxv3EwJ6h6RpUUV1CN/tLzlS5/EuobjPtL82MPWlu0fdC
+PqDYtIiCuHklte//o5MyWOMJwO32yOLKlr+xLUeQDfhQtszF5Y1QKgK1VovlFnE7iSj4R7oPUSt
TrDv6U0g6TXxeDAnlZ9ObHb3Cc2CXszXShcNenQy6p+qJKaO7fpFfQMO3NYYETpo/64JOLU6ZS+K
oGb5E6+hcR+oBToIUyTL9vw8y++rLEo0kZljGW3HQwG9p7yxH1eWH5zwjgoShp4uOttwNPSa6Z12
HfNxCLYEq2Bucpenj2xKsgZmFEK2FxUIWUg4CWY+xPmK9qitoW254SuSaGQZsqO/cOxmeeOD0zZ5
n2lUp3PXZHFETG+UIjz3dVkNxh+toQQVGr9YRRZbb5lA79xfHHTpDl2UAYiiv2aqhRMqamefavcP
TaISpiMAS1jaMbHtVtjwPX06c4hh7Wp4y1Xg/goNWbvFE8heO5W1Y3ov/O+q2VARkjJDFp6N+Ejf
qXp9GEJrtoPwzL/dPdJ/y0XiWzzKCDzPIYl62S8NlzQ+lRXd94s2VjQwlGpNrbQZeCc5TY6n/+pO
kVT4yUoiJ39659wE/jSWRA2LdTkqEo/dZ7JmZR/tHG0cNAiwiFmuzIkpmARvM5qqUvGHTmCyzK0m
1x9kD8azsj+ENml5p2cQmFTkVBOWFGKl1qb8gQWu9Dsq5rPaZ/fx78vM8laYobCQ5ieLhP4sfhBH
TiXkynZbQet9QZ2tr8YNSJjXxZBouOHrYc+GTVbbHQtTn3V1B24ZyTgvrLRKRJJoHCwhii1/K5Fd
COmVNc40uSgxgt46ulHnx3/cvgNGkDVgdYcKQYL+QOOOeYlAIVA+KR9eFMm4pcztyJ5jYPxSAq0Z
pXod2lANT9Uvwl/a4cu3VSD+ipyvLuQU466kgEczzBNTi357mey7crrr4a/5CoN6/2OvMvYvkhgD
yDOqlRatQhD1x2IJ/wPbdEpMkMA6iBKuYYSzwgFzcqEqMj5EqVEHWbD1apWF3cDoVkwIDnd9E7FT
cFDgf7QyEYQgtaviVDbBfahqfOS34hVNDOdRC0EAPgN41Fi/yyL4LcZGa4VZ+B7qD/y9/cRdNV++
2nmxpACYZ5wtbdOq+vfCaOjINiLMfJhLXmOHQ3FD6NlUyUC5od9o5clV6Giw6FiudZ7Fy5ECuKOx
uRiK34Uem4fc69VxexSiUJHByilmYXtShfej/jZKrIkRrzfZdnNeWaV1n+TTu4N0f4xMYpci8lgY
8TmeBnx1X9i+vWYN/j5xl1Bs5rfUW7e8nMlOQzQcmSTmzSCpoKxAvZ3hPLVT++abwMfk3O0i2gf5
irTGMk+6xlp7g7ESOddK/rOu8mA7k2Z0LcZ09rOtBj5QrC56lSSjik/HM0Hb4Kwoz960neHF5Oe8
Br5gGYXj9VdSTS8wxVO6DI0PnVn78dvZlTdfo0M+jB6zkc9zHAIDhhScxI7gkoWYvY1cMRDJ4bEl
ukcF3VY/8T/KHx3OGNhKxkF8Kj8IvvnqwzNc12JOaH8v+gjz9od134stHRmACsHxzf1wHL3u0Xru
jMJTCbp+79/If/o2qHbArOvrSBZ4BnzuWnt2+v9QZ7H8DEjXRjcNWW4bAlnETqgi3WoZpFJCG1Yd
OAzEYAbYzOhMTHqjChgPBhdFg1nnMLlYFN6Pvtx4/JNioxn2RbJf1yjdP48HT0dw2pU+iqkkY1gF
MAfAlbZZXYG0krDOcz/y3AiKgmlBSbNHkqwLKvlXGwQhRyI4zW400p7tVVKpXdxEpjXJYxdcKuzn
XpoLBAmSYwxc40abceGwpuGxsnabsvg78fum/k1LQaQ2kE5+qsNQTULPZ4RK/gTKiyowuaf8l+He
MAiiY6E7sS5A5DFHTVcX4WYmosR7X7Qa3EeWm24RfjnD76Ca5pF7zaqcPh/e20+5Y5D+rTve8nF4
9V+BCRkQ1v5+odVO/aZDA7j7xGdsSW2m7fZzQpgqiKocl3ZIUIrQ3EM+SL+N7TSvni41JLwDnRa1
S9GwHPlvTX91aDRRuPDNEN8cjjy0/LTeISLkXz0M7DIXoJIFqs/xyBY7/XXJhjskZmbbfksBmgZw
9pPByxzinHg7pV/USfborvwaN28K7Lz4BDp8q1CrZtJzVkstEOypEx74OSFWuNZcQPAp20xjDWuR
1LKcJYerjM59ZgRR4zgyn2CnoAms4jtcvDgSk+lUhZs0iQ8j6P00SP1oEIsp8ra/4fayeYp9u+AR
JKmnild43BtRHrfzEh6vv4+rxBcgm/fup2SBfppr/RZhmXHjJk1nMHeO8zmioOvWzbNa7+XEauyy
W+ZRbUs4CNlqYZe4Sb4MA10Ur2wWQzyr5vkP7O6EOSbYEobWMbeYGEMlJNASol9XKmTj9J0F+Laj
vwT0g/of3KqgaOCdZXRwwuEKT8diyOaLNwFMBYpwSQaBt4+eHCqPfNPNBQW3rkTV+3zi5BxcCn1n
//Ng+B2eR4M/fgv2cOUYAtfmeS0nSIvfSC3MxOBgtBNDcafHcfS/nwMaylOmfLhyBGRojwjw4b0Y
rUEaX9w4+28l5zJ9iSioLdWoVE1Qwu2IxJjuFsQAqmcmD/aY5fI1GU167avHWQE6C7QI19K2HCj4
G2ABtZMJpppoFLkZesSa2y2doyjkyTU59ux7x5t3kWu/8YP9Pa77AOrWFboSHMGrovVR/G8dHIef
wC0Uu2iy88hdbruwmqqgEROiduC/umRvUFmcTdnTweXZcSmATnlsxblhkQlaMCvllBI5voSAu81e
qAkPhY4F0RYJ0E4ZTXYu7L592SZQlYBrBkMD+sN0ffcUzyrcfWQ591dbPXW1q5DnZYsXUOyQRnpp
YSFCkMFR7HyX4N/ZYVH8JuA0lBO6vKXk/40zM3DMGwKgUfhWzlUf30m/FaavI7z5GRk4cXrSsg8e
Yppu1fmYF4O0W/m5kS8p4KR95nkBNTYaqlxByhG4BR0dIm9x79DL+ujRU0Gkqf2rwSbLUPl/ixUM
KhvT0Gbqjx/Po+7pxuYUORrNk4fulfjf5WORXDqMcG9UBLa1OBhRDywJ7GKm4bHyw+TSOGbP51a0
QwFES6HXtTJJeXWSWKMyjLAdl7S2/trb1Mvg5ENlBaBwAZAYrKaFSa4LRHsw1DvtqvY94EEEdDKv
yKH7UoDMiwmbVkQKKYsRYRz2q9jHwGcSAP/yLsOb3L54f0J/40blz4sJjTpD/12JzhMP1BMeP3Fg
DrtLfw7YNfKTmrb9sVa1/F/E6tcwCPFK6l7uSUScuWLkpbsS0a17U/APt7Kjtxy/K+Rer2jepW1w
S0vRPjW0tH1L/dSZ4Jjx2MSJ0o+xgatDKUiIil91frJx1dy1BGSKay8VwPl/68J3oGP2U8jMbBEB
IOUxlX0Oo8Rc6n3UPOwcizHqVC1jKwgKdJ10b1QqddXzZEUlvNK+RiFeDozpt1t7LvsbeBY7g07J
U+WE5GPKX4oe4SOwGtc+K8GmIRIghB2yHap5Ko9WTywDHWBVDUE9bRiONoNkCVrf7R1QhQ1gDvdn
TfP0/HqrHJecEusWPXJKBGQ1W8+r+EwAGhDPhmUfoWa7CZcIYE5UjqjH5LpZsJy8g3AqgqOqDP6j
D2UBYcBMNCq+woIf0fUeMNaIrnSTZKlvLgIIyglOkCqQlumS83ZhR3rHdjd4FWYvENH/wcfRi2Rm
4uWMFLZjgAbSlGcIIUlz+cHY7mPRteP0gIs5t/rILLkx9V9RJdCpEO7gmbWf2Z0kC4cOhSixQA4D
JVLFYx6fxNZpUJuAEFWb0lYW3qz9QtjK9PnjF4qDCt1kK2mxzueXDhaQZwFgxmp9c5y3u9gmY/nx
9TW8n4xfvTP3b+bYENpmYjQ/oo17rf2vXFcQNHgs+kwzidlQn01bLD0CeYLHrIu7cglEIkJm5ciH
94lYYCGwwHbJ/c3VG0Ubc71yjaQ761QFd4JktzkZl71L3xnsrm1AIr1eGoTrkLAsvxqQJOd0Qq8A
0XN3EA2084NAK6KWR2xIAFc93dk0tlv/mC5le/8a6VOeFCAvKdTdnxsPyaKzcdl3bIBuFuuVP+dA
E6T7ieIvdlrD+yncA2DSRaIGXMGDVIVhll7rLl74iBfC5uKdtAcDeroXUAyiradYBgsKv088L25f
tIdikCEc4yKJrfhv6uCvWfPppucj+DndWkc4Q+MULQA7OovV3A64eu8DE//M7Fz6++m7RBxNAX3p
scjkz+5pmX7w0TnqbBxoLPXvpm2iXT7Il3hxKYM4dIsaatqAPs5LEJg9MkyHN6CxXSEfzJCwmMXZ
aQnfb46QAxsUXOhvFFfE7Q+xYyS8jzdnMHQd0ZfYDojgtEwULZ2aMRCUk2XpW5msd+mvxjR+xpr7
XsQU+ZBa+ycVnDqmz5MpcBNLuC7pwiMzI7YJLI1DalcvW9gDyle7iI4oMgtmZrW+GurYJwTjFuiJ
tkmUI6H+D5mbCgkXh8gkhCjE1Sr/PnWkOpQJ7op+dWAUg0L8yalKDNx3wL23smd8CT/jc1VQgnwb
a6KzPpbQD3wDQwFuWfHvcVAe7L3GvtvGrAM1tnCiZj8aD76gaAfXtWK1JbQUPXjOodBFiAxaKbMm
wmUKNrBfjd7UYhkGW/LpaB6OGGgD81BR5imwX2rgWUgMHudANaJ2bnyA8MljE7HVCz2XuzLtSSqB
ru+hjINX5G0zxMgWygFucBIXXRZGWORnHOap/htcAAz9LJA3sfa82WSM+uxOOG/degqG75hlNMzR
aipR1EybUkGSnf/s5LUzx1H+IEiSB+0ww2mbqqIWU5SrTTto1rqQVgobNSlTH3gp+gc4XKt7muCY
7RlPrkSCgMdaAoN1Xll0FfjjfMzHqYWLNFmTnmAWO30gJfIDaYQA4UuADas8/QUzU+RuZCt9fCza
BmUsG9cGZxtBt8kn1DdTWnZyZdLNbkxtDZXWAg5OTe2OYWOsyxlc/vlDpPwa+VkEC4zSNFOMSRrE
4ab+UdmwEwmgOEEXJdn+1NNbG3h/QlhssqRoZs+rccYFRgq1VVLXnmCoEY93Ni3sWTDkRohiYnJo
4/0SDSeUH72y56vdOTwbwMXMbOcih+W2IlAym2dKsy9+lK2ZZLdbPTkXnDK1GcmjqNZK/Uyo8WeJ
Uma2H1SXUataNWw69/R8HTAJhtF/OxMys2yzg/s+qIyrRefRAtRvGQ7gfGrG4iip7D0sVzldYDtB
ukxkb+5AmV7nWXAnx6Djv/l9hsouQdSE43bMp5eSkVAmggyGFkkutKWwDb1MRG+pse+tPR1XohCn
CF6+mHOU0HiApQYMmHhYp4eaeyqYGr3ufPyZ2zPnpJLOe9nMpV3G/cKDQVCcQi1cbtqipC5LiSjF
DCZYOQmhTXgI+5ulaWo3BurqYye6KicnDRlkl4J5ab5KTJBcolqVMmjWSHnI3EXyqTZHeP4GRMgM
YPJWAOPIsZf7l0gjqtY20Av9H6TC/5x4yFvO+z/o4r52hgzUs+ewdPgFTyOpFEYY5NymaubqmkVH
d89FrDeldtZ9ee4AzoelnxDGMKteY0SJPbL2JPeaYac3SSCQg7hutEkEjNxOx5y/KhQt8+kt3seR
6MTzXukNX7APlQh07P2ygrst1Jr1cieXFka/0rfqcD7XtYyr12rU7e0JIB8mvcfk0bwBHupvrAJV
zz6lX3u9/hgmv5JIGp0CNUN6O7uVJVFGrK06A9I5CcQgtgEtjyv7pg1so/6qerAdtxVnWSzv/2Ds
/OS1nNi0fAlaF4FEsrIA+uoLMtL2rzUprT2u9oqsHkPuXa2woyRZ/f48P7+uUREE96fukwQgGGN5
JLibh/3It3SeNGn3nyA6vX9pRoeVYS8rRBx4CSpSJFeTzvrK/Myb8/ltG1E4M+ZwfTM4riDYHWw9
TJNYPd3Gj1gW5mpwmNZiIkDR7S3ONzL+u1CJhZptCJEh2km65kVvrufoaxK8EQ3/hehl9DLSBeIx
WXFW2+EwNQ+mqVXhIu6k3NzVGhnYPwsyfqaOe2vLa1VKhT1Uxe2LXtw0vz5BwZu+eBaYWMjsRA0F
+sM3HO5KsLKxqGJOpeyQVvSWaDOJfL6wAVQiX+sSuVoUdQekLXKge6/iPN2VHDb8w4wY7UExaaQr
llohnWdz+EeT/WiLNy3+8+YdmH23/8nk/FEcbAJBJ57OTFalyOsXvf26mP0BSeuT4sivSjQoZBlj
gbHWapBwCOqXGpqc0NJuCivV39EI6BTV2MX2n0+TFUetR/6RUEldHZ7UHs5wIrRvHKMZ6JerYAc2
Cn4uhWxfzccG2XYr4LJIRgmhqAfm0SmqQBtgUmGu7685/oAQOj8CSYWGkUZkhdTfL5iCg9SHTSvt
uFe69el/INmEzpVARiH5jkKenc7ONkGw3d8WjnSp1t3WYihpIMO1rdtiykzMSOCzAYfkCPD2NuPi
aXPZ8S0AdYYTHKpFxHhUNeWaXZHjZ6gbLWezB7iFBC4LiwjDMi1fqxLzPK6opEINimaMnPiBQXWv
HVzpK1T0XGtr2SIhpLk1AC42s4CIOLSZLharOi3Ug+OyCF7BNeguNMQ2s+zp8EUjC+xGGOFU0sBQ
ByNyP7YzhqPcYHI4uMpU8uJF5rmMrqdaBTMDPxMN7l1NvREJkhAuQeFBcMgCo9YBT3VHxo2nBsOI
gDBkZMe2AqHo6XU7M59+hPPlTYDuoua8E+8VGpetLS4Z+fVJ071pb2nDb3/Ci8zR9VPzOmMdKQHc
tLu2AI3kDfqvtvxDU+cD0muw4iMcSAB/1JVgY9qoycwR4PuDUXw2kDLBCNuQUMGXJ/jmKtNRSTC+
wy46Lh9+tQRRwFeeW8tQVA4TKZRSwkFn2mMt6xdMCewQv9N5wNItKRAaKZDoUO/bvFTS98y4X+lM
uwwOjLBcLCfgzieH7yl8MI7hA7pj9UOUAcmqIVvvJ40RelKjrHwmFU4BPv3+drYK6gAO+DDHk1vT
tEt6cdLtMAIbDE1KzdbeQWNv1gYCayavCh8o0ZVJQ2VW39BHle4+ZNrVI9TgYgqXBM7iTkmqMQ5t
nsK4UJ/0RMu492OjCx5IWJ8Iy7Dr0uZ1nBeBB4s/A0hGUYrS4HGin83o+KMdrpyUTZf0P+XbIPH7
kB2xxcTSSFVm/Qpg+bRwnNf5JqQ7tgW/WSkw+Z+U3fGMwhHmr03DgU2/c/jiB/mNFqlgKlO0w6OC
gzFA3iI/45U8CYS+/BroUhy2GKloqRRtjjLkvrB3L4a9VueYvotEHMGpedCtoa0un1S76JnHL27Q
+/ZsM5VfI7EJfMlvTfKUun9ASLsc4UfbnO1CV6+kl5VcmYc9fdqCVLRrQa94Z2DrG/w8LCH1Zlzh
nNjgZjcyRRf0O5HaEQXvBGYJM9p2l2MpzwRXt6l++4WFGYJr4lcohbRetGqC7gCy4Mj+7eiGIgDZ
ZzFW6Kdpff0mImZD0aRIoV2H2eCLLmesx9ynHDASquSLkKkFe0snDGvMVf4Y2wtWPwgs79XhtrZH
6uWbe/zjl9y6S2RLEXTRc9cLVeky6te9BRqunRYwe47gL1Hkg7QbK6NaAHquXWJX+aLkK88TtQhx
xpP1kpDeUHFlrcZahoS0dJ0fpbvrDj2fFANr9VVYB6/KN71DbCrPQ2pUS0DudEXevX320gAeASTI
pco5mhnOEiiAPthISydm2JFAmYIS3LJS/BJLbJGHLiZwDmHDEqiE7nRt93JyKlWoYbg7oYpMr7+6
3KUuFvtwEUgcAYUXul8Y/US0SDy8av5t6C9paD3lBT6n/sVUYnKU1+nvZBLJaoFz7ry0Gbc41LT+
2BBykF7FVP5dyrpycxI2Zh2mFJGOQDWB7ZAQACEt/+NHY+1EauYIuGEpWryEhklNRLgN9KtY8Qdp
kFcOVbscEB3+HZpV88v+e2NFPaaC4LsdKsaentWow5ldk3HCmtmBKTctQXZ5bupdbsyXWkAK+3YQ
IL4Qxg1gJLgGJeG22lLdUlb5E3ehWmNZi319lkOJdJdhYBGv+L+J0b/qUH+ifqqTNSSjwtTifoKo
rTtDDCJczxksP1FkOEenp+++hGwd886t/DtGhBr4BzKpujGC2QVeSD3oEyxB0qLsIzdBBUqAjtHS
gd1vfubajgPSLskrDyxO6QJ4WxTUFrJI86myx6QfjfqJ0VulfHpaWRe8I6Lg3bzz1dUcjMvhu6xD
ob6pfdBym8MpVYfkrn1rjUcjdA3/ih16Srltqcji9XujvZtUazFKfbe7NjjXwTLeK2ITf6qn1k2y
91Nn5AIzRgae1K1tlcF33kSWP14qFCxSfnYL+vsB8wR6I8niPcZbBZDY10tSvPb40KVM6vgZvwiD
3rm6YG3QpdXh7OBlUfRhcSraPxNY0S4LwayKyGt3AHmIHzfU4KoIpIRZ+9tbA0zpySTxUU+cnyLr
adgE3Lvitga1nhqUEZsm204Q1eNBdsFwNd/3DJon63kKqLMcSIapVzJ6xPqwCb5uSCDuhDXkI0sz
YBG6LbT3W7xIh2Hxuy3U4jSvbjV/s/wmXkgrVIKA/zGyddp9V+cQWF2e3uHlBaTy+yUurUwJhveJ
jeEJKD/ArIXFpuLHyHMSwXe13O4RLYe5kwPujvdHaOxGA258otAGhi+0TnHimFCigUTHWyJtNlqc
CHp+J5pxcwYZOeAZfyeUFxAV20QY0/6yirTaUeLYgjGPMJMqq7Jn6jjjVGY93U6fgjpy0vQwZEnv
oUkorf0AzglpOKoNEpYgGi8PEaL/lVnS+tx6jw+VxSimhY+MOT3uhbN6R4pjbmF+8Qjp7UnRf/I8
declvlBIc8AXIz6wsj5kgnm0sXnj2KXMRnqWMRKgv/nYGe12zojynyQgxyf+5bHxq9fZwNMJDzoj
ZqZq+dxQm84ikAnT9/WbWR2xJVK0M+rhSOGIyG93M1HE0FuStXeaRuUdS75L3clkJOmmFPW5bNky
fcQc79XP+2QA7f73tZS2gv6LFZXXGxowpbpz/XJ+okghZJsXyuoZDaRcULXZFIoeEB23skl7ZutN
MJYxLalcFN3k6veEhZgdQVL6FQQTZyqX9GPZ7Q1qoFISDZ4q5lXkSic09Q2Wpr0odwQsXJGP3al4
HHWqumwPDR4vmVtv+F5zCY67D165kFna6OEju6St/OY97Zq++Cy0gdZRlspbZLLDzVJvExGQhgIF
dF3OEwLMq8PmrippqbCcW7VEupDhR5t9U+aHb/FDGeuTUSzIh4HCdH/EZAA9rl0ugRjAkhPHifpP
567nhj3WBVPCNw8yY/OkCvZVc5ThtTw3IHkVxveqoK5Tz6+XKdCVH8zX0nsuQLc0Z+0/osKoqycY
Z0B4wtwcR9oooDzKUvCc11Xy1Dq/d8nvbEUK5Zxg1w9SjXnBevWZPWopotSQa/LOAYqPV//girvm
GUC5azwKlbDJ8vs9AoHygkVv+/kWMLQj0oG7H4Wut1caZDA2vnuGXL7ZF2KYY5PHUEvkJf9/c6HS
lyFNUeuHBWvnhYEL5WKGEGN1sgde6ZH4Obxjbhz5tSkvOKmP4wQdmt1wrqCNPiZPW+/kxFFpF8E1
aBu5aNy3yJtl522vN4SOzuKQCHrGaj8DbjwaiEif50635Yf/d4ac9m6qbpKJ/f+FkVGcEEFoN3cD
HISL7OSeRdEZM24ZW8ZPWkt3Z8QltXbErFxav3ZCDxK3HY1oj+GxMHnR/6esEYy0ZBwnkbGh7MY4
2TnrJqOGEFS/tNvOBObgQK0SIK9xe/jG5556DlGg/k2iRArDhYMY6jA4ALPD0p1YbiBLa6Do/m5S
omFRXbhp9RflffnzA4BlyibVcBWdBMplpDhprbpZPKkfMZpgvQsP6p4MrtNbFO2F/cy0M0aFRaBg
oNPpWL6CFUu0NyyW2xGoo7MRqkkoCnqbRqawqqg4D0EW4gWOcbokx0AhI9pDyOdzNBO2nO1V4HHR
p95MkJqiYLjPL+CZ6ZIpXjY+ftGcueUSQV3DReLWbfxGh354mAlTBAi81wGJD/Yt9AejP/50hbUW
RH66u+msc96ZzTXEL+tBY27b6cdY3ifdQl8t4Ic9Wnp//t1DC7RZckxllgaDzeuZqJASmJZYVuIS
nIBgDYHCOtJREnlgpsJMXlW+o5uAJgiY07MaPuWd3G9bQmAIVuhLvni28G1D0cN7ERjo5TSddoBb
hYC+SEXX8UHLt8ptB2iPpks5Gw/g+vi3EebvSLFHOCBGagF2RuH3GSUKIYgJrnZPnjlKPUUIrIgt
Hbr5f9F+ybTkDz9R0mzqiUDDFjUAp4gf+z1vEX1Mcm9IJkYwLzFeqo2kuGTpV3F72pc23OiSvBMo
GCRioWotud+uRWiFxw1uUTG16AKtriqkUyJGh5JP3+fmZNQ4+4wPacAN+ba4/2YLCutysKgPQW8+
+/I7CtOrQq2BzD5W0rh71cPSapXFCPhlfagehPfGv81pKsdwmfKVzcpsA2Fv/Ni1GG03BA7kHdvI
JrrDk77fqjnrQXGYM0HNw6JPNYYBtRJn4wXNLTssP3MEG4CWZIt0/AJ8GDCNbtR95rBst/kehaZ0
2365YjXJelCyf+LVfozQl3Cjc1Ot9FtP4lgcJm+IGisy2LYjhoebxwefTC+AQQAsuMxLeqcuTpxv
QcpoixHuFKxoqzv1GG0aQ3soFN/OgG1BJ9QNLUCCE/rcx5VV9+vLygsS+dC0XVHRCISw4aMf/y1W
/073IvtfzNNbP5uYiFHoC/+2GEql8Jx8Tcv4YbPWlNBtiaHZH0ra0dpCKm//3ywvGBj+m1OPb5CS
pCN28VlN4lon4ttq1D0rNfLrA+eZtlEh5DhLqjTn+NfnorYfZi/UCBuqHDivnQ0c0EZ3QGq6LWyH
14ytRuWUFwchATVKegsXGgSc0nHCKGiXRXEMnoehCSTJrYq2uI0FxK0FmTnfChzMwzTSdDJ4RTzX
Vjm0z9+EdySwjuqxySZk5eNow3XRAu9sQ0IHSqFoR8dD5Ulx6TZ0D3Vh6cgjCCEQGmBIPcbTPenJ
eSCOi0kPUeFscUXk9w1dTXo5H5+QPX4X5C2QUNLt2bf8liDG0b4mvGitRyNua6b/3r55rPEQSRrC
wOGQlBcQ7pAm8Anob4/v1cxliAVg3o4jM0otFllfGvYLhOzw7fEnkSVbBHI3+gtWdqGh8/wT1GEg
88qkHUsCwu8ZvdWepApMIEV/BxH1MPdl1nSATMNiFNE/tHD76xnBLHTDknGj57MyiUUu77nW2TDO
8LrMGKXB76tVDVTX8ZHyun19C1Y02prr3Osn7Tb4y7UmwXvL1TvEs8NWg1brCKkjFuImPFmslFTj
Y80Lk4BC8kZlvbh9ERiCnB66fyd0Kh0ZNfwr0Zxfg/uVHpbqU8wwDPzyl5G6jkoTP5OdoUHJfsbj
61v/iFMkIy8SFRpx9hOt8VK+G+EulVPF+jv7awa7YrnWf681BMKgaKo6YgB2xYh+fk2/vWS6aO5M
RE1D/iYv8UVtbGvKjy2lMWg5ZsggWZ5D2G23WoOPpr8OtZLWbIZActQYGZ9AbIlQunFBaqDa6sbA
b/bEixQ+qNrrMAghxH+vk76OpSdnh20VYxzfg3r87DpjeW6GVOidgMPAGctDe1zJc/S2wCGKQHnR
BSYZgJ8Si2bUcb9lzuCiS5RYowfbZLi/Wdh0RL9Z8noC+81uQFe/81oxCS6n7x23UErb3lBLjg2E
7+QzhuggMrOqUw68SA0UyqgQ9qMzwwA9iDTbe7xUfmdLfBfn3QAT1UIg54b2pkeMmYRTV9hhkZfO
mdA2vFxBm1PhrzhgyDqzTkeANqQNpHIZY6o+7+uj+I8HEPY/4xOj10b+pSjm8mnbo3Iqw4TwZtb7
mTfCj4lZnz1ChnQFS241jYRiebJemO8o+RdXOjIpXq3MSuM1vhK6PyooRqJhz+1pFQPczijZxO2D
iM+LQL3vwrQhmvmJVcHPl4Pa6+h2qZXYeX/Pu4/hbRxlYAkscT1YFkdC67UIwYEWhM9DBeQ9ihu9
iJqV1QHV1xKZukDJsuNonB0jkJXpxRQtMzDj8a/rE+9aeIUgl3H/sp1T1HyxdwZsL6pbZq2d+IMw
CQ30nMi+xEgtUH+WV1xtdWr03pPOx8IJ26b7P3nl2UTRUa4aLkcLOg6ehgo7YGJATPKpkcbfKTpG
z/FKGtDmYyPY4iY0HD7AYtYt9VP+GIFrt9wy1xpISEYtbWE0m5dvafIEi+FtZHUkYcSTXl1GbkCv
YFUzdOG+G3X+JNBVvvLL3iqcs81rNHPsxYdrpFQGOQLLY6RcTrNzSPylnigv+4Ouuw6yUJ0654qO
6ndZwYm6g9OW6bLQPe1LvmLNMJqp0gRlVuJ0tEm1t4hkCbm/sqZRZW5165bz5VxRyjKU8DyAqLgf
vTE+dkiNWZ2WcPgwQNmbDIKLHkg8PsaBpLxumb9wNldofWC8OQFaxJ3qg0O8XOA2/r5L7hMd4W/z
ImNLS00K4u8KcPkA7Rm+COoFvVNm6jhOL4qi75D0gsA+xdL82mTeGmTvz1hz2QInsm3K6L5pKvLQ
bqMU0AQ6rnWik5PW9TGRcYmRL33vW4t1+AHIJB/zdsY8fxeTytPUqXXtXlY/Hdcks+FnBs/Ipttb
RE9Ntzb8jMKfTjiKHVfzeiX+PF7ZIX6UyhF60H5L3Khuaana6dxJEuqtTjf6/psqwMaHkNWNwsCY
Qzn6oWozBodexdwID+YQPlPxqAeaaQMjh5aNKPzlwgQ7vsXAn4y2Lw3cGQZDAYvOW27p538NJm8e
Q2JPHiN/KE7wZZA25kt57SGb1I7ZaiU290hIKBfaiFJMt7WtXf2uoUHwP2o/o6ftC8PkOoTtJgyw
5rTAG5Bdg1tkPYyrVrD6SE16VgVMOFN3dkwJNP3jQEy4t+i3XKr320O1Pn45ulCW2CbjAfYlhc6d
ZfSqMFyAfXAZ7DnScObUq9/v6Mp7QbjQDRUGTA7ZIkgTojJBhGCBwz5yOcCBy+A2Unk1PPjw1cRy
7dpN3aGMw7vtdIxX/azEiCV8R5Oaexvq34Gx15gk5SmuaneiBntLZteSCZtwtNkbctrUq/PzaK+H
h6MQCL8iVhDzKA9davXWBOBkqIVf8wjMH2yzGQYHPaorqLyck1DTDW26fyayjoLcP+9O5LknJvsC
57ZjbBA4S6zBZYWbdmRqTWnruxIXfbUbEXewzorGZgtb/mrLVXaix16IlscF/G1HaKit5Euy/gc/
D9QEeD2UYd6ii+H2pQIT6zEkTvNvVYxudsnPyLWiWDVPS1UvYcrHY+Yj6mbI9MbElyj4ni1O+BT8
NvCju2iKyU71FrKDpVXLBQ71Wk/7FmAPm/8lL/QX1I/VXdrkxV/C/0CTMu7NHvJ82BFapPdxefhz
EuuxkTTnkaOFTspz8bLDLB4q1viE3HAB3+x9NoxUpS+zq81f1lkv3lt2NkYR9pEz543+jVu1u/Hy
nQpaKrcq4jEdrtUE/1ppD9FhIuYLhLdd2qoKICe5bi0Y96uZcCk+pBaKHIrN37coxtfKglqwsYoR
MywRf4vBBhoYcX/DzOkybzzRfPHIaRbtxyhXRhCJmS9pOVUiHsvlpurZree+JWFFJ53yJo8SngY3
1t82NZMwIPaThPZeuCUGGHG7rv5tWm4atBhhT5uDaAHA6ui5lwMItlbAYiWj+FGgTl9NQFp4NxIx
1I98jRLinks4Qfl9BYaddKvRWNfVS6Ge0gf8LFOhdaUhBw0pnKbTCVquv8oWXUjAG8Oe5oLLXw5j
07mGN7Mk2rmvP3+zi+EY0rB5uPkhPqVaodeJ6naI/EbtPNnjkqDXOpPIPhSKt6AjOWYbn7IlAbd5
s2K9q6cQY+ziXH/bzOoW8Z5zr7z5/DgEK7Ylv/G+BV+YhkL14c/Wby8WDWZKoFYdWvPCDD0jGUGr
7MYPM0NX9l8zf8LjXSLceMJL5aEM0wO80EjKq8a13QVi1D4Oz5VhBHomXDCJ+WZDijvmYsFkGokF
hxhSKTNnqngTX2ASCuoKibZVXn6/8lu1V51o39AW+3I03djvm8fb560nMU+uSJUZZa2od3EKR8Yq
3BNBcbk7dzuPwFgWStjAflV+pVsccu5f/yzqgT/H8H/dCDEqpoQqNFrZNJs/adGnmHqF9rt6YljM
7e3q7hFBDwx8fbPYvytNxTteM0+VipoQfzRNukM5rKNE7yQ3o9a9oHJE0tw8TnQeeNlqMtjNXxcr
wkHUb7NL7qgOdPsfEOe0YzYvtU24pztroz2pCgKTFFAsdSWLC5C4qRm5wsAUrYZ2RgNp9SIz+NGQ
3JilbPcAwLEnB4E5saaQl3t+xoxr8pRINd9/pY8FakINoNZ3ScKV1q2VZYSrIoCI8BiPe5KLLoMe
c0mGilEhZYi3ofxHpAm/Rf8qOXpb50mi2jgJs4qNZpLIOWBZEkYUS6uBKVolZ4cUh1mPkBxta8HR
2odJ8n/bcVrh4sb9i6wO8NiPBV1gvyaWlzza6F/pi/nwhSJhU1Xm/uSjDx4IHJPUfvuhm6bLOVaJ
fAKltBRacsc/X4y7kb+v/mGDr3jtpHawKVz/8aNaX42gJ1nH0c0Ju14swaAStRwpyfyvFYV7ir4K
xVYKtoDt883AKhxqZ42kJ1Koq4xUbkfhDMRjMisYN1IQ1M+dKxjEBDxrwVLaJt8MQbEE/WTBHm00
7UYlwZc5+S4m38xvaDWYOR1Bm/QT9O5LR5mVW/i2CRNOSWXAx3hWlJjLNmYhJDwwGAyZTLjiyFDj
LYmx2KENIFTHK2/I+ysHPvvLW50+u5NrhWtTAySF5I7UCD5gCBywZJbtvNBYHEI8wiQq+pe95uzY
NKxe5F0w9Rba3jQOKDyV6AYAJP5DlAm7dwFdDQNU6IW+zCRSkV5AR8qBkAoSLcJjwUhyv/ALzSAL
/jnG6rvccr7JTT/HDTug8xzdVnplsiCfpddKRx5x7VptPiUsrVURr+1sg5au/GWmkTzWdh5jMOIE
LTgOWt2+K291MGl0LjrW13id6zd2lL+moJlrFmJg4O5yy6aM83EosI0j2ewdtietLGnh5jvPMm62
+FZLs3uB7Js16jGE3pArcxqdEwQqDr2rXarc7YpA7BYy1fqo0xgYDOIr6lE5mW0Jw4goYh+5XOi9
LsqImTAT1505GKpOONEkNdkU5fgZjtJvmH7ewSqyS8DSRHkuukVviEE06zBcZnYFoWStLljofhyE
fVt+sUfwiHadLAFoW1p4Qx/87C98wxer28O5vKnzH1XGH8nCGfkcvzgi53G8SRKs06kbmZ++9as5
P33iRhTZRcqIJzeGTAlndLJeBrVwfPmzPe9rkUDyJy3tQgjR5XDTP83E9Mi+og2krYyG6qLNGuM8
dHLAwKXYIOQBZi/ngUP14MdBe73OF2JFQ875SsXww2JqzibZXDeAAh30wCQxngAgQV3OS5pW9Gh6
EJSs7IcWbUaUIwDW/3FYxROOuLAM8u8mrpaNzdPWB5lBI4A9T24bKYCWWlE3KCfffNX/X+qU0evt
LikYrzDEbhkxOFYsp7vs3NHAafl//x2dU1gsTdvrFjAclHFKJDu1MNev3SUn81lxxJ6XSKgsqa3i
2twoPfkxxU3zqfizej8dlRDSpGneenXNJW1htMxrALfRt4+e87iBH+HbKtNRMZ8ChEYgNMOgGiE+
aH3IVoi2QE6xiimGkXRuSq/SZoiGCF7dO8qkA3YXweY4X3jbtyfJYpbZdqptZnW5W52d8OPuXgKS
TeUeM73KATKkDbNjV22bfuPBMBp8LlHP9b/SOAfaorE1ase0cAgNflQ28O5o3mshRNEvy/tcWKbI
ys5w7r1KyptDiFrMYjXl6hpZfyjO8BYeF0//7stD06UrdQGjTkjljcH3bTbSrdywtcv4rdWa7h53
B8K7mv65WW3bC1etKZqtll9Jpzk79X5OzmGtRULG9cP/fQqy5wWY8ohGOEU1Fud41rBU3sfsBsXZ
A4HVKijHsFbJWJNOOufCVBJH0PlhA8AMsQ4YtEinVWSkpSM2PACkLmac0VXDFoIYPIxyYKKtDsts
IwoNu5ZHnL8m0pNXZ6vMNVHg6R+6XOc5ouZyV1u7SNZitYtR/23Gy7kDRz0yucxZccCbuHk45YE5
3XJ2xLcyMWfMxRypGMO24SgTvsZHW6hz4ZCPhewBEXk95JbIv8/7ZujlLoJkgsmnnhkeoQ+Z/5Iv
7H3uZq/qbNJWT5NRezSqwUuxfWrgRXwrb8j2Xs1/AVwxK5ivHSWF1JqLQ8mmTlI4ZomaGDdtU3BW
7/h9yHfay/e0KcGFkg8pvC038/Ep4yQ2wNHjH3EiAOEgG/Lq6g0IdVNTuSWJ7HP3leGIxnuewo5g
4yY8bH7vznEVuBSu0nM8NFP/UGHtRUooIx/xFne4fMMuWkEB7TQwS/VcC3of/uhfiqDghFnMQR+T
V8PwM9+GFVgd42KLb2bg4cQIzVm18DJ2iZtp4/i7QaSB2O/HEdncVfSSTCgXpMX3FnKA76om9hjr
rZl9rLTtXBBPmT4YzI1f3V8F0aCr6akT9Jn5hB13OlgDfF9T2ZKj827IqkR/fsFwSf1Pp7KpTd2h
UGjfz/baREqOe4kZ0p8pVE4MgXzPXGE2CUUMoRKqb5OTNkGeRuhTMjH6BtUqqZr90mNq8ZP+Wx6g
ZbNK8jVrtGIFnHemA8jSSHGMsEQYPDJ3ZlQ/uujTORTbSj9pmeNPIHVz1hv4Z1/7yq7XFDjDi1uI
Am/dRStTQSAJ0L0cPjXTOr9ksyTe/0zPhVnT1tEnCY3mLgfeVydfzq2DGgD2qNO+cPr5XAFdF7Dm
EvxljlJmWQqLR/cEfknpHVzCc2JCLOrEC8Zc/KUh8V/tiluTwQ1+sq0rAdb0cno2YuDuObAN46cg
CVgb0VfYAvU3c9q0RB5M6pPc0iC7CXk8ZNV2gvHn+mB1ylTSg3D/XsFGb6BnL0jNTfefo4gLRuvp
bKj2MhdjaXGsmrzAajfTwoD665y+nbz9xWE7SeCcalM1XHdDoMfJvIh1KZS1dRNb+2KAWDhN+7m8
/f5mAZOqsXjC40yvHP5uszfkpS5ohCCtgej+2en1m/bw0if6mpW3fwQPJq8P6WBEZ6iX8WZX2FH/
PJ6vTiW2M8kq4QqjCPBPdX6ofboVtIcK8j8OLC6xmUIksWQ0NotQ5CXzG+APO5f63Xz9Y3IwdfTp
FxwyH74JLb5JIX9AB7UDoKjPmtj/XWCuDPpI6/8WGP+Y4322gVqY1vH5W1uRLrYZ11fg/egf62/h
LBwZUEaZRzmCSrH6Mb9IRw29IHo/tZxfOC1ImdHRVR+w1TvLug8NJl5WpJBi46wYePzyIaT4LtlB
c0RRw9tcW8kEFeddM54SFLmoaNBvWQGydw2WupBFXUSGqJ66wNoT0DVF7xVyDLKLJSrDOBV1pDHG
2hh8cmchWqyhGBv+quLS/0qNsRiL6lR8MQBkF7CWHc1HGB0FNMGZ5oe39mWjFSreUaBPHTN5cN90
5ClKRGonyz6VGPfxSixOv1Y7mcsDTWsjT1/WDQa47MjxZCiX1VUwnLNLxdyTqAmtuoXEiLgE108Z
4eJh1L+4QrmlklT3DG0IwXAdbCr4n4AaR4USFgkltr+itwEW7dsD1+fQjbYpcqxSbaszxG0/k8as
BQIGAVxoro2LgUz5GwRoC8T5trT7ZTcKhzjMTCtyqt+wGGFqPnrKcGIs1E2H2wbw6BXLN14PgX16
9w2NBaqYiabAojYHAn7v6VQjp5cx5o3GUtnCWL3kXtMlY77sT+2fArtHsnZBwQN46bVm5CCOMxPM
MqVsFXwXIMRHjcjk79x+m4lfPQjdXx8EE81Hxwzu3rwKo1V0PPHQwl9+cXbPK0uTJ63qF78pcsWh
Yhu18xNG9Oyt67XwTVBuGNz6Ru1lOtNa/pMBmUO6AfewQorUd0/qDB2jVjFa6WQMM2d01p4rzdOL
eoJi755K/gvdm3/dK0b8OJk9X41pJQ4gV7GZJgwxzNsvIjGlzRy5h1TIy+F3tQm22qNHwUdgG+C2
HkX+9rlkgsUjMd/3stY714xVzAFoQC1xnPN/RYqhZQXi9RoUlFEgNz3WG9A3zdieYthkLrPrr/42
kqhpHBK15htTZNN6FO+AqYc5zKTMF1I8E9GIXzRzj9zRSwGYzcAXeB86m+z98Hf0kd2hEtphhJ47
rBbnUcVeFILXYlO6LdL8LGM90GnBxdM4nm1zXzJafBiBdXWX+IhD/p6Hi02yAH/hYw+c/+2N0zS3
a3Nq7i4BaU7WZVGe5f/6yO2Z9OFPqrQ/b5MtNZ4Ae1W9HLrw0sPraLT2SnoaFc9YstJh0eNGfLia
W4paXpaqtkHvuRhT+BN0cByuZusQXV6KEFwtZL3LGBw7S+TVHgs2pMXelX97A4/lzd7+ddlIBqMz
ahcRQaSdH0+khOwsZuBUlghPK0Qnnit0vXS2eWcj2YnNnCZTONp2rEoaWTLzMsL7HHTUWZYaJkH1
yt6scj3xeOvvH4kjzxcUF0Vt4wLn4GOg84utkTHRU4TtWhpdRQIdK2FqxLIYQfAMCGcHhei+PNP8
/J7TzIifVwgZR6mqkrVBX/EZpwYdaHxQbvGT8UTFMc5A7WdAI89SZp39qW6kghD06tUIQ9EOJrNb
X0GFa6XH69msgc2wLcnDgZQSWhAo3EI7Q5Xi8tbZHW4fk1CEZyCdOU9FT2lRUrBpErX5CdMnHfo5
w1o7TDfRPtTtAx5HZGXL8ChQi+dhSqhMzfkXRIP6PQRknPmKxAJXhrmWDC28p1Hk+5DSnprvQrpG
mqtDj7cCENrkxV9/oMFZXsk0wLqUzvm2kTFvGxK9P+uVSnDLR7qHIvzNst+3NN5Y1bLm3udOgS6V
zou3IHv+BEcY2zU0ElGcQWatG2rHGn2ELgBRQdfmMEtrtgDJpyf4SoqihpeHios1IPRlANwqmOu4
+vmFY8jqTGFdIus1ofSYt7jIPtpNHhzqJSA0oYm+bbaDKEZrjuIcBHIYrJEx3JwGPZjGUJRiiiwZ
2/eh7f9wmAwxO76ppL3AQUgrL90wBpqsNcrU1okkZeMN4qGSSUz/Nh7qAIBB5c/5QIqu4BNhza/1
tA6YIm5M/RBRTcurYTXW4Cqz4o8izL2zIcjXBD8cjtb+vZXJ3wexmIp1F3+BAFSti9nQKbgbT8R8
XzW+YUsN/tbRF5ZvDVPp5E9pwlh6L7ZYoSL6ZKgPw7CZ1El0RVga56D/cJdhbmD42FCx0Tm1RRQX
+MD4jfvF/dtRCpDuP019C78NP4RL+85vMDKz/QTtY4F6s5LiDEhDG5IONf2vrMZNUYrNvoVRFYGt
N7iLRKToAj7/aG7AcZcEl68RtJuw+89YwEEK0hwP3NPPiFGKR0TVl9LwJcNNUZno7Be/UGc0gtid
9Ep7h0tDzGv+/GX4iiho40QCFMEPIWT6x3dExY2KI7464HRs6CkLQim+tPjSe1ke+p8FkdNDiji9
cxj5EnSgvMnsFIwkdYtnVPxoxN5AeAnkxGBTLODNz59sShTKhWvZKNqwENywH38jQG471RbOJD39
2Rtbc5Rw3+kPkjd6yoBvSO/swZO+5Lh9nfXa/D4m7HozUYJ+sRB/csDI4sIVFuT4M6+C9O2UJY92
pOT2rDOR2p3Y5eH7gC0ie4hGJeobmaibo9YsmRan2AjJAwVL+ec2zKSrzxzWHuhp6eZzczXVqhIf
Qxtvn1+RAJOOUxHp5sqaejGF+2TV6giJi9UcyGEUUFznyO5ZLrAcvLJSahY8+9zTehYnhueaKJMt
aSZH0UD/lI6sEPf5ASrp5fGa08xFXyCyimfRGsbSDKWHIVCkWV3FBV7ywH8Fec0BD76TSWTPWyHh
xG2dTGI5qNPbVEFwGk9yV7lTZdcqOT7+e2UnyDfqAcJu7O/hvaQyLnEpAUQabJxIKU/z/Nc2RqO1
zBto4HSGeQakMbg9k4uNoPXjSNcoX0HupkINUpN06Nvnx3jfODbk5qYIJJ7W/6xq576RLfQET+8b
KyPi0sov/JsKtMOMiYknGB7pzmrhk0+5D10V6Jg9XX7k4jCInBjYphZb29SDNUymdo/mtSN1il2h
2I/Kf/C8i85j0DrlUC5uvR49S4lfMRQHkUuMHotyTl7KzcbwUvNkHUza+YrkIvcw2SDHCtS6Ty5X
QFrhfrkurbDD0WZo7OuurHLwGdlPixbdc8XisKvC9Hq2ux0eolRP03k+ZETubkNghUB+WPLgwBUe
bsYqvak79XjMXY9AT4cT+F5RdOTccGdLQvcWPrkPZOvqrS4rw3McthtQSdqnFnBPCLBAFYYe7u7W
VT/nB0+AL6vgZ0zKYp5hTXYj59Mbiqasuhzi2MFCM6c54+tHAEALcGF+iAZErthQNxm+AznNGuOg
kXo8qBceNkGFi6CdzmyJL/DeNbB8Bfjk+lOxTYmUuBHXUpy5KTfZMzh9QK6+jCh6fjKADQtl659t
XkIwfWHGsXnOCLd4q3YsN9Srru+m+Zlz07F9dVjMXRKkqCDU5aCYa90oZa4FCXuaTxt1s3JLhLPB
/f45bY2P2KwfTqcfFq4oojSN5AvoycSgDvFx1THiRu8vtXCTUpO13qR6CqsihBc5DLtE/eeQ75G1
SIDAfP4cc7mo5+0layIpQ49WoZZ1nY7I83XJagaxJmy2mB46eVM0E+/cKCLNL6vgRXs1uj+ffk3l
PfnugkfcuQoKrEN2F+9Xio8BmUQk68fISFk/y/lW4rEjO1TtTeW7bq1HUXbFzsiwhTia4z1bwR7/
EAilpsrM8DF65y72tl1oBd8cVFbr/8sn+R+xdv8ymdNkB63Ie0nSO+Xy7tunn6Il/KI3qwzJLarH
agghhNtm47Ij1rUcq5Tm6RkidakIDISn0xFUQKjBFWnGoRzzZ3xRVOF1HMzsomz4X7CNwwSXxG1w
/5OVOzBkEXSPO8pKYQ697Q2cBWZOpt3jk5kQslru98IzyF3DmFebeiOxA9IOW5x3k8Pm9e1MpkJg
6v++Gt3OzHqVdy3D3ck+i2EDZvjqsKxe4FawHMxdYUw2WoYo4L6gfmHP7MK6V+iV9+lWFH27meYI
it7e0b81Yc03u/GSM3kgMVaJTlElFrD1uUtFoIsNoWSk/0bvi47ZTyZFMiR7eaUvOcX0ToeUNkr0
oHjqfexvMnpyK5lqyx3IG1ktV85pJvcV3U4Wt5wC6swkxQJEj4tedRok496DIDiNvi3DqRRtCtM2
FTbjiv36D4D5fucfWXs/+AI2y+TVoyMTGhZ3pgOlDvfePQg6Vzfeque99L+nziSxlV0g3m4kYp+1
EOVWyOv3xuStWqFJzEahxmKDVDN31Zz60e/9+YKdZZqGKF2zM8WrpH/JjUiQ+ysoAYinVCmuSEpe
7zmsCGSsGR2Ql5ZiG/1zEC+fSpEcZZQMq73HhR3BqTpPxYolHZuN5U93+RTAop90tzdYTXAiEikV
Sqi/NLr0vH4jJlh7yijME+ptgV+cZwa16zwMRE2fz0Y2Y6M4veXwo8DIvK7aRxFqwW4PEX3LGVux
uWTlr/9PNLHgqCiI/FsYe12iF2eukUHgrJ+6acZoSM/RpiKaaCoow3OrAkyK0PCIhPzErYTMa08X
mzKl+s2H3y5k7TQXoT3ZBXBNy23aUHJj6NJLtplsnuX8YMBRLFwYVuKGttj0Pqp77m+V1BQfc0y7
WlH57p8OFF8VACBaDD5+j1DW8TS5Jn/aAMfRRIGqleCL3GKsdXfRMZf5PXqdNmBkPMJAHY4RimX/
9BBQ85TOT/P5LVOp8bWFfxR4SjUJ+kxGSFgLD5laDA8+KWb/O/xnIi3cGjXX86BbhAUsccAs2kEK
3S63vAvg16hTCYR1hJkfeCz+e2rlj8osaxrWhYz7RUZ5SVYU4mkfna1gUTi3fVfhRoRP6UKJoVEg
JK8BdzggvXY+UODbR/CuDM4LGNy/HEt55QTfhnI/wclnWr43mU3ijWZFShR+oBnfQOACuP4GdEUf
0ZE95CnLLaAbZa311N1ZHCbywJAOyQDyHW1FmekqygW46J0b3xM4SceBobEciRLQmaCgUUBxb/1Q
UUZeM4qnO45DWgT7upc5bXC7a/MFPrR2w44u5jlP6SGid62NMum87RxxkuENH8sO6yxn6YkdXLOh
i0ysM15yGiYl1XdZk766mWTGpz7EOE2E5pHPKcMOp4BrJfkbK2ciotM4GTXVOZop30BpD/rrup8g
HUcJiH9LsnIp96FFEBSPtH9Q3zY8XN76rSU6sqz9i8lrWKbWl0jX9laTZxMS3AoaFh8FqboJMHm5
ulb7Gq0V3A+94L866axUZtkuytGQiQdfILNISjM/Y2xh2xagJkHoI1Xh4MxJ5cui/Pp3MdcycRa+
GudoovY7X1Ph3Xaq497r2rt8fgeXLvcqcF/kSF84m1dUofzdfHpTONIeqTLxGSJ3qiK+brTnRU+L
PqrklHN9TQIA+LG2k9A2CUL34VFuRpqmLtG0SlwxXqPE7y0zbAh6UKGchcBGa2iJvVqtvZZFHuO4
9yYDlXqNtBNJdEB9LOIbLpMEw9sg55LDC86G1GEv13OzXFQ+8fkSNzICD7SOxaN9Jjx4MTf59+89
63u6FgrJsC6LbSWChH+C8bzh9Dl/k5mggeUdC5Vubrd3Vilga4T8Gr5DRNknqZ/skZjyaYFsSRE+
kqY/00IDreeNVjQ5owH37vyaZ4aTeeJJrFVxIIu7sZFgEPlcHs4PmvOS5D7UwIsYq163l+A4ldv/
wkN0ATkZpIO5I3xm1o7/uJ+KMrpzmlrycTzwaHl4OdO3gT9j9Lbirs/HSsbUZgnerYpZdFP45C39
LEwChKlMAvcOFkqoDtRX2Pfy2bDN/0vkTTN7ivs59jCC5hWRxgTkrV1LcLrvZjRomcGZdF/1J9jB
sDZYtGPIZQ7XPrK1zj7pV1V5RHlRv3TTuid80G+jw7s8V+FYVF+V/cSEY37ndj+yYKyGrPBZi6DG
I5owEbODWPiTf1+1gYz1MtND3svmy/Ts4stGQrR5FXnH00O33OkPxjtVuA3l7AO9Me1yOMGb6WMY
UYHpIuq2U677IJ1itpvcl4+3WSqDN9jfK2NJ4cmzAvOBTIYs8djjuybO/oe0s4emN4fbVA6Qbij7
ZdQifgBSGIzZnVUX7MXesmAwOCDa2WbwesEmAdUWjftw4vEyQRhs49hsXMxr1htQ23MY6zd/V6Zb
9ABpf3hZQuYFRXwUk8FVkrr6bfaIP1P09fo2kQd4TrsKS9kO9uCp9Nw3gxsPUmXE3coikX2i4pV/
bx3gKW1rwC2CadudAQqQxSH7YwQEZ174AGWdnhAytH54aqA0KB5chMRsvyTZc0ABRk+heFSvk17p
0DuhpkkatyMVFq1QmDRruFb+eN0lT6IF0GQV6plSkQZ1SX8gJzYuqQc2NDOAfVQeT7BAsgJ59Z8q
j707X2ifeCvhzlJm3a/My9uAUqEtrFb7yAfzwad66hgZjH/ggSyxHZLlioB2d+9oHp3GPi5rZ3yD
GU/wsCt8OiNDV+X1uqZdA7TVHB286aQ3+9laZNHJ38D3c3gZu1itIoznd8kuHeshSXVH/rEpLRSu
lUXNU2UfvZ93/TTPwJdXjbjqFbtzc1sHlV2r9/tljXQFaN0pxUoK/x8zrhWyf3VJBwgjHy0wYZX5
Rs+JoXh6ufh+2lZREh/6gEOy2Mwpjo29U60J9qFlv+dCYu67DP/NEL0iL5wEh4G0Un5n7D26xpt6
rpFoVhS1hKGlxdCFKXozafGt5SgZatVlBDyVhVTKj4q8BlrlRU0fPar6UT5zFlzZzPjnKU9OSkuo
R5Da4B9mmyfOY5ahGcQz7Y5kzGApxpp0+lf73KKLaqv3L2zGwZd7ErwtWEKnmPfeRKVZ4wA5G49l
p0p1LONcxT5RU6XMNOeD7ZJL3+NIyW907za0TNSEJyoagurbTzVGPFAZZYWmqH+/gGzqwlal+pZN
ks4eLvA6+9hCiHuNQ/Vd+sq6WriRTpy0DIdOb/e8XyrEnofjm98Qqwab3DzhbaBONsMqlQKGgH9l
tQ+Op0FwXHLBgCdB3faQi6j+9Ur2mVzaLDUBz5vG1F6k8uV0E39rbFNdoZ1QC1VN3tl64vhbjzb9
ovrBXWejyPFr34azjm5VNUiU7YWSikEcQS+Ac0o7f97U2ztraZS+zjL5WfXsFMfPxhcLAnLeSN3Y
L4zcxDk5KPFDAh0sB5Adwp5PRD6VPqWY3YunL4A1oQXW4JMsWiZM8/k8KShr9qVynUzPRd7mfcWA
nQ1eGtTcwx+zC0crWSr6ifUvEdhjhwhHHRf0Zrl73ae+3M9uChAUmE0wc7q7pmrusfXoUnsxGisl
IxdcyOyjYpKuTPsRfpPgzRywEaBjfMx+LB3Kgm+8QfD+f4kY0HSIde2iO3PU6nFs11yiOaXjlve0
N5BSUIICrRglEl1ZZyQYXvwmprwKYr0CFNZfdKTjacr7F6rAQtXtuVvk5GvWZ9tmO5uTxEoLyLa4
X3H+IS6zN6ClNYXw3oh1H6fEZdQ9n5ad7CIhZrQKsEv05Nf8Z/zEw0Q0GtFIhn2agsN+uKH959o9
LsXUJCwqh33KZa3WyocSyCw/QXbBlOhwKDHuB0QU9yW9X/DB4lBMt7DMyU6hiLt3dNZXCVQsGFh9
0RWGz26/QLblFwuwBvJtjBVEgH5jzFcG8eyM62T5ANQjUaJ+8dRh/quPFswfgMkW59dXSLTdgFYY
6xh30dBqcAUyrY8w7V0eQD8sJCfwydYVCGOjrzBv7mMT88n1ZT+gvgOlLzVio0an29WJgEM6DoIX
FiSX/wAko27+VAT2dSYCI/SCShZrMjJSW1FwMW3yBETt3sPxb7FKk3HIY7Qz4ShXkkDNTEFI3Thq
Kf0PxN7fsnHCBqAIHkVJtQeeTu/gVfA342Q440L/tELupdzKKm854Viouaot/UjVk9nnsdmrWgid
FMoDNHTJ1rmEWh6R24t3/54ubd3XWAJ3XOvRVayvYt6qyiPZhvlLtTuNPiAxJ7GDtlSVp01m8nud
5/deV0UENQa09dy0cosZI821hBDMGYoC0Iv9wWuyCVQa9FKS8p0Dfegsx4rCHVqtREDXP/MrKtHl
4JEQeCgjqKjo+p/PiGjfQErPg9asM0dUougXdrQLYnmZ0aYsf+OOQYYtCGBjv7rjYiWc3EOUxYtY
qbOyUUCL8T0wsPqCI74DNKBV7COFkC2+gDspe8iOtsaw8vpo8tBfPh3TxSDZyGID+0NR1Ug+hOkQ
Rmp3WAqj6m4Iny76PiHDugUuUXS0H3gI4dWLDeBhc7/NG3v3Nd5bV5aC8V+vKAEquRAgnEfHm5/Z
NpjWXNw6C2IMzkHDgLLsgaVwVTpG7ML+el0r6WK2toKxeOMQAIXQbk6Qp2NMkP91zW5wMkohaIf/
QkEeH51ekhbCASrc0sI4YHok7ipDHyg2rkpYMUcJQVBUQOyBhMgOWIgwHeLngPCI0p6HWogWQs4P
6FiEirvlkP/3DwOy1ja5KKF44udRu4vc1PaLt1br5kbOmZvv1hI0IXuyOxtMX/Lr6di2x7PoPgI7
qn1FE2Eb5yKgX/F72C/Tgls1NcxYHW1gciibUFm80VnWbQgNCZH1mORAIALzni/T6lPhw7OmkbQH
zkFKnUBG4KSUmbOwByf6HcATLJygzF2LQhsim51NmFX1R+11Tw/I2nrX2Xp2tRxUNCEe1pP4ghtF
w3/hydpYzRZXFFWbIgYToSGNen3ASdx5ttqkjQa9VEWt0+KwdR4zAqSQwIRK/ALmODHtsdD1exON
M2YhbI7hyNaP56FfJeBljo0fFZwAjrlsbcSn64DX9q7Fx3t+ylntZRc3QNxvKjr2VYc7Cnaks4b1
jJ1QnthQ8mYzkdYence7YTYbqZSK4Kfmt20JL4XjMkb+bpkF+ubeRqhV/PodIvizNgZUthY2z7ng
8skMjDAlwVUcbJNXvuFnWvX7tc2C1FcTXwyL8sHLSA1iv53Dbb9SmChotXhiALQl2l3tuo/9oykr
pH4SoLgHy/S14IcQOamHsqfabqg/Q+FKfV1VatqAmHBkz07vqrOM8Z2XZ10dwpeMI5g6X3P0+4c9
8JlWQfmb8oparJYDI0pAGKeI7chmvIrP4oXZ67JhXNvlgEDviWGWPxcnM29J7tVP7qRbViY3f99n
rbraBdUEPtR44Wn19OWcdMZI5Nc8Ly0SuRHrLGGrDCOMCAFr9v4m+DodlUHnAKYYpjkDxFsi8uWs
mYNQpTDS6Rzuukl7sNU34ZCTvogrN/jeVYRfBZCRvAwTeHXpPiS23DZdqxMsJjiBLiP7F7i+Ia44
k0s4dgNNs2oLFUhgljP5qer4h6b7QxHV7vsNYQUtzDNmGn86c+IgKPgIoDmeohWvZiVPj7ynqIgo
xWItgWs5QbPiXPiiko5dZXBzOGhIKDoWmYeREPPGdg261yl0wzDM1nd0LorHPQpKyyl0aLc+wJnu
8BFr8nxK74fp03wn6hdcCH/UO5GQa9X9gp6/iZ6l+6nJlJ8iQo/2jZUfHp/GQ8O0BL+fzSJLG9ym
C1afKaGpMP88lBCMtSo1ehKgy0P0vvBK4o6T0b/mBLlHMEXzMl3YsqzFUqbTdWpdUiUdG2XA7pNq
N/5iPtz3dTCIJ1EoyuzejQTHVz87MlCa/garrN7apZtYCJfwSt3/Ztz8Bfj5tCVaXo1JUPJCpqvM
ugMYwJbGtwmh1N2xcPlJ9UVpONj3AtBva2fosOiypFIwu8da5Yc+ssDhzFrnQo/7QoyWJeuj4d7z
/9vKPKR8yjb8RBsNJ/Yx4kmIWPBOUrqp/KuG/l4EBNmT4pwKXYaQkKI8h5uFNlvKIykxNV6UhvnD
bcaOQbpoUGzg+Wex0SyyR5b6HM0qsQtZ0rnYQGQz5rFZ7wYtFfo6RmUjdij3AF6B72aK91aXfnPQ
kcxxMCVLaF2tJQThVitYwf6lzvCCK3O1XFwF+1j2/ga/m1eToHtH7gt3eOBg5S2X5U/jb72gelsf
WdCMpIWm7BWJ9J50CXu08OEF2XbOP6W1A7QP1TB1TRMW07lMGBcwjVm7eftM7tXO+3+STdNY0pjZ
DeADlPl1OltXbd6YhztPdtvTOEFTP/A1m1ppU7psAlgOpVj8BjMGOimQ60VRKn2v6Dtxy5YqLksg
vrQ1Sr+Rs1BFbTm7T4Nojeov70pnxsTQy3T9JUG0OLV0EslejXqrd8lIT3SiwrSmPXap5yOnivhB
m1DSYIp+hQK/FKk4BEpuwCpsm7TeldFOC11AdnuJfes4f54vOHuXuOPcFge8WRnr/vGBFwG4DvNw
+piV3S5iKL/AXfcxCpbMYFmVc/9XQNnn9i24uxM8dp8BGTU4/xCl+qnXlLLft0KRx657x8bZntOI
tFszEoXGKPD+mdW8IRejC00x4YZt8SLSiihzNPZKA6aB9NumwviYuRQkyXYkyhuSGaEBmeDncMYx
XX2PffKWkooRsDXDULTa9KL5MuT32U1NQFEho2Qy1und9JFTx52pKeRAfwLooaQDtu6VyUMXEg6m
BdBWGgC5gJy5Jn0ZkxjwehglVtB26F8RMJdJqB3kh3Yk89twYj6mMM/LG8BgpsrxL9BxoxvnPPB6
h19MM0h/e8INbEJjDnUhVuBAXGTi3MsExTgvqMozOQydOH/FAbuYbPKTVsEq7Bzo5Q8DtqqGuN8P
abVIGRWzIpeKTWdQiXgoeCoG3ITMfYgQq0e0QnphYKQzHAGfKEeDvkAjVaTAn7MHJyeMv8RPNsEa
FyG4hkkD+HNWC4I5Uy0bv64kye5VBF+kaRomxIqFTITU795RjRE0beYpKAmmW9LDfGAPHGurKsyX
Wi6b88MKgZLzmSS8Lyx3vFYL1m8zDAr5+fnekqDjmmjkR8WJXF8BT/eAcDlGayRza3dWGcSUwF2J
ieksKnJJeQ5TrbtTzkVwdANCqR8o/jO5IpYHhdfwaRjPkOoNdUOQa8oXUAcA8Lzb4Ni1AaEmTOLg
7yemlj604Qy8Q2VoJ6OkPZ/GCaudj+NzRKkR94uXWJMhLJHMD4nJEGKFsVG2aw4Rw2LASc5s6vgQ
VIygJDopzh6h81jcl3nZ7OupN0PmmHCwKi8eZXA5XXJjLV/GDVcLdaflaCZfY60rEZMqqewcGzZn
vv6D3SoEwB8Cu7zQ76cLkRZ4SVLRtCBabwbMy6yUzzE+9rgWnDofgqXMR2DUHkuJrXuLdGsLxN39
SjmmcHqAMR0Hup/625mKPf6p54qjbu1HUSxegwdq3Tn25TjCZdjLBN77UVkCU6vFYS6FTTrFY3dW
s7m8rUX4yaPpSScS79MW3trfu9s4c9oY6+i0fguP9FtG/pTlyukNVJYKRE3D+R2SfNN9pVg+LNN+
klGU1ntGTgDtsOM87+NX5K+lYcXDyEn5CZEgGuYHxAUzoMMisdxB8eUxBVf0PLPoK7Ll/3UCFSOT
GGsPZX3mmeF48c/IamS/raSuteAvkYstSEJKgWsCBikwexbp8seSz3dGpip89hbDzsA0OEyv0hap
MYHTCk5NgNxS62oDcL1fHU3vNiSTYHDDwuYZh5fWyzohM+v0mnn5YDTuGjLmn+gBm3792VjlpS5X
HLoZfmxnka1VHra9pBMqhHAUUkJ9hNHnCrVPSMdoS2wdSsg95BjeR4zgCxnz0N6jOPpmm7e5gWdA
MUYAtr/4CQWRnyOnFaZ8BtZ1e/NRnSSzns2RBBE1JP9LaV2Ed3+JdTRzAt+aQoKpwqsuFCtFvZqm
FzAV5mlioCy4PBm04SkQlYltmdFxqbA07dBLIgzZmHYtefS1uD6fNmHjBKsynEM8jA/M83swczdF
ghC/iaPF8dpt+Q3GO7wb9TQwjlDEs7n/j1S8Rmcvid326XUxyByVk+5M0qlAjMDXaiBvhfse/N6E
/ctXBksud/C15RmhYSRg1q1A61mFOC+nb4YAc/CYX31AiMpx8KvofIBiX5XkG5rZ7+NDBLz1/vWa
KSw3EaY6lRMTM6yT7TY9DL8g7oHINA67pjOpkFQhgHUpKvp41juH+TT8KyOCKZbb2QuTvdap3iOg
PGj6uDRVzhlNCV33xi3jguQFQ0ufAirtYDfNFC+TYGo5+yBk6nfy8mJ+EdcKeWi3MaxDejmepugE
sMnwfs5szuMKg0QLIQ8YMf4lMpROQ1isg2zx1j8EERJLdoo692ZWKGELqGcTXNw2NHr8THw4dP1O
k1Z+vXUU3dCnaY6t+IpaTKcKQdK0ULI8YUCeu/ES7ZTNVF7TX2n9Vpr3UFMlZyf/pHLW4jEmyoAz
CmjpoLMnGQcS2JTOvsECMznQaISqJJbvHWPNHSbnuxmuWxz/MgSverztbR0fXxHVdMt7+C3lVO/E
CQSDNy8lVFkRE07NSXZ/uZf/iBISLl7qjLkhY5avw9W3nIrs0HQffvD4bGXQtKEsvuXi38Y3Y4lz
fLn8mgafSC/Yx6svZ8j6A82bEpVaJ36X+77tH41aVb478sp9DgnVd0Nie+nMvVqUqkZxa/bdQfo9
AQFWdSQ9whvN+zfm+ulCEcQtjpI5yW2eCOO3jwbwYTahSSK2N29VIZrocsQJS5Fw3HB4PE2VnqKl
9HqNHUEPqCA7qDILm60nGo0AkblmWGqfSN9J8eJlMMjB/fiogL8RkxZX9QdAYEoXNe7BUAcd0wZp
GiPjZYqaEnkX0IhBpaNZUaXYmmQdoL0pgoXo8TAv5NGNa0LCmDKPgk2fisLVAKxUGXkMDcFUzKe/
cva6KO0vIR8wvwkabPHdutfzYylhcBIt+RSWbk65VDCdS8tUN59yiSPxcbaAlUumc9+pInjXWSk5
UeSa75rLVfp55fndb+LzPQcAD45SqcIY/tnLkB0BL7ESCSlVI5fzLEMYwz1U92zsARnFCJyu/Nhw
sXczFu0rL3GZ+aCrcV3ey8/hXO7agLIF1xI/z+xPLlvoMjJHDwpk6pKIJmIWJ0wGvItjJh8PUjEh
9/z1BcxQpzBL8su8XDAOWpNIkdlQJFxODR775eDWbEn0+7/Ifr4bqDGzM3iB/jkoIfPD3/2+/Wsj
2o0zD5o26PTjOmA1wKDw3rZejN16MLMx5Xzy2pxfQBWoVhTeaeiwi9CDxXx4DnpCKHQjz96gAZ2W
rl4dIbQ4COTXpMQbI+s92xCt4pJ/rX8SrFclCSaN8pGO8s4fO4Y2llslnLNrApSCLV3JImzR10Ju
oaEN9vEAAli2+XHPUwOojKQ+RUXvLr6c6oLiR3zNJlASZUSeb8J2JnSv1VZbpY9xu2tcjihH+0sv
+cId/9yti1JpkGCHht0AjkvEaAkrxaIQl7/eKyocxTJARdVFJrMbTG9xj1eeha88JfPmmf5+zOOj
QDuT9/rc+BUzJ5bZHrHzo2fK9CBfu8mkpGP7JtIiv0eCUKIYjmUkdVz3IVVfRFaPRzX9qfx7tFKG
jYND40zyqDR0xyZto4uGrTnyUgt5D1yob2ZrYSNoYSmEcb2IWrfZueuv8O73XOYomPH5ESPmudgS
ncaNLfaWmOYM1u2PjyA32pZ2f74D6mMoU200Ot6t9JCDmL1ON7lK9GkReUi/foYtkYjSkSneqACm
mIPy3jpaqrSjojwP38GMm2GCw7hxb2AfjVKZpk2d9zu7no/0r+HtKXbaLgj7VB5ueZNSVeYBbG9t
J88JU7fGT3Z2r2WuESF0TnaBaELhgYT48bwoUTQ9awR2K81JeOSY2k3AX+/s9d5SBtW4sAfOjoaV
q9moKNM5WPO/0Wv+qsV0EF7KtyjpYR476rS3T3nXBnaC2MYPCgpt8DrzB8cyQO7fnqCN4Z+wrH8A
BFWW/UyBwD/B98d76yL2zvJz2TI3eUGI5B002CS7TkNPTCmhzLrsdjKlXuhU9Qg5Pt/vQMi/hFtq
mf9dSsVRERpvqx8bwx/SsvNK49uYIf4lQljxXa1545nZdTvh3alBkr/I7QjuHQM1knYtUmD2XOHH
Ubp8tJQGhy8l+T37JGoVbzsY2a3f+dcZErujyYBqdyEZIB67Em8urRod7gmcDR1VeMlMbbUxMifk
g0qlE4VaV43JCTFz61cs5lW84WYoYA46FS56HlloV53//H8dt+Zx1rP8xNJWFmUBts5CD8z8AeNS
PmR/vZ0z1qz0VcvBZZlv7mqDCsv0XGlFdC4B9np9Y2gVNJMIu/HrYgHH68Iehq4nLbUZXm95ATFF
ac+H1lSuasfTWC91mxdBMUp6nJcH+X3Vt+kElvvdRdfQeFoyf0oagZfFiS8JhZIWeFiPp14P2ul4
Jqcy/UL0IPnvIlLToAqtSTSfzh/HAwGp8VZA+Etd/PsfDzhDlgjR7vYcXVUX786uDJa6cVdZIszO
lKTIlWZZgFC2OJxr/w3bJUKz6mJQDxtnYsEiu31IwA0P2x13ZjGQYlQq6HP6xFSKLwwr6ENZb6lk
m77wFQOgZyjQbhKOQH5rTqS+Ve5CDykfa7CF7An072fSi6TcMXDo6oHU9OhkrrTWlvpaQNu7OsT9
803f9PQtAkynA+swR8Ed6vGOaTlD+tCxGjlF4vB9hOhj1xMhyR4W2CogsP90PEIeG1kqxqqCLdkK
eBK05HzxWC7ui6DJrrcov9q5mbfuPaMR4ZnY14jijfdalvaSf9ytuZouTZ9NgKipOl/nHGXFZZVl
VwvQqMErsTHHfu3HpO3+eFexRhiUutxCQNm5p0+6tuqTZFf1azxSxQKLKvV1vgbGJtsChGHPsPsJ
uHtGwWBy3Fp49n8PneAxWcJlGPzwUD/V4DU1lA21IInTbcyRMa64L2jX22aCJdCY3zfq8KgpWcPg
mzJSjnpYh3FNgNPBtHUV5hCvrit6FjpnbMhPd4rOdpOh7YBf4L09uE16j9xuDWjYAel6iTOqPkcQ
FxCGPIlLrPTIVOWOchX6PjCDlg8SWWPKHa95WAqEoOUOSWV7iVA29VJJZfvv34r3V+Oq3J23Gw1d
HZ/xhYKl12dLSitfkUt0UluqTQqNEYGKwmAbLS7lmT7ridQBv8w21fksflGK0Qz2+VLUoaFwkEbF
LxuFpIl/+GWZwHTnCeGFIMMTVgzZtgFxF3ArFZCHkUfOkMbpGmngzUtAcDTp7rE6IgOqFup606aK
LJ6lIW90ubf4KcRJ1TfwwxrNBuWQyrW/9HtaXHLMZe0CgV6b8s2rJOSw9STCeBKC2IrYB5wB50Sx
fEsmQOCSdGrS9vKmNWotduNuWbxnUYpFU5MV1sG0MFJjuMKJRnUlLMBfhKfP+yXUAFmMN4QD+he3
g1dJWdkpORxyHiw0M1Vkh2FZ0qi87hgJ/Icnw4UjFqkkNk570Jb0Ioj7sQcFy3Ef2DFLGugoG/i6
6f09A/0+Z1bC+sN4EiiM2yuha2iK69Spafkjc64C+lo+MJ38R6PNZIAtaYtidmxFZylkWeqTGQ/e
GZnRddRHLl1rkXVQBKkPdi+CxsxkERUWG0e7XF8/YNo9ppkMt/KOPARqwbW4UpK8OHn05wPSNz6G
9W0vX8e+BeiGf1glY5oq+9trrb4qiJnVqltcUaHdZGbUsv8WP+iQpPmQcuHq4AWQr9WnniAEwOsN
dT3SwZVU/AVNruMq+XzCfa+G10UuTQgjFNqRkE0sQk9NlV0P+q/+EAC75YPVCJ4a995trSbdFopZ
L2AQcQt3mL1w/cz3DwgOudESbOAgI21V3JnsO8P20s6SLR/+UL918hjeiq72C+kyeqK1v/0Afyo+
N1lO4q0t+R7hWkj144Z5q4q+YXiPNZ6Iw1Os/ztepyiA5C7TtAsXePUuGhZppN2m0lbbdEBhMd6R
9FyJZCLrczfVxRWw1yNg9C+YTNvoyDVHD40kw9YO/46dLjVvbFQOFiKnvCeE+8F64zLR83iGlxcs
n9UvdycGWBmnIy7Z6ymq86sb6fUALdOv1+JU6hNrKPI13vbzWsw6GbZcLls8I85mgwfRE7ogx+Pa
KSo2Go7Qyd8zLFBBtrWtX4KyozPaD0s5fvFPUbSzf1qa5Czx0wupgXNJmQMfYmWKdrk2FzrfQ1Su
NDdokI4XwWKOc2tjrVBuwkHxcBu++rks0bQzB1U3JN+7dXcYAQ6iZ5r78ukZpSdRv/jv0VdYB1EK
b0oTAF0dX9UOLoUuJx+z05ZictjvnSVxGuCOdWnfDw4y+ARCjSBK6lhSyrWTLPNdX+zZvlWvRH00
BeYlkvk2SJ8ay8KmejPTfEHhbrxZxTYFnQWM/zA8UpCoEHkFzXUOxF2j6mZVpaT4Ng+BTRW9tp10
am+u1YdAl3i718d9P16Mf3MO7OI8xb6fVnQiyxZyyt8pUDjO0Y8rBpx0nR/yCh6RpHHthqN65vh/
HmCECYhyFOX7BjjF8yH0xz8DdNBR+aiCyUKfT9b/BS73ZJ3dad/QQz95sQsQSFcc7kEGy4Z3cY2h
DDDxa2Vu3KfmKuMIDsJ268O1vMsPrMzEDmMAWeGfy/HkChZ3KOktXkxDZ8Uz4/j1G+eVcgQvucDT
m5hXkA1AjC5s35wgyeLZT+PyPaZb1muSLm3u1j9LrtHltR6yX3Viy6ICnCsAR1Jbx/kNBTD5fV/P
1t5GvGYJiz4cfPrPkVmxNVTueyiIPFWBBOPwBc7sDpwCiLfRMDJlPB7g50O0AbNweGAlCgL2SSdl
1vtyOourtZywAX+ziF/J8q1nONLYPVl4I3usTmugfgD1hthlzUvUD0jfKL+Gl8wlXfRmJ7LpLPm2
S17xdUmIqKboTFf16/tW7GXEsuMGBfsJtc2X19rWiuTpc8EaOAKf3h4K4C18JnBe73m8bsPowUgF
uF7CRJ+syNksvPoihNLTL4WhKXLI/mFVagrp9IxCBaF4fQkbaufcUkq27VnKLwRPqr2ywzr2RMQ4
XLrDBVemqgX7yKpsS+oYVhPJVCGa7UB/MrRq0o9QEOFRqaLDpfCi8YIEOlBpRYg+mDn3WbzM2Nei
O8aXYWqygmNnMWoVgtqEcNSXWxe7WN7ROoznfLAfoAgcEQGpADxbaeitldByef5JOGCIGMmwa+nK
/bVnZo14QVXrwOBW1UQmvfsW3FS+6j+PBma7rkl4Jq6B+jwkmtABdZagpqFMGVQjZjAbX2A0zY4b
YEk0hIysKJeVAwm91f9PAdNpRfSuShv+1YMwIHq0G/YjzTYQtvzNjh9IbcCxqqsQSMdYh3oXidRy
vUB/PoHWAZwlvOyTAiHUJBJQFXka1MdEAmT5ODZQMJAbZLqfBnj4Z+FQSIDCCxwaq+qq0Emp2T8b
WO8e0rC8+nf/UloTSF10PiB9LhhtYIsw8Gx+uL0CWNxQwLtG5gtRGpSmQU5wo/ny+Gx4CtB081Lk
FpIMJwc7B83XaZYdkP1M3mtvQ+Mnexqe/qEn2rmITnTd1rfx+MhtA5ZC5nFcYTmoJVDXouj7WGwv
TTQ1EOh5OAJl//suBdJ9Wp4RFe8PBZs97Kq3PW/JPSVFd3SP4PDQ6F8GJjKPjmjBBTjPZbt58Lno
GoBQxCD60dm8G5B7zp+Bzkrq0JvGQo4y8IkVDs63UXahblpCDrEOkUExyVqNmjYD7CrI0JY8tt7l
y2r6DUO4CjOy3V5g0WU91f7FSHaeosJZQMcfBeUqxMVZYpUZOpG9hJ8mkAXGbUy145gHOUzCLkLi
dEcYJXBW9kL/D1Didltn1TpDOGPeDr3UUAwS7ZjEkItK00DY8LWnkpOtd9DTLczXd4OcYxk0WUjJ
FSECFOy1sH0H2eOKUZlNGuAgh5hyRSxrOXGc5inL70EYdhCzLJA7OGkOBwH02LikmX+/O+VZmTMu
BEvG7E8S7vGAaIYXC8WN5kVpmPbk3VekYx1/2KKMRgLvK48753J5FXOcMLRAUjBC1GFdztGX3hmr
io4RKqCRvPgnE1TAuFoLmdlIS/oEHg/vcVGMD7XkUH976n662Xrh5sVp7HeFJAhbgQ+UKvHl6VEz
minuGlLrdkJeJW5/gO6vexaW1WU1P9C+ZmsyDvZfq1ogzoCOT7pagXTPbqNNA4IpFHmf15phV4SD
/SZ9OGqKGlwz5qoviOXSZ/e4BJ4M93CNikjXpP55XOv2Ugl2UDLrpWaAuHDe8NkCXWtB6G79Jll6
ey4eHrwZNiIF1bpSQaHHEp4kAb4eyftoZLc6WOND6Trqw1XdzMGhIukbEmdXMF+uWuEKCSvdxpBP
cfVR8/MU9mS4z2U3jUre7WufeXM34X2taav1G25VyH9sWdoDEp552P4E7V9QTAW+2jplaGRV3uxn
7Ni2ud8zsIo9+KSFmkhJLIJzEUxdvmjWs8jDl/JbUkDFgb2wqY6bK0unBE/+W780xm2FvFTs7n/V
35F8GK0HgLzEvE/z3PzBEbS1sXZrupLrr4S8LpOv73C8GUK/zchQ2d+65ELBi4ozpO+pjoxYTpeV
W7HXNIv4C+Njonk2EVu19Z88NahMljvEYg9pB9B9slv3H9baZ/PO+ANXfsTpC0gVsNZiGPuRs17V
UExjkTMkcxDzLcW5JGGVqvdESULBeVBt6dGXWBAVPSVIBVk/lBmVq0S0nZFC6vXzfg+gKGdzZqY7
B+pLjvbuX4/N5TP7sgO4mIiKPq3VHX9RboVVlL4nJyTs5aUzl1zhd97WyACC0a1yx36GpTucKJs1
iGU0ao3eYA/aanFYD9sYhFLmimWVNYf4fzNk8TejCr1EncQImifNcAUNgSuRP2hvbMDBA91mbEK9
skmFO4eJFk1nWm1Qirsupp5X5Uvl2u0T6I8Pn+2ZwvK8ScmkheFwPTQrCKZzRKPul787RYIB2ap3
B9jOFf7pXI7EsdTnXL/NJRD0x6KOF7S8H1mr8yxyKoHp10WG5A6Uvb3drPXtxdKO/V+MtF+ypv2v
BWZWfcHVqaYKTjizLzdy//dgbk3C6nau9sCEgU/a69rAcwk9je1nTGRJe/aChwxhoqdMAvYnklUe
waIePAmOvu5wcz6SV9VE6SD96H/VO4LTvmXnp7O6xdbnHMTY7EzT7eZp2qOc9hOROP6Xx8KBJDW9
q5gYrepxHGGXUQKZgXaIl6a4apmuDdid4s+hC3aSVXIs8H+MhNRbMOsy+L5/RkTsIfwrSl9GZEsV
fiRRON5wTqDrBisj8Htlqan0RuiygoDIAoU1eh0/xP4c3ac6RvwRHMM9eta4Yz9x6grfOjlGJCIu
x+kLN3qtqgbvUavfNu6wmniD1fImp/dLf4MQrnopu8T5a30ANpM9LdQpTeYydi5COngCo8p61qdA
p3CkpZYZ5scdeGCj/DgDUBpbXyMVKMonDASkySKyxgSeyYkDJ4GI2k7ITfy+WMr1MsZ4YoZ/OPpK
IaCwqyH9H32xfb70Va1EMbCRAw2pIEkvOAG+yTBAJ4wfAqinymSMcW/2512H05JfsncO6y0klF2y
w9fIba6h4YZU8sXfJ2vI4kkbk+Rc6ZKxJbfpqgAGnDTMGHovyk2sqLLg4QF1k92RWZzUT1+mN7ot
T8oT/Tgu4GTw/ZlkuYui1+6SLJ7Z97+nHmhKE+5+b8fSPMRM3Grbc+pSUjTCrpCQ4wakzXE1ksPs
UYSKeWJ35QxmeGpFO8PrSv/160H5V80o5WSFKGACJjKl0ZAXcYEckq6wEwcpMT26lJAcEajT5b8n
08kTRNpbLsB7U9Gd7zyAQHF/jDV7dz6Xmcq0s1YAOfHBJCSgE5QuXkgzLgDFsz0X/C4fiuoKmtiK
Flu8uL/ESvd7zI2zMgsTElYE3rdBTt8HTMUlGtiCbBbYnhTUAL38w4wljBnrYsdPx7YMivs92EFT
NcW2CZwAAsWoLJYtMEERKZcveti+qdvl3KJwWoSfP88MBtppSWsDicBCRy9I30ABYE63+0+6CU+i
XgYumOVTYF5FYWnMIpUV6iWHzdk4PReZ5XlIIsB/lSzKuaDMnzVR+tsW1mZQe6KWHIDiw+77blkm
+HVh6IjMTVn1bO+EZEpnfyybhhuQBV1z4kZ/xQH3D/V1PVqZItEyMebSx0uzsv9ln49hxv9NodwQ
wsLpzUeivmAxRQaiFeqQp3vwjxZ9a7XizYlXU6QdKUr17BS+Id+HsMhrRht0/wYOeXW1rtCeWARt
bOq5NUS5wDG75GBbusb4dKJIgNqh6RlBgRPc2YlbYdicgH6LEbpU11wG+ejQb3m69eDV4nR9nGkt
wYhLTtGBdnd+z66m6ag8OL7XdYqHLXFN1SwunHwR9gi31vy/jqGiETuIU5eRCtwcYBo9NWl/z1+m
GvP7tjU95LpshXh1ma+mTAXNeKBmmByHY4WpacMPpB9ESUEiuaXlQb7rHpmakSuYdV2X20aruqnV
5skhLrt5uz8MlCpSeULt9pKQp/4nzoVkvvNobKmyCB0nrcJvft7yuirMIPEgt2ZS3wBIwRQ7kRCV
8+o1IqKIfLtfn49cWK+76axMl6iV4Qp8kp4MLEL2tl5xL/6jYotf6+ujMJuq2QkzPU3QItS0szj4
sHDFf6jtGbqUcv+mO0aNQudvrj+TTQ7vpoDEHcZAG7f1JbU7EwfgVgPgxjIDIXcYGY4VNF2AA4pb
KDcdY9sPuVawvjjl72EuRBZNrlcm6kZeH4nsB1YS918IfsnG4lXD5W+Gzem+/MlgjtUKpOgzRJKq
wrTv5X/NBQv9Ba7BXOAsaL1GAGWMJNrRL4NLpSjCoLULHrRMXlSPYWaYhT8gdMPixCFFZN7/KlZl
KN8u+c76CMLWU3vgSxZ4xef3bfc1BiEN9IkktjJSvRGkHUyE52zm3GdiWoakfqC32QryX6UBCETw
esU9VIfJuGMqihwjQ9IakVgAUfvrD/9VONNJ6J/8VV1AuRjmx+DNKd2QJ6ytjweJusi7GevKZFei
Fo09HLomaEjd1QbkXwr3kAGgbgdQFSVGy73l9NRcbBmvGs8elPXn26k9GToEhaM3hTwm03MNEqk3
WiEt9KueFeUtHrqUKiBfRblh4x7zCJwhSxZVEXLMGRCL+ptab6juA1sVHpxJP5RbAuCIXYg2Eetr
yhBU2Z/2nZsWt3gO5Bs3xu0D/kgzOg4CUML4ZP17UoHE/2dpHC1uEpy4DppBDRxIPPeiOhzcjAH+
KA7tl90dROSH5mvZ/XJ/eCixb95IluwONo0W4jc2cf/4ed41s/jNzWXF6mXjzW3CKVB3mhvZUjI2
KfVAKY0nLger+0uA1gv9BahVsBfoeaC9Jcfxz+OU7/nUftLVRISF5HtduATp+U0BlVzKVPyZYv1A
A2EIKrXFdX1+i819AK6/QX5gGQHnwCVobMcTvTqeUTa8ihDStM3sMTUq5nCQ7qycgl5HD8pc27oh
Vt4A5NqsBhQLMRl+R5dF6EBURYKiSwnYsy+qt4yFNbfwV/Qt+YLJuf9KgbAYDolsB/dnyyjVsp31
uWosFuAdHjJVncYrKePJA+vsKiBJV8HPBaGT2M72GoZ5WHDKbS+OzdMq5b6tHZG1NRY2++TTymBE
yEV/BvwCEELZRieazcspkwzjf5eq9I99EFClK5ELWN5834pEOZyusOc2UhDJFeE6Al/cNyr+/bEh
Uz8N/OMlly3GB/H2AAgLoNfyoHfCoWiH0rDBvrY0NjKJ1pPFQ3edAVjw77IGtwBsfjvGkwSXUuvQ
hYZWdRirIM+hYzvUycMIfeONPyemj/VwdhL4HpabY9XG9L37P6NxTHXHKyMogVLtPVJjN8Xfz7Sh
Hqz0wOEqyaJcVIgeoH/MuY4qQhuFofi1KNM7MWSs8gY4iz0d5IzFJWvzh6Irv/TSoZ9aH/pr2JqN
PSQG9HhcGs59enpMq2mFJzB7iJjT0SynricbeMWO/MrdaKp6A2RIj13XA/2lVmy0LZvV3O4LHa+Y
K5kW5V6QdkIHvGPDf0n5YwcUkjw9jAlyGWr2xuLV0ddI0QtjDRsUIBJg1Yy+i6CXtx9cFeLr7p5l
pDRqwuRHAj613oukKvC1iwB1Qssyd3Y0D//axvOl7QfeniYOulLAEit0+kbwYASXJBbLig2BB1WC
0n1X0pdxLll1EzPUAjSvruKs3ZVhK4AXLMXt7dMwO73M0xZjCZ6UlrTIsA56wbeSSzyLuuSP43yt
WYE2EMi521ZXRUTgtA7uhJiFh3YESf4HhLedeBCfkeYhi5xe9Vx9Hfo0hgzOT0okwuMatMfkA+rv
xjXX8hatZE0EWYHQcP/6pYA3ljeVTT6O/SWF3sotTyk7c79kiCGwRB7IOz7OPhs2ujzLGXYchKrI
/LWfzDLB+vmzFjkGlONv5bh/jVIdz9dkejjRTNTA3Hd9E7wKN2gAWCubw+iPLZObbaJbcWT3bM3K
RsqKgDAKVAfnDr/Kgk2OlSh/kHC/EbswQq7riqNvEd1Hc2rSqU8+rtzpNFsz3riOXNHla1c+F0K6
cy4tuYg/40r3Ksn6+VkGszksIWasPtQxyY6bHCUg5F5CoPLXjypdfSA/sF/gm5Gqo1VRuK93GJIS
/V19WuyzHcVI22rfo0Q794aKfeYfI5DU4+NV49UxObvKOGIWBqGUYG7hKosHgEVEoCcbLIE5G2av
IYH/r7N2BKSRNoo8yuH6oiBZ0De4TG479Q3aC5rh9V0zpVzGcvJVNTh+M9jZfpzzUB5me8xXYe/O
VkW7crA/0xohxndPBHZnO3QpNx1j7QWI9eZo2hjai29hp7IRdbU+cNR9ERSL0T+mWbor63oYPqmN
dzJ6HpJdgiNekif3vDevuRUeKRzGnee8vmtxiObsdtkWgd2Lgi8jNlMT6CVA7/0TQK+tM88lNcap
e4cfaNp93CCRbt+K2MAEf7EIo5PsMxp13AqEX95rGw6juwos5X4Hyj4gKS1luny66brLmv8ULwBZ
Dxz16fyoRxwTs+C1zvFvh36q8r/bmUf8DIcMC61nHol++AMitqCco/OBhTqczfQlwoEAOw2Mmdh4
QccIQtRT/u0wQvLvrJMUHSS3MLTsz9/PNBCmYzjODi4ax7v29iNAo7yfNEKhx0PKE88ycbM3BAxE
KVAncnBKQYRa64kqRAzuH6Dx4Mx4xipXRcxmJ43Gx5/7Kho7yVUEF3SD5Qw3G2CmqxbKqdwmfoyC
C4omY0fYwQ9rQ0Q37G6Tn29oleLNWNa/JXUA1EQnbSmfqTvscZeWLxURN/7SJ0n6a+cznDxxycqc
EMp8pP26Zr/CG7bd8bwDQMlTKlcsr/Mlq2ToNaG6Jp/foohIeJ+xtDoieSOMwQHkgtt2Wu+yOOlL
aafzT7N50ev95zh+GWFbpaGrs0oYu/e4sqdzuPao7Dz2/ee/2Jj8HdmrA2YyjBWyzroS4r+PaulF
iXNLw4R6//AaWDunJMYU5WMrobBh4vFxJrDZQpJleKH+ZsY0WJ1bQ/GuKX9kLrJNi34LK9mCoyHF
oPL5Tg+Ih/SkPNaT6hMTXdmupTLln0NFPXNDQv5lYkxrLQowKuGH9s6/gIIKLxRNCcKvuC7c7DI2
A/LJsHa35S5OXPazDtfFpUi3hveWh/lVYapw+oHElKDhWGqb/tsP2dgvwezuMoHSIvD7+64FYfrN
AJNhpigSQ99qRFIbz4VOtAj6zRWiBdmmrruxlOaQuwQHTNGBMN75KppSDvkFHYDcDUxHR8aRPGAY
aTplsSCuL3glK0g+LLIv9lRwzhx1WaGYTF29RngW3RjNTBNa0Mtyp9JpD9HpxAgtAAUqsHuiW+mO
4NRqqFk9LaPk/1c/DYbSFnS/UQ4l9NiReJ1jDQUB6tUl2tSlalNT68DzDG0mbnLk9bcoLLaVnLuP
S9R+hcTxfy+egQFpY6L6wofhLDbrh45SZK2UU1ik+9EYBMbDgjTyhCsdA/e4LcUjuAv8jyEjD4u+
pJX3YsDUK1xaKOF2aOiv7Wo9LskMp5wbPNeJS6E0KyXsWNzxD131hhIRe8QtmVZfixRBlV9rRGrW
/Jb7neUmXWM1XZ23+N2RDKW89Qw/9SC7r7jMZ54Wotzk0Dv+d8eCa3uYRw2jzddvYPKatPInAZxb
sK+JKNQ12ERi/Dhy50rXqBS27JMS9zwHlK7ApOvEvOT0zywKGBrJ1/hJrsa9uUJvcMuE/SrKt5Wh
AGYNzJMypqpCYH2jLfWYshikID35LZfe6/znyaoYN2ZF6BhNJItxecyGyhEizUj8sNxHOOk9FF05
mNA8A2caM8MB1NcREFvvVWnEoa4iDHBxD/xB6avd5K4U8Ca2rI0sdXts8Dyz61Nv5bHgt2oqLpnZ
epdhpP6aXVyQFvgBg8dtat4G2z3Bf0h3qAyoSKxOQA0Heas5zfDmFUh7P4f2cVDKaekW/flk1cwr
EKlIL93Bf7XH1dRsnZbiOJCmcz50e6w0RmW4p7EbnbBBp8QoDOu++IaDpePowi8vzP95n4+Z6iHx
TbnTA6UBjXqMX611pU2JhU8JeIdwjQtn459aZpw8rnnCzLtZ3XxSQI6gtxB5xDmEsyNBGihAD+E0
2sbPevWv84eN7cGFz1M9QbyLdx+glPiiKKcIFSjIX3rZuZpszzbfqXLCxn+fgp6eQodPQDvubb5k
hWdyBlvh6Eqs10TvnMOoADYbqP62BGAhGg5MYrGu5bJLFpI9UgwO3NfFYsBo3NslfNQTB2jP8VUV
4EKBCiS8pkP1Chv19ppqZwg2R1cBhiPmq3hGuoxG9ZyX4ucmOT0vYYx/x3ijWeZv0l7JRBrxXGsg
keInnISS9j4nO5EU7H/87ct1jbPOnEIEMmxw0XPt6X2UYoQHFoa85roSe4bHHzJQU4Og/p1Kv5Ja
FUbb70MkeuDAildy5DTtZOW0VuPAX1icGIT8BCZrle1Zm0npsr9Kkrc+sUx5+MFkadvKbpnRB+Sl
/L532HU2OTLs7kwHamC9CGZRlOLfHDPU2eIuo75HEvBo3/Kr7rypf+R4MEZW5MsCLcRE0xA2vr/1
fLZgkkLWAkK1bKp2DcuyZYyPrBEuJE0jCWUXHsOViCVV0O4NzT9ntsX5y0AwgsCttnV210s7B/SK
U37VSNezn5BCTKID+Dh/Zt4FtHJTKiph4XQ2m82mes9rxW4CWA+YtG9n+Q6+e/4xAJIo5EJ7NtCq
qcx83zXHu54yM63pJi7t1O9O0ZQeNAE7SjD0WhWPfF8aQfwR8cs6syApiPgFx4bBzz0iaUdG6ihW
WdBWJ2SPGMPGHFlGNS2pr87wVxslzhm/MZqdPtgkYZAx65zH4EjQ5jjBgD7/1LXE6wNQNlKl3Uq5
cBlsCDDsxx3gC+u/frM0/HE/np5b5eVbfQ61LNhuJtx4opcj2cbKAne3mGHa8ayG6mhj/nSgayNI
GxuNd+oq3ilw8+Dm/E0cRseEbzKY9zFym5ds2Hc/TxHMVHaseRWOrR8lVQiswWfd6uytPkxIM7hg
WmPtLNgrkP7JpFraRU6Oe3Hcsrm3Uc2fJoxscj0HfpAwb1uKBhN4k6msVOHDW0B+LjHA9pTC4cms
In8pgCDvPfUXMY/ryOl6Rxc6rD2xz8NdqifKfEterkyEkVRTnRvGJ2MVNkrhC/jghH6UZNInpXsc
/jMhMy7TvFv+fEDA3p+ZBg/o2osYxGPHJHBixQR0wmvi308EffZlBDch+9tChhXFL7z4rfeKlnCo
0AoaOmYZSPzkNg5dldZYGTzEgDO+dmw8KCTdMz0081Tm68ZI79mYXUAn7hmTJoKb8psyF72IgsPO
HUkdIiPGIGGt+xFTyYlmmFXa1LXFoQTEZc+lMtOvX7bMFiqHqjJEl9egGB+jXdxhaf9/j8B8Rt/a
p53bM6ddjeeui8MW/MUNHjiNKnSqme7hPEvqHDQsTw6hWytlIxNH93KnuL40rZIE8Bb2rCTgLJZN
IT54VBT2hAbn0K1tUk7CFYntgXUCI787++R4Y7YoSKbgS3NFy/H1FJ/s6gX66ccBpeAgou1S+WxE
wCf0FizSODM70sEGyBp9FxWF9h/W8GssnUSceQu066iFtM4tPJaVaTKaMeA1U3pKG4PTWFkddjfH
wcRYm2BVOF8dCyHWyS8R9XIDlefeFzUMsY5JnEaN7e1PLAzEnA3eZymZptTr54b2mcNfrhZy2tun
XCzi97x2yZgdiTF6+VLvPBWkz7u6h9b+RS2/6K+7hNQFut9LGvDE1npq2HPT9QoJ7+b7Z1cn43mx
Eani9tUD0cdf9PjAyc0Dy3KvFpbC0DuYGu0mn1+zd/jZ6B+6MthDataZLU5jd4FMZSE5/37aqS1J
90EgLBxnkAt8NB/MdpPrPJ5iEuPWHB+SuPkWpiUA2DDdcoJ9XnnFAzLrPpSBx+Bdf9hi2xlnbwWa
x2aT3zP66Ppg1OIJuhZGx1bb1/OCR9rpfXaJZtALa4LjBbDq8dX/GkYV4UXu3BIGysVArfH1rQHg
/29yi5tpwMz6emkLP4qnqUd5y7X/0PE+uDp3Yug/qMRKfmviRHG06gttgzw07E89BwGdRzAGj9Wn
Y81OZontIaWtA52tRx5X2fsSQtTKV3XnJgi8qX/zq+q7Rr9roqP6icwAwxaUVdF1CfeqYPL+PHbA
QuDlpJ1ItwCzJe0x7O0Y5KT5ir1N+p566n+CxnnI0Si3KZMtqC+IImxE6ZvQEunY9xftWwXjqpYs
eTwe6V2HIVoUJH958BsMd8SBFXuCdDlHFqqmiLYnay5GZCmY4HJTZqh2qNz3MeMVGM13FqHcw79w
8GsjdYsnjnXOH7gOu7+2yFQ1F/gw9Gtoq3y8lBwBfH2T+g9WfRid1gFgA5fK+bAatQ16XwxsaVmD
YDGN2ghcN5ffrn37NSwnOoDegT5g3UDuYV7k59kZ/23w8OJqoam2/qqNc3q4iy8O1xG4/p7HzIsL
0dUY2fM2tnjM4xPrrTRgdV4oTI7eM9j63NPwn1r3Jomt9EzDHv8bPVGdo6dCW7giUyYRSkMM+y7K
wvK8t2A4itF0HjAuicecfPVNEzRXaYIPwcEBtQs/9+KJawtsaoWYBnNhA67MVf6QS169rgZgWm6Z
rfQzE1Cd6z15otiOjMUIwd3LLldtDpr905pGQPGeuTTaH22vOxCzysKTrnhfuMhAOwP7nEZUOzLo
TgOjgcXO3QOVMGjd/kdw67ymGXeg7FeStf7UejXVvIQlVRr6Owuj4hq8ONZtOzO6OcpnKjmb2HL8
3SJa7Y/Dlqv/SgtgryIPbumu3W3lW85/gyu5UodWTK9lTv+ts2t6F3mwEIpeyYoGYYYW3InokCYe
ARA0kZGQ5j0Je+nnt6woYq+ceFZKOrRLDIZUDe9gIFFJCRPu9HZmEbQvo0ZsSzrXAfpXUsP+CXoD
3BQIUI0LQmIMIq20AnRKXwTYn3Dx8MOsCtBaZkVR6DjlcKq0VARHi86HN3e6hS3RMdqETA6sAg9Y
XqLqptWyTGyMowGgVcHmwThU/v5MOkLCVj1f48lqPv9Pret3QR3iJiDXJ4E/qH2YDQLCC9IneLv1
87jhGeiz4ZXWLbc8VzZtJ7BEoAu5EbQLD+HA8Zif6BGLy0p3BzzqdIC8ML0/njr9bCJGykl6wPhL
qgD0Z+acD6qrS0Kh8bg+DKd3gUSu/3oBe1Ow8pTNqnI4sCosPKXBhVzv05T0MOvaRwvwOHX+vV0t
+jsLhSZdPUQQwMbiiqLSTy4mXNeGxw+H23yJNUkHYltvnNnOKzp+feLCYOWVW2GyA9QXDm65C4gO
Tn0tuKX4CSJnAors49dGVjkIYjrc9XW3UMvlvmij4xmgNToLofI2/Pn2kuD0GGk2v5pDMDTL8kSu
VbaQ2OU4goqmT5q8sZegJF2KvcwHVbOUybVXc3fIAy13/v6I94zgD4VPfO39tftgTrnfJOqTj8xu
T/3BHtvEC+6aWxadfL1IbXy8LlNfmTsLoLw9WMs/Y+KVuzHZ5woFof0aArjbaRCr2BtCNATkeewh
/zulHG13gA395dcSaz6k3Eq23QJvke552H+VrsrFYMLtUCbguNdeZDPQRLRVCuMU/FjO9YCslg83
VJgUKl7xm2oMdKdOfPrvgOYMAVMdxOskAHRMCk8bzJEoaYsJVTjUa9LrrKH8VsIN/lyGzKOEQyPy
fyBZi+OLFeqfc/CRW1zegxY8j93JsLaARZapGKQc8bUahG1F1s95Das2LXW1TIq0trJMg7Rz0FGp
eP995MJQgz0Wbjtzg0RfrLiA9Yyn0s5IharfwzfDxHstRvYeKd9YqtIlLr9CudP0NHFn7AOAikeW
HvEqBnetC0I8vRBSeV1LTA21wzYLcfhRzu0xY143ZJ4y/V/hzpwP4kRM18usZWE8dll695kTsydT
foDv+/4W/MQ04NJnpQ4LupRYdtqMUmfnSvq+Uy6rGNwaAxZSyjFzgRtAZQPPg8G5wVwo5H4RXoD/
49+dJ0cAP2XWJ8B4vE4Bx72scwDv51K6mHUhXpMpnOefsiyuHDL3l/se+K9Oz+1C8rBp1gdGF7QT
RTXhSoC8XNir+yJRS7ULoc6VnvuEoRghsPmIFQkzzpKG042D8lyf8hr3JD7lEQgd7BU2LFOsH5md
hTQbhQY4WyYnWrGZ+vgR6I9UglBUj3wkucDVD9v4DsEOcewYgEBptC/ybGucGKjEz3mlHtPo07GP
OR+QfXGpT8SU47CmrG6r+sryLl+Si1o41d507vI/l5UxWPhLrP/pdfwJgTIeqAApqSsGfWRVp5Xv
w0VOgT0UZF/fHTU5VbtqdknVO2KTvtJro4kcnzH2Y0s3G9k5RGWrF1TIjyuqWRDAvB79HVJAQGc9
Pld/c1TCfIRn2E3P7DHtow/8hc9JrfXADK+0gMqomC/q6Wco/aYZVArPBpjLI9GFxJaQ8o0SqNCT
E+DCuzRQvwqkQGkITSor4cFtH1Fp1uMTS1KWLf8GDdnp1hALItmtcRCgnKJP7PN2vPbxL4xP34V3
dEroYNPFreHXiWSOvNCy5zUJhPkSJqjcAi4bQ3YYwr/YePJEq6HrOMSzkKe6w3pyJwMqVZhy2khW
JAkQXZXdhWvRD8et/hpUx849uRb0OpKBX6TjvX4pfHdTUpbbWSHYIBoSe/Acf+S+J6mClBUWWkqh
MxCAcqENFgE82JIQ6hm+gg+pSo5WbZesFKxvk8SwHwODCv4MWgXaPZVAZ5wzUZcuVf/oaFVB0ITG
/QrGWmtSru+uuNsXThRYjboVBwE89Nxvu+mRTDHCzPWGcpqlrjlLhygLowGmcjliRyqF3RzwTdII
3s1Eproc4bQtVk7QycD1nQyRq897IEOIXZ7Hcj/45WcILzAdaKLiTDD63uZV1KQ5K3dpK7UY4lx7
RJmjrgUxWFPxveY5+LqMfdwr/g9wpnAuqK/kTXkpmKwKLZAr+GJ3+dHuy0YTqrTpPnX5Yi9/nJzv
VdxkXj+SwGGVibLB4mi4jFyklCl8fq+mwXf2AWb1iFX3wfh9MZjFv4jf5IEqLD7Q7cuDBHnNvImK
amVUxxtYLMbXgHaD5YBLTNUUwzuPu7TPZIh3DlxsHcEftiVGeHiKMfxCuDCuXoBrLS3pc7pv+oEL
TtDfq0qGHm22WP3a9Xzg/WzKVDSafqL/pBmUV4GdzVlodfRfqR+pUK6RvOHYhkNxu9XZBra/S9yN
tch4Opbn++tybn3iUg32gc5fhCHgSaUQJsUSxx451tVNd39ELVWlBceOMX3mWLCKOMDHmXSzGheL
LMw5m8SHclEmxcQdox8ZJ32ZTLVap12CqnqK3ERNFGh6sw9OtouICashlQPo4IGouNsvorQjRjdm
3DprVZi6kd5/TYWQawqDUE3ITx3Xn7HrxksO74TAcfOEwFi/TehGvhWqxFczEuQqz6ZkmVpk9cYY
a3+u31JKx0B5XTgTXVUH9fYNvTj3UCySQHeMtByNvq64k1sqDpNVPOquq97SMOOOFJFG/3NKSX6m
HQPQ7DyynCTKTYCPHeGsX7E1X18tThYufazVGYop+0p9kgB9x8a7BFBORuAYphA3cxZNgffu8YyW
uWT2uV6D5KiT3ASbLZhnHgPgsAx9ovN6JZyAPP/w1hX2DX4n6scfLbmXpnP/C0DP5jgwD7k/J76O
jG36LrZzGfXjlN1D7ilvZP6wIfGawLYPoDW0CgrzHYL04pgQ2DTHG24u5uqhnmZ7yUCRVyLWZWMQ
dcoY2eWCpO/JLjqVIzBNwYYFYEMamJM4Cq/z/H44MqB06Y1I7rchpIZYa+CF6VS82gwc9fPeRHYi
C743hnA+dwTb6Ri1hrAmwPq6lGLOgOb+rVNYdpVBSxkQ5owacEb3NRa9/l2r4dus/xRTcF07YpDK
T0pLLHrHAx0lMIdCPt3/jUiLp5uJrS/L+0C6DwU5AaWEgCSkp7mJFUC8L5L5Cs9DkEwkbIY+Rvi2
smCF/8rDKkGrmmgMHmsyRt0YwF974kKfoWOoLdAFi0DH7WCX1K10kxh0U4gwvN7H19K/SX+mMPGH
3XmGuNzlEcSDffS6XbrYxgJOeuXxNPdQIpufZ1Jhc1stq+n5lfqkwtdsrhLWB6FyZZU0yuKr/DNj
dyoGQpbXFW9KWmZ80kCb6anaWmFp4P5AMOZpO5SIx7QlkSRdxHh2LRGr/+mM1LHc5/0YusL2oU3p
cW929Xjb+4RNw1bHWPB5dnyNEaPQdYCN+oiCWjT6bholQtPVeYr+c0jIPz3x5LFZx1oVHQqgDg7b
MGIUcOKP6tVa4L3JjYTSh02RDbT1wQjrnkf4QOhsaIhgQAMQ15zNOKVzOn5a+MQZEyOSI014u3nS
gK0TeR6ca23I3z4tnVBByJra55oe5YX+xyY7Fh9AS8HbMqf1TUdAHJ7IK8gVrkbpU6jA4Impn6fH
4SB04AJymvf5qq3iWGXLmuLzoKjdgcHeestRAWx82etP8UQGggCOnnq0qllKyuciM2hsN/rQgPnP
LqgXtuwlSxOSH0oBGDDPv2/ahdoXVaKZqenrzBD/wgohjQGZ/RqR757TW4IFZaL6yiDpZPwQ/aJ4
X0u3vpT+0dsgNaZPH1PJlXOfAJn+h5MPPkzivvwrmKl+GN2a78VgdBaG6gvuoltOz8ZnX3hZblQe
xkQ2C2xwebJPlHv3e2BDHxJZvOyfDqgcLI59eNhLt8x5tCrsaQVz5fti1M7prtFWHz4+tg67GY0N
61BNYrBMxKCvV/IubSgB50Wzfe8nq2yMMMRo1UncfDR2+FKjsm/9ir2v0yjLURP8Fb7DPWi0AOde
AbuT7XTiBzTCaHDdVLujQLTWWe+M7gmJjmGSqLsoS00zDThrS+jQFCcFLBUCb6eU0SSj1eswCD4r
7g/OCwodOuBP1b6Z0sOPZSt3IXiy3ZwF2tudQWc/kt6ppOVf4pT9UHRu+s3BgbUDCqsmW5bMHml8
SzED+2Fxy89wuk82zyQaVJZDN7x21tWhpkq1baX12kM81cJVp9WKaWg55V/h2fRsDD9GyoRc1OxZ
o7yQ2zmrzKWqlChMg/3Q4gLTbuMbv6ZJUhY75USkRGH7q8k3jWU1FPJMYQsUmjfAXnNZ1j+OSrw2
dxVZb8TdkO5pBdDlWlvVpITxAO/1GzctkP2SjepxOZoqjLDWDeeURb2ANKzSiK2NyZZXmmEBjZHn
jf2aBXWY86BSpZ7mYCWUCnFt4LemNMXOR4L5xd9Ae2OoCs1SGweNUHIuyB0RYC+zxsjLfeClWwSt
hY0emvd60nw9JYFxr68l+0VevGfopQShDZZYpDqbEEIYqPo41aychBT6zG/1LYvU57Z13F42GxCx
fx3PS2gjz7mJ7rL6dxUvisFlHcUq7dpJ1rKL4UrjxaEf2bTaC1U1WBHLxcDPQsRtgrQc6B50sEGZ
j/IByriEDPOF6Lk8n5jBs3RAeKNTBjUKZ5s+fdIHY4a2ilMDW4YnmRgDMhQCmMNhpSQC/eQbSD2Q
tukd3YGpBhJZdDxgIAPPM1lJ+ZzTsKRBJ5SGA4kIYDNk0EZuCj9+u03CPuqggy1QL7VeiCCKdZN/
Vis0+Tw3v2kKHz5t5nCaHyoLic97UgwPubAEBPQITT+JVrwGa0wp93r0FEcYZktEHTZdd/tyZrk9
ksWaWf+AMlT1DrPMdFrx/nSN+4gIjdjyHRMtpH1StUGs1e5t30P9owcg/buQs0knRjeJvujbngxB
X2JsPw8O9qv3tkgMU70ppMXWhWdKkvuw8uNQskJVlkhginEJEpGB7bqECxYUVwvRFQR4MZxZwNZb
U8G5JQQobqT642yAmxlU2fWwE6egBYQb67lEg4yiM9muVtifO7aj+dEY1juzVjjueYf9KL1ucU76
tEKU7Us0XP9GBwaY+Za/LIIiMrvRv8idNfin53x+qq7M+6V77sdL1z2g1YqwYfy06o1BAbSly80+
Ns3lbSGCiJFh3UTlK1fP0ZrEvIObVjkAEPngg57pP3KOTlBk0w0qTcELVRKptN+6qHKuKBqi9DyA
Dkp4Y+tACOx1mP5FWKCo5RNs/LbZ8vvnzwW1kw1wVAZrXn1SxN6PU0iKYhVn93qP2dUwqAX2aSR7
UjwNqQVD+0E20tWOFMoy6owT/ujhcd+StxlJn0L4yskGh77Q5R/BSGtFs3chfuLOSM0buasWEjIe
6BJ5heLmSHS0kdEFcSaDhTNId1jmFHM++3dLdw9xUHbiefGhf2AFqBcRhL95mCqv5DdUfX7fGTjT
xhMaBH0Wm+9eYEEbLkyxKrGO1wiXEB1Ywv0QHZk1TtjN7leurGS/Du9FPR6BFRTwGF9RR4K4QCmM
5OMg4nQZHLPCXk8ShXAnEsonjbyAsw1AQ1EtoIbPZ/poB1yieTCOGLhdcpM9J/T9FLNeYmrJs8rg
JzRXClJaIE3YGf9dS+DQ/R9DS2OvzXlOvuIT7Req35HqJfWkqoABMhub9SFOU2MlEE3MuPB1GIan
LoYLCrpnilxsL0dqmWSIdafFna9zvzN07MW66zJx9Kn3Dbwpu9DlGegLNIPPgExpUifripkUuqKz
CLmQpzzM80JRidkyCG7t0aS5PCQVAGR42cGAIpF83C3qVsC4R920DATjmauALwQybchWSUIOZdBR
LU5ztrBaMYezq2A8K5KDmluR+xG7WCQmD52seY2r+jHWUsxr/qZ6EFFJVVW+jtFyV21wzuDeRE98
nYkHToWBHfb793veEXFFIkFiFNHXPTJb1R3k7f7skvxbZvZS046pzLeF2Rt26ypDqn4uhiSAq/kt
l2ZaIstq81y5huRKT11XxWNGgm55A66CjAXR2oKBx//NemZZiVNSukzgDr2g1SJx2yydSXKOTv4n
WAs7bdtLfG2t3LYYFTw2/raRAHNG+2H36xWmBYuGcV/Zuw0BZAfUQpYdPWjwrZiiLCao4465LwvU
Aj+o/euX4nDORuA2ffJiSk5pIf9usTODS+YohoWokT1Ax4I/5/YqihQ8wKMKQTWFdAWjbhrH1Y9e
N1fpi0VJkWg3hlynOixS2mbJJCvsQNaP15xc3kYqGvWcS67qL9iRBrq6Y0HeZ78j9I4fy3aov3VC
vHDT3c2GUYJdxNaTKCTc+tHQBoe1dA8+OtoTLZcN8NkCDUgYaVIN37S0Nhol2g8dT0/ckvpFHU2f
MfaDTDpPNsRngjnfvdz19PtBxXJZNGfUw9NxF+zd0w70/fEdJcc43zc6d2hhCVqsqSkYyhmSor33
KiKZXA+Im0iHoGflXbGzeSnIdpn8PWBfakShp/IoXrPSpzz1UWtyAfFuIYO7FxKj2uf6Tv9uULx5
tsRYwA3LQd9Kt6V6XT+iSDqFdio224FQHvgewrroFFXD1VyCMLlBuQ+PUZRYYSaon6bEDZRsEpmM
4CQNd7XVWY0hC8rb+eBkgyGJ7YCBLiB9PcQsrTOX382IZio2uPX3vYw1SsV8LA7OksKUUwOSD70p
YbLMVX7+Ptmm8zBdTK/+7NT+hN29xQNSkNXNH5O597PXHhC/AMOvHeJMC0zjRgEKBFoHmXtkojly
NkgfoBvaHYGp28lYvuaLs3M1HjgdueAEkoF2uc1iYcAZCnTfGcUPv+Eatnf1amkSCRs6S4gS25tr
TYF4w+uY9jXFBWod0bAbMrmHrXa8CclNXfKVopq1j8ZtQLiDrosRlcZqlYchWi9wedBH9Xg2kD5f
T5wZ2f7OPgjIK8Dnu0eLgzQWj/kh6TAafJWZHVjr1xr8fQZST+5f3OypksDIZzW2Kezf4kMqvbFs
WXs3FYui+M3RvzuUKbjvo23y7kM69Avp6cV5+r2QFzfImW0GLvGigaVihGMqBOIRNUQCg3CVJLUM
BOi8VRaWqZPaMXWr+wFniM393CGBhELcOnjNPwbnxOQr+ny50Z44NCHXhl7lhoFgNFFaPCOIcTKP
ltee3b8TQRvPydER+0ZLzFE2RHF+OchjdmKMX9qSc3VraZ827kk+cu8miHO+T1sg72UetBMRgQN2
Zs6DSVr2oC3c896dwlAA21aDBsY5Ik7V50E7GrV5eBFcuKcaKj8rc/E66benxz/dCX5GNtOzP6OQ
WgvdYLeWsDujETcXdVNlWQYKXQCguXM4xuDCxBtvnwY3oX1Hi2S0pEaQJN3xvLzSZGfEgI3XoFQM
UwPAqJDaxNECKhQH7TWR2dX1Mx0uIuAi0eKlsCa+VtEM4eWl4q1LAW34uoeDNF028M+1TQQXCE6w
p5eo5kifGv9R/WQdaG5CwQmQN5RmrSXuiiUMLP0rBnNuGbvk5HsqEKP1Vz0ZDXhb3lximtIzmW/I
CHItqMwGUSHapCPsAgU5SXmP9m1POf9mKg7JIGQLsI4jboNMESmAosBfC6eOwa+xueKG4Wsh+q02
6bXdkbgXAaFX4FtdCKSwEc2ISoSuTXdS2jYyp9dDwsd5GZEhmRE2oyG4y9CV3UKpzDrulHDt9rK2
nfsS/pMc++bibU9JxWBa0yFT3xsJvRteX6GaltdaTHzywnK3prBH1tytO+stdOFh06Ge1SgzVNsf
hdZoazSGt4sU4DQLwAgPhYrqhIi3Mw1sZI3GnwGvK9UkHE1/IXk7xPmFzfKQ4l8+Xi+oAj7qLl4B
SNVdgko/979pOEzrX355oUjquhuS4bUVlGXoezZHNWIJmWfwAAqRAVZhE+aLzdVd/f4yschInqTa
X+UgmBk1HEcoC/I18lKkDP4ENYe0YOD8maMWIivHKXM2f1J/yU6aRxE7dUNAZy6J7DOLg6AHUXbj
0rWjz+o4BgMZOgZ7j0Xs2uF+L0StuFZTPrRnfeiNg7gyeoY65sj+XkDwFvrhf5R2CVtI499KuSZN
bHPXI/ei8vhQkMKxpbmIdkf63BKVf1R3niyKh1AF5uQG9R/bkGAaEGRyymhthfS3wdpAWcQ20RwQ
ghtJ9NUl9FGGRbslbjqHwnN6F3Rd2NOz89ij2c1XO9dW+4Xsez1f4TpACZ2fWUoMtb5Var1fOP+A
UjgkXZM2hAWBy+SPsG1BW7QBW30I4cQ4xHjbaqC1jli27c7Zn4XPtWIVGexMNzVg21KTOJ0yEuPj
8o4njOsjR2+Tbk6rRNzEGE07HQcTsJklYzmwaHi+R8xkJvr6nafXDYQQD9pfVPV7IphHW+iCAK66
bvLufmj+CsSeG/3UxuQ1rjNSHKzqxmB1FffCje0pgCj1BKZoDjIMkflBuw4kIYD3vr5GLjRkyNTI
AmCV2GuxqEIIaCN1L8crgkcbkNwyBKqGDPHqVqVcRb2Os8YpInNRM+2arFyLAfSwSXfUAhb8nT6D
nbPlkXoEZ1u+ET5BmXG0+62Gt13tnJs/e+CZNVKX/4ijOU6LpX/jeLxG0fMq0/+kCXiY2yZEUb28
lkPp2K86Ysbzx89iUn3WHiPHmoEef0QqBFiD3Ch3DTBNUxvSWuwIIyhG3DcEG6xuyeItaYXcp9Oe
lPhRojPMrcDTWY5Ywj3E/Kxbmoo02+XMeFzDxRr16Pvl/kKCc8gGtbAqlMo60tQJWKXCPmjVgWDA
8loUjwbgGDNPzhv/YjwsQofMH+R6Y7hEKFDuCNfMBA4zn7ZiMT0V7JP5ikyRmKrHBV64oD0D+JcS
SS0SiJ+JM731Z3HtydO4igONkxzHvjK26mhfphU6z/avfsG9QJKrn4OSiKIUbqxfH9TSSOgtlWN+
SOAte6ZXUN5ZtR8igbpSR8etPsRo+2R9A8rDbV3TogprAjTecNS9GktEuAkPSIWI+HCwdweY3TyY
zScWKXy2s3LiAVR83ZEdALlsYKWxSSWIbzHUbHkroZVerx4WDISD/CWV2aVFAqGMS6ePMCXNdk3B
OmfNO8OUkYOkwLYGeogVfIBmNQt7o5HkkDvVhQpVjF5A+uffOQ+7hUo0Wyq54PHnC5NE7Ec0EwGg
aVoaO70weYcOsKvxZF/8+U6wk4Pte9atkLeeOOfcF3yGHzsRyQwrGZfUPZ/m3D7lYIcx6eUGgqFR
IFbZPnLG3tfrTdqhteGz8tPe+UtEeviOIUi7wJuZrBHfGNnmKGU5cEgFjWwb7uDT1hrgvAXdRSMg
r0fFSRYbrdr61cj5Y9Vh+d+Eyf7C8NoPz+33WQnu69Kr+ck5F4kVSHgHZyYyudd5+XA836T605V+
Sdee0PC8NeMXeFP1k7Pd9VmOBTS6bZeTMrbUHYJ5+74tP7rTy93BK0/BXkceQVSQtzAMhdxgrqQT
Sv3oO2fbxLDpmyBgvxy+mwSp6VQUUDis/vXtFNxLH9oYDCJ98sqMDDS8Lx8uqaGY00zIfLEP7exM
H/7C+EWiCdAyfvA+cOXu+TjMwlKq5Jf/ukrF7cC2F8uNWJdxBRM1MczSCizoNAi+cG5wI5wkf8AL
VSjcJ/MwztLcqM5q2pbgx6RcyNYi9xT/CH9e9chQgzcZMSZBn8NOFiVX5668/o0I0Pwt5yEz+TIB
az0pvRKDNfrgebbk6yD3DPLGHgBX0Ml1X03okc7y06341dSoZjbt4mZ0b5GOzkEBqwQgm69xAq9J
OOlDD4DTH555kTMT7wgJ55ZysyOumMyaV4BJmL04OcEAX5eRnXtZmY2TUDqy+j5SAh2ckvhiZfu4
wnW7dXhuMMBOELg3DcmLIzU8KKVtE6QZe7+vdTGaZsaDj6iT00yLfQv7/+8jcao+vElISxsbPZ6C
LdB7Mtfh2QMxGbPRNHKh3QJKEK7DnxVylZb5+Z3EcEpRxL1BSm+7sm+x6eFdiQz8aCawXkSuBtou
J6MOOxUb0VUCWfGpFD1t0igU8Ih5Sa0xo5kJFoHisGq9aYkaqQvo8WyaNXpSJfO2M10rp2zVzuif
knEJ04gS/2m5dpXALYOfJ/mv8RQhuIeOZvdRXavrO5FrXM/gXvdVzuM2NCwg5Vdx+40+0G3Mp671
pAmNZ36Ow257+lixQSuhOg+mvM+EYKpenjZHLJt5uKsAxWrXUMpGxLeW/bQPzri60fQ3gSC273NG
ElAxzalD7wb+QtG+CySc5Q/S7RryJh3STNEXqHIQGPT9/WZv42bDk9M9jvA+BF6ghDlHrDvMA4+P
cxSOJRcGAEleXQwaxCo0hT0j4fvZ3MupImc+30TcEadS4feBqPGw2Sv0wUDSZJzWzFuySTZbscqm
fzhfxp0n48hgfq0ko+OzADTAa9BK6YP1vL5Bk/GHGH4qGv0e+Fq0AWGbP1RKoBCLV/YJvx2kTvkG
W2gKA1IMpIW1oNitBIWeRmLC099PzCywuWXHkvp85saRpTeXKsaJYAXOrkZS5hXnC4Qzre7vrGjh
cBDodq0XpJRsK8n7e60ZJekzFp8RxRCpjh2pdWjI2CaDkctS0xfMSrXsuvxmcaN3nveb85EKP5uZ
Qol+/lmIkLnAQDIN2J+0d4a+Xm5HJONKFbBoCq18TYEATYpaoELbcV04uJbG7BKito8GDkG/QGwc
Z6l7CbcCnHwjrlX6WdPEFHFIYlnyffgU82Tz0fkGyHA4lzTkpqcog38rPWJFCT2KSZwYz9L1oKYG
XuFnP0CYVT/80mG2gUYHsFH8z6odPbAzcPFQAEDRMo/7/BRymKCkFYBcJFQpHhvGA6U7ZPrXxhMZ
9ulR2/nOAuzMFb7QS9iyJYWoNichDZNYQbEz7rKftC9viGGeNtOlfY2e8B81CLJISdyd22PpSt+k
ThR2Q85sFjhkcauL1yEuQW6IohVKRWBS1PV/Ut5rMkT3Nfjk2PJq+K+P2ivZBH8bD5gGL7aI0Rnp
P03lizurrOTb5PNhffqWhzyrQ4ErUTc1axQXryrRa2My8N4Wsc1X9mnW7UBg3BmQAdi6fbO0zMmV
q697x0wcY3rPPovYV4t7nwGvKks/X34t7Ypvic9aYiPvLJ+xn+eLW78Bjzp9XsQmVgB7h9eYknAW
3c641Le7OqZy68eZ4SILzA5x8g3Yf1vchUzaWAGwaDsMeULUc2TnLLZ2hAbwr2x4fL+IX3RxSf+R
j+kO7nzatJLeBuFLGDSVmX3n9i1WJpw2EnybmtRPVbpLVZLeQ2HUHlFz12Vx5nvkkR1Q5GQj0SOO
svfpU8j4stv2jfW2XqlwrX247kaaghWB9gEJzD7LV9oz+V5yBWDnzW8G4fvECyoZZjKCNtnZg/XB
8NkUxOVqkWFtn1IY2nzJEl911VNNKOUyY9Itlx6vL3R5bYdX5YaXck5oum36sBTkkMM0YH9Ef6Gd
toNqg3s+kreT9BXHJjS0ZPXYrlUH6WtJyXSGWVsGkxWwe9yPOWjpFp5x8W1LsE0XeGlTmZjtx4y9
c7ioIKUJTd1SAW3CCUo4okq0aai2Cu+LdAhExYdWutJ1XwGOgwgrk7LYoE13rcPNe2synP3HhJUN
UztC3ZNbzyK8zsJrC98XTTljX7v/GeQJsBEnBND8+D8nZMjWk1sOyUIovdsKNvgzijsqqGBVaiNt
J4nDl6BtgquqXwCTp3QNldoVYfYfgt2LNnWn6g16yE/Rk/aJGKVpycVc+ouSLGq0Ifl7Dc7agp+5
CJDnO5AeBDBNfRC6U/qPW5j377atEOeAjFZtLdHGkLdF7dz+ClM7f0TEAG2GgtRiRa+ewQGV1aZS
5XM6fKmKBtAdvX/2yL37VINtnbBqKnzNh6LYbZYa7bC1DIWo04V1e7CdOWD5z8LTzGTmZCKnxKnp
5JkOFqLjWLlI635wheGDpMjU5cqEp/0xw75g39qcCDGk7sh0vNsLfW+AG2fEkEVHjq0NM61NOr+u
HAw17sq+6olb/kUuPZ/fn4rC1K9yAX+pONP4Ov3uItbDXxAYt2Zk5rdfb4bYerFO54H5HWjY2SS5
R5KoEJOxt8Pn725szmS2ck3zagAGM10T7n+nLRfG4xVbEqPMmo1bkLe4uhAYg/0dMaQBl5Brzj0s
4IJFRXoASAoXh83hVxc5376XcNDfA4q9Uy/hj/dUR5eVG3ZZXmtrB8bgamFI24Z6dzFY4L5D8gJy
dVexS0vFC3biE5Avz3Fe/5rhn0B0fmoiR0ygxwKE1PXvABcuUIhipC3llZkVV+4/BbDzD2N3bQDu
ZlE58tv1vtx89un57b+/NxoYC5pzUoXyNDcjedk1zH8g0UvzjPjum41aBpL8T/AvDBW1JQt+Xf8K
3jCHmQWC6E54MIKPZfY7GS4mQUQifAtTYEcd9Mb00HSlrZ8QhKtwXy+I7JqMf0MWAbNj0euJQg56
fnxzaSCRPKsDGYTDlc7aqVzRRHvI0v2UP3BiHufs+vUnvgsL5dvW5KVqPuqVgZmsm/dFMFNlD1bL
qWqCDAPIg2DPK195cuKoOIlSBbYiFWnEoGN4rKAdvsK87qTbgp2dVvL2hbcRWX0q9bB0wIPq8fVw
dOx1iwriHuLFDeQYBuppOC5LYhSp7dHdX9aoUypyb9k2aarACoZlBZ+OjVM6qpasC/KLawtVi+Od
oJFoxCw8cjD+VJuePOrkxDB4p8COfUsIjSbYer0N2/Ro9CTC2LUhw2LoKYJEfv96IsQj4xWmY38s
ZwEHEjG9hjfrkV+OkaaV0dqmN6dGWDOlO6QMVAms/MC9wDa/ea5Cu71zFWZ/+1ohIkhaY4Y7ragH
5r7lQlXRyvdpN2t0Kx/h0Y5Zl4ylILlTTDp4t+89iuIL2Y5w8oT/LhPwkgOY/c4mORybRu7AUx9B
oW+A0NJY2rU/Kznwg2D20PxHJdN0rqU+vqVLzR7QooKaxDQCoi8VGLJjzBpTC0QdyDnUcNJG1Q42
npk3m7wQC36CSqt0zhqC8hq/lTYe72HUTZHxeI/cSvKqDWVWBGxFcyl9va9WIm9AfxnKF2iaPWjM
0eSonNgweDo+oK75Fcusl9pKEfkVd+0cn7dn0ltsFwwISB9qfR5ZJVwuON7kjEoDvA3lTEIF82cC
OL14vfpKPlrECLRqCrYTsF+0hJnOhsd8VvT20co0YGZxPf0qcaM4jj2OOJxGTwodOhwL25MXEbMH
lBrHPhUnGydsYOTVi5yTCZB9ntc/TzmxRIxxE3X1qS2SJvfoq/AWYfjCKB4uT8C0kRedmT/AmYax
48PB4nbn4vDFCuLR+FwQytuyhkbihi1aCy7RodYJ6TObdBQeBiDlytKl+Zkc5VeqXWqBnlz6R7B7
NedjvXxRnDY4m448R2cp0eyu+a/qZ0G6eP3KWJMD8hmy5YqUOISPwyI6qGttfz+KkBhl8Usr0Ys7
fPV3tUBE1ra7ODLG/Z2/kvRzDrMdlDQ8ueDIe9OUCcd8UxQzPr43RolWA11xwCOhDhY1G6Exziup
ljWJ+j42S76J1C2cQ7CP73uZ2KJeIniPQZO9iLOHXZI1925uWca9VDfWMuoPHo7Ei087Do1oDhC0
S1M7jBzvM3yfGvxBEhyuLsVvvcAJovxQeSqpEnTIBbLE3vp5lzaVPdLv7ku6CRAlHov6tmItbcu6
rqbEOVXwN0tueApu2L3Ni/qxCncz5b2pWjxruRMBdeL3FBM1NhHbSSxtpIqbugYmQ5hTtJ0u183s
JVwpw+VkoI8+ABSPrYz5fIwCQXQapGXYRCLDCYENGKnEgWquGtissX71IZn/N3OU2AYOCLEcizd8
fi1LNZ2s4XQGE/n+hUT0lgBtMNDKiCRAhXpN4ZC7OFY7o+8Ykv90kxLc+9JNSH7Se1EmqNOoqA9b
HnHQPkb2qVO+37UozF3ALr8LAUt9lnthBMs67M9QPeZ9JjCD9B8ZPCfbvgmuKMJGjfLZ9T+PiDuR
+advLzN2r97pJsd6KoY+LbB9S1La1oJJ1nQqa3V8lepKsSexgxUoxn9df3WT0NzkBzfhYO0ZqHnF
mcIKn73T6s+8jx71k3fO5RUfKJMHduuCVX3FXVflOMS854+zwDT0ox8Hg3cXQOtOA3JEH3uOeqGg
2V8TLw9p/WO/5vxd7/VO98lvU3j27Iw2U+A3on7aTmUPyT89SYMdfQYaOSGGnSCkqwTcmQTMHH7X
z0KWA/Dy6W8m3jUfUwkTA3BGLahkKuhe3EG7sPZqeAkXDV6KimLjdE5mzJ77kM7GGRFOXZaYoJzT
9f8eFzvz6FddWWDYnOKa6l1Ys9wZ7mqqznEkQfiIypXO0IIgOKPlY/L9FAwr+wmAceln2vZZosAW
lS8zTpdjJQR5rkgbGLS8kgb93/7gkXPGt0O/y2e4OG4c5vGJp+3KR4B+Nla/IP4JYprNBE2W2JxI
+t9Ow+njWmjyBKRDVUUj3CcdsUvxTu2T1LT0QWLwXLn5OID1m4/K4FCHRThbEUvqD69QdO9Uh4dS
yDW+Vloa6tCCIJeK8asTtkgfmixJY125XmBfaUxTqFYP7h/eLCp1QyLaKYzWK+Gw40UDQ9LzkI3s
pcr88JE3//oLsjI2hm4h52J/khTA/NJi37Zo52MIFqyWmwsoM2iXWcUdjCADs1M+pNEukk0uvwoS
Oa5jnE0N0Ad36t3AYGci8PE4lRBplrCf5Zn7IdZLo61LZ077nv7wxAobLyoSGzA+IlkszOPA8GKq
5teDKyzoNrRJsvBSZuDaQ4xU3KE6ZexZdgRe661rwq4pE8krZmi1aXTnM5C+SLXJwiYSPa1RdsFA
iRi4115Ts8cgRJIfDMNUhR4pSNZ1XpF6BzhQCw5nYRgfGQP7WmFmpXNg1bDWnOtuR7gQG6LwSkcI
eHF6AyLBgXRFcW3/8IRG7sF5AVeGtJx59qMPKlXrc1/ox97EoGGN41Fs95f11JOFUZ9m2xYxJbMl
kteTcuB8BbNm46n3NnUhjIbjgKoDxVKq2sIqFERQtq7qODUZOGCIrvZlZdYqaxz4UDMFcaVpK/oz
lS3qYq+RP0ITNEJtnSrppKlAiO8mWk+S6h7sz5lVGleDYzSyM7UBKUh0+0VWTTfrDKY7sy1/lm3w
7RQ1xw67cZoloOu+9prhg7etA71JluN6UlJ6As0fRZupbhgmhrUo4FcTRISjn4d7ck4n68CvXrWG
6ekPodsEuUSULRJBDAREUB1t140TYyTDrJ+v2AWsbUI5eFQ98ZxzejGs30x/myR8uYJIe5FKnxr3
VFoX1Bdw+CdM8NEPhC2sBhrRuwPHq43g8zVAz6JrBBqqAUaQuW6dYWAq6QSDw8Qd8wFCTMHJ23BZ
7Xw6BBFetGD/yxhvKT82p2xtWpkFxY3yfH0XdXFXQgc8LzvWIsoSoFeXr6HjeUV2iEBA8fHYoqb6
b4tuupon29tvhRyVqVbnPUtdLP1L9QTOtiz7W0iExkeJXUNnzTGIVnY+NwoUIIFZ60P7UKErIpIT
HRKFvXMp/SLO3Okqm9KBwlB8VaGVy91VO8b5Z6IReId2jPclfjjCjQf9KNv3poJlZhe2EkbwSjMk
1GBLS1jxbqUTdjnqxHNeEe8WdlyQ/eJkrDYDiRu+yxolhET6LnfRxkb4LEzx9Hp0xKptUmn0XJoL
1tF0Tt5Gt7CLd4tEZ+cmg2LQ5lksseCD1WGgUriAnmoT2BdXtqYOM6gAkltCFthQnLXANc5DIjbw
2HPJ40mtk8bpU/Z2OyDTC36prBFB0BJgMnjtQtnqEbn/RXJFkUuIjDLwHKYrGnB13pvk/KpjcgL+
OJXC9HrbQjeptzhpOVelPSPg3wBSAuC0S/7YNEnnhGTMSfcnbXrqZ0KbUAER77oA+7TnaLF1f3So
Ee8iSRCCL1JRMlj+SW5B1xpeNEeUCnL2+MER56aHdd2CCcMltkzMggI5UiPeptREeNoOWpfB8gHW
nwoQHnRlvODUxR8mm8lkz9Dqgki4DdMJREFZJsyC7obqOjdG06JxovfyYb1RHN6q4Mr5QIY/7O1l
IlyFVWeW77wD7iQ8kX5maP5ilaHD1SZ3sngiOtuo3QQoodXHv8vLNdxmUnh/ImdR/Xb7EWfybq98
EycPSTpwRDsCTAewQyty7ywB/N4Y7/KPk8cZx8i3Tkijdd1TI8j9H28B9PgKUp83ZDjAmUJ/4TTP
8LEKtQNQqEx+QoBxMoigzglsgq8BHzoSka6I1nax7cXEI1ed9+Cvq9JJMktm7WA0bRBftErh/FDp
EwW9hVCuQTLsPTlJIAUN+b1Ire/u6KinWyufXVXpYnI0ABdeJCGvwaoqzEpuAEUEvZ5lM/5g3IM0
YU87YsJ1Dr5gNX/JxVxZC3d7x8aHrx8wL50kEG0Cl4BjcE3wvlpFP7dTsqBIUsu9Agna5Se3BHkR
Js6/EM2ml+sZdaL4+Pnk5tDT6TpuemLmq5pFJ3Da/qVw7hQkviocIvJYXFDLnb7T2kLq8ryDJqXR
9Dh6JLm00TBo9AsmIRezx09OqWb0UfeFeW+NKxIgXSBgQYrUdlTWgN/4Gnn0MB/WGvbQyzkW8ISH
pSviJzzMo3ADnm/DZOpNX/ySbZ8Wr+bBmIqYCZNZgbLAJ6OF7RL3N8nQuGn5zTpxEa4o3yv0pffn
FvyiGSfO7MNf4pLg/F9VY+my6lJCrE4PRB2HZPmu51UyweiIe0dL0QxXvaKTkcBM1s4YyIZZSi1+
f6Zg5CHKhoBO4tXBLx45l+9nJ1I6ZWz9kub5Myy5Tmb6IOxDb7uZ4/ZnrE9yzq7rF+JiYZw5B1Ui
+2AC4qtm6NT5jd8YNVos8NNfy2ddy9QBuwkbKhMeDvSlUd6f16sYuxVCXAE1Cb6DgHuM+nIshbXa
UX7s5iz93MHWMXc6jFblgIy+surLeJgggYNG9ekH0yy0PmJkuznogBSIawsLxlYK2Z4H8iLM/nn/
jJBFPRVppph56TETML3KUT9xmvpyxBdadFlhpDlTs+/eQyj7DdIn6rDkbqklF2AvmVrCiypPT4sS
Wg0kAnQtWJUSfJDfFyXqVaTbgNQAduXgjJtFuiP2BZD6sM+BuT1XOR2ALvDjWScz4wjVT/P8I+Ha
3dZqrFsEZCRvmp7f6sw3h4tYDHT+vVash686dR/Blt41W5UT6cdR8w9PI0GG4OfvEb59MJeWEwUD
UjTlA+1o7+oVlCXWdBj7fTIqwmyzW+SUzWVNV/GSvM15Jd2uEq6Gx6YjbkBu/XBJEOXJCbTixCK5
9yP26URUa4tAS3/THbYjebulhR9z9w/nfAdaKbUpndmPN9ElrVw6WT4t58RMpnBcJhtpUhRDecLY
VJM//TmgsUA36qhhVyevF4/b8XYkZMfl1Y7Std4J0wzGhtSYc5G5J1skoUhqhYnMUc/6BXkoNaAW
89p23rJypMiEQwC7W+ifltMU+j3G6JFwkCkrFkAHkeT2KBMEPz5Ock6UgADQuKxYIGT+M7CPxs76
Mbb8ihRWDvr7kp3QUUZBBBUvjK+pB1JDmKIh7cSbgNcruek+Cw8cEy5aAXf0Q/Dv6L1XieBR1/La
1YFPcbGNwqklOh9lG7dvjGLHaQeggTNgxvCdfy9ig99KYxbqMebko1ZKWfmDpIhLuiQW9AEJJSZx
PemUsCmv3T/dL4cwsYLoQTVzxszU2siJl3DN99Je/s3yAkM+6j3wFLRX11fd6jjK26YRjeGLoLXs
rPEA4AGYZoJoja20G0R0HS5cD5VpIOu4rGIyF+zruQE2sHcTj6vus1GgauqyPnIpzZC8rb9q5s9m
a2giXvvCWKWkHScCn7dCQijLz/V/WlWuNsorTD6XG0KhKTrdF+wZxUVtM6/vK4XTXQefexZ4MIhH
UGIuDYwMolxijFSOF8mbt3pT/rWeHu86KXL5ROP/IjvG3S5qJEDMu9KUsywYW9K7TJlfibt/TcVc
gBcGg8nQcLETl2R5bkgTfSZUKNA2nVWr7Appa9RV3eG+o1OYz08QkjRX/5aF7zFhX1CWM+Re0vIC
bhgSQlLpPC1UkjmU0iL2Rwa6wEIrbb3n24hB0fprbwug+vYhpNYDi05eXoRXNXQxkVrGNL0Vpt9O
akyD1cF1nnbHo1ogKig6eMCdgyVyVM0mNhC7ljmCtwK6SOdIPyZnFHnSopf4KKha1rDZqzIajQv1
gn9YDVtRTdyUggCdYyFscT/SIYrNcBmtIEnoJpAbZLSdLEcxIEi5ruP5PYk4Q6pkE2xdSr9CcQtn
lEwtesELEP12rgDrysXgYrN2CKa4bOTu6FMArm+aGp3EO8Ipv/yVU6nfyw3s1IiR9FdU48UddV/p
aHzqsJ2UNM7KQY9i95S78lvldVdHz5JCZFJZeVi1NhgJXr4H2en6DmUe2OaNDjaHjSnBteeWC1SI
g3Hppln6tTkClqbDaYF67WGhIFT0qsz0HqVTbmJ0Lk9lzxYAsEAQSaz5pOJYhbbTYp5w8iTyPBzc
ETr+bF1PTQoXva3XkG+MdsQXLclCRlHVb3Zxb94S82sYrNGiFTTtiDCTNHbXOhpuNT9TLmFJGQOU
rcfUviVxBLoGHofQFjvEjKvrMrpx0hfBnf3nnlBdyoHpbaV4Zd4XJwK7kny9/0IQsTi0xRRIs3A4
JIJUoJimnQn7OO2u5p+MdhK5/2lvltOxWvod2bkUm+zrZHCZQ+NOgqTAy2oc2IcP9NpsPOvNRzI3
oGbXoDu2kcmSgUB/hKsPJC1Gjwq9hhk0lAPx56nCi05N0rss2N2q3/TcnBuAEuklPdF4erbRzupa
nhz2DZCGeV8EO22wetO0UwrYO5glFmNqDaU9puBJWFZOn92nUHPjR2wPDLmEeRL5FnO15Yoqdwtf
BQq1hKT0xBx4amBNCFntnWABrKolBM3HEkB5ITmcAMSgV+yXGSHWUCpyVcVch5bOx2qJzkhjybc5
VXRZDZ10/WpvbFQFN/UJpVb7yKJOPwJvtaO45GUC3pTliIG6UKfZMU11zRdltcy9c+utvt47hOSu
ZVxPOlDRDh2q1LFDP6BuquASteuPJKGuBuu/LTG/FrzysXIBFvHxGE+uBJ2XdnbwroP/1HM/eYE4
+f0vWdBr2We4yp2RP+OX4k0zg8H0cXQHZupsiqqDPiqAp4jnqO5/Us6o5YCWWZlhpeDpoVk9QVED
aatWrSWwnSQRij/lwaEEcwUmBI2tHrNykxxSKneRjpDNDC4dyPeKJcFQFkvrUIgIjY9eVwioyv4V
RaTachpEWbKrDTKuautb+vU5v4T+j+pNi93nyaiQbnmVqk4TmLVcOFTt61/4i9yr3r2jUSv9RfNn
BVo4ZDfQLujE4tp87GRNcOMqlxg+BBK9fC+UwEuYNnqWIXC/2V9TlYEu93sjGQYpVPBFAqhTqMqB
lwVubkBv9oof+Fbw1YGCP0tT4AbHXt1matMDi8+YMa6FXVu/vEF39xT7NAoz+ErO70Zycu45jMGV
pIf7JNSt0NDrOnSdLDJYnmFSjg8KJYGKRFmQrJ4fc/SG2VPSq57IIDgtlK9dlTfm08OoFTvS6awM
T2rknegBoPYJhZ1GreQPbVwTLU/H+kVs38Bl1jQ57X4KGPtvOUKEbyj0owm2ko6hzyRzZ4N0ignM
C+T4k43coMq+oZM2tH0HXFxHbZJ/HzeHb0Y4fswdKE+k+CFWJH1miz+kuFjkXUdpz5xyEQi0JCF0
nbD5HAZT93aS9D45Ps2dA3h+bFU5cfflVQkT7gHLzLyu5KBqUtPHKXJWuCa6uguMu5PRwZ+h1ERD
DE711pkOvxZh1+MFkHMOEcIvcOvhE5bq3xdZod4bzjk+KLfOh056xsGl9O7zKk7iuHkEgnLu5Dkc
StpplbWaL6zKksEQoNEEsr2PNjt9ULsJzCOmQyhiBBZ45LDH5ZSEPQ8/teiIz3ClgmNw69IzZCy3
TAqiOnusFsTqMBrvklwopp2/LfHpIVwobaYXDYZWqGdMBN89XRdLkU5ZfQ68/vITIzG/RHhofV4w
guSM7WEhMbSnGMxo/0c3U9JAOpLFyQppN/UJNoXiRdzewDajuGoni8NY5wf5zpBGrqhCtYLKH7Rg
QK0XsSzmBOqQgJVpoVsaLavd/v+Jy7drFpbL6Fkd7GBBXZua8zMNmlFo9X8H4oPAsFUNKuAbpQME
JvkJMlwWWbja9KIFXrya2B7By7BnlpkF7OqHglkh8UxgInS8IZ0+pBMptSqodH2/ZD7dEsyxV2R8
PR/52GDfYe7qRwWeg+BVWGLsLJUadT6Wy1LEzT8JWP1uW0NED9Q+TnObPLa/CJl3AOxjdIbZmfoZ
qqlzi+mCylXYaSEztSoV6PbwHerZxNX1IqGiMbkhBHZ7t40E7LFIvBp/AvrxmMTJ4HczpWZrCfQ3
PmYRvxC15DbMwSiBWx4SLpAXZuWrfpKQpgcJJnbJGxor/SiCgaE4mz7Xz4Lqsjdf0fHQdYq2QLCV
5Ifpjc1XdPXZ1jcNq6EJNMD9Uet4n3c0Sy8hxe/WqAYxP0hByDEpp8DxpupGbB6hLfJEguO/jdwW
fPWJm8cTsiMnNq3pgi6iB+pw9tfE8UdVJH3QSEiJgTdtSf7p4SihxOcLeEae0E2eME77+eQvDF5k
EAhAIJl0WAKwV6IAdYRj9WmmVNWFSS14bw8VpQd+e0mllQOhQ4xHnKusXm0LCC4SYC5I+h1EsSpl
eYAd1eBVu5KvUr5F40VhyIi6PLnXlA44KO8Oak08xAp1X3bsuVxCcpIU2zo3+9d9BM0E1EtmgX2k
Ts6a9dpNjQrBaLevW703rxzBuTr+ODqqQdhpM03mQ7MBvS3MlfGoWn/tbxd8AZDQRtUwPuAZc88K
jw7dcrwq/XMYkpVdcDoy51jRlh43n62nW217Gb8GpubhVt+BmfOcJkpDq1csubr8gG3QycTp8tAh
ZSK3oMnNgkZNfTTo0hnvrfmkK7WXxNn/ppg9ae9kMF75QcIA36puv0pP++gB/9sjS4mXDlpmQdL2
1hf0nJXXxzSvRXEL9WMhzXDxSOnUXZNty7ApWjys2m7u0HU6WYJyMxXoT5RCAx1f793KlmtQG7+j
CoMMaMKp1lsUbWI/5m1tKek1XXfMyZ2qmoBb7gHQBl598U5SK+k8b5QQSEeE4smh6uT7Fl+RnzG7
zD9/BEuW/30ykll6dxZqVQyDWYTGqfN6M/l3hGUSScD3ZsAVlIMZps0JaR19J5PyoSaFXH9lfxHj
TyeNxNS0pmlgLUX8LgyWXbBfVX+/Kg+v735mWWBkqSXai0WDqLQKRVUy8GkeHGuJNNhXyVGB4z9O
SFUNLY8T/FisVryWRRrXhEfCKzfXbcXIc/PT37M4cg99w7vT6FIJGs65Z8NSu53qi+lUMCYZATZt
xZ8BOYo+r1ypm0knJBUgFxcRPoHBUbCjhh+bLFxi6YmlsVBqRIUrvza5WmwY2zkHByLiClXUrvGk
1nUrHYnK/qYEs5ao9MIRpeUEpm4alMe5VeRTdKRgSbwTBf0dJoBMAg02cGpzvgvQUzmMPMtCXLEd
lCBdSeq3Y/SrvHgO+heI26uWSlHPAOq8IRbi94nBBxZJOOuCbrw3cV5OXaKNy4awj2yVCjhD7+5u
veN1kC/YJA1ynpAtAjnqUHbVoYYny2yqSDtZakfoKtuCJfqSj73KwVELwZJpRwCLHNaulMLqTvw0
DdJ5507lsyI77oKxgW97C5V7Abg0att0BMsK+TlMyV6DuC084DUdKlQNXr3YxNRd/3clgEyECvBC
03V9tTr+sraAiS+Zf8N+VPmHvnTSKM4dHlszzmaxl3rX9v+q/+RQgY0KM8vZccYL5z+y/IoLV+1x
sDjegO8sr2DRHvdHgHfBegMyrxFa36pMHSSqAeBuE70tO9PG0jeqQbVmZ4Jn4is3qRBnJse2xDUn
PngAVJ0ftqqZpwItunSTQTbu/SMhfimXCSNpdy+guHYE/eVwwefzVBpKdMsn5w+oVT2MgtSKSGUk
E5sM32gyFBCgttvnDlvDGd01G/w361JiVw771shfxmZB+KLLyj7EXYKMJlCGowKE5NCH26CYsqIc
2R6he/m40dXXneOIozuot0eRPyEcBC1NdDqtHDeC/B/KLmAbFXyfnvEaZ6StXyCKMzF0z+Q/zV6K
9sYQtOvpDoznUeXbKmit87WC/nxxMrmFO1Yl81WNrw1RS3mO4dBRYRF2MlB8+zCq6VEHUn0Yo/Lv
EcivjoWap9JtogbUUGlpAPIN6E/BXx5X465c1rOTrCeQxTPKsyvrHq8UTI5Sb6mpmcOSNidNg7KM
mlH6UE3Vz4rvy6KmhyAzR14JuX4LwiS0NFeu4o/vp8Jwig2CpfK/7ecnWTTVbuOaUUFgdACvr3nw
uiBUQZTFOovcTcX6A40/KiNeLS/8DKD1a1knoqx8OX8SV552af/braA1I1LpxayzWvqxzZZ/m6Go
Ll2KZAwcbAaTlb+HjW3othoWGIYP6uh45JMNLGB8IFXPluD8fPUYITJJKjMsomNxCysJ8w3pXQtA
PKMZFge2mpCkUBLOlXOzdKmfQ5EsYfhSL3ZQbUGBvw55KT/tK3ZMzr7Do3O2t5cXJDsh6uZKwSo3
ClplNa4m/skRmfxRSU7RvHUt5Lw9rw5mL+hT1wu/do5oy/DM6bzci+hpoBe61NkelN/e5YOTU8yh
M5mChy0iwGKxdjb9KAtSPh0MqgRwST4iSzLxn2TboWUjvohpJJ6j9WrzOOAobxWQBBK6Fxx9KZK6
9QoIg9byPK2zkppjjI30/4DhezPugwBsvoldYyyzwYfLJR+JnM2g1jC3Z9t1BcwjpTgGtrniaGdH
Qu15LDoQppgI/svOHTdbjHP3EVaDTAltMt3tBmMyRHoAo1NYtXtrNZimrBKAqRaDNARLSMPFe/fX
iVnMGDNjjdUXSfTzrHLwGWwB2MHUWluupRcT8ECu8Saev3B/Go8lvyNRgzUFxFr1ZjQKnCVBQLqF
otXRrGahedMAW3APGhc4rmIdS2NLOylgS5tvQxKw9iBM61T98tRzjuiQwBlxH7TEXbTHWNyl+Id2
cj2J/RbJjoCz26LD6WS3al62NoQ4HJFtJRsxY5jnpOhsie19LSE8Ay/wBPFfgHCH8sLmuw3w3/6u
eesATZtuf/84kPIhw3MK7ruvaD/ss4XqyqKcKd24mZdStMy8BWNtuBwNF4x5ZGAW3WQ4Rs0gBMy9
W2fXNutmkNbOelshZyJ2SrfHbMK3qW4rMyyn2R0Oz7GbO5imvlGL6XQonw+coVqkFzBoZZnP9IMY
4Zc6h2Jpwq3CnKZXdHG3fKE9BhgRGHQkVSyb1wneSnQRZHEizdsU2Au22NXCwK/5xVIJJucuoFas
XkHUDF3DRyUQ80Gp5CGU21k1AOtbr83ZfqJBrAJ/J8qesoTYpqSGkpdsX0Uhbx8C5uZbogAvnLA4
3MC8Tq/zFzQktw4UJukocjUblKqIK59uM0f5D4NcKCjpRTMRzqtDzfZb48zg14IvhYz5ZCg7qf4d
MHjVkbVf1Yg3iIZRMgSi0f/NqkgGKLBYTTLL2naVhqmvyCpQpTLz6NCX6+T4FxgCebs55Wjz8ubC
tj96XTZg7bSfoXadugtBdS6zAg8vHgr4Ab17ipm5OJhVIsWf+IHYmmfOmobikKd73avB11aXGVwI
PPi1I8pa2Tm9fMcbndjqO9U8bIrG4wgDib4pZb/ib2jz/tePTkEDugdaF1saZxlMHPWLbP8pKsgC
ltbT7pHafPiOJAN8JoHFsQlioayYmVVteeEVM6CpcwPKosR0sm6TJMftpk+j22pgfiqPfqlHe6b8
Ty5qSknuG6dV7hC7JXU3ZEBDxOIWN4iTfKwxOmX9nVuFYJ47SEY8yIwMsVlht3t4CGg5DWlJ8Y3B
hHZaMtIP19HberMmQ0gX1DW741tTggYa2O74fYAnjjw/9D7K6s5RzV6T5cicvBcra+rBeRsVZV9W
nphVnCwjVNkbVRjQk9ZVydCYncCFn9a5NTiItlb7R0BcwPo1lxHlO/8w01SMvrIr9G+i8z6f4Qnk
CfcTP//rLX7u2MQfim9i/GkQw06vAu9zoSJ9Mjbh7ycrbMKHCH6lEpuwHZqCUcKW5V+7vSu9xBD3
6iAav7hij3PcgP0BaZCGtiVlpKaqxDO6PFv8YFhvPqlRkDfZW5bCKWUd44rzX3F+pwD9uUlPTyGA
nncCV1P+kWCUWq9vof/x8cNOBWaBceQsyaI8L94jMz5oHXj8yA7bcGVMQYQt2kfUREzqDl7+Aopu
pekaGHho0yE7VAx7tB1KprYFkqGKUM93XlCBtRIUEJJC+E4arJSTvE+xlXY0szbLuHmoVR5TxmFt
xvE/YRRK4QGbJevLatEgl/+3DzKS2oIB38lax3dpSVvq7YQxk4xCLiOWa0gurfLY2galyy3a39lI
mOhK4B1WiX9MAsIRDs9FqDBB24QuEE241nuViKCcGJeKCiauvIsAXerkEt4vzbaKOOhNcnXdksLj
p+lvEkzQ7laCphFmD07Ns1O/ZjjKVdxIWJbwIKoEe6SuRdwT53RJ4wn5zX/50Ag1zhspQ/I20IYH
HmXi+QE72P6H/ny0EQCB2/CX4ab19VHnKeIDN0KBXp2rBlw3EcITbNHawsH4Ehbny64sQErxIB94
rJKDZYYNVaY+Ucdq7coOcoeorOfmnZHB1x4T1YkCteJOhVO5vwmyhHI1RaNJk2OSMR45fd8jk/vI
p69ozbiTOr9d3nrOQBSR00rYD2sgfG3bCrzwYhGTa+cQrqFnccGuVwVNxLWrpui8GfWu1Ul4Olub
OF+OgsQ1cJkfRRJoln65NkgGVWO9D0XKQErSi9FSEtnfJrO6ypGC8MbAnwvZyQny3kzQ1WiXkk7p
2BLtFo3+ULzZ69PxjclVRreqKNP2a76wzMb6nuU9PyCutQtpXjbmjHQ0zPXTBypw2VZaXD/qgnML
H/kd5ekKCDkUe4JZrxvPyrKQ2l2iSTwctdWdkPmicoGEOCABSDRvE/fonmtZZGKugPgPAO9QDaDE
Y0vGZnoYkSbB7tELTtrR2hgoVceAroJUo2IpOcvKr9cPx7fhI3jTL4tp26LuCkfVyUjBldQvlFxU
BSkeEVXZWXne5LsNukE7t1hVI5y9GLj592oe8Z3k92BEASpJpI6DUfI8bCKsIkyIO3oGhgqH/qkY
RTFc6gXRE4WaRmSUftQO4iwG5GzgJPo3T0eokeKqoxi6iTJML8m8FOvjffW1NleM6/aBNqjOrR0w
k1I978NcpMuYh//pUXHK7VPK9FjNMq8Beni1S0po5Xls3z8g78eg0j3ZDEW/qg2kPv/SbEv3VQBp
Rzny9A9kyDj+o6xdLLc2XxiiyY/Jul4J2pz7auqwNFHjIajLjLRJAfh562MDkQwdmuKMbqzS192S
DldldwLkDf9x6B6h8zwQw+1CTAYeN0ak/cGzSmoZOelOgZRFug0y37B2IOEiGSscjUv5E4/zyMuM
3VjQHGsXPExPhyPKuZ0MfNMNUtLdCVJT+CZ4yDJWR1aRkRdd+YgLLRljuz4soKtbsFrJCxxd44/S
Wz3K/vRVsPpVYuVIWeexW5akiw7TJ5oMjxmqmkxNLKKYhdYq48J01yNnRoLVK7AyvB59mpjHNCAA
4hmzTNRaP+EvGUj4o5Av5qRXqb1QCgnwEexucJIRhYZ8ou9H4zAcfDz+4SOwbjsKNG9buX1p5i+y
0bc3nnh7WwU2lSXy080qk6HpPWlX1j2P2Ub4Lq0sfXt8Cw8R8Eudov1o+DOslhUGL67Q7Gnlmzu2
IzQ7r0Zr0wQC0yTVgf/sTL40CmG4ean4Nl5zoIJlgWKCFYErOt/jSiV9FKP/qYIhkOpPhT/gD0As
g/9I2PQcQAfgieIeK3LoW1IF0VzN5qPmX90jiGqLWuLqBVJNuIHh/69T3Sv0j7klY0LhgZgiI/Ad
fylpqd5DnBhVObEaWT5eBth7HHyjBV4WchT8OIXxsvINdPgFJNItz1rETT+l+5WrpguZ2xLoCm3s
OYyBU1N9pkbs1MRpuB+0sUkdR/sjBoDD+xdUet78v1tSesGMbYf9WcnbCq5iejtRxV6ovPs3jT2b
fM85AD4zgz23TUOWzIthcWzNA2WiEP66dUHF06aQ2RcT91dXZDbh5a+GC0QVJRi+A8ZILpWVPIT/
i+aNZa5WKr8Y0WCwlk48kf7etC3qd6aA4FYqYBnfH+Qut7lWcbhk4qY+Sa6rrwFzvHgpZVXvmWk/
3TVRcXpqna5yOlhyl0j07BG0cizO3cMxZxPfdAJdDz/PxDpgWN/ZPkbl3laY3qQ9jrFrHVgZpFQH
nbHTfY3ULlFf34YRIBXoRYeM/u1V8p/9HlhGqYkAMUuKZJlyWygUYniXscM/l/br4IB3/Ng7DgQ+
4h93ZIerpo+upH6uSzj27L/2YhlOjgARZMHNPFRRomo+N05zFfIqx7Y08bZgZkB6/+TIwsaNnJbb
j52tRvHVJlQV58kTbO5s/3mlZA6JnjYAZO4/2T6T9LTCCyy0PnDQ/wRwNZAozkvsL3rISgLvZ27U
RYaRVInAeJjTN6GNZBACy5v/rE7aQ7sBkE77ea5Cb90HE10yI1s5auw40+ZtONg0vgwJc/kWjHLz
zfgMW7EjkBvoTVTW2qQI0YjIkroU9xrHfnLLuHEC+NrklE9kLQWr140YLVBsaCZAy5PejKXquWnP
pCoODGg6Vj92ZjD2eTgh2da9yiHLYzduuJtk4QvDvmlEY4rVy15fTpjMs4uQGTTX/oKx0s1w2+op
rfuuHiQkpIM+5NVl0aZXg7cg3Rgv1ViYMy0nxc1oZjUJ4aP66lVJrK6ayHOuSrKDuwV3T312b8al
78/JVc1Dq1TMU445QJZGAZpKTYNXbbMHoCG5n1asQRjy8mB0+fDmb3+2Ng66FX9lfQ6n8t28gCN7
EC8TqG0lZuksgUzoxSDSdcM6H0M3L4Sem3S5hJY33NOB8Kx+ajgt2LxvX9MPg2E/OwpNXp8ZuLDI
W93DbqwII8lgjTlw1rr7Au5DRNoQCetgf1sUkEeBQQo6Jiw/M1uH+bs6KM4TCrlM6LgXRjPtJene
uqmNc9z9OsHgw37vO7YzYmgV6tVtTgadj97WOCXzac0xFvBwi3aMDofIdVxzJo2GnVyoufHz970c
1k0YVk07hVmDvf0QX47mDR/3wXaIae/2T2vOHnxyfJm5ypAhVYReCSHvkIuAUYL9PyMZ0gHN7nXp
KTyXf+oYc1m3ANZj4SqKYLT1CF5f6t0hRKIL5M9OaGZqGc2gXCXPX3ix2dDaXM9nKIEvEhkjfIWl
6981KekiSzSO8hzylVNn9FhPWa2gV+k/mtni3eB/SBfBwWpY/3BTsBRbSgcN8qL5wyaT4aqS07Kb
+cLAP99BKUaEJXZKRycYMaywyW2GDxaBgFMj/YljGBsok/tgYIW2gZy6qbiAc3lV6pKkM1pWibKf
ODTyMWQzVagMI6UB3Ko4huVHjtsprulg+yjUYKuPFhC8Z8xR7JSzLLvLbY3w29RmN3Fj66jC67eT
KD2W8LCiPaMunXuXy/lbvxXp+kPofvGU7OE4BFeggvzksDCHxR+INYy3b+NTz/ATWtPNVcKTdgrE
fg0bpYUqxhgRfeV2QO9c+6pcAtKiME+iEypF8wkcPZmN3BS40fldS/wGYy0bI6IBQ3fabgr9EXvi
fjuJ2xg0SRMf49s49sINJHby04XUl/JbJfUbIZI1CMR/59wI/eHdOmKE/eIN/RWCkQpBlpMa2iIe
8L3Wmi4vD72FIZ66BUQvVRKxbUWN44YoEYsTf9oIzznvQemZRDCatNr1HFOb9SEj7NMrLZVOwGJW
HjT8Q1quMHZLgXGAgMshUwRSwd9cg/oXN1jamogyrZbyHTTfg0fh4bubU8mPJY+9wl02XPO630Nv
E5eP0DSdQGYDdqJgIxnfNxZ/9pLwWWMwUG7R/+E/WCZX5A889ViyRPdSk0ybXB45Po1xkTjjQqhE
9Th/cXiVaY/5sQefzHO/CiZrALmSKxHUPO7HoWXTfE8ST5tr5pxx6R9Zf33oHnRbElZiZbbedKt2
WxDt2LeogWvOsQX+1Fy5fs5/dbY4jkmomksU+u0Skruz5tvaOUgzZ6uyZiipwgRtpWqAhXA73c5m
BhrOvTkSMGnBlUkF3TsOrh43ir7m4pduiUAMSLfkfcFKRhXu4EPUYgP+yFvdWNTtkAFLu842cg7j
/n/tNHyyWwkqjy1JUDoaisU541/r/PD2FHkjzKR9A3ot7I3Ah7jjY+qgWy45vzeqnCy81RJwjrAG
jrtlugs+1HwKh7qqVhvt4hqXFor8jK56IJHN60qCWpg0m4aC3BrAqkdIthsnjGsZmRr/PmwjbZnU
/4EEgyPWBVIpvJQpJqRYjeSnAk7HcWbFW/6mW8mNrxptl1VOfVmbFJdunm9h8Qhc3Aw4zNA4sJJ+
VuFC5Mw30vaQ0zbWnZlCQe8PUnae93nFDm/TjhUmok8KciA3KpoXgTV1DVA3R+copi0WCJnTXIT9
/4KI/RqF/9kGm+6quDmo1UUYz8oN38MWq/elizHNWjfHYQ1M6YuWjaegoLduhsixogdB+Xgs75AS
Fjo+bZ2Om1/XIK4ZNMsv+LDEh687OImm+6qxhgFF8Ov6A0UUD8nw4kmenB/TMmYigEhbLSSMVRvv
3nfQmbKYgAJQEXmKrOnsS3GInY/yLgvD1BMPRPEeurefC2WqTmFsWC/sDMZk84t3qdr8hUZlULlN
Q4JnCbNiW4IHowMTI2w42vYd/7v1+0i6XO/coHVPcWJ7GvGyQaQFiDLqsydxZ8VWXXR9yeUtlqTc
U3NV4WCzk4fEq8JCIND0sjO2ti5wxBQhsLINp0km3EZHsD+irzXZNT4jzSwmEpnbzbSymgrGJ9qE
A92IxzNSsgnAYxW1Ibx0rHxAyNT/oe3CnC9324tjqLpbdjQI9LSrEahphgIIvD7yIx/YciZmpIVJ
ZjE3+ZDbxL8mveyI12Ltcq+XVg2zE+l6rjmoVrMDiLsgJusK9iTcUFcAssuwJ3xfEdcvLwz/H8gd
JaXVs4HDH46A0CRaVBqTfYyEBFgfE2gnEnIapb7S7iIeac8/JuQkLLLn6wQxmF7ZsP0Tdvwu/Rqs
Rfx7cod/PkQTAZUljgM+bCXhYQjVnPaSW2G+cEb/k9ljrhciHJoM8Rrp7c0fKu5TWH78jtail+cE
OkJk75ZhZgLvf57885Op/FIhSis8CrdCT2HDRCPSMDq3KMrxKI3FhUH8g2z92Q3w+dy1YQKAxk8e
nR6wa01qkWT3j9S1PKO+k0jHyJv4+DCu9C8vZg9PeSj78prYwT7dvOth6zP+AG3tBu3w1TTIUL69
+hOygEszq3MFxNRDYkbrvbmYoDDsRkjlX49Mwe4MeDaLBoupAdKHLb2E30KzCbYYLy2ivbXGoDt+
7PDHJ7MHxMbWWL3Tx9R7QcCCHrK8QJi/r3W8RUr0DLrfxgsiR3bAs9w2MjsZsGUx7gxvM6O45l/v
dHHSmT6V9zrXBS8Urf5elgkF2MdYVkdU6NICXGpBwSfzvrtL4H7l1o2PciYCIgrJwSWVogn/7LWK
2CEInhQ1j7wFTkqwWJeUmhyHoJVSfWtiMFBWboQfGxds1S/oW8tKaSQMEecsih4f3ndlBNq88TqA
02w88ru2wbcxEQLpu0z0RtyHLskk+nzrsHqSxhJZamvpvqekqCiTYbtGuActXTCxWNC/9SiZ5VAn
fyUrwE/oqR5MHhXJdCRa/Z2EUvA8K3X/v2Hy3SVTVh4Zd/2UUjCqwlJih4sCYlIbARy5osus7npm
62V0qux5JySXtiVnY4O8LsMWUADs5SewuW4Am3W0tbpUJydZG/Q1SsmarG4EoJfbCwtZ/5wOxQgI
jWLeD3o5ViugW7e+/S1k9rsVkGbmvOAB0Im388s2juEH0ZRqqOVoeElvRL0btp8CWM8yv0H/f9DS
bM1/zQcbFEE24XXbK0aQRt9KFe7GUje62zwbaZRktqa0jeGFt82hweiJb/NFq9W2nxXrtJE+NH03
18+nrHGc/A/eTXrgaUEbi32wMlsBDqJ3JDs3s0q/S+sXZexTCW6YWFa871S4xzsmV/Q9JK08TVJ8
Ua7/YdXe38kISLTMz7AmrM6pBhMZxSwZdcuMcE62gExgNgSihDnAgFUQXFryFTV0+j9NU5LphmOO
oxbOopT0Uy/KLiQVt9ll8WLQyyCQ7JlG8efwTLDClSxyQtOspNLp8CZn/w+H/ironJVW7MWx2JBl
Nt2vXXKpNKQkXHLWGTf0r2S2gVdqoXI6flMziu5UXe40S6bo9grP/WRQDBLMsxpXmVW+GckwLQ+P
IFGEe2ax5v/mMYcc9cuywlhxxjB+bTgDjfSgCTVQqFTofdG1A1P0pen4XL31mRajdk3PhIXtwteT
6zgBPHZ0lnap0Tw2bvH2w6I16YnSBp+Oc2g3UFIJrqy19jLisXCMfRNOCodjHkBycL7YRbHmfWya
91VSkRhD9tleteH4yeNSVhicY6tJGWmr0miMfe0aj9L3Qx0U1IrK73inyJHCkVhdC5V+ZWYWkd5V
au9i0l6BT5TivSJWJJEPUaKObiIy8wUIT+Sa3Pgn34yEvACPkSt7xDus4qwCFA+Yv/6kqoOjz7rH
j3WH/OjSlVKN9MY1VQVRuabmCEk+zTcHhvi4oPMA2gtAEKdENHtyyxe77HUTGl6ZVdh6sN/zaYeI
pGWxqzCbZdW8sQxxTBL6DKQv6pDFpQ5o+KLeXLFIN4+B8XbDVJOZKyKR8j0s4KJ/t81Ds0x9xYBP
8K07tDWnMSQvzdrvoDMDwFHbxi6doPq1zjrcngh//Jbfbqnb6ak1rvbgCcQf2MAEPx1Et0GpLJW/
sdwFr3BEzWw2jgPAlLd4WFvxlvvx2ZTM6YV64o+8cqtCpSvq6gF1e742KmgFRhQOg556tYKLbM56
LbpZpsE8hKD302oaRSltQj08OdQ6ffp8GyAc2bK3ZOUdlsVWyd8Ei3bETKHzL8LXO7gL948yTcY5
qJA4c+H3YZMlQyOEVP1NrMBAbOtKFIcMAunSnr18d+M76H3mVRF8Sk6b3W51Ixk57aRBJBmkdVnQ
bgjjpm0HBIAer0QvnzyI+x7NS6sLmr/0QKOh3RT1WLYraJKyVdj19exUnn5XpXZcKFl3kHNhEnk0
Jocxu3HQ9UmPWMAlFVT/PpwdrwrpL/PxFS3x53Qmmdy5Se1ncUAHvPVckw1DbJdifL0HPAkhFGo5
91fAcLzKTnWeYl3r1JrBs99uigC2ZA4lB7E5rGlWvq2N5gqXndM+GRd7l3yh5ZRpWI3+5xVXlK47
Ai+voQgcFTaC9NchYxzOcSx+TfJLTgRQ8o3SLPdvOngv095MLJzRedsF1V5fQeXgAaVCg7K7Tawy
WJPTtx8+i7F6EKKYchu9nQcZMRfuANtQjwd5DOJ1FG2qvLc/6H/Saflisqpsj+DMhDqLZBIaEz/+
pR/2ZT5tKtzhNpJkZiD241y6uF270fn91ypKDJTC0kdgTA+ZGQlunPbVc/Y3u8Vo70/BpyhzQFz6
IQ+4t39yX0SHfVNdWntIzP6GdZYLxqlVsUWUdZh5X4dRdX4BdNhZfTyVmOw8KFvSAj7P0kJLtcaY
sHP8QtieXicluJB9x3ih304EU9Jr7oNZEbGjNNT1uvUS4VxfY93gcEFNvEsPbzFmzjqQs+CJIhm3
MBDYfu2q6awFlZV0n+ibHnI/rMPBP1Oyxgq+0K3T4EULUsxoFSpBd4QLfvhR67/8kFl1kmQYtTS8
5Ig0Kxv8vzxC+7FbUPXxc+/FSjalLD2qlBA/XVBcsEVU/CBpjqW0VTBGMkrdnNXxuYkp8YAoUb1L
cPE74SeNqJuNmZ9urG2Sdi5asfFs/7GRuD/tHLRpYyzWwFB67jBPEB3Udeb6Loi7EKW0tubvaca5
yDXSd1cX2/cdpHb48igo3EAQQwsH7V8MvWwsputk8eMql7TLqPnTLXpVPMHA3gBtoN6CJ/ibKVvh
wee1DINswjRjKYUkbGXKWaS4pe3iG1Zx12TlJwZwvP6Pf5Sbh1tDgGccI7bSjJ6OwglTamK/cQkf
R6P8yHkz3I0awEn1osnaE+wM4/VYJpSoBMaUY+C6nuQJDVPSPHndw9pkQw6yjTRSMvnMx+1Mk1GB
ixOCB9s+5cJakQeNRIoj1TyGYG+eq0+hecyhNUT7BJoRWsWqkip8e/i3P7Xx3ohXRBn80a3zzoSE
fu/YVwcRtUW4e6lRH7ULN48t2uCN4kJJ8KeQOjZNguBGezCP2m9VHXC2RdSIsKdut47+tpd/xfeu
t0EpDpXIoV5QHkE/QB6SLy/EQ3/O8WL0PZo4/e+P6XHO4u8MQXDixr8PTXbOZlnUTVTcIqc8QtRR
mMO0JSyERbMFnC0vpwnyioTXKrUMseDa7sg5OzjpIZzvHd2IHlBiBdlhlUv29gOkCk0azEB+BS9w
3ykc/Q7XY2pwho3mxm5OcAeCWIYDl6kKKSVeqPFWACtnJu4rc+fEAIos5NL3san97IBAJ3Dkkera
J83Q2Lov1KD6Vr4fy9SuLoTDZaFTCm/qKqBqy5Pvi1pw1pSeFn3yI/wl2jJohDIbY0ROpKjuYRdZ
BtjiNI5K9WmwD12EWDqXF+BGDKN266J9LKiZvX55iRL2GS0SfatfEbhbIcRqYQOojtwpH5YIpe8n
RcSyMMEfrHVg17QBg/18LSd9MUv6TbJngGW7MyVpCAjQZg/RRnAVfKDaU99ODvTGdX8Nl0EQhnns
FMBB2QISia4iHlSEmEXdxq6jHYdz+3mStBQTQ2nDFSeO952yNb1vw9vZ1phEFz4mgTNGuVDuYr9A
2ZCt+wl1nQzW64TVKLCszDkltCJ6t5cSDvP3O79pguUiS9rmnafpq8TJZxwCYs2gZNlocjWIqB5V
ziyYQOYhj4xd7w90r6WasrNu00uy+Wc0V67JkhygpX9iI8UpRP9l3i/M1meR1UQ400ScKaCkUABr
KSWhabYET7npP3VysKzkL4T+qlQZDkwvo3hsu7pitzQdVuHui4Y1gNdCXmwmRvO5iRgnAIMg0PVD
mnnkG27eo3dXoMBWajZE8BIoORmi84jnQ8ZFJQrKkJOWgbNYrCB5wx7uZppHqZFz1j12RivfKO2y
cRBXA8e/FOk2ZWbWkU3GGJZThGn/3xSbpWsihP9NiZdyPb9vVKQM9UxHTMTvasK7eUdjCQ/uYE9H
17DAX/dYSid5ItktPYp2jJPL7sv/SF874UYmxfw2UoE63r3eKkILkBpI3O/knDKo19thjvaWk7ev
zpPfAoJPJ0Posv5X7Kj5uWzb/mSH35CtgCuGX4JtoVDfhJg2/rXlozrib2jg22lIV7rrymMgWRFr
jxhXOI0Nd/LjYlsgAE+fkTqeVz9qBFhOzuW7OWSt0at+6zMzFK5QflqZT8HXgMJ5C7sG4fYnVfzL
zHtg40ADWCHUUtHqNPIAnjMoVF23sVpqWWvVVtycF2JuPTrWZ1SItZS28rei448NNGxH2Vd5B1k6
7a+6v1FubxFtkqwT4Jw4+Rzde20F4N4SqjUMfDAQIyIpAXI31MBTcM4WOzUStcI7oM1DcKvfuqWV
aCGulIEVYwUBGJBHxPmJNcumTid+VfYO0+aMoc//0UOnDqgYoywkuZxlnWGFTc/GD0RDER1N2Rv5
xqivVGzYTyTzchztpwWy5q4P9l3MUSweFevaVRUDRTZrVu9HN4boGUT9hfAfmHfbOGz40/Al2vXj
plYl+qtPXHuG9kznCRg5Q6a0qOzzbdc4Zw30aRoXClQzOF/mpNLG5IeRDUoi+Les6ix0bj7f6Rby
VX4CxWkm//b/YoLslTFZcpvMTgiVnMnI4K6rGJ3rXI5rFmtet6OEvQag/oCtKQ/ISHraQt3ve5X9
/fSv+4u4K6sSnd70Xo+LvHtlmwaNfJwiKztA5etPEAO5Tx61iNSLeHQKpltRfvOn9WqIAW91DCXz
iiNcfZm8mUzuhmBe2vxA1GMzuoFswNd0r+Owz97coWUuCulaELRqm/xYP/eU3Fs1eLEOJkRz5I5F
mkzMVfy4ndb3QyTeGIeNlIhMCpfomfGtyYSC0hGnv70eqnKnz+XVR6ZUgENbFNvn4l9t9/9ZCSp/
20siMAJfrR/01HRQF0cfn46pzp5BYQ3Qks33i7TuFYx1gCZAStSjk3aQGzcMwflWEmnNjS9KOnbL
5VRYiF/nPQcj9Af+hJsW21xuRmkMZ1sFcFieaXXRCtBT9xv2Ux96eCou58UzAUOJYptd6Xe9XDyn
hoL1fC8ufQICOfdb3Rt0Ovp9nGVfeJ802wmECWTvNy8FvYxDRnhd6wDQ5nRhSyeQA9JY83GlaAEz
qoi+UJLqqIOO0MYSEv3F+9VUkh697jeZyQQuj4TKj5HEDHtyLbzW9hfEicKppCGSRWzmzok2PK9s
dZO88V2DWGb1fwR31BlJScUirMq+8zu9b6v57rpuhq2con5chUO9VhPPx8OdxFKmcGWFlsOPpSok
UoX25K3o4zk4wIgMCQwDhVaJFgEvJRwIcjkql4FPonTX+JQTfSzAZ1E9R7z86dEtN6XeIXOaWsSA
7giE2C64BE0xg7hTTmEvvBmq0YcqS0Abhm6GrXzBScVWhtdhwpzIhJHjuMCeihSh8+LlxEzDti0u
XIyy3lfTUix5dWD/5Uhj7qcfn15x6I/Etom+lPlEhXFI/tvQyfHCwkQfZir5Zu9jG08kaweRNc9K
K/bUZ5y9+O+bszovAAcueq9FCHfzw4B9wi82BYfI+di9apP3sa9WYBjGTyl5g8DtP4YrsLf1kQE5
IV0aLgkXi9zDS9xOr2y32t9BE2+9y1zf2lGsqDef51FnRd98GHb0Mx/pRZYbaJz5WS1q1i/jUwev
lNt/CbzvFwcd5E8QFN2y+WklpUV7ZepmTMLcM1qM7uA5xZzyJaWoP8HY95hRTY1A0SLigjoakyIL
b8ggcecx9bmkbgwRycVM7WDHmWQwCJA5bvWq2cl5JfOcCyoUCiBamheE0Z5TJhPgKDpwqprvzV9w
ZirfD3aB1tJnsI4e2+5gP4yak2YhActP4UkK6FotnoANp1pwnpelhCXmdV/oqUSYDXV/+DjekoNY
J+xaqoV7ND5bbikI1tIa5FVNRgCO0Z2cEiRqzSKt+JewvjgpjnSxedaB5IgSAYBYgp6w/h5rrMM8
UtvLbu9T6cyFP0LXw8iPudXcXZ+96yhPVpO3tZQmlSGLunq0c1l6VGbcGmjwSI8605UIvyFsh3jt
Bxm3xQc4TdBLTxB5XZszqybuPOxv/EIQ001zmceV0NKqGb9t2Xd/BPVWUg1U3aLCcpTo/xAgxp71
2YywSJdpL/YBMS2u8frpntKm1Dwuj4MH3PDLOW9OVOGT+QOyCj9OOIn8d4CJm3CEVAlYmzevuZrK
Fj5Qe3zwEGYYcLLIHwlfyaom5gQWVbn3YCHKvGUmJ1t00iW7Gzp5aVi7Ps1Ul+4iRi9Y1wRBY2CW
TC/1YB2TlHK35fIFCSOU66oyC04JULfbvSIOhSCtRYTJ2K+v+FSP4ddPAC2UpmGj9M4GWkAV//94
ss2Krmer6wxYIeltZQDrJeVFh6Exeq50McTtb3OeHzMLxC+w5VtkjfLWo4LB9C5OBxxXy02x7yJO
SFUyCYPTVhIIMXphLrEu/+cDIrCGjumgoTViRtAb7mJZhQMENSln+FGx6YNFPZlwQiH5wBUa31e0
qF+dK5KQAoppCsgKEeK/11qUMsVP1wGktb/oq9P7aEt2vIFHL0JcYDSxZig3ekQ8yFq8lK2BtldV
RB8BJJHDhfJ+2XsnY81crhHEWojgZWnpuJ26iCF9lZl1fKe4K2iUNe+z09toXsypgEnaBzxmzsLr
k0+ZXz1hC4TZpvhECQ3Ak0BSJZfeLJTaAHKvs/BHXFCR0J6NYVitv2qu0NppO6S38LRpuxQzRAgT
5fK5AErZ1AhFFaALUZMZw5KHn7SASBVjuzAVKj4xK+7s0l8p/wFs5MfgnJpD7c/ZZvKm4WGuryo3
55Rxm/oqsiH9bUrCJiMYfTiwP82fCLuOffW77c3E+laPBff1x70MvD+G2PuN2RCa3kO5TV5ZoiCw
cEcro2aOdPvnw/35+mz2en/+iva94Ip19FlbGE8gncf2jr/ud49RFcwi5ar9QmmfyOUvIufMZm/b
pXYL2bxIv07X0yBBfbr0h8P3EoHzXJf8l1Th1nSdkT8RS6lIe/I3DbKorQeBLT5HP5jdCKE/AEXM
haM5cYz8TCHMSKRgR3QByGV8RU9aWlkwRH84ITky9guCfTfmVLEVfL/ewWWZRjZYPzQ5qSQg1RCi
2KeRLNKp1GoUM5ygtS9X4LlYZZV/HpPE89gwKURIeEnduZwsWDWNrucnSN83Jd4fl3AJY3L+H1df
5fXcy6Bo7QHbf4OfnTuhdZTLZlvJoaDib57rwOvlX4A9Lhaxp7De7u1coElkMNvTifKY6cC/Bkcb
fmeUycKwAVvItC+OSpX86jD0mfElW5VibkyDJzQvlOEDW5/vO9qGu0UmUHBorlSk1idz840lWthA
xjCrARaWlPts26UfzjNEsqJVW6v7pO9F3hv143Z/HLBAzRCC6YE8HpatzMed6JmINbLv1KwHH5bo
twIVtA5x+tfxCLXjs4d1C/5SNLdK1Uui+WWGUpDda1NQL0TbUT/RYLcB0jGizabZzEtHoyNP97a+
iBEKHv0tkxusiPqHy+tl9MqYNqC8yya49o0RBz0duA4iLzZhuVrF7U7eUwlJYJSkg9tVDdyYC9yX
2kTCzzMsu9U3Ufoy4Gd2HNnRbVBzodqgkXGyjGuhl085NXeURUOzlHc80Jwe3r0o6Q2JbY+XXBcZ
GexMLWLBvztFrKzxI3v4itN/lmR/r0UG/hx7zzcv9Cwh96G9IC4yGsUQbOy63vIIq7nM5cQm4vs3
+YbEW9gz6vD7Iub1prCXz6tzxrY7BzV3oflIsIAKjwksNtx+Jb15Bwo1WFtG8atn9xu3F5MB8zRc
q78sxYP95UZGfevsMTMIuOmVxXHfy8PnXVa19skn8hUXb2d722O3nLVm1MJBoICNgigE0d1qrm3D
uO82eQnjvuNZeCodb1iMmQrulLNTBAfwh0yOmmv/xGw7/EcM61QwlPW4iIRAon+/SnJKiJmW1vTN
cFgFBOWMszs6d1S6MARqujUGM1YUgsHSB749zdIfEYc5Ir8XWnWzybG3fojHZJWqFrrY4bJwT9JZ
7oXHGOf55NiLmjSdkrhx0f5gslXiZj82YKbvifWx1SfulJiX+PSoTfHLMf8AemwMugl8pnmhX3gT
Z1nQbwzC5U0m2F5mGhqDA/4QQSf/zZ7VsmJOYNEATY5o68lWdo3DmgWSNh3funX36tczUWsagd8/
uRpvy/LVmAG+ZiZIjlx7U+XPmFAbnvb8GVVkx1y4iu6XJYSkCAMR80UkP/eCO+o08dkh99I251sq
CGCEx5tGZU6b+XVaxgIe7Oi2usohmwtQbNmG3NEzmxrh+3vz+IlvgdzQRCSMpUTp66QuurxbvNU/
u7QsPG+WyPJ9SzRktzrFj/sx8yPka39JyLNyJTkgKQuL+dAe4P0yAh6R3Ih7YhamTkS7qtNcVV56
I4ZcBQwuDEJkKSuze+ygMULNM1cTHDdh4K9jqp5TCD5SIxJDb/IN41gBpij4eZCyHWI2snU9fMAu
Am5rTUwwn7WSUk1C7ID+KfjS5jYW8AF2QKw5UbsVJoA6sEZHmy8XMUMt8TXUUylz59M3IvBRSsmJ
z6PjeV6UGtDWA4ggqh3YCr1WvwPWrdlG4EG2rmYPy/kwOFyW7x9v/y63Dfk0jGMs3Ib5gkfj+sHf
02WJKOsrqlNiB0e08N/DMMnZJfEJ0HburWkU79JhCl4znIJBNm/4JOzJ8ZhHizcQlQYpX41RPWGI
fz3covYFeIlxBRxKNMfVFWRMTvhZT1Bz8aiG3FvWgMOBUQu4ut6Snw2mEKC3FHUGHXd6Fi2hnBGQ
zSgyGeLshHMZg/bpKKaMYFichscWCXjHijK4UYvPZZMEbtZ2YmA4zvEzOHzzTlGyf4ioc4xlQ3Fs
pyGtxUJtSwJr792J0rK4wwiWE7NoRJuSvDapQCyNjLr5q/QwOudj9/y++LmP/TaVk44Wv4QvYd1U
7TO81PcIuw/oYFToFg3j1xk5neiyJZWBQNYsp0bEII9FoCSfv9+VGQ5f8ri4KHKO7fvV7DdBlBCP
x8OGx22744T2B9IgbjZs7XvZ6xx574Cknv6q0qa6K29F/coOqw80qYH0zG6cQl51vtYhmaLRm69G
8ta8fjegL6h8wKE+k+EXozMqNPLmpcEPDKaIzfHHLU0jhc72BrlAgY87o2KyqiMd3t/wO9HS7JMC
GkLdNc9o5lZrBlcX4pJrY8C4UU6BOl5qIh89t9YHmO+lURh11JSxZN9ML90wjx6e1PKHa3ELysA6
NRTvknexbcFgZsV/BYC3NwFgFBwzW5FhDQMKkM0U9qGcuVPDxiR11pEQ4eh7kJ0/KENnncsyNY68
E9ke1Vff1DA2AelnvyhngV3AS8XT6/IAht2Fh+xc28wIf+chn0ppineSdTGCM4tYvsPess8yES3+
VHN9toF8pY8XnsDiIfrL/+OJcVlDARXe17fv2+Iof9w+T/j/HuJ11DsnkIttHWUfmeiRt/9ndKnA
cNsABPJUM3DFdRcGIGFXksMe74sbvXciw4B47UU3Cs+Z+Xv5FMHv7vYla0XRPTMWtZ8Db7HA9RAy
xUtPZ2vVFt/iOLF5712qCksUvGixUk7KUYrIkeUpF2KSxjZKbk4a3jNDpMivfa0nyQ+P3eddQlIf
kcQ1k9Nl1AAcGT6JSpJ0GOorzuT+xdhhzdGLVgvkepB5bAfcHY76DJje1RPAMZmy5I7Pdzz4+2ON
o+fs1wuwBdkZO3D1NIoW7O6pPXGXZ5wQyQ3KVma8DYteeD58Lq6eT/pPfFUQkOMJPVlFWFGlLwLo
+GCp5zjf49Dsw+be8A6wUhdKXB7jm8kI6j1jJXhseS1NjXfz9eDR9yC4GM0UPXQLzzAkAlGKLS/Y
Li1jLlG+vazsK8+KMfjZ+m2fwQPBaVKeDV6x8Dh5lO/NDjC3/G0Kq7fybTwspWtWrrESxTh2tF8n
rqDaqN0vyzBOY7qEYBi7b6Ff15IR7RH+mydWpWOKa90BB/6heAGGZ9NP0XTrLRWTkJFwor+ccjLG
/1z06zcO9smOgKqn5mdg2q9wKQbf7DSCcmqdlB+q2HK/j2qPaOuT0vCzfeSAJMuwWQkGLaPZ0kJG
uPRdyhFaYrxS3/2GZTbSz7TlPHV2IAN3m6qVmRoIQBs4kleJAB4dcqB2j+ngDXtjL5gy6Tgzc1qy
dxUa0DUMK2EfsSA+TxMx9ub24ko+flwsat+wUT2ZN3EoxcQdJp2PVUjRYRIu9qCrMzJ2c4uWiplf
OIKGgkXxZ/dPpfEaKJdlSMyucz4BJgAJRB+swHwvOfwyK2XLP0QYAeoQMW8CSStUYW6e09KRqVsj
SNNkai6oD6Kpzk9afc0iisz5C8dZaG5sGTU++XAvkd2UNOIMZMl15MK5vg/DLfgUzQrXKGQp0txx
MFudG2PIMVFW0RhqcP0rcoPXa2+hWbRw7z003ZfYJI6pUFzlTZ3UG8tZMtadj9diOpVRUiLJLPNr
S4zKPXvy+PustKqy2IoHkESN8kO32N4016qxbTaPRtkXOHwJVbJySeXXWlYT1eooPeecQlg30eEU
2AdNZ+N2iQVpynBu1Oh5J25AL+vqX6rORI+hQHqH4U8og8vxowK1xF7k7sYQ1yypRlAEehUFYLjV
c9makZy72TFqFw93M3IOuPqn/D4TMyYiKatHPTSY7ZU9f/AGJJO/TdgCIsRst9HzyzCHiCXKGKr/
hDjWPzojw7Bmy1LhJtHybkE5xu8ejd3QV2wwcL/A8NV/FxP3bJmQEludGRXwCXI6FejO2zqagcrT
qE5zP6ugP/RSrBEoOQRB1Dd9OsYEWJKuS7TfTBGgkdlb13RCAxD65FL+AQoXKQuNNrRkkP6M/jpP
1gdJcjaBJOS7z3ATc2DWhBWxFPQ3aoE6ZJe5/ucn6L3qaMJLXskET2vF/GqIL+kZCZNx/aTU8Sbi
xB1PtnVxvL0ivV/yJ/vTGt+ddY3mFo+XNizU4j4c7QwnHLKU9ICiX5pntYx24rekX2v3DplSOmn4
NdqwV/QPYgdx2ZYiQXgCLLDItIS1g6Lpw2/U6a6DqH/du7RRRmR4spDqw1PVY7tO/k0jvkbRvovP
3uKL/JrY9SX5AuFSS94d6u+KANsujS1x3BxTIvBSd0qd0l3QkZdBe8djwTApxWGO4XBr7XCi9s/d
rYFnHbwXpfEfWAprcRhzUUksUoEaJEDEyo4iMrrvRtuE5lVfrHgtaMLlGcCvWXu/OGbg0Y1rg+iT
6e3kPCh/9LyNlfEzvaKbphxCACD1EPcF6wV5r9ecRaNJ8StGQxzm/dygNLCKq/uI9MZ0OKt9vRCL
mN830urMoRYGv/sqeA1c1xTWSXrlLrrcBj32jwW6VymBGCkRkSoUQM+15oFscdoqFpYswCbFqZZM
GyL0ahPB0/S+tczyjXwtzm5tEsvmxSR7c03WBvGDhsJifyFkQ0G6WF1SvZpbgzk61d1eMR0v2TPW
iRYdEL7yZ7G1ECOjXRMamhatA3NDxTuX7ARZPfwz4xbdzhjrPpWpDFHgTbrzlMsKqoufLvpYYOqA
h0l//dtj44wpuMRNEHLHh/97SAiZQIT6FAdJGhf7rTeDJI5KjTri6n8Sr2m7e0D77NQtnNjz5teI
2oFYU5c2UIjT9WGIb6Rv6CdSzESJHbAbDXA8KhtxXiQv51g0I/lZql6oby39ogqjT4N2muzua2jq
pSFNx+Z/CALRl0plMXn8JONUkw+oDs/+EY8ddDH/CHUxsATuYg+q6K9jlLj5lnzQiK/W6MZm88OO
eHF+M703CyYubND6Okddt3JOGzMlOUl1xONU1ZvD81sfPKkb3sC6ectUYR+q9Dtf17+K1/X9ZZh6
FmB3WieUrpYL2vCGNok6uCYJEU2nZxQIh7UkLMvTvSFWI/HpvrDNbdrKkZgqfrj7H4Af5LzaZVPN
clIptNDN0GaIgALMlrD+xCmndIjM+gYRoROU1U9lVWdWkWJSRxwrrwj7NNmDj77QiXmgP7hnt8Sx
OnS1XFwJ8XT+Ym6QxCQs7rNH0EkFyKQVBIKike15viB7RWGwE/pprokTy6eU9gqSJwNYywW4YxoN
3cFcX3ollVaLI39+VBRAIi0AfyFbdh60urUT/uvCiJZ7Z5UFDecJ1g5Z7PjYWUQpqygwwqlwhTwx
OyKrKTeg3dk2dSHst8kn09D3oD88CGZrN5ckjc4lLJBnV6eZ6FW1f/OWaTeax0NAPauCUHyiz49h
Wrbi619bS+XtC6JW75HNJ3ufKmdlSgB18CR2j5Ej8Jpy7z3STAgzERiLmZNBkUImkkl9+V8KQTMN
l4gSwTX4f3eI0c8veTWNhfry6iXjPxEQmwcAawUmoJPtXi5qTlSYeTdCoh+wp1ENK8xzQbjBwFVS
MER8XT28WP7y/Lk0nrRAfhjiP7or6P7jAlHPgFd72sL2OXoWsEdV/Exwg3KIJsEflZhnqgnkw3Wo
u3Qxx1+S2lWbCyxr4ywLVMyActs3qFpJ716fNyljA6HD8dkR09UGc0dbFqgAJ/k4a2zesRrsnqf1
zQLjbgrfSBnKBZvyehyPH6qgSBsWM2tJEkvpJJeu0FyCmrT5/NANB9J0rZpV/GnBhzVYiFW7/mBM
TldNfTUVhBr7S5qXu7NBO9SChQvpsj5DuxqN90cHyJ1QV+TS6lJ3ShPPBmxl3uLHcd8p6e+NcKSa
WM5MTa2bERYU9d8eiZl7TDq/P5NUNLL8LFUjOh9DH503p1Ym09en7wfkJH9YEwKRDHQoUpCVq8BX
I9tnTYYvb1+JP+zXOk0KVwLzwiCSi00gR7rWbvQdH8yCjFKneaXnO5DnZ8UlJkjrsuUuXjqd5pqK
W/kYaKe4OLo+LV1yRT4ZCFWomDiowUvJtgYGto9hWm8675H80qdyKFW8gBnAo03SklR2Za5frE2p
QpKA5m3kXnD69Ru0hsAwNZgvMEPv8VgTp3HQvxZEBPGgOHvcKJQytQzJ1R1lphIpGKlYSChji/8P
DEaVAFm2L0M97xFz9CZFiK4brj32K8MTZhQUSIirWpW7oNFkcb5yvZKYCLbE22Qv7ytOBgl7/eFR
uSpprMifxwp+iseccmvAoVaT8u6fQbhym+D0ptupkFkao2zLfhp56RB1ABAVsnPwrUlSPcysozh7
jvE2V/Rml1PWGbL7jSotENcYtZInqywl3wecjOPLHzdM1Gxdx600urggq4J/2yQhpvD1Es3PfvNl
/m+nWS3vcE3DeskGcG0K0ICzI2ptm9HOaTxpw3p5+hOvFLWTkTuGSKzZIaOkmL5jvyY0DOOKhZor
iwdm1VAUtfhDq9wSgXg+eyIbFHaL7TRlJ1lltha/fZwmBPlARy1T3baEXn/4tmZPxYwmTjx7uuhG
FVn71tu1qfL+8AhXPU847EJxDoJwuZEGevr9lD7b+opW4ArOQcX6kuAOyZalqNUoc+UmU0jyJdvv
q773HNUvrEflJlYrKSwMJ0Pf6QtkOBFJMKv3M+O3He766V5DiLWVavMuHVyGCP1aIrelmrqCKV1P
mm/Z09UrEZMYFZDkRcSM7iRywiPHujwcSfSSISTfcG6E6yBBNG733UGdggABA9wNco9ErkwSdDIy
VliNNgikqu07ZS6T6DLp0cWI6y0kEdhJiVmvBoCRD3l/TMYUqvQzkf7vrtUuKh6aG3dfMMx/Izcj
DXQDfVcn25xkveg3ec8Rb1TXZV2mQUL+MDr7mNbLBMQiv7hfQu/IoQCBUlsveRpXZpb5Q0Ggeyff
OB3h202Ksab/NXzfs2Jx6spQSniYBIvIblIUmgI04kD3m7nPcAQ/J0zbko+9vm4WD0rf+/Enzw4N
uLIB4eZR5D2vrUjiY/MZK6togNwyK9yDvy/Ke6My59SfBryL0mighGLH0pQ80DrSTM/p2IW6TN6q
2ytbeGZY16a1fxhPvNs/YkfiNB5p0mE90l91DeBMzWO8PKLRMRMc1hVqJku9ahCMs+4UPt4mFMRb
c78yYTCfvqX+fJZI46DQZgqcjzfe4PFbd7Bb+m/F01DtN9knvJ8P7TPMRMxr+XslO5BvHUckvLky
ALa9sq0DYP8nUH2OQ+ZqjOKg4FiyxukvCjPfAQhZ80Qc/acYbHzSrgu/uWBP7JB6Ss97u11eKw6f
WZ+N1p+ScfN22M8BuFeH5TjOEGoqFN/u7x3+RmqN331h6ZaVttwIBeT3M+67cpwUc5MX8Pe1zcq7
jqAUIDYFhGe9cb99Ps3qBIf3nH7AtBsN9CuuNI37gbE/mLGH/he+rW4PwJ8owX3b72T21QGcEXwa
0P63TnX4OrLANRNeYC8kgT7GJW5EpYQP7j6kPctFiPBqPi3/6vh42kUcRU3jtErPEUEwBUnqrlsK
5e1hUcRK0kGk0GmSZ7KbL/9xC7miYlLvfQibjQCoNPOWrFwG6+ujrKh2mKfgjqSERA5I1iT+Xx+X
6RBpSrm/jLHS2Y1O3tvnJlVRh1fCQqL0f+iTcu1ViSYeCsJBpBb7nxQa3U8iQbVmXno04AQWjcGi
16BL292RxuUkJMC2oNVaRdq2vs+ZmTpwosX7YDo+a+okgMdfCt5gnDl1F/gbVE0Bnh0u85I6G/SK
RNHH439jsdtZxdg6kWnUfhSE2uIy6SX16GoavYNycagO15pXxptzZhSyQcobsXCL8tZlVpYCCCKn
eGTPsru4RqSh0Mgx1ow2YlEunakEnOH69g56gL8pc1nsfWRKgLCNGLAdDi/nGvn/Ac+9CgeiqCOR
4XbBhN5zWJJBxCFkTldEVDtHxgzDvqNZloOzAPT6WkXozdh1hnLVAuusDlJ6q2oY6Ws5V1FfvMAT
AeZ2LTlayLYAXJO4Tbj39NTsIdiBuKx+PFNShpcdoG70yaNYFbLr4DLS5yuV2SZgi+6mJblLmq62
+gzwCmi3gxhmH1DJ27SW737DBMwMvFysL5c9KQyKlr8v2QnHxNpNooE7P6Sgpek9nnhLek3wwz4c
RUnPfIfvG/XMHI9RROD1fi9nkkcCsb0xWu0haruG7pPEhFcnAXjdWn7qi+nqQm88YRenDz6iLdxE
s6ZpamVmaZ5Q5Qq1/YoUSnLit894U9MslXsCJ/IcTBDzUSxvdxE5FKiqVwqo8t2PJjbYMMFvvYD3
gJ5wLsUFYxmhytyp2Kp5dizJ7xMpKMioxtr/aA3qCECg+tDe56yimFOokdTHS8mcyVzKw8TzKrlr
ziDWss9NflO5CX0ubAhUBaKZP1hlN/0Dz1st8O7s64vlbGNCG3MMk7Ut6cPuBBOHpW1pXc/FwBph
IR2LRJ4mBcfL6Z7NAzRDiRIHtOK0nwglEuyVf7a/pWDGx34FHl+92hzQhlPWhV019myM/16SsWR+
taceKYziuCHslIwAcfUHZjpWE70jj6Imz/x82RDUoPYUhRT6q7BC3tRvOBzVdmKsMXe9vqIyZDqx
+9YPwjO7HGk1/ghq+uHqcAkbGbkVYpaGgbwj2Dum1iPCi43RjUzONORB4T+Zdv14R7g4ZqXDG4fd
3E841E6cBbAjLeeYC5j1L3TQhHK692+EPYHInGlG4ZlJR06nb4NKHYRYMM4WwFI69BBEI0kVjLbu
1dMZmv6FXRCdnael1XmvuWe85Ra9EBW8D0e39phmxOrNiD3/ezeJFh1GxETnDgCz3KTVc+O82wfR
EmXNM1qPhVKMsj2RQ7635DsjsHU6K4XiEFYmyrC1VM0YDAno0aj8P6M95/xIMK53wkh3Ji3jh2kV
FHRlVs2LxCpHpFw3E+9kE1bTBfDtP/M0JicWh5gFQVx3CnRfwQezbFhs+7Vz5p7LL+EKuFW7nMva
L6pfYefnxH0fSOMyW78O5hIwdZ4gUhf3QE1WBUPa24rH7bGxq0cy3TQdRxKJ81C4hl2pvy3v0E8l
+DuJQd5fPVwAHmL+smTmDzGC3zOrnDMd0Srw0bfjQOaNwXRpOiUKVqhN8/UhECWsf6vycKh3FJ/Y
nJPo4u2I3DctPq4E/IQH4aIy9EM4k+CgozIgHZRQZutFW3zcgnkZoBDBqvbT7X2SIptyrVIcFPb1
19bUaH6MUG9Ek7Y+4HFt27xlbo0DseVVBJGuObgdDEhLPpn5o1n0nCys9S1lOeboAAjCpMJJxIAT
5L0uzXr6R6o8S5QVnmar2Dz+U9I1jhx2TAxVKbnDpfwXZ8bGFIZR4Ur6nKc1/NhcSNs6CSwOQwUQ
G8x6/Mf5yRS5sKjXYG2BF/jt3UFufd4y0WVhO7oHe7fByzbCS8VMgkpOFikdic95341DSYMs1Db7
1moobQJU5QdMJ+yXfk+52irSI0UFc2th0L2t3cp6z1gRPQBi+FbWQeeAbzDUJXlPBlXRuQ8qp3rc
ap6dj+c4jDsmnTd82zr0jpWlUR2Ka+XEWGoZhRuCNFj632rdvnzS9A/c9Aq2Y+uqV2c4fFekmHpr
Jii4+iMRupmsqIvmndColwAR6/dP6LDRyJa0Dj7tKfxKv367K9s4V0pchq2c7z+x/pRbT8FrvDtf
+4ufneid4Go7mFxCIs9jCNpsbBcSSyGm+FcpVOppqjgAVyXwrm2TqsTMY+4s6t07iJP6brN8z3hq
UrWedlbtjj1gWvpBzekTq5FdSigSZEkQokxPYgwQGhpZVmFJRmd09LaXSuPCvOEMU0jM0vkh+uES
X8QPtHa4yyVnWJzLbPNeMqOg7dYyS4kx9oml8DKDONU62CUgwQoaEbUi9h/ZKqEqDgn6d8YpbHw1
foVgoWLHI9/LFRlAplCRgBG8xqbgmblY7Ikd6P0zsEdt2VfAFNnlndlq5K8COovVZgc2072R/FQV
iF22zQnCWFfg8Cdwx0OA7dto9qUKzvCjhJgQrfb4xSUhc+ULBiCSjIER84kW4HdrQMm0Ffm7JdUe
rqrFclwhFnyV7uspx96OcQBUwAJ0LZ9JSE0xHvhN+0EKwEDzujehCNM0cAPhOZioaF/F8dGGa4ea
C6uzqclN9RwU8NwV7SH92R8xoqunyr+FwdpLSDHznMRIajcPrCbsejZ4Is8qYuxuLUCW6DLySNmR
HZhDJm7H5B6KHDw9VL0YxLOvTdUBYKkkbQZF2Z5r5xBknGadJwWsnsaaNxU+sbe9nXazvYxBB03O
iAFCrz6mxiI0RFUYOIfalkipRUtvA09txbZZSRZR+VmvBuGHkEnnoOpbWA+RFGVTopO3jabTGKxw
A3PyiMrzoxAAh4WlVc4IAUV2Hcp99eXMJiAONe8ILl7UCEFZi5PtxzJxyZefwozZhRl8TKL1PxTr
XYItbcT1xwjoWyGSKZXNf6oD0IjitvbKe3lBOho75yF5wLDdCN3X18cPRzdpnUVb/ODCkaEh6d++
FBcEFTwDfln95uq1V3DPzZTX1mbc4J9Yhqf9Jtz0kCcnNOTDGmYR4lo0++MJB0ud0nj4ocj1BOFH
oxnRhUsE2zgHS2tMyBxiEcw/+HyNsnztV+POaoh/KQa3UTwJ6r0jyb82gc7tKykCWjA9A71yQ1cL
H+Atjwpkhrt3fhfSandub8kmEIO9u17o7JiwjwBvJRchhsMc72TPfA/ujSo5B0DiKDWUu1P8+YG2
lQB/wBNlTxuZnuM4NnX3Ga3yEogJft8r+QgJbUtjVo1bDtTcTVh6s1c10gHJ53fvSdYOmRcPVfdL
EgPKF7XHlf6ucgn1Lzn3Mn1BTYwBahgNYwUBwVwV13wjG5rl2bc8vXXHLe/rvne5t3ROTNvBWd90
AHH4hXbwAzOAhymCXNRFU2ubcHUyXnlYpgXXEoeK6uioa1f3oOFVUxNFrs7SZf9TX+Ax9rnqXu8z
gm5IgIv1Rchi0HH1aXZB2ut1Fs+O2zLY5e3VNHx0AbS3cBtFrYlWp8wi3iJQpnYLD9nPOH3iwJbV
W6z1JDjxq+0rGbknRdJ+NzQchTisidY37SFvY1nQzhP4By7WmE02lJmt/dD5srqtBoBMFebzZJeL
t/YqpuzvJENG5vYKgZ+6U1dJ9nER19szYySKzEMotzq7oGI1ghh9ua7ghTXGOuMm0Xe19EiVXuW4
bz8ckX4QoQj7m/DpVDO/VKpf+aL+JgBLFc/IHfig3Y8HfQJ9CN8cbZgBUG0SlN7kl273upMIPxCk
y8XPMunDzh+8K4sAca8f5RCAA/zmH+X3G3dsLfaUYDUqmZh3p5Wr0ZnajAdKPBEw8m3sbSRCMmNF
jGhDUyvR94TC306iegLojvhqqi8UIMT+ZLzoG1gSeRfhLrQklaOp7ZSWQafP6Ztg7cEWPSvpZl3E
54YXEI+63k1DmwrvKXNVyTU/TYRUDNH9hIeNwISjTHVvJnurkr+RLwuFsh8VnKK1m+G1hOBblk1l
zHO04Un8Q0+oJEs7nU7GUAYlx0yGH+CPDNMbKIVG9OIQcLQAaWl7t47Qnq++m500aOuQf6fOBcxX
SeQ5+qBkgbOMSQa6AdZMH2cQOrfD4DZUBbf9BJu6VBQa52JwhxB+lOQ3nnVE4+md12YcIaA83iMB
555T9ysXMW0cOEVtBPCSntFWe8I8/Iy28DntNF7Eza7LfTAMXPXGSYpHaxl6fhKBajSlrmvEEjer
gKOWbssrb/5RE2xQxLpbyuF/TFpM1KtCO7fP52Stewv+CuVn4BzAB4DuxYXcu9ReFVSLeBxf+Vtx
C9+2qAB00GJpTUvun0NlAWJ+95q6WUUHghizFamyfI8+AMtnUddIaMAXfktSHi3SA3FOOYG611fM
B4S0dV3qkqP/46XjO5qFUwOujiPZjeieVAe5l8QA6hxAKVsWAouEzDka3pxR+sflnw/A7Rvd5kKg
iRrIgfprd0gyU4V+1Tn4E6O+SC1hpdPmkNerGu2qNY7xEyydSt3s6jGiGYVZu3EDdUBuJbHglRIu
icb2xqspJ4eFj5MnJivIAwBau84Pry1ckL0o86wH2G1bBfRpniIMeXtrhnRpbXhiY6/bauDj8QBM
fxawtBrN+LTcmyro5rP9D6Ed0Na72bAxRdwAyQQHq7WHBMiYRMjqHx+1Y9uY/RRrKutOMqOAWb3L
k6ikboJvVABdFrKiNIgQMa7a5kph8r9Kp7QmSrPU0MMmnk/q6CWR9lqvfqrfcRq0J0UajTPikRHK
C6C1YLLjnEnin3UrlflTBp0ydeXeTQfEcoXX/TfwWY9KkdUq/074BQ3yCeN004HjSQ0yVG6Is3Y+
qldPiKmagYQ8DQY53tksQEDUbpzGs9Dzn0ESJSHAJbUPFQcFBOIGXc602FCzJYNMkAJyoXmyutPj
rpoOpIqY3oAUqjoM3NWH8U5jBDSYsCToCMI2VAL+E84W4aETkfC51qjClq0lRki6aEUHibgvJcYk
Ynwc3Pv48xm4TtywsT3tasPF3xvNNZ5rVgsXLKW6ddOl0GoJ0+cuivAA2L1VRCaIbQSuG4ZJbNfY
aas0FWA18/dG2F7ZBOzhwYBWwY4X5m5szL4le+13YrAJzfW2/mSXIwxFgj+LJKPESQimB/uhmQNP
ojLUp/6nAnoEfmUPhFLanDwlSbbzr3zeKUVwYkhX/HeCo0sWMMzUxtMdKPf3fjPSSviUm23/920e
1ln/1pq7Hd+oTDmhyBS8YndoGUm3APbkv39j/9RF0JDOCG0vEUX+rZ0FFRmnBnQZZgyNCYCiDIQ9
CfSXmGltWA/2kMmkHsFSbS1ppbMoQf3Uo7pTGg1j40qEXCw50p5IyAnudip3ikcyA3bjK5PSXbFR
yWjPcStdjqKh/0UX3RSqOJUCFu0tFTbQN25NiYrdcHCTQdZbFrxVgjWw0kL5VVzKn66UGyR3d2bq
jWUzsM3XxC+m9aLjyQyM4+mefRIkNPS4eebRO/0XPHzSeozar6lh+CKaZ+r3hrSJWO4glhSU8gnj
VmTnp/QAmr2LONphj6depUCN0oCdZDmwg5VYDxvKOjnqU0m+rrZM8dnbOXfVvdmWf1ciCSbq35gm
RYN0UCRbyGXeYk9MeElJEDF2Pr10QDlIRoiRNoClCnXwky3+SsGk6UuSI/Oe/MAZBQ8QuAJsT9aU
0IBDJuJXiLWY1Fg4YIOPASa5bPx2tmHYPizaLZb+GQYluTGcZxHzGvHEbH3deyP4uxbqH099smDp
nle5GOkGb9SBaqsUrbQ5IglyFky2K4b6Wxx8ER1G0wGjewNE0RItYLA4VPwqSn4M5idvY48aD2h8
0EEsfqyClgRciM5hMbcwluiKDQJDG74HyD5oHOhcLRV9NHBL1dG/Gsh3LpwCX/XPjWda+AKRVRQ1
ORhZ9efu/ZplMm2Q/feZ3IaKJ9pKKfYuQx9txpvLdGOKcjXTETOccTBQtXMa3sdOU9SxBkHBDC4W
X8ECeIYqKZHWpIZK4rDN8lNz+iZC5FXPy1RbYGAePx0Ho6LKGIXyQAMckwbT0BYJkgHsnhpPSSQk
jFCZNBxrWgsoFIG9ibw/DRaVyS9MnTr7R/8sXAbfQm4IDZmcrNx9TjmazbCanyZshGY1Q4QdmMBB
9RbjyANMAPqYxCiKszc3ZoxbTAxnXds+x6z/Kt1Ta5GZ6bEC0xqjswN0oln1Vl9rBEIIFC0KD8QI
+E1zEQ29sn49i1uxityYBbRh2IGQdRF0NvHc4Cwr3FIljl/Pt3vi+9N6P1RDuC4F56vlEMZYv31b
NejjxsI2YU71zua57VhsCqOIWWJWgMjjj4DBsNi/bHJiqnGrQeZ5a9jkT3MKsGTzgReEKpISv6H9
xYOPVVA9yTuWLGz5YYZKeRCVmqOPq/pWVy0mtVU99V+aisc8YZLFsfNua6yAiaj83iBtwDHoWU7S
eOvO7831n8KeIk/UusU9sHAGEdicCO0gWam7EhnDXWoFSSogIAPysN2/rE/k/BnMyG8uXiCWlUq/
wvfFQf51+i6oBrhKZKM4lQ1SrHgszKyf2zBzqLI6gsZC4fMlAQwddfKxCcrv4s/57q5xTuxA9vNo
NmRDi4i4pKI36drA+EHEgYG17dw0dRaS/gOGi7eMlO0NASp70PSr529RqC3N7ppJpFZg6iOuSj1r
KPN6Mq+9G41dZKsxs722r9AqAcVKnyWhsrplWqod0wK0VYNdtT7WCnRR7VtjZ9wyIgb+jpoQnWgS
a2LVvrQQwiTurPU/PO/FhSufNbuNlkdUq+htdb1vYLRbLp8fgTUTNj7RdUrRna8V3FiN7+FWSz8f
/LzBAdUT9WE1sD+1qRlcbsqbnzEwBWqqLjLcFl8KYMK5bhIyKw14MrT914oYgW38KZglMV/0uMu0
sP3JhT/q5aBUoVhBZlZQxwaDtjP5HTj0pjzLNn/QxgV3+Gzt3dsd6yrz+HtjWrHWOytD41MqoEZl
+sT1x+Qcj/+0Mu7u+evcjwBsrCganAp3fjhQv+2Oyu9dM/sSps9qd2YdaDJpugs2bPC4p7pXgmW3
17doR8j4Oq8/QhZestIwsyZmkYPxOrfZjDrIW+22QQ7ch57KbEXUNrPmD4FCRE6enEC87Z0P8tcb
j0eSBTuBQLJfeFBqhuFsj9VXlWeF4XCvxkCBBOLM2jE23FGv6D7xDYsC+EheRc4XiSa43kDgYTSy
AhhooEGAsqBce8IyG+QHHSg26+2dfG97gC8JEz6tvy15ivVSh/51xACI/VgbsdStXbaRFXWCKtki
Q/k4KaKJp88E/mr98haYHSKL+9fOlCn3RHumrZEwgeVuqk6Nm9trpGUZ8ELYrCMtGU5uwrszzPEg
g8LaqUKDc9jvKRO68/92VgAeSxsB2rMCoEkpL9UPSCSVCmlhK50kcEa7SG7MzMdxfSJyiqPQYx2m
ojrFV8c8whCIlSya8hKFQhoRmjV4XkIuZ5oO7njsh+oSyC3MdZHWA+R29jjY3ZsyxjNoYC1TcnaZ
lufP4L8hoi7CS+DPOUfZspXKZdLUsntkiINGmdrs4sfzWDEniMEePAl0D/BCvmuzIGmhHqAVqqge
SkwjqaUIfLbG1v+zPnlI1h62NmMNZKlN116gK+k8p+yjQRfNROyRYxF+HahJbFJau8vD/jqGlLtc
U1htHYtwDUyI3Iln6IfgSjwkst4pi1ci47by2YJzcbDS+y6V3hM269N3jCan+DSRmqfwFsCGLCio
6qF8Empls2rJJANsQB6dP/8tR9w+mm/0YRGcfDkxMyzRsIXjhH3Zn+ZEsIEQZpljP90ua19iwqoL
nYKX46hvTL8LyVXPlaHNn0A2XD7/Kb+1Rz0YvxtRQYwiAuVqBUJZyewUpW2NO8mp+6/r9yPJWaka
Nz9R8SqUAOuVcyCY2BX/YJbCfE4/MQawaUVFx4w94xkUOCVdYDvMzOo6+9tzJZ9IvWKzNX4iLppK
Dt7kNQfAb7y3xSCohvhm/xO9KI5JRDBLxkiOFvwwy5O6VB1qE/iv6qZYJEXTEgBfc8LF0cHHQLiK
ZP2RmID+icG8AaRNrnw2BAHEDYxWxoAXxBKH/BKO/uvR7JyhV45vwj0mYF9vzocYE0TNqyr9fGw0
3mLhCZBMblIuI55Rw5mta/apU+oNcVm6dU0m0PXIyCr+T4md1KqwOM+HGqZN3FHwmcB2FZuGoyRq
txrb21aHOTffJSSEimSr2LFwWypRwMiRWAr/HgN7l1gtRO9PuRw22ABkLB1OlALEpgzItxaqNi6a
6ezBRyUecEvJ45d9JSFnDm+7S3LlinFDxueRWvQHcCIrTV/L0yHGVi3RZqB5hpf7f8L68f0GVHtY
8jHzSp5U9YSdfqvdFrQjFDNLh34o1hQChiu2tvFHRVEvEMpDLPnS1yoh4kdvl9m+NppkXVuwJXG7
BrYcaALcJaCoFVT2SfBuUD6noBz83Pmlr0YyDzi+CsUhq12zueQe03MWBZhyTYjSjPWuka5BzDmx
Y3elBs4ibE2zwE2fii0XQOcZSh0P7EHnSvrYmWZc4dSn5KKBBdHt2xi98UzUjlBhbtUn3W0RtRVp
EIQ8MAtjMdthAIzJM6iQD57ijSyLm2j3Fv/SVGlAa0V8etv/lZSiiGsfiOkUzAPl7Fpw54pDCHe2
lgaprsOYGLn/39XrIkBvjqdgA4q6myOUzQoxRd9EWnjn+/V7UldTfta8In5yiNMzE/Rn8DQRfW5N
xDWVb2ee0zEPkAIzAUaQuRqUflP/u9jUNhuibxBGn25AaxLMA80OXryEGsz0Y/FnR/FsrNWoBTV/
GQEn1GhntlQ6v6wT6nw4tjjYm91cqzPImygb0Wuw3GaOAGf9XMlatzYocVwsYM6GdPLobPuYPnmT
bn14+IHdTIxCnK/Y4Bbx6KzV5v4EIK08MtM8t9UAMyHvdb+lfbDnMzudEpgie6uwmqt/qZRiqYDJ
X8dkkuzgfenGOatZTfMVZQ/zutjRsEevfQ12wbIDSkzpLBg02kCMJAdwJ56yDE56uWWxyh99v3SX
fnRFeAIx8ujds6xKjkoeQQ4/fdHk4zlGOQGMpVpULoNBN+NzMCfVUFZn+MCHS8pYqwMQfqIGETGz
rQ7a2XtzwOuwhhBSENKQlcghVxik08bz9NEv2El5em7WF8vGinitMmTqWZDdV0Ryn7PiqXTDQyC5
Y5eXTCvgShXk00lnosaPY5OSwla2SNmuxrpxgQneOUkHPAJyVoLZ5gfo/g5ibhqiJplmdYT974tp
LQLzICBAqZ2Y96jZRyijQpBe2OZ1seunXgyzwmFIpFlxSZzmZJueYJEDbNIBTx7I9FeVsE8EUA2J
aa3xYOif2WDiVmAqMCmMkrOj0ZCT22pns5hvPzJyrVn1xTKpVIYSDRc4c2CqTmb/doC3sD2JCgHK
bQIB+fCZIUVEDGUqaJvA6UKY6rEXt60B02kVdYoikpmQA1JVx5/Jg3Ihk7+CrAago6Vga6BXpWkj
mvpVmpecFn1wJEoDIr72z/c9bhQ6uxL3caQbkF3Hn6a6rsqxiGvJ5mcQaequAczwMKABrtIfzJcQ
3Y0W0rx8LA8ElwywKqFky9sKHgVYeAqGszTvSx8ZqkwDKj7W35puKRfH5/pOK6gPKn5Yox4k3+gI
DIl6TJbWx+VUdvLv4ehLKOqRTtPbGL4M4wuuAsTjhi8kkgRFsNreSP1r/m4miSqNaZti3mL10aig
QwlKeqwRjwavBwTXJ6nvIhfwnBgYVczdsv3kInJ5Hhb3L8wsJ8C5pF6XG6M+kGLlUYJtNTdjZEFe
RTnLx/cz7fjlbx0B72Z/qJn9Y8uCEmwdBt9O7KUbeogW8rBg0Ncvi0NrUv3VnP+NxYNy0z4qlYCa
5jvVISsQRQOLoNfhYNOwE/IFM0zyp3Nxbpz2EIzPinPzTPKSoaT5fDjdbxobE8sVgZkRBaGczTtm
QebYLbFF1cRGcVVcldnokz24j2Uv/RbVxzHfyiPS12z6UTDcmYHyavh5kbAOXnlNQq9OGecOh8GE
gMArevJy6kkuWC+W1R9E6V6SNQ9FoaK0ZqmjJ4LFMT9WVDH5p1jNPLquc7+yGr/StNWa4/5vsNRP
jRQbAGgGLGFfBP11X5SuYE39S7zqq6hF2pbsDpCFttQ9zC8Yn0uKPySvu8oLp1Z7y3Fe6vhqGj2m
qBHjUc4cHvWn3kMIw3Bznnsc9SS1exk4FT3MXt4cPi9R4PYDtEyxO6wWqXoubdw+I++NZvCISk8N
JQgcMnunOGmVtBLdiFpGfl1j9k/YCf8DEp/OnVbQiIK2Hmk+u9YL0XAADlV9VSHsoueUO3Eisx7Q
hgoFHrt3YJX0YjBqheJM6KPix1RtgjfFYCCRDLCbUX6f31bVJHVraGY6jwMOp/II2k2/vFvC++Ce
lXjIVfDDqzM6wIXJx7QOmvK+jCxLnx4CsAAyoApiI6EbWUBTPfuX7DQRls5b7YHWgqwXchBxmXJr
ce/gicybJLABsm+GxnQRjKvGE/EZ9pWWkKpcsy+uCSrVD3B3qCzaA6gAXKHAu2F4xfEf7vDeXwDb
3hl4LOlY9kvrB+2znkUe8/ZFbp0BoABPF86XImEF8XIQmLQLDPOQOrp/musWXnzMmNzsDuJfYvgd
cLvHV2uWT0SLKBMU4kNw7bf8CcEFGnCBC3K2SFaSxDq7JcoSNnaImKP3vK+Akc3OaYWARb7iEx/f
ut8qtJk0UWFD0B0rVljUJ1teSLy4q3hYL1GrpeF1oIOp51f+iQyHq4kcjjKMy6cBDzi7hZwwsp78
8JdGbQI6pT/ky2IFAyhHU6+sCiRV49izq2JZSnbwSKJjOjOxbsBxgE7pNUQxJna1eXfh6tKFBUIA
uDklF2n5zzqFb+oRHnHRYDeWyWQY8QwteOAJw95w5MDzi57PW3ejQwyzYQZMGP2+yekrE91+SRKw
KX27V4Jr8bAWpBOjv9wv5XxOx/VMbrtrlTdkQ1Uot7VjskxeyWQhn4KppOi+U0cH9oNm73Ca9n7m
dcdzky84gGd83J2JHA8X+PgOV42zEB4X2/3DYTJ+wuSyaVkZCpUKGCkFe77KqR8qdd+O0X3rER7K
Q8oqy7pX2BAtu3PwcuKLuOD0tUEzuVHpJ0mw6tH5O4YH4/JaoLhtmJuqju+av9Dp3KjVqbDsFKLg
+VMJAM4Wew/J/NoFV+qwAetAizaOkOj97FkTG4WOpgXgfDkptE+lM9VRZ5wJqN5B53z/mTh/M+jN
2M8wQN+6Qmt/wVSjseBVsQJxqS/UTNEpKmtMDBklgCHTXFKxib/xYLmVjDBJMxRsrc8yYNuWfIoS
2SpCxlU60U8/IJ9NphhqpzjatUICJTTUyGTPrTs6mVGmkt/mLU+Yu9H3sV25IVcUWArqRBEZ2mYg
kZIjVJ6IS6MmEPe79uESI0NqJPO+GeLRIJDV1IWHwlBtcaUwlI5CaI/p6K6l9nr09iIKmkPLwxNt
zjJR6C81RADSEx509BklcJNlm59zTdK94FQ2IZXgwzs6/LvhOiYDL8M/WKl87eliRHrS2Tp6cHa7
sc+An9ytt9QQ9idmDfN+SovD9mvGC+GXdG4wsVB5+D7n8c2uchnCKxADUw4f8laLMmR0Ha/ZfSfq
f0qstbQcwHuQdXqZtg0B9aF9nGbgx83Q7w8W339vCxIjPfnQ+WBh807q+hFrp3PK7uN2ATyX5+Mp
QMOaiOLSzKuS7U8YvsO9PX/fNcVy+9SGSYEBVp4pG2On+WYXlRCfHv9OO5rhcfAdfuLlige9a1D2
29BXCebINpLRfNyqS7UkhoUsoclSXwKIM921Ogo2uj6K9KVla3F1UFZKM1B19v2EbOiyh/fa/2gO
3aRh9VLjNrPUr/DOsdSYkouymHiUZ+g8KQEWrWjdSSITdJhSJ/sm6ZBVl2JVPwqXVUiwjHZaCvuO
ItMXuM5d29CtvnW3TTrARgjMiCFYNHTWFBr6P78QB5aPRQ04ncaN+EvkulaKwew/igUv9I609qMq
LqN/d/sf3ItuWhT2E87MH992BBGYFpOxPlZn93BXQn2ZBsZohIkOEc/5J56oUmudgoA1S3OG9WNo
FbPwtcUvUOmgabzAKQqebNirYigi+vfzacDQQYV7hnT6vT6J4AxNeSQpTb9y8cYAngEW2q3JMVhp
kxoHlXP0hGja31MbBq3BfPngDvqH6IMbDBPwgpXb4mC76Vac6chAM+dqXisgN3N3j5M44g2bUl3i
5WLXG1DKTFnYa+oSBuYt/NjWXUhIC0MZ9IvNNKrOMMVXgij5jexjZDxhxOZJfz4Zlx5buJnob6jA
V8oBCyJou9SXZgd+YqXRTsM8Ql2b425Xvx0y6+R+hF+DKKkU2IEU2DkjzAbRToIMBZ42nNmE3Dya
0AN/zj3qBhatLkMlrdHI+mGNxqd7Di8GdI00QCSoKiLFr5KOJFQpnk0YrNZH2m0i2lvjKi5lbLrh
oHwgkYe0fxDGpV8mxeuOi2kk4oBhX/YSTuyuugY8yBjZlvw11GwsZN37p3ABQHhPH3Dd5qvc+WxW
IJwpVvpcG/80K16V+2/GgtIMnwgG3GJq/17fz5sXR9Nf8mhGRVw0vOibbJq+CRiWBXZMnEYyUBOp
Uw9YFnMrSo2D9lbdK3Wdn9RW7oFVHwcvyv8gSNd5faLLCfFEESZrDT42Sp+AqOJr+UmCKssYWS3Y
FTnncIdT9c29XB9prPAUCOjxIPfVSBI7AEe4xA/fWw3DNNpOIr2qi03utAj4NwfW7umVL9yLZihk
+FTONqlCUgDnGiIIqIJoIEPxWWk4MoBFV4vhb9lCjPH8NAh5F2UFJbD+o1Of85Al/Wb1xb/1CSDR
1MygwIv2gfcO+P8UVlao2jaWy1ru5NZjJji/zNCkCG0bCO3jkBqo3Lodb0d72vLGs/2TKrCw+C/9
vFck+edmh20B6NcuPeeX61kitS325W7kqgHMBr5Dp0bXN1XYrdGoD1LL6buc9q9TysRK+UM45KAF
Xe9ztDWRcRST4jMjuuvAGhyDS8EFcX2hYNVrKrCJoa+24ZiE9/ujVVAaRPSc/RWBPXNx40iNIh08
6+W+gaavqO2DZ2PF7PzzwJPnBnTbX/fT1UpfLENJ2k38eC5xMY2VB7HhAi2e5XULy166KpeN/MEg
ESTq5kIyyPCmOC3z2SlAg5c8pTu0c5L1h9eJumc8v5utQeABRJez/moKVtRq/Bcxq8GBcn1h7PII
ZlLtG/e3hWnzDOPcowkdeiuoy7bJebJwADH2WvtiMwYXyqSwS2NXmTEo0zx8T3rbM+fQPFpmHqyT
K9yxrj4zs/YjVYlDiAggRzcO7YVJP+h0KopgN1fCCn8FjioUM6gYTApzcRwXaFmxBtjDWeVurKr3
1mVJZv+zQxadHX4EcmxHfRep3vnjYgIZ2NU4QWXByEcH5dGnofUdcNjvDI6ibEXZ8q4pDVmZ5VD1
dsY72t86SQGrdUUSVAsKsPDr08bsVluyhWSnT7d5kPvB1MMKXHsxW/U9W+8R6aKtkBCdiRTCi81Q
9FoiarZiKubvqJhEyCTKlSEP0n70z7+L7B9oglu9OJKuBoKN1FHl5Hji7xLOclWxV60atlZbwUKL
BzZ8+fy7Mxd8FicYY+k6HNsQZQhwqlAbsQQ/QdZ+n4fYUVssFJTllvpIuDjuQUo71fISlujCidTq
Ry+Uir7DSUhCC4lqq9ydB29zrDjqzWDS+SapReTV1PhN8PCNuWOc0bfTaS627cQShielDilg9BBd
8iyobPWe3MrOtxtvH/f4ySVKHg+tXPyzZHXZfo9+sbVlCGER0kPczoWov9q8LKuKGHsWJyuYZ1kF
66eBLIUAFi+Ap/ZdwYMAqolBT/PY2pJRDAjlUfaE034hB1ea0ZcHY0IOfoP1BLh6KY+JIIKylVW9
5njmFObrpXDW3ff9mK2egKgTUaxgu+czK94SNpeTbRKf+wuuz903ujKOPdnK1PoXa4Fu97vNZARk
gax8R3vPPQJwYf3/oS9JtpzA1dVF+7tPGQrqyX5/p0TXN2dYmR/htSTgeMm4pYP+HXEu6v2cE6zY
errV6ZbYVvSe/sdVtPf5i/oInGbmKF/qgYT2B/R/FUFlYRmeaUXozd0yQoXmfrXdH++v+c1eBrpD
eLuh5+T1EOI7aNiDp6KqoCG2vRgbyzdDKY4Z/wk6P5Q1ukgapRcZstRE65clYjFzZhd8WWUaSR53
75ieTwBn3w02NNJwOO/qgleqvCasuBMJUuDbevN4eGT3KQYka04ujCZpFRZX8T8Wox2CpdfGsiBz
dDxQBZD7U2yLlrQmUbLyG3T+mDvqC6WDlEDW9eZHPgwU6Hbiri4K5B6+irfy6oJT1kFtuJ/mAcp5
cUa3dZKlD2SRob46ZYzbOTw2iTnJPn2oLQJVAgIpM7vyfVGdM5J/7Er6IT+vqMBQmC7kUphpqzLa
+jdMLWS6hJyUUyIhuM8NGUcmsnUtFK99SV4Ss3QE5UEhJWgit4ZdCIkDW5M+hk+LBq6Hwprn6Xpm
0zk/GBTjDhWIZW3YLUBD8Sat2jcA8VFSX5ZBN0fgDTCBRur8311xC8Z7oYAsmnJwYbX6oYY28QS1
DcqvWj9nHwB+jdeVOZKxR0+kQQU3bpwk9hG9Sv9egs9rn1ulNK6fFlNPKnZCERpVdsGX131qQVQl
/4756Vav4gKHwxFPfhEpUQ0loA16pLTPcxlf1Z9M2m7v2okCCAamnj9xP4FfTAM4Wmd4fzbOnc0R
3xJrW0MEtRET2LdnTpyUIbmkPP06MffO3zhHvjOWoLQpnGGNz9LUaaIPds0vShVwzEKlm9sqMdR0
x6vRUXJkXn5eNWPMQL3laIAZi3RHBczBlUBASRCb6B1Q9Ju60AMHpvV7Cg0lAsXgBdbL472A/bxn
aKAm1vpBkeEO2Z3p/dytyuFY0k/bjYtHCFe2eHTvTqk0b9fs/60ZenGAEBS+UGl2uPDu95umTOKS
i/QeGZ3TjkiRWTZPLdL0pC9x5OghUr+CpeBorue8aKujAbY93wVW5PPfYb0Vf5w+aqv0pxwWzjCT
5En9zJ+RjbRIHzTKwVOXDl/A29nklQURgy9jfo0VceNG/BgBfv/68bdyv/aZuAZzsntJvPROaeO+
D05O5HsLF4dAdsDV85cLelcp23i6kkwDa55SJIqgTRuAe/+3mPZG8hNAqoGVgRlqsVLCcSzZCneE
x8Jjs3iJFJaDnuMUIAORFvJESjGLmRSXhfZlRVzlTkGQQj/y8Srw3Qvnl7EveurMckTkIZmnOlb6
x3+SG7YqsoPJMI4wLuBy4GmkU4fes3z/etGCCGcQkVDoVNt/049IUkcFmyc2EiWd1417DXH5r281
GKwgikQZshissZvNV4maNdwk5tNDvj2E7IGrobk01mrRz6cxYj2iPIBWGYMZnguLIH8TwFT7a5eu
OgvP2WQfirFqHtJS8ewANDdKBDGD02Rja73ZuwZtHuOqbXzlnIr9tXfsvruZewXVEqDPjiOlLwTZ
rmML9cxWdXvBFI1bn2qmkSJin1ntDBDn9TwFH+/YtYvnatRB92qGL4C4l+oK4XOePDQW0lFhoM2n
LFaxn9OwvXHg1/040fnXMizBfcqaH6CIHIKpo4XTUW28jhF83wWl0f8I9JIupJXz+qQiOGRsEe8E
OR5xa9Vlu0VKGCPwAUX4MKSNn0jXnUDIKOzan1drFVtTOUih2/68unhd9p/0otSlU1pP1m795WGY
JWlqCvo412jR1F6b4bBlUYdEhOozVtR9fbDLqrIM4tFnq5UzWsTsW3F+TkleltPTFeP4+Kdlk+Jd
Y+ZZ4gzSajjR+mdrUnGnKbrPP++maoW+Wa8OEcGMeybL+sDZYYeeQqYlRowmbfZcJKnHvssxkq+W
ifxvIs+v0xgLB6XkgYv8lYdszsXoU+AmWY3rkhGTEW8naT6r4i3MMBEZb1bzfyq1qTYvAg2f8xiF
kKawMucG7QacrdCEAPvE9SzOSbi1HVuhMzHoKgwn4585IEKBTG+suCYc//Y3DGaXBs4iRTTi+J55
1kYsQAoNEFVuUFLWfKFFStg+55CB+ZaJ+YK+tc52kMhsSGBaQQGc+bxDLkcNtRoDEDXBLrzficrF
KMPQ+WilUXDbRF/1ZxV2Cx8KD+TuVO04ng5i3QFA2/QX+PrzSVR3C34CX6TY1tA0U8DqTWvtuO6C
UHSd9EbTVZQOjfZh6cDXEtcKMdKf2CLqHkI2gNv4caZi4dhpDmBSSui/GePGfl1NKaWgvp3b9JXf
yeSYqWI03m6LxVgn3C8RpoCfvA8lBGuw/nWfxvDBzuKbCGUkyTTKSajo6LGrGytAl8ZE2X4EjFA6
vosbQgrGseX5oBso9gh0l8dmhEWdkXun8gyQi6cGRdxbHy3G+ksnbRqsUZqv/8SwNfj04V3Z2FrK
Pvl6tJdRi0BVpNKyWb+3TU/dKjJ00oJjJo/r/z0lPAOKrlmekd7lcqvSUTmjbFTI8eEqSGk0mksO
+xr0Wp2ex8Fi7x3b0EIjb/vP6ks/lryKcYWc0JiawGOuineNHdUzhc9UHyX1m9lipHvZTxq8n96f
xwrIovlmMBliKoXa0IxyHl5Bs8GJIBtg2RWMinTHxvduM9nlvnrPff5O7CLLlL9ADMeP0LwODlIi
XwnXd1gzjq0xFbFpdzxDz0/UXAhnVbPFgcmW1GwzMSEq1iNFY6XfgF98Le1SfacnLrsztwT6UqjQ
uNQSeu7SRKptthRK42LHbzk/W2owz2RWISDRHm33KGjemRNvDodSZ7ngHMtq1+ozujRUYYihR/BJ
XGkeMHDarY5j4T16T6fkh0c1o9w6qBMeqQs4OBKNYXEaIkpPuouMWzRI+qDVZCJ7mA+/wuw+vuEU
2ovStw41lgQg5oSMsp3jAJ5dTAMy44Hcg+4OxBno0oZ+je3qgekl2DTDMBko1NYtaqSGIaaU8DLW
EP5czTqHkzZXm1joNm3FvJlrYKI+2IJ8HRP931oesYC791O1PylXUGuY52h0glTWUpZbVn90LLCl
d4az7PbkckC3kyuIqFL7/DXMUZu0c2ReaHoq3NdC6Lll1L4JnUkwG5mtGrnJqFPRF2f8IjbX659M
Rfdexdw+s/shiTZBuW6WE2Xs637w1ltCkRtnjzyZZ0y3J/Kg3iIQ6YhXjHgBb3yPMSJn3Hq6svJ/
9z4gzLz+qG23eSzPOO20iQmNfcsnwQpnpeR4+1L1AU2qvwuYkyCNjFhMJYdUYeGlqgReV12VZeLg
mox0Y9gdk2H4bFakM0KLLq+sx06Fm+uQDBJF0dDNwtnebW/HoEYmll4qKYdjMAJy3RmdVMX6vg3M
hIoumBs9R6BfAvNc6AF3dizgrNwDu5jBVPEwytQu9B56V+Msxtu0A6xrZqzzpqnrYh7r84QVBb+t
nxxO9XjQwb4dibr2VgaeuM8kUXBT71c2VRZl5ZXsPH9w2qu/nD1fieGdDzoywH2w0jDGMwnFEzrT
T6ivErSrA68zqSnNxUCNW1OeJ+sjALK2VlNC4LLpF2FozGpUQVABAR7suIWamVGhokMgsC8Rh0bg
dIcrJJMXpTCWhMLERZ3V97aMrnRU+7M7WXSxZ9JTAORlCGicdWzkkUguFeGnsVGVWpFZXE6vyPex
mAbP2hal7u3gn0J9T2nOmVAg5O+Kvc4L9sIXnYIcHfscCGsv8oCv0g+PRh2PjUe5e96YV6TKVnVA
ecJUJn0+wGrfmv5LOZSLfMsGpvzMpLTtxdrjvt4/pxhmvLfnnhZpmq2z3MHNp+0VFMfDdrWZEhro
7WKYBfVIjpgLV4+pwV4Zqbl0e3ch/Husa7cOVPleXjWg+XryNdvQimEZfZ9IK7ZseIZDFbI5SvgC
U33OPV3z6Pd2vvAtBtbcOm+XMqPidQlTs5pF+yBf+5Fd3QgIJ9NlUpcdR/2CSHqOIFLL6+drNE1v
mQ4T6rjuwy8Xxa5qK0hEZIneoZmEvFBECWc0+eb1YeHJ7hExliqs+602f0djLTHmjSm7AePeHIxL
An32+r7/p46z0zlc5RowhM7Guy2X8xebHIxDDjhW6PlnH+vX6eBc4mBCDqtZCQRZ2boJ/XItE3wL
Usp8VnIB3X9GkZvQZFiMbxylrTaL9KQfUI5+MQxRIHfaVAF0r8kW5aeQ+WezM/fvztr0qAaLDylT
uWc6OlnKgPvG1+EjHpAjF9L1GfBnzMguIkTw5STEOoAIvcGy+cHLwz6IpkAXYtj1JaZL8pWfcrOC
/N+EWll7ZiylK1+DIxv2Axu9IBe/ppsg34dc52mTdX3xfZEbu7tKsP/NwSKUFGNq4ndVynkbmMWv
hcs8gmd5Ox9oQyrjzLhyrjBcBFED+4yEhWuvdQk1IwothoepOSL3QeIxN6+Ridj6zQFZDN3QGk2h
b9fr/Ot0Lhhry3z/t47GSpkZvMMZPm/7Vrr/SfKq6dG/C3zDiagW8Y215+qWD932bEzMnxNFHrok
F7Gq1fh//fBZGwK2T0i1AVs9h+Xm5Z/H+BBz8jrgHPG3b5y5CVTmWtwAvt4UTlU2ShVJGL5jGo6U
O6d06mUxxHcgZetizjZjRBOVpb4MuNFJCyQaAu1cExmVEyzL/ITMI6cQSrLD/xLPty20Gz9999/W
vXCanbCzydQD0YiQPRZwNLp79PYlYyn2a1l8zupQeZgKzU1wyCkOkeANHFxf3v9JiyWOGmkkmH1D
ix8vLR+PQ9/Gkgv1wgdpc4WzeFBVjcA+TC6+1jRGYENeyQzBT4zK+wgG1wbDdfJHog3q/e6kB4Je
emh/183nyBOlwzuk9TFJM2tzuAbO2hAsj8VTB1P+t3MolHsdcXrJfDR++fbofGLB7+os/2Z/fEHN
IcyIk10dZRflSp2zlTkAjZrpOJTQZ2ynNqAi0S6b4M4Hg3nEexJ8XuUB+9Q5UCCXMevmnffeBgZB
Z3xpYgjNpdbLz1RODCglb/Z5F/o9t6HYOM2HBMq3LHANS2DPT4QfAmO4elvD0LYiyIldQJCZN2rg
/0iZ1QQCa955H/UgvLuEEOiZrgE6tIgDiM0joE05wq6v1X/y0KZ/edb9KzQ+5GmavN+FwMKVDmwS
MbiCkmrM/1E5/HnLrSb2jRkOXENSdzyac0DMocvfkhamRRRAxGlTdTrr48cM4z4qMUdTIg+W3D3/
wyrT0+JVIhFWCEWh/SsLDY9wJSNoBW9ItWB/v2lTcXTrM7fpSXeXIYAdhvzAsZZudw+N7tSfelh/
DlDvUi11fSWyqX3qQccB1272+uQP2r4Cf50rt9SFpXA42xt5gXC4zFgyayKaSDD2fPBeijXOQ6Vj
a9+Kd6livWP2DdSkaNdxn8vbZepXNG2X6Wb8I4tdW58MuO2ZuEBszUDRFtRQKHngiBXXhKjh19OO
78dpgFuc7dBX2/kLLUXLfewLFokCGO1/8cOSJV5p4X9lzsmE5yyfDhbpz0p1vHyDZlpGZmMc+KwB
2hYluUewPhA0bWGwSnD7nGGW11BMqjc5yBfzKgw4ZvKn84luPWWlpddPc/K2jCOmRcb22YtMLRsR
QqFGvGy90ooKdDS8a+6JEWer8IxC0uFmSTgY5jcSSdhP8IUaMy1I9t6V20nii5x+4sU+n9VW02jC
WP26xMcG1Z6YnqgDBsHmqHNheiGtVufdtlzBJoxKs2hfiWJuoqLUOZn6zLEsYoBkdbEoNecVlrK+
NJ8vtBP6mu5EqGlmEdwU3oMRCWM89l8Dtg0Yz+tpqZ0N5gCmW8alm3IBkScBG55W6yMvcwuPXPWl
amZO9+3PEDigRoSh8EFdimESO+o7ZXnbz9LzpTYHE5Kemaia9xJcz4QArKutmPKTKtGeBpirMFWI
WEtll/yWNJdi9V77LtakfUaGictWTw703cKblg4nALerBZ4ITfAAk/xX+0O1SDTG5IrUK3vEjeXV
fpQwz5F0okW58mp15ZOTfsvriD+Q0Jmi58M7tSgxjPT/qQPhYvhhc7v2PzA1QD7orDNEzMaX92o+
UAshdE8bbbss4AWN0xDzZ4Qam+Gp9BzyVLt67+7PUCFlfeIf1aU7Lgfhyhap62GryaFMeSH261dX
kqHCur5+iD6qnifciWOOtySegPPW+u7EYbcesCF3YH32v8m25U4ZjaPMkhro/69seAUUbY5pxQYO
rO9V42cEguo07qI9mBWiie2E4zqdvKJdGLon10t8+YKhQ+pnePV4C68V6jyDFZxMyerAXwWrB7M3
Tm+4ZbyeKnh2+TRNGHGnRZ5RwKbrF5ByUY5xPXBQB8zwk97QdIhGYSuNt16VShM4StQBsGqulIef
fSbxPW3CWlyEX5t1LE+nWhfLXMSCtmItUTS0BN6sB67RTTn+P5vV7TaoKOyTKILNfhKshfgS0EVd
luetYIyHnkx9wOpolSG9+UqLr3PsDh0w6o88uFN88K8UWxrBCQhFXeI5J6JIhGcoUCYHbtvLbQCc
yXuvKq8ADifKLNy0L1xvlNN3ZX/hGmlbfbI79wCrdXY4Z1FY31MCsT+T8YFEYKlklH5FXMwpKsyM
6z8K3EWEZrmfVqWqTvZOj7raIAD+B0ERomB4ZRlI00O2EJTRd1LRH9TYHtQfanB8bgKDtnBNHM9k
m/om7aqdsqqExc3FjaP/T1DPcAru0d4IAB7y68DuuC40zMXFVZnJWjQxVQQwn+1nuKADvoBKSzET
XfzGSXLL4i+7dRjGcvaDEiiupnuxQOKFH2ygSVwo7GiQpdsusJEbcp91HnhdnecWguA0jEaTR6gk
WuHLs0UsWcmU7e6WAENYr1Iao53UMMmuW4Kh1JQy3h+yNikRpq/05C3iNnsa0sb75M4MZI7vCDMu
cqWOoUMbLpl6e+PeS3VgbcP2qMYK3E0oHBKvHnsODIvzJxuP4ZzL734Z8dtWWd/H+bw+qde+RD8v
CGRLfYNGxsOa5P2BYh/pgvmT8SdnI7XS3EE9dmsjXZO8DnRurS+JmTyTFOsAk6QSe43pK1pFAn1x
S88S90VsgSoD8B9WDHWAV+cvI9tmWu5FZqZafWSQSnR8WX1jTrxHYP5xbgA44SMbMELVS6deq3U0
PQV34pi+qkPau+rCT+vD8A74IoQig8h8dfCL99pzXkE36JRLs6cB/rVA2uDkq5EJscGO5OjnTTUJ
agxHRMxllwV1H+FKKLXWfD4Gy9jsTRxbOSIXqP4HMJcxNmpyKlR7qS/7khMo/EqitmZjhGDQ5sEk
eUNnZFkWcHaTYUu0rblTmPypD39yixK7Pqoi/cfT8WdR4uQFbaPpaGQIg4Y6lmO7oIWMzIiW/UcG
l9Uc2P7X3LFkkZErotEhQHFnuyvD0vQVpcCScNJ/imYIl+qhbffu+PDUDhETTN2zpubEoii7kNQB
JLxKC3q7lt7ODhCgAfxmyGqCxR0Y/epgk4YMyL8f3Ukbd58ng4+wsenvEdYwJ/ijMe+x+J8vwLHg
OBll/FDsKzybWOYoTza26JIIuoMWrBFZKp4/nwLc7V6DuviCJjtoTns8LsYvgqiXMsZvhzXqvtTr
kKq2Ihb1847dmZAo02e3Xj8JD2G79vOOkEYjExL99Ii2MAHjVtKX6CmEkGsKKUGhrk04EvYdR7gV
pioGG5NzHYtvbLNUGsTyPE8NIs37tySNP5/X6cppu6FHXBSJshuL+1teE6qYTvm0hXAcW+l8dWCn
QB3RVbpR+aUBX5jr+GI8dG1PrZawj2WmcDp+ofyy+kbC5ycSYyYTzggMC3y58QiTbxxKLrNV1Fgm
DHP1kiMrzp2usULsbUlURmxx959Sz3FTM5rd9z5cA4JKlvViYooG1cu/peig48dWNssbO7kIBp9v
TXB00D4O4D5lgA9JWs2yYzOVjQF1xE2qaBZEjqGQFLZuL41dhsxz7ZxZyKs/qzFWzz2gooB028KM
OK05hWQ7p4IK2Nkqou/Dctb+HuVEd/eFxWCdrIL2L/MMYBMzuWc3/orLc4B83iZm+p2qHphCuhrX
Af4uNA0xi90ApqlcyHXSawmz7mSIsiJPKR/oVwk8CeB4FL3z1VNGsa779Q/ULFu1TGgu4xlxwyzR
cVNtFxxGK/qdQEn27nROnNUYQtAsqO47p9cw5TSc41iqRnLrHm+e8zDDaWQXKYd/T5vxCCnH3XM0
UtJQBusEDdc6NqqfX+AANeqOWP44YSIFFj7msVsKezsqRWj8zxMFKjlxdkXti9trEV6xWR7HFuaw
ukC7makqawkqtX7WjRkIcSFEpwe23F9pF0iOQTbvgI6Zq3+7T8qCSuLaTQCnsOmqAryHSTA4F99M
AKBXrvMvf8yvktV90H0oJ/XhfURcbZFemx9NMgL17umPMcRyaxFcnAe3iX+xnY/etGLtD7khXmEW
v3D/ZoAaXXh2+6nslLKfGsjbuPKl2obgg8QCNf4T1qCBxFqz2jMb7set3YjMrqnvAKDcNQ7kLawM
jx3GOYIZ1HD22Cq6I7kdW8AkLIak/94XzY+GyPQGO6PMf6zWiAGpj9yjMyrUFbrZROXJIKgJzN/t
7zbVdrqmXdZSP43eoDma+QE52x0dyb5LaYqrbdUOruHk/yCm78fKfRVnCPVqm0sAGsjha3yEacSV
XGZCrUngzP+lMCZBOm6OiMDlEk32oJiFZp0LZGG0e17QZu1IPBKV/QGnG/tMbNbaTM3dks8oeJBX
LcDLP8jzYzzy7Y4BqcYnlIkA3v8ntoRmLj2cOGpMlbI5FkdsHymlPNXAkSUzXP9fuKBrJDqVzo5u
y+fbqcSPe94DVdCRpvNhwSzVTzastqftvqW0lH3AD+B5U3RN27otIlcuCnIie2pI5KXf+/Mbzwgd
soVP+hEs1qF0VrmC0M7dlkE/a7I4Dnf4Sw7kjG3excOZNJUdOxw0oiijrXxbLk0sOlL9CVcOYE/g
GHv4jtd37bbbiyWg9j+gU9fC42hTTBTDCNhf9sSdlCpWjSOvqxjbMPCo4MDsCpTrHiVoWelk6QQQ
w3ynZA3Rf4l8SYY64/wXz4fmNpy2Jx/Vx9kQ/zXW/jVDqoQAQ8YVmtTWJIXGaF1lAZsTo10QYbyL
RaG2i3Zz5P2IPoNopSrTUCv4rVI+kjulecCc3pMMHRrgkesgoR278Rj/vl96jP43BaQp0IXffrIY
W6f9B4jeGQfIHH3/7e6HpuSfaJsIhk0CmbFDoUAJYGG7zI5Dk3BiQTNVVfo75gMY/EWCDjH6g58E
BqAQ03aiv1t9HS414zNE9+OqSlECkKNvahYR+AhpEMf/vcfNhGbnTvSa6EKiJU0swvgCDChd+umk
Bk9MBoF/ZJcyho37AwmGpk5OssI/I6V4LcPmhNvtqyWiN+Kss6Z6T32vrMFQQqJdnAtksgPyY5e3
HotptztoLK5BBNELPJDTaJREiJGt6vivjDWvZXzSwJykqXNAqcEjG9GrDtz5szwIlqErWKO/HyDM
gLBkXQ+Im4+vT+uieehaARwajBWeC5X815SFCUCPGepLV44vTUG0MzMbUMIP4ZIoZefYntx6erCi
fn1yDQ1IABNqKQQlplH1AHJA1jHXljwcq6kBhpeRKd1zH4VvZVrlOp5NLmMGaZ+MdzS4JmorFRoJ
Gacgq5VaT7LoEQPOb6s+NVKiGxXrouzKCEc4BqwX1NQdGzE1zNhDhyzRBOdNH/X2Mk4AH9DxT9k4
H37l0acwEL+f8uS/nr6zo9SXFHmG4iT64BFMf3S1wWO9K8NTDh3jJw4CwQLyKqwXeovdr2nf6T7n
PyYD5z0y8XCt+FZ0fspFJx7WIOsjn5p60ozCfTlhmtN9xxl53wWU0gJnq/6A3qox3bH9z63I3nM0
EZW9r0P7LoK5u3GccQbUHTbzWxQultYSJvLohweAjlvtnsQTU9xrwjrCFDSLoazLlvchWsjCtUZh
0CDDiwxoy/SRClljNhgEv3NCSKS4pXnC+rzA02CNqFtqnusbjnZHBARCRB7VeiDHFeL3uk15aUbY
HazN5ByEcjUPWT4PKB1i02Aljb6o/hzUAeSPgboxe9Gyp9IvbL5hlzQ4e60qwS+uddj8G97fjdKM
ecYzGV+zNMZFH7S9yVTJOK1kUNysi5AFpWhRJsDt7/+BdWVyMvP/Ga0Hi9wXS68ITmb9cff8aO13
3a4qANcW8sRFcQzQN6oio46zEUfoZiP3Q3qrd8jqEcqCwqGH4dpvFfjFmwNEAyI/1bpRZs+ueT8V
Ywen0qVbU25do5n84pDjpg90EAfZnuS/nyC2ESXzznhVPJQ2U7ZeY2ONWHKoQxYrrhJSzAEb0ETF
WnRA221WMMkl8nlkmunv0yy1b+sF8jQHeID64T4pv3zwZ6Lo1UkzXRMojebVkSONb8NUjx9h+oys
9TvNugqE26KupoJDYtSHlH47njzDyBDaUhNAY8jNorcBqWsR2rRkpq/KjtzEqpRtPAEbsFd+y4Sm
RpsCRyrVT+FQxDgN5bDP5kRBmCmnv8qdEQzhUlwaJJnlwf0INpMlml946ZRvYTOLYufadqE3F8V3
sNvtweqxBJk7Br9vYAPyKcTCxxVqKzYmwz9JnEDHN5Gp1g6Xa2r+221nsxZRtjc69v/LRVqLP279
9KHq3FK0vvi4Ia0xOXEh3H2JDUdNIEOVJ+Gf+R8us8/7EElp9toeZXtv/rkQEo8a/hLAcb+56dQW
JrmW8q5FG/T230SPbBRKfbXQSRDpMSYfBbyfOMpy016gV1psxVLRffLQokyTtn8nIRipF0YcsIWl
jgyICNw18+1+Z51XOgIoH8Ykwh/zisIugAdVpnRdc609VGT0TFzA/WpLaIxAIEwI6EHnMJcUSPrV
IPbRqT7YN70DlfV0DJV6SoZgF0ZZJwrmKXuz0wtH5/koRCUa5omeUb5dJ3i4bmOLPl8Xyr7kj3I0
dqAxy0MZvR/vD9z8VzY2WMWGB7bSIZcjXevn2orzZ5sVJ+VP4ZSmVZnvDEq6ljGR/DcsCWroNaK/
/foh9ppYrJ1G2qKCesULs3dyKILzI9+CWPGAERnz+KobAcX3PX8VcgNPD0oiYFDF9p5Qceo5BI00
OPfaincRSTF9/0X2zkSppHhoDyjIaoxPbXAgsWem5Rs4PiMk0ghff7uZonL1fHL7S0QCcCOdVBLy
C4R+NS0SflEB4LBVmQCow/cBkKfh8UHdGEuPBSCs8XLuitmQFxr4tfHm/A/2l9DNzTqUtY31y7Ur
ZJ1jRoO7+TihXv2lq5seEkKqH5FrrUiG1oRd4BuI/AdgX2pEq8Su0RWVpFahESJsqFyKhufOP+9f
+sIQFVUMM0BetVz5MnZyQ4Elwdiy7PMd+2TifclM8J9Y+Ww3LClaI9IswVbiiH0s0yUg1OKu+odt
dSActdJpypbu0kye7f6s0rKdmOZcSI2WdN9gDjAH+8l8Wa7fx6rgamPRGOAHmiWBQiG2DMhby/hi
OXwap/QVLXX3YZP+on6kiI2tlF1peztIKcV4F9uW0hp9wsNFggo5USGvnp4HxN+4t24wxLEAdwW3
7kHOL+8tFaBnVoDAGNZx36K9EBxmNaP1K2eeqyfB/gYwAeds5VqyP2wnrtBZNBAo+IiZfQ0iSny7
Q93jTJ7wTnnmUPnaCBfFgSH8msQprrAeJoUpk8hRvua+bgIIww1Ipqi6Fdrjsj0qpTAC72u1/3Nd
F5JNRcjqPhApo2JPaewKBYiOhoP2T6rWCmyJhEaZgoxWeq+HcLRbNWX/i5KObtaOCjo/6UwmKRt2
Kkb8acXhQF3zeJWWuIsJ+MoW2TSx83FuiLYabW7ou3Kl4Le6f7zUWWUvDO+TZ5Dppa2C3iuwyjan
skOrEQ2is1bXTBAW/0ZNQyyro/ixQjW5rRQxiMKvOzR48+5Qda/M45ep4HINchGSjrNsRPc13RrI
jV0NbBDo496LVgsadN4bONDh1kuFkt0WcguiVM7JdeuE8o0tZxroun/5NOKKUzcm69w7LJtL8kgU
VpUvbPfqi0MUABAxCsBqiupvXOwLlzpJpglq9+hOx4ZaRuKmAjUyTyuxpEXfMJ3aQcAXXu01WaaW
wGSLee7I+Di+cyW23B5GHC8ehG92NftLnAMyY2ZpPB5tCbWK4i8/+7vb7OwBxBPqFF6wTPoEVCDr
1BSS4ZXLyd2YvBrUDnYVyVfHgGq0c4re3GzjDLBvrFxpezPZUmPX5NirTZ4EzHEAjjWfty1lbPE/
ZBnTEZXzjroO7BvENzftwgWcVSm+tO8pifuTFwZh+2ds+88yCEDgkOWse94kYrkD8TwdWO5waORo
oA8lEpkOXYHOesio9s4N4n8OTEyLqvjutK8o4YGUx1J48VGOYMLUXFmebltXqOvaqq623JQ2lHXh
F9eHBaK/SOErIlYh5O2VRuReMrtzDozfsV77YhIG+6gVgvwVP0c8LiJxQ4ZQxmwVh3di3OnoqGwz
Oo/ENRD+43lnm0FMpoNC99kzPGt+nCmz0GUzqTuIBnB2Fh/OrNUKXKtak5fnwXcNUXCj+YCcVGAL
ZJ3BEIF69XA3P3LjJuYVw7nLRAXtrGrHgQqZnsFr8rvxkzdIOoKmK+JWm66RI7rd/Vb4yq3RodT1
/G0JQR5kXkdxMnj7b8tvZPZkafdfASk03xUZl6KyNv8RWT1O17oDLaP5DO3C99Oy/CwMmJW7Qp+n
DzWTUKl7aL79wKZTvPsa3R7cFE4TCCZM7nOMh3I3Zj7gjFVziYbXNXrYMjZbz4s+pfo43PkG35Gn
UZrTpTJ9OL3O1QkCSPiGJsGIs0f/QF43Dr5kx6irQL27Yisjn6Azcm/5uoq1quYFYs2Zf077UwEL
KnT3JIG+f0mkC18F/HzLIEF/LTi+op5C81PgZvUWzCokZ2tSIjyoiOMfwi/ZoXyB8TiNd+x9IEML
JmFCSBd9zbpoP4DPD1J1i0JJxNg27ld/KRskCpczghf8GuyCNdSHzYTqYACz0gq8EAufk5iC1hGS
8DMWMXM3bNMebgLG/nm30hS2z78NDhP191QArcQ/D8tyKDvNRyrvCtw/JftKyqUsZ0LzdON0o+M8
TQHGSI0xkqWKnupV8v3/1GW8H5Mw37Uf+anHbZ3X+da7BXWSusfDzeVQVGBAKxiHdvi90R3gZmcN
YhqLY4ws3/0B/Bc+CEYgOMS7QChRa1V0qkf5AJ0zzWIe3kNTa4KZD2U0NVB8nKD+jUsYXh56PAMG
MZaa0/ssSNzhogD3YFdYbxaRrMM9HBU/zUHVTqMcYDBQhG6Glrl+Ra/k4niTGU0JlBOaEyOlIsJo
jlFE93Ug5n80s6u+FkD0UIzBCrh/jk9P5a1C/6iHhcQPT43xpb/DTxOjELzskhTceXiuj87/YVh5
tMEP4l9cDXcXIcCZ3M0Q+oO6cqEPoHZVZr6vR4eETq4a7vorazXi1l7OopWbCLpz8KtiQv2gruJp
yhfaRTfseOLEhLcJ4WrwGTv1W1CjLlV+XCcf1Z0R5Y+CAqq6rW2dw4BXb7DG8hn0yWgYOrnsTEON
rfDPkNiIQrKml1FYrk14kU4lMAKLeT2sKKpjW0nx+QXsyaxcyQRuSWr3omx5kh5hhz+R4on4V+3B
1AdDVLCF7C9t9FcrHb1ff9BH80hv3cjaKMfAc4MGEsNzlPTBmYS1oYf460vmx7HluD3c/OSz5adg
CYLEhs8Rdo3u8QPOS+lfQZ0oFWUCk2fMilBKHkB9AHiZaVHeQU/D5jRLd4omS5Reo/Gh+KHq2tWN
Eq3o1esrXsNs2WQoMZQf7kQ0zxK++Jg7UWsz3Msn5Y2hrjwtVd9VkTNTtMazWZgBs22+KL0xJzSM
9wHGyHKMmgSOizMU0KU092YQrpUXIBVCia1nn3nZ5GeWmrS9W/Zu+1xUneIygxMKMd6hrKz2O+2r
+45yIXRHQqUb6682V9LJBJ2hiz0g5ekXnVTi9rdT3Ljfm8KIRYGUUzMldlPx5XLVJBgVS8KhaKsS
a373hXdQa+wPfWiXyVYLIUFRus9yAAwNl4MMlQioW8oStoJ5wawITEon15rrX3KWJf82dhNaYw0y
oH86pTkPcHQRaVbfL0U7HlpG4eS8OGxuipjNq/56yBgszm1KFT2jjzzzx6m6mcRvGPmLQu9MgLiz
LQM4Ewwar/L/TqCYvP8Y+6owgzweVqcbbnS/i9CefKi7gesSGRTXfI5l5zNd3xj/4KKHDFwwp6jq
iyAWxGgdP+XKTVfi8IBmdLURROaDnlnh7GkmtrqrDiBIuFkFb0f6oDPY/JfLge3OF5zDd0Hp+w31
SEzsLYfhlIff2wTFUebTArHY7Hnk2bO+alQFhpL1J8ZFzmGqIsMCqgwtVScYPHkNmC9Hf6/qJqe3
RkY4DDWOBbAP1KuRSWd4x1Q96Sjbzbxvhb7sj5mrsNfwqJjvusSop5N4Lv/iRXzzaWyR1E2CWOph
Ae8aTTG4b5rcYbNZk+HRTX6kofBrMEcAwRx87VFGKL8Y6hE0FhXgzbp/YUA13pS3r1Nvy8yAZrM2
sYoUz+CMDOzoD7avoHAHZc3XbOoJvGTRxPhYkEiwt6JGFNOyD4x1jr5558kJxB6f+fAFXp4eAIL8
OIuBqUQGKGyQW32zObQe6PTgTwzC1PSuaispS6UQYJldkmDRPTTVf2PdS1wg3PAQr0/vjZDy7mCk
Lr/YNxpdANMAkz68w+XquqzZvywinhXLt5dK33oWkOpzGIpEFuNqPTlpozW544lzoNtVrspe6g6D
mSf4knIuM+OPsTCX3irW7sjiCt78685NapOcM6PQw3IzowkVjzor3yWr80wakV2slT3PlC29YmYB
afTe9Ih9dZkES6bAFZw4r3xvhp/bAiTMRFwtNJ2FnVrUmSJCQo2Iy2hmFkbylwg2kjOmaWsUlNMS
zFbdIAsv7fN+//tHBkQaC+aEMQBtD8kYg84txMVHZXaA6lTQQ+TXSZU6hwCDWy/HCrqa+AO8Qhjr
tdE5SYCJvgUg5JWDjSIgNT5P1M4usTYJNh5P1qg1CijQ39AAIyZLErXWq8HVT4Ep8eWnjIS0bH73
+5pYKJ+G5pU57ssv4R+/Kpa8DIqH0jj6J6m8xA8wIdDnkDbBu7lLTIORpFEoRPziZkDSdyey46jE
YT64YpcZdgvEClY11fpU0PLDQeCKW76qEeagBzaBb9KrgER7Kr15XCf/9gfUA0SqTuFHwWn92VPZ
Hq6DJkMnMv0Qt90brCRVqvcISQZFMFKz9ob/ErWXOFP+dx74/o9VW2WuhThXQdLdSCxgFaQGO5lp
rFWxP5vDboZkrvbDKuDiX3xH9Bscug8VLjkW4zZqj4lrcEmmliqo99bZchYFJUVloZseqyDZ/rEa
PpLhbemp/d08OS5X+6H17g9VYUOP4d3mahDPXtYInIXq9dD4MDzWpchRnBnFrrdsAti+1q9EUh5/
k7NLwhrFcykIJ4FZFmRu/C5bANqoEGUZbKGaNzhber/DMLdHZI+xIh34AFHBXigSD4B780fFNUU0
clYFYXEZCiNPi0BbxZUYze9jOuJIOGmVdS7Sp+q1VzPmC8G/wLzI7UIme9WTIxEtfvqwAUo8raGe
UNc/D01SSy8FTDYhPtRIVy73dKUE60q7qallELdPZe47k/SxVVk4ARDBkOsiIX24xkmwnxlpnIm7
/aruvyW9xyAdiUdjD1mxDdxVukspW3yihklDpooNZX1frrlWImuWwTiJxs7pmaZ+QnEGOTsxtSBz
YcTLmegDkdy59MMLktLTCXFJeuoTzkZ61u9YHtoIVj2fXYpjs2Xa1u+1JDfMogJR35jxpqi5v8ti
7vrbEtTm2cbgOpY0F0TFwubD9csZ5ZEkySQiAi8SqqjuYTYcsrR41tTPqCwohPuCzGICmuJkzkvT
RbxrfhuJwxEGmMJwsIWeLdRvIIhWhFc409dpSOR0lyYTfHdQfyvRp3SA39ZxBs8Px3lQZFBvA/he
XtlBWUNtDAfrzzBj3374Y3zGhAN1cmJwL0kOF9icPGEGPy9Nu6btVqEaMmqiUeVq/RdaRj20AFel
/s7VrPW377Roqnx+Faf8CtUyIxav7uU15keyDMatH8CL7tA7yc2EDUA4n5uXIHXottUStfSDVlnx
li0GwpANCK8Yw3phJb5bKfM336km8ovFGP9ZsmzwlPbx3t+jXuMfg7gBd/Q0rgARPsPpucleCgOr
eTDQHlKAqgOCPS7047Eli5wSakZcUBQjPpbZEF8caqPJUsxq+VtTFEXT4E3NZIwW9l0FTgdh+9Jn
za4bA1v8ZDx/5cN9h55FtLx1xwrB8gzYC10k9QcygNMtTpLUPUDVSZf3WZT32P3qjQJ31e63qYr9
CQCQhFD3cnEQRnwoBTPizTRtFDDfKDVdc1XwqttsCzbOy9XC5XozY9Ja86bQCaxkpe4xXhwhuOKA
jk0R7KLfSkuMEzZOci5bq/frjtJ4nrMXZy2/xom+maGenLRK5HI4wlkVusEVwfwXQatZlBWRba0v
AgXvV/jaK5wyv4Piy1pNRQP1XOZqKCdrM8mJ5JGHBg/PgjX3FH1Vub8seTWc3FlQHBZAEcO3Uieg
dcJqi98dQ+LCjGqptZFIodV+ZbYSIMqzk1k7Mc46lnRuFO64NuRZCOn97F714FIalLNYhVKl7Gfl
xeO885QBS41YXiApdWujwF+APY/TgcuTnTOYiWN+M9ZMntBMN1TeicFmqrqPkVHIC0FZdkSopvyA
JBHTFWNoYM11nLCOBmvaHRJeX3pl6v3QNcV9V7j8imHmmvPsQwfp3wjCBYa90Fy3TQJTbpUNVYYY
W0otUaFanbz6NCvRPCDrW6UeTUhxeMuD4PYUPj53NlHbY3RAcp4CDir1GaKfTz+8yPLn0G+1sMPN
CyyL3u4o1hjBfnQh9efV7RGCfTLAJz3cAnFnqyWfmY/hgdqcwZVV9jasOtnhUV7d0KPqmDvvv0nK
TXXSZEv4cMYh2bj+iWUSMHQFvUG+7PavCaELMZhNoKOblJlUwQqAO0wLfsV/zvBZL4BY0GhDH2NX
5+yajU2IyXAoA6ahVSFoiLc1mTi9yH1XloOCflcY9rzcrZqbI0QWcRv6L0EjY4ktDHk2TPeCvgwj
c0z6ZC+unejlkruEua1PhMJPUhOB43ZhSb7xelH6Cvi9QJOo7O189Gp8rEx8Qf3boVltMdYyd3uA
7A/TIdlefGRR36xnNbD/7n0ZEM/serMcfVXabl5w/BhBBVrl+Df8xZaL+t9Uh1zzvlNA42hJrMGK
8IypDrt7pM/qa21RBe4qo0r7H4WggF7FdO+a49GnQn/4VC0N1dJbn5UPWVTjrh1BBBXTHxgs5Hov
k28ITAlG8Yo0ePUCasGFOiuyqi9GL/wzA+bHdPO3wAl/mATs3Ts2+43zUzuaRlPGNMGUEqAgCG1m
4/5tQjRBVEMeNDOTpzraU94W1Z/QFXUP0RKLpYE21nCI9MLTly4zXI1DBbkU0SQFF8gCkvjQNTCd
ZmhFJcTBJd6HS0qRTPaWOvvsrDDBAWc8268g32y/pAbOaRVzbr1Bn/Tp9GjT92E7fifE9aUl5wcW
TJvZ1TToduo9ZeXqmAoH2ExYrdP9+g/LeKOsr4UyAFQpbIwkcd59A2R9gRWt3IkzPyD3wj2OKLpF
4NUiEWzyyK+rBos73ho5WMCkplrbos7VpoZEV4ffz5d6BCLqQf2iOrGidpc7htIWzWFXk8wuFXLe
th/BrXwoekFRVlEvBTTxkXCaBNOWKAaCEjBfiurKXDLhfmQkUar5jRB8eQOCeVkQ/PitwTy9KrQl
ncE4dYrDo+7St8aQfKFpVddUsHSSkoq7zRyMWBqRDHuLX4J24M5NF2IezQUTrvCtXuI20Rad3ZMz
K+ed9BudQfuakICAto73UZuXTu+fcXxMjwImqfXgRDNdnYEsXVqB39ZYneowL31EUkiWczKtoQ7n
X8B9A9r35V/E2HZNCFGfTUQ8M4tWuiquu4KCgDwhK1FCe79sgrUNnJmQIcmpWbaveEvZZM2XSaEZ
mTvMOE7578rhjiYR+Fc0GDNCEpJMOAn2A96tcs4VvYrcTpZMJBz4Ysup74qM0JTujX4s5HcK2LK4
S4PKhC3JsMQaL/5OZjqs+ZGDpeaeygL92DsR8BZprOVTakekVFHdzY56fOzq20RaVi0CJtZA/VZ4
ISxTTmunTsBPqZO2rjgTpGFwkMOTxnj8zd63kEQ50V1axp1tIwNsDYEuXkXW6Lq27F6LvnRxDSdO
FAxYkif/+JzZJCExcZw0JUWsLs6L0ML+oJFRBmEMoGjBzLC5PQgOk07GbR8v9mYi3PpwXs/jV9n5
ISOIcHB2mR6exZDldxHym3K3z8OoOnqyP+TeWqqY20qj+1U9cw9trnLkU59Q6Fa4dfwbt7fKO33j
PGOHBnN3/Y+c7GUr67OI/ScVkyNV7R6yAztlynkhfuvA3Eb74LrkRMUGeQjYITT7MpDI/dh1HrtW
6SUqt5YlHyIRAlMV0drC+VLj5TpDYsn0Yq+591ekX6nQEBCRc4HrBAk45jlzs0EFP4v8OcNQim+/
qftRhIy9e3HQU9N9t4REWfiZ9EtrOCl0rzcAeUH4jb1A19XUfINHHIuGEWGtwgtYSXmWKiLeVLPG
obUMrnpIOMJwLsHXo1c6oa/NXo9rj+WQov0ldR90MfFUOHFXCtMPHW1FZLQLDLpFfdvFUo0ufzWm
/u6uzq6sPKfji+4szbQIkiG4tUT1T8bGkwmMkg/EzrAwD+HqkGDackXCGnVCZSzGm5k+cMxV+9lP
5gs2DBLKunlW1mEtcBOusESHCPdrJxvtMk2svq3n1wJUi4MvApSIZDzvlASe0RadCR4A8Ytj/RXi
hF4zSKzHmcx3UTHmWoNGN7o9VJ8+8KRXCDGleadtlYr87QLv5tEZtVFogFwgPoPArfBc17XMwvF9
oJPftC3Pym/de02U+W9sxEfP6VoUTh1IpuXyrvsdwKzxOlDFJK8tVVCKCDzH4olX47g6Qr+/JIwx
M+ZgbirJwn8TIIV7yj78EZjZ7NSi+fdCZ1CZsFC09zzvB92Cf5+GiUEqFO4ipPzHMNwi72w/oHDu
NoMcoPjNbiTM7ldx2H4488FomSVRztCDe1/Hui6rnbI+HOgXmGhYnn2MKagxvxsCQAyv4rom0nc6
5d7rBIqF5LaiG3J97owfijNLkRYx8PeIS6njffothOjPTfMr2SBwR5vTQ30ROtL1IXwrol9P6WHy
Cc8jNAf1Zr4ziTXVfOvHaphWkmZBCTWSAd92/VoKopoyHA8lsEjIkSHQ4nvqL1b87FegT/QNjx9W
20phYDW3veqeM1SgHtFFw469cQfmUSV5fGuPTmpXAuXMtd2JALjdq0oO9sY8d8em829EeHmQa/4N
+PsIrKI3cCuXhM4ikdtBMppRXq8r3Zb8NncG3DtAzZBS31I4rab9gR6M+yE9HZqRc2pskYrwS/K1
LT3xZfwZW9eQCJR8jqptyTV6jCIqzlfYJzvXMKz1xrTf+uo7Kww8llnGJQ99Smt1G7rOSi4H6srL
bFaYfj6CXsLFmbfTQ+SGAEgIkTuq9iLt/9o6QZJNTJvZDXKmg/X/mtpQHGZm1itAlC8Mcv2ig7b6
c6F/GquVVZE5Yjo0TO6oSka38aaG1BoV37nbVyixFunFiXk+LK5w1R5ZIrec7YWWXeQq56mWFGBN
pVLDKRG6x/f92Fu/JoNiDcoZUKMf2W7PV54me8/kJXydqw8fuGEqfjHfEwPipzVHDHEsSi6alnOQ
syroitTtK92e+k77NbmiP1WPejjK9rnT/1+p4MWxAMTzfmvD5qJfb3ixO1boa4+crtC8Z7gZYALX
D5+uzcoo1P5J/UMSqfhkyVRjlMfK4G3v/PqJck9ogqlYPamY0tl+8BmCnsXW9g+ia1AxjJzyUQme
zdED5e/HRb91sZirVS6URhV9yESAIlwtqFvRrSrkMgLfc0YN6vAubROf3TcrjveTjAVKRjoH3Gjs
eoLvTulZZX9fguROeOHsREWVqXfMbt2bJqbPwG0wG6VE1QHlKQ8NCz2CjsEc5KSU0bA5WyuS4C/d
88hTunvf0p+ICrXtlxq9vl/YeTgBLFQnBQjfRfaxQovezlNbb5yZZ5fdUZ4OsRc6IxUCRbIZI6sV
p68c9j6bo22VOBF5fljfEcNvv96i0eYiOoBfdjcxutX9bo9M7+ehLwPnvzO/n5fdFb19Kr2nlPkC
kTo8BPWMkEHp0LtqGMHJQHozXiN8JqrttcoMv3OzdC8pI8zgEGQgOrjDlz+OmL8QOEFuzG7GFGWY
Vlt9s5ep0AzTxV84q5AG0aBZdk28Bks+hP6So5woAMaxnZh7OX89QhvXlGZo4csxzlCnm+KzaxQP
yDOqpwfBsQcDwwSPgGwlUzOaX/eQxUnzCiZwcevr3VCVsVbEsSymhFy31kx1STGxqX5IMlasdiUj
G9huH5Ptr4/ztvgX3406KB15Wv7pKLSpXYAuCp5MLTwY9vwO5olYpcDHvNRIO2Ev4Mj2lpsntMzT
glcwQWk0+aQzPBlH7qUanGDOg0PkORdUE/s4+bY9mNUWxnV024I85uA9VLaibbfo0VUsst/VO8aC
rpwe80MJIRN6QkEaVD/gU6pZ+9G38LXPdzX45hIU370HtXKbh2NuY9kMuD2CBf0GsRaCMqPYeYW3
2iRW1G6kiTBC1JsHDUgU3Ryi+GwUb+XYeiFnbRbSuxwz656dey/wLVn36/jToBT6F8mxjVcJIqNA
Cef7uCrxZFwoYKWOm/cn1ooeNqKsa5aO9CAke4DCG+HFfbN+mXaeb3T+OgA9iij8yGbKuVTAOo5c
rnNDNvRfj0QVf6k5I0pVCGYiAdHOnpdW467FtajGg8ea/2MooYQJ3Soab8t8hzhlEndjvHt5ob92
IqheDp44ImqP7SJG2zh4FSNFxW3I+uBr+JjojA1dWUVV1u0e+5TBziMSoyBRrRLhlMpXIAiDXq26
H0juota+Nl44z4TQMY+YZ+IbVFvrjPsVALdgLlAIWptAveJz+YpZHBcx1mN9p94rVjszie5mxgXU
vUWSrwckKIHqn2B/1R8aRloqsUjOJ6j3EfbyHIgEZXfq5r4cr/ooPbChv1rNi1ETUYgu4lWO3N5k
W/w3Agrpjsl8SAgIEmVaN1/RNJHeNb5J02mhZHnwFYulRTlKRB2s83aIClSIEROOBm6o/xnX+RGK
woo4aqIp05jNrWspj7acIiK+rZg4SRu/bbd2wlNCgWoGU1SLishw71C6Nq9XyHsvHfFn1k6wQKzJ
msBU55te5kggm58BWnaCXo5D+xwGWaU+n6iOe23sflDscSlnIX6t9H4s4W/iqeFeqcV1bS3bnuV4
yAyuH4UJzfng40L/rT61TZHPLvZHr0EdWzNGga6bQzrzqi2ki9900nbjMwH1Sy5OIzQHfmgQ3EvC
pSgeBdkpHQqZ0MjHNyldguPzPlvobNQZfppz7n/ghWD8TT4fUOrb6Pv7Qx0IgJxIfO1SxJAfJGrP
RIpfU+SbPIIdKLLMLee+p8WwEGiUmT4LUWN2EfOZHSK/gGq7YMXFyvisjcek/YTbWFsFI6XwMNLL
Weh9GBi0k9DdWJFEhCtq0QmZ/feXlKaeN/l7+TLEVtZZQhnu1cQxoFm5sfXYNHDUhWdrO9RULmos
yYzMNYiud3dojc4RVS2u4xM8MgCfGaoOGGn6HsV1/jF+6LB36CaBFG3ZiwV1DThXUxqNoybYz7WS
bZOVMVxVMcxg5FW7y5t1QI37XGZQUMXDwV2KqRS+j/uwXDqdbxGEY9sUHQpAPpAJpgP/KO7M9mT8
/B/NFCiv71B+qt5+z+uMfQZTdn1ee7NstuKtyZy/MpHtXnkQo8mIZyPMswD10O9XAZ8lFOMed4k3
LPX+x87etgAwnqPxI4KaDql8t6YGr9tqC+ghQRRM17JWFq44LWuPxRrpuqh/o5yXjBaT1EL/qyWF
DU+Nqv6uRx1jIMwNusGe+Q4i10ob4LU0tAoEgJfrbC2/flUHqZ5s2Eu3moWMgwE4ZWmzWx9+R5Kk
HG1XtR8hG8jbq8Ezrg6WIuOPkPsDXT1pz+D04upjVoXxBGNKmEjboN1+3S0vHuuRb2L0jHLYsL7P
fKFc+6k3kSkulJgmcFLmuwdU716JK4FsOfejSK8ToQD2bpvSIbeItKX1K4mEcn/e4G7G7fj7dNq5
soVXuB1w4xWKHo4rXJ4GwtDEvHRSFjQqo1UuEKyf1Y1BmGpIbZIGgKv2+yQ9P5B9JLSbdZVhdOkn
Dhoff10d+vt/6ZZsoOhqAJJAlz5mPFaieULCudilZM878RMHwjNNhAKTg2jDwGY47ub/34DeDnFh
lkWFttAqOZOdTVCRs1LhuLzw9umWNfSoJtbdx0eXpDyvIyl1l1M9d+TFzCT80dDL5bKaDEJ2XkD1
ABbiOusF2W3Xknim86Qutn6GFDi1sgtbcISIAy1FzW5qjmsBB/mXWMVAicA0J6NsjdxhunJxqEYr
DbirEoANBtAXIqLzCqslVLkKKF8p3LE99AYx+oSoaXFJsKrPF3rQya3CXwDThrygz6xlkmwZ3j3e
jIPHxc+5dVLftfskDwflT6Wx5EP5pxjfIqoGhYFqqwSBnf9qUcvaIjf7jH3VJdbDIp/szUyFkO0x
bi0vU/iUiq2VmkUbhH8CgGdx5wzjIAYg+H2P93QimD4GzDoqDFebuOCjxjX80m4ezfFrkeAHjHlA
T7wCSArfyTelt2IBv+Ji6iuSf1JkxkLjSaI/ibzrKCGjUFBKXwGG1wWWpDZkQdPjEPuY1MWcbClS
lfsYCbj2uwU9va4l/ZFBuQtjGzs6vAwgGUo+oslqdAKfecFFTy/CZFIFd0s3+BS8IvecmS+5Bx/v
nz1K4iTJHARg6uaaU5LQOh917UOR9Y9B4rPeRDgJsxhW0s9uSiOijV0GhWlwznyDMDetViVnFDCc
RCroznR9DVZXIBL2CayZmDJZ/9kGayXkOMw13Qmj8NhZbZS5Ts2bnqrtPiiNas4areXFH7EL7Zs0
PCgIe6LJtwZIvQV3RMKes4RRl0jAv3lI7Ge32WfLaENVHLL17Z+HKgGrZXoI8fh3EGi2YUoxPDJy
hmSgKbCzay6gvq4Tn5kNcGnQN177WPtoxaEJ7kA7xeeceaP+nbcwMdISES0yeHOTtpSQgQbjFgaX
IDXfEB3ZKzG2CbLzvlJ+b0HMHvBG6pEekQ+FV8ueoIi/RrYcdroKPuciDfO4Kj94+25wNse5zJ14
y1V+CONCj9Yw1tcTs6I8+B5530A6rvTogbdps00RNzVe3pToPkyRY9ess7xbkUQUvDNDdy1hxdDB
VIAi27EOvufeJTYfseWSv8HSD1lu/DNrOYSyJmrHGlZeOMzKLzKUHbAPRmqJFPKGyxDwGrNErSwj
nkwlCoRotwtUkw9b6uRRVhfaAPjKjCiibo1zm/UmZTDmaya4OFsqg9uog5gHYDx6utk03GHhxXQe
UZClSK5cPYDGSQNNHxMJNQy6FIZz9pqpURuKwRIxP0FbWhPwdqmZOlLo+sBz0n2oOCpJb/c0tWG5
stR3QRbeRZ8xlI49oYmYzwD5rkL5007RasYhaRNHaixqvfjm1hk9IIPtDyZJXB5xtc8rhwx+wmHL
FhoxBcFtjT+M2LJHiYyNy+WiHZ6sWa5m2JbGTZ0wfnkKJdNnifiod3yWOCiTqwZFGGsj9hP1iQkv
ko4VERSaVIzYIlE7kDRaIE3sA5+Mjrzy0wGvwdXGqmwX3/ied8U6ArEX8XdZST3bjcOFd7s6HjkD
dFtUD8IHn4li/hin4HWk1MKGxPFVhhgF9n5uqdf418ElWhzwSrN00KmPS0/LcHm1mdFb/A/v5XeD
9rVdRx/uy++Sm8NR4WuvMG8q9r0tnriMwkokkdB0jwQ695kssRFsKauN9C2RhyoSzspfG7ROLv6u
eP2I5Cejn9MIybVj51R1DWfFcVDaEIBFtgd9UHl2AQ5LYvoK3+gPVZ7DgBzgrgFu4EpN8Xfc34L3
5xo16JicFgDCvuE527l4+mJLqYUBPR0KAiX/4MyOZxlpwknYakA4/hedWIVTuZn0XgRt+rb9rdQz
VHPBPBaffZzsHeSO+1gqmuuEK7ccdM83RuRXY40fDf93w84c4nLCnBVCAGD9jD41OvApOhcWfTVN
CYRe4WhqEI8vXAcTizjPXOFX9BgtFPfPWjnZkNA5lHRVc8JhJ0qq6H8uFxQ+khHgEJDrO/V5tXnQ
ClEEdBLYMGyZxrEEZIoJrcQEE6LE3MZHDz6BUE5HZ35gj3kDSKTBx8M6nyQXuRBf66dhPBcwcp2h
/QGKC8SNhA3yCVFtS3hQ71z7X/FO2P4d1OaivZBoRONNy6GAzLFdvhvcrStLlMFJiMIBulxyzGXz
lpjiCvYB5kCjPSijVBRDhELrRNxu+6ZFGDURp14fsw8PV1zdjn+zEFhtcGlibvCf0YjeA8xt08wg
r8kSNUXeeTlV4Nl7+abnMRcD0FQQ1tAtZBhYb8Ji/2OT9EIf1zSuzudhBf1t3ZGQyni5EEY8IyqN
G0LqfnPv6kb5mNx5ZuuMbe3VgdKekQQpDJXD8WUIRZBpiE28+kTq3cWUY9mkVLFlOXIq6bQksG4C
CFuTusd3alQWtYNnXDDqGnG8f4Q1I/g2/2P5y4hlbqE8vlReKtLDZ87zg2Q6xP1qdUjdWN9zCBan
8sApLOSZjKelv+3uspJC6onfd8aCP/XcJxLOyEv5we159lGwZJ/yZajFozKJEzWi2TtyOiPQl+VD
8v7TCCAXJjYahedpNLb4JTUMDhWCUz1Y8zhWw6yySGyZENH3GwC07xdXS+ICo8TgcvvtxpbjBtHj
5WWpoCEm7hCi/7Sx+vyZhS9iI3a+XH53XZ3mWH1LcXeU0aPu6DnLx/f8MLoSQ12lS8haSdis2A7I
TuDKCQU4W7b1cSCeEMUfMPLdiHqLToI3XF6PD2+/YqSY9kL/GwgGnmNdQNAqr0nlkNz3zuIPhGu4
ZdDpja/q6VVDkgED4k4bplU1mj2Vg/GWRrv+EGuSTVrK8qUBHRj+53+XCT4W6otq3Ipw37R3MRxB
05QVtgNIKFczfLEm6rffhlSZb7FdpzhcsQY/UIakOeMh3GUZiG7m1hB3I5ltLb3x+6V6d4XCenIH
boPiUepMb2iKHeX3DNojqbkPIj9yv3D2yB5wQauzohKl5nyTftD7Dbj8bQOmCC97FD4eD5/Gptg4
SORu1vxFxS/sy7FGHlEAMuhAX9bHbFTC7lk4CZMql01gfpzjVoGqwQAb7pMx9vspflF1tuA0chde
y4H+MTq5CA7vAynouEyggenmM897f38P2NNRR8kRFn6+xOO4HcBAOQ+fux0toJyKv58/S4GTC/HB
Bzm016QHrjUMTGewEHDMnv/PzUmeTFNy3RQ97ODsezpCyZmN7QvANdoMBY6Bi/66tM8dohRukqH/
APOlUGeLY7kLFnCzkaI+xz9exiAWF4fxFDfFp9bGkm0QhtNTIOzL1rE8ifS3qZX7bdVEAugqjch0
yubnIRavJKN+Q6SfbShIwcvb40zKZVF6HYqOk9JM5eGBwBZZ+Wi3+JsfLFN9lXcEjX3CI5o0M/Bw
a1J/nJVEAaws7gL+mxl8QhZCLM0lJuLOhpz1Wl9qf2nLj5neOymMhwcHl/RGol40u8jMZzc2E38Y
mFfQO/4I6THPWDILbqZFZe6RqwMJIgMCmMcELmmgqDcqrQtsQD+PNM25ofQpM3eb1wXvL8l94UZS
n8SSxyFCGpvyQblFc8ZvthB6zK4isoNqT2td4PUoy0ti4euMohQfU26OnS3DaNunXn74iwJpgi+H
DzVcHlu24nTxNzLzgz+Pf+Z8XmwjDSYxHalLtJrkrdY6o0LxABo7i1Ws8xFi2FnG6C2RJaxyNKWv
kD5ECI0Pm+f7xArOD4xFH020F9ARwX8kuCE8bWKEx42MyL/Z2FpwMnN3SyG0TnZZ1eQVnEWVjRT3
VWOaaMkdwrYq0dUZagUpHteOHC6kc5iQPa5v+ZG3U00yBdV7FILTYf1g+nQnlnAhNHuXmWgiT2d+
UWJMMrh7d5czGWiIl/OF/ND90inAMqNIIGAvfP71W7tZQ6fN83ck0DU1puPMEzYWyFJCBWKaAaZO
rxNEBokqYrCe9w6uA8RdMAfSpsef/0NXvGx7xq3tN8J2fr41peVkWkw3LGunrFGJiTtOmSJSdvqu
6sLPqGkLstpRIveAgUXJJZ7ygXoBSQya1eWmmKjxbN9k9W3Rq4uqipUejSon44kkb4FvZF2DNtKQ
g8xgSUGCHQe3w1c6beaehErxWe+lUzH1kIyORDxPnpmmMwVEsaDW8geKEW8AFgNaZBooRlHEFqbb
pnXY/vW7aS9jWvDbSMn9xd9uUhpQpCQ8GiDqLJyG48o+m6mvFx4MR4pkSA/mrS77CFyxmJevGqOM
2s6K1JZApMVCwxdk/1PMbaXHmMnrgjqKGZ/EB8h6A7WmJKRzKpvo39W0KJm3ZtORswYxrDa1j/ZJ
NNNYzl0NIpHjGVdoJHv7p99BYkYpy/+4X7ufFVSqmHJB9+LlB38CFXCaY9FiNtVcOptLyhfNUY7X
wtfwYJMCgxa+MvOVcxqjjUvzexPqBcxUgnWIa3Bg5tt5MMQZG/oBNsNZniVcQ1UnX6izNog8jiDu
nUxLL2WK2fF+S0O7Q5kPbuYyprC5sfHyaBiK946lRwcuYjks6XgD7V7MvTtaYTfeyO0kUx56oTP8
BCvn642Icvpd1yeV8jsZYQLeeLLsSqwFKd6eWRBkgHJ0Ur+jo/GyK1M1TcsI7LuzyI1AOEBkVHMo
AF6SBczad8eauVeorywrGPZCRF7KdXqKG7Bh41navFR9I8r/QyLKNCVTioEpp+3mrpNbGJ9RNZHM
yiqSb1c9C/kRAOx9112C1N0MN5UrV0pcB03xil/VzVU4A52pOsFCMRIbj3ONFQEpn2ma387G+y26
Fkn37oQ3RwLbAflIa0uEEqZXFzy+dmv1RbDXqCLzBT2oTmojNyWJF5rIRmbRdYJhy22pSRGEETek
M0Prvlzuc2f3b8Fu7fz4btoCuWfWQ13Cb+tIBv0c73vLRjyPa2y3kJJxCPgpkIsuYr312v6HSjUi
hZLSgtIAXkzf1CnofcHgfRST3qFRkarVvi1XRkUrE5hp25LMYTZonZQ14cbahwbJ29kHU55CeXmK
yA1El+WZDzl7krPipkYl87y4LiWnH9Qf4cOK6zvOLeClxZH91n3RncA2hwuemGaitp0v9wrlNEzW
7tryucf0q4BoPZGFIXPNFn47ll5+LzGEEVJ1xU7xsab7NnkSgINxc5+gisT0TzL2t8XBqxouyDlV
mU9qAvZTzWwf4L90jFg2Tl/QC/LezRxsXObkVmGaHQECjuGGQ2pn12yALDygE7Q7OyVtO9aHtjcf
rZIzczjm72eMfS4X4dLcQVz1F4HAAYAgmvjW9GRzzkRyER/qdeHl6XWvCmqXFY4wRqLSbKAdeMlM
KpciBHhwb2FdmKpHxFk+WexsK3sc92AkxXFXV7AIeGlIQCDieBcCPJHv+iBr/cmVY0f+3851hwCn
K/cqlFkoAJ5QHtiyoV8ymu9s8DFVfDcFLghc/IKKlvwN34t1+/+YHFrK2vuvqtxrkWDTR/bICFPz
WzM/u4QltHPmaKHi/YZH+xvck/g7Oj4JT8NuTE9lVfruRZisk8f0eifMO8rS5fMPw5lGe1+k0syF
0ADenEWsVoKadCVj4rqj4uSAwISTZPdkKxgFLe/kV1uZtNUbbqMExPz+QDgCffVaCnvcgss/tW0R
KPiCsKbMYjwrWfP9+XMJ1aemGXaLllFrM93UjhWN5i5mrB3kSOWLsTelPIl0X90XpNCFs3kJ1k0v
b9DRgNlK6r0SgDffvR2q6/wHY4BqVR9dc1fUMTC+pe1N9GjreJNkhN+gdwrVNL7qy1hIkSYxEJze
C8tZskeC/httIxBfOJLBXiBnS8DgHRKwoaXNA8KJ+KGBUTnkXc+Ry2MDhFxUMwwa9mHFRDGX7Aml
MnXEXYz7nlqC+8TDOMTQN/NtqFhXFHV97X3pRcVtxZQDs+dsoJjg4qFP04oIXfZFV3V3vcnx+B/X
amBh8OtPwRtgdHD/4YitSBARbpC2g5ZewjvsbmskN39S2+dSiEDVelVRZSLAlh373tWRtCVj3bp3
RBsaF+tAMh0EUFjo6wT3qst09qtQ8nUFY3FOngJ3j+ORorEhXXSt7P3xG/DWdW09UatGjXHd9jsX
af53m6cQIEXEeVO4VuyZuEjnjls3Z5/A03KB8NkQgGJ9421hiUCzvx7i9IeO5+0mLdAftluRNUwr
ZxE65RUWMK5npOq1FmZS12cYeU9slOjt7IBYF3VPcHRtoVjJPQYEP+dKkbXGohXHy6ZEW9+9H0qU
oU0H1CvkVMy4PQq0k/WUUvprcXIbQnxc3jR50t6NQJShCLAmOeLfoyOxl9mu38MvSzEsEolOt7CZ
+DnSJV5LdM5Jg4Hz8mNSVTsRZ2AlPr/4rc0kcACwY+8Uwmams+AtG4lZ5A3QFQ4qzFAyIkyUhhb4
WULUPP+BUfvT3SCyuz4B4h8PDGoSXecJBaWb7pZgbD6BOZAPV0S223Ga3ye0cuDITPsKCP/NCglw
5KP6G/FGycQMmCrfVW5BPB/wLfrBZ8QfzobgyliVTm4oOJF2jaFLWbrlI3v3c/dZzK/Kij54oBvT
rfOY5CkK0p5NPK7wjj27B54/28jQ3id6vbKlU1pmPDQTgyJSJnSM6iatZ7+S2SwumFH68lKuiL/7
hib0aZ5HbayMNd9oIZFZXPIxh0nGuwp+v8OPA2eySj7N7jvI8ihReu9L3L51bNk7B3iUqcHBtG89
hhlmjYLoBTjt4+MKt3pt15ZG6rHHISUVzLzAKoSq9aX9skWcME7MuHG/76vNCM0zwJYFTu4PxCit
0H6CpwHoZL+Jcoa/Q4DthXkjxh7WhKlPmVMb2czD6FBruPBONMlPnLu7BV66/9oP0ons+8DmxzTm
YOKq7eZJqxi6lS9IPlHXVaqrpjup5JieH+hu3pbGF3PaMDpVi5C/b9SLZg+MKR18vz/OPDYgF/2M
7JReYv5DJMIrwmSbRLx9WdqQaYTTFqwW96RTEQEookPd3sQb1xmkD+mL3IMO52aposfSMFboxHGa
y9nT0jVkcYIFWB59RjZIiTxd5Jkz7CcKg9k2Zwn6iYdPAUAcuA6fkjCQ7JwfFxb3+nRUsPVODqOT
w5D1FcWGg9VPektVKZaceKmQdbVLBO6SPuMGqjvDvx4Kloni3UqfbQZV16A22Llm5owW8zzHh1d8
CfaIBj454jLjem9jp5yvYm99vhJo8953c1etHgi6aKgDpVcAuk/J7m8WO+rJCYnZN4TIlNV4QJKp
BlDg8kFh3AKj70+y9S38xePQVpS9LrLTsFs82H35cWgWfkLq69lb6Lgy1Hu2ceSeYcN4KXMhG/cV
Tytp4+6prgLHic5hNkzcHhpvqHLlJRPC6EzX+7qNmWc/jWqBsTSXLr3zuDYNvUxazaRiCI2yEOxp
0YhmujuPBWtBm+U+z9AzogFH1L74M4BiCIZaxI2U1SS9x883KFBNbSKpiPPZc3+oYHPii8LUQyas
RRhXOt4ZRvR5yqJKw7o2al0yKF14lGQTY7HSKmOgFPYtm6amEZlPPM2OTE26VoKGBe5bSz84lFq1
hQijQTE2epLMbJS4jiviDltpRCYuFald52mlGKZOppMm0b6wuBTvuzM9Ij5wXZNB5Ghplu3Z2H6b
IWm9LPWsRO61oyREENdaBB5UMZ92eboaWkpp5Cm9/2cKxUvvO/APt1vaXrrwTZZe5meNyiQkfVN+
OAjO8Bh1FyYdZsXk0iOxRi1n1b97SQMTIR7r9DD1pdLe9FqWwNZpQp9Zuxjdj8dHjFhBUoXK4Ajm
Dw/0GUG3WxTGcrTyRzLUNSkaHKpbaza54+WNSCHfQYG7Rg1BUMTB04z9y+pIaTKrc8I3UNMPLE4m
CguFr9aFkt+I/qc9gt3EXbE+sXHxszX+/zyL7hj2xjXxeMVpdnpyUE+T1uqOynUcH5kZHGNA4RjF
GbAfjbdoih7aiHXi0g+VloT+MUF3IYVCY5gdEzBrBM1O9qW9xHgeB2UFkwgrAMIRoiD0yTwfzqP2
Ob/Pus21/C0z/eby4npKveukdHZOfJP0opTPLGEexNfe1lVi/qLh4ez+lLfkvWgL0O7Db7TbZn7l
YvcWAXGVssd3HrZcuiLCbstlku+ewaibv8bTrPJhqGRuOBjxnkk6rnNsfWBO3761c0tpCMLW1hYq
bDmCZ+SNYYShxG1NCHLrlX1ZMkxD5Ln9LK+FZb2jXUAsGZ9zFqEjb+5TZlZJP462op4sIIjEyhrG
x6nYovXzVXmjlH9OwjjNEIhp5AfDsfnea2fpd8gz6PLoW+t6taeINZxRzi6rttWTnXVkSJYVwRI2
LpM+6VLj7pwTld3BtF4cOvhE66lUkF0B835XZ2CyOQbQAPZRz2+Sti8x3M+F6F+dwCO2vkiKevl3
dsl6kvF2n0MXAEIR9R0On4bVOlNMW5GxjZr83JzruFxG2zXUAOmkJ1uy17g/sE9xa97iRFFLF+9q
PYPojehegnoAkM6jO8mtsVtt3FURjO8Hl1PIfJY3ZQKjJSVNdBGgHO4k85lx3gNUWXJ1F+EeeMVe
uxQAEGToCnhEdYJMuFj3X/oZz0E7QNj+XWjggwMAHXfCAjH75wDv1uMofqwcYukvMZzbrlKop9DA
ZyOw1gRlXVqJ1nAo26Vp+iHAbg4zcNFJTuPmQ4pYYe42piTEAlAl+12hfUZ7TKihncyMngPVTTLA
HtBkLjBT3xx2rjx+Q+8XN2sOAYdiySaizTtXnaZVwWmyOpFkxUjn1XppODnjsznAfzZQ8+E4MTHJ
YDsrPrOWCo7hDxeRrdsQI6uTjRJAIZcyNa2M3D3gsE72edLK3eLlJpDkUmQR9bo9Qdg3TADc3sPh
icQvzLzBTA3NW6p0/ZRS1YxzrvNF7JloQW4rIhelKkR9PswruKKrczfpFaUC9S0mGXAcSjXuLdrw
PK9M1+90V3tn15rbw/tpdXUadI134JNMYrqURTfSSTcP1yo0RzUFe4z5M5Yv3hqvz2Jhi0Wk/m17
Gjtd9ChRx/QwEJt/K6z4HSzGsIAmieRlYM5Kckyi/EMAm+O4nCcQ+SPA1ZTHX3fy+3bmNJywPm9f
txDgts4mnDR0rH0V8idZVt0sNPU3/pFKLuv7e0LbhMk36kGtoRwljm9d73VWRDVODziS5uxDEBGm
I7uZ01VfK0SjTHdUvGf9epeMQCIQtYTmBsWOT5LDwgPkA3kXvOOQUcs1ehyVKx94G3T/DiF0o0b1
nkIkKv4EK/pu+EGY3PjCkc9brIhiqymyraX9QP0P+uucTZVy+4s7g36UcqbPL4JS31iZnvddFVjQ
c9ekUDoK5MNWl0JH81YejtJD+aXAeR3cJucR4/HOXGabl7cQRQVnWs14lx4RhlmC/wUf6Sc7MCom
tsDaMikleRzsIDdt0sePF/HVq7/Jeh0GnBXi4cP6IrM9F79K71Xgmj5yTT1CrxrXdWmNaERx+Lqs
ekzF5yh0qlOtnw3w/68lmpYQsq5XMFpmgoV8jGrg8lMtdUDiPJgn45xxPG7t4y9NL9o3lG6+SWiE
3aFr9dAMKDMci/njWTRD8LJ5tgom/tACtM0bUMs7IjAudp6sBwAtjTdvey9Nsmk0EqJUNGDup+Ri
WFEoFTyFHNHfSxiCW3+SuWaimQsyuUr7MfvR+9YoybORBg46nL0tbkbcUz4ghY22I4IX2xSDNFYe
CKyOeSYjGOx2mGhNQoGjXVI2PVJGaAbYftWLipCXf9IbtbfyOQLC3U8ecEF1o1ykf8v8L6Rg5sWE
IeNbJ4vDiLVAr9GTBtH2t22ywZf2fX5fOG0ug3o8ncM1M1uuaog+mvdpceacUisaBVa80lelVhQP
3e0a848M9RxHEAEWBWJ9WyU7ii/ucO7dtN3jXalf6zGZZHg3ciNxIF8PLxfE07ntDdilzq05VcH2
IWH0Mw==
%%% protect end_protected
