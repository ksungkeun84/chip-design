library IEEE,DWARE;
use IEEE.std_logic_1164.all;
use DWARE.DWpackages.all;
use DWARE.DW_Foundation_comp_arith.all;

entity DW_fp_div_seq_inst is
    generic (
	 inst_sig_width : POSITIVE := 23;
	 inst_exp_width : POSITIVE := 8;
	 inst_ieee_compliance : INTEGER := 0;
	 inst_num_cyc : POSITIVE := 4;
	 inst_rst_mode : INTEGER := 0;
	 inst_input_mode : INTEGER := 1;
	 inst_output_mode : INTEGER := 1;
	 inst_early_start : INTEGER := 0;
	 inst_internal_reg : INTEGER := 1
	 );
    port (
	 inst_a : in std_logic_vector(inst_sig_width+inst_exp_width downto 0);
	 inst_b : in std_logic_vector(inst_sig_width+inst_exp_width downto 0);
	 inst_rnd : in std_logic_vector(2 downto 0);
	 inst_clk : in std_logic;
	 inst_rst_n : in std_logic;
	 inst_start : in std_logic;
	 z_inst : out std_logic_vector(inst_sig_width+inst_exp_width downto 0);
	 status_inst : out std_logic_vector(7 downto 0);
	 complete_inst : out std_logic
	 );
end DW_fp_div_seq_inst;


architecture inst of DW_fp_div_seq_inst is

begin

    -- Instance of DW_fp_div_seq
    U1 : DW_fp_div_seq
	generic map (
		sig_width => inst_sig_width,
		exp_width => inst_exp_width,
		ieee_compliance => inst_ieee_compliance,
		num_cyc => inst_num_cyc,
		rst_mode => inst_rst_mode,
		input_mode => inst_input_mode,
		output_mode => inst_output_mode,
		early_start => inst_early_start,
		internal_reg => inst_internal_reg
		)
	port map (
		a => inst_a,
		b => inst_b,
		rnd => inst_rnd,
		clk => inst_clk,
		rst_n => inst_rst_n,
		start => inst_start,
		z => z_inst,
		status => status_inst,
		complete => complete_inst
		);


end inst;

-- pragma translate_off
configuration DW_fp_div_seq_inst_cfg_inst of DW_fp_div_seq_inst is
for inst
end for; -- inst
end DW_fp_div_seq_inst_cfg_inst;
-- pragma translate_on
