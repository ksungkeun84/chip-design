%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
LNAJoirHnGsDKLmdF1QI1TfmnyYrQbuauKpM0r51UoXsQC7P0RvR0TzNa+te5JOENGCW1fXrFK/2
3s0nmbJalkame116pv5xhwWRtCN/R5sgB5tgvxAkE6SSSKuAaESrprPmAefwt6qJ9UGOp5oXFJSh
34sunBukVQ+1p5mhrGXMxJQBjaFpv2UiRsnqxaeunyEWcGxE0jXS4F48vJH2nP9RjbUZqKc4kBBC
6C8LEL3rrb+ecrStCcplJTk76ctViaEXFEe8PoFhOhbg78F7D5Jw1XzE7ZO0gUZTh2//tMsq5hB5
ef5jA8dRnEF+EeiGs69SOLRe8mlkacjCWkZKTA==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
J+bilnW8L6/fj0Niu9OvzoHCTgnQ8GzQ/dpXLourDs49A6JjR0zozdc6q0oNJJsDy5bvt18r22Cz
GC5TCpq/YMqZGxUfbvIBs0iJl4PLjCi7xd0uL6UxX0QcSt7lax37/C/NDP9T0+SPWbq0y9l1Svt9
VvWOY4YNE+q7YKAH7GtvbwwQWjs4MtuR37pjY7ZffF0ir1Hy/smwmJ7sNqNiydZO4TQOFAN/CIxx
LwwO/pyEwGFx/8nBg6nGSZSStEZ5E6IbJQlm3a8IV7RHhWwfRH1cqi3MEfP6wXm7pHydrnFdooRT
APDYbEiQ/mfvOrqjj8uC/FUGO14bosBbvIqX0WfGMGZNBg3CvhWpxego2KPcJC3NXq0DNP2czKFt
RcUzfwwAQjPTVZTSCjGGtSdDAyh/5ijhZHwAHXLOm7/zPDj+lPU4DrnleKp/ZbwMMfH6RU1jCLrb
Gl46h2plelfRpSfAsTIoXMJrTyUar+6xrzWLbNwXIymjLvMZ41gOKIVguB7vEGG02jJO+Oh2Q0aF
Mq0TMTSMUwSyD+T9xJSe3bfr1Vhv5sN5HO9PAVX6mepMtyN6+2nTbBXZ3MDq2gxZQr9nZi5DFgOu
FBNDkM3I8mcjws2A9IZegt2bNhLHTuTVjgypVgenhMAHgXt2sAiJenj253Hp5xBqRXj9ccHITmcm
jAqZspVekAob+zj9rNwlk7iDr7JoQZ1ey8XJfDE4/jDI8OmtYEVqafM888YcTeEwEvs5xFmNYVx9
5LjIpvKzvhc5tGMQKh47xbpWDQQVFpkaDVgjlDLyAxH3DUi8XfSq2ljR86uVcZBe1/hKuwLc+4mK
Jvjzgisihn1YAZTquXIXXn2XM+WJ63Md+obD4XDfUVesGRlmpdQ92dPU/VW16SQqnUMnYSbAczjY
/Z6wifQefldYh8G7h4PI9yojxvYmR4YWSybE2KmWYrIMncw1lyH4oGwFG5upiOvs28EjmhOrm1yy
pZHPWptmCfdalFKV/oMneTt86D5444Vzcpu9iZDQjp5fHErYBL8vu2eYbH2kPXXY1OWnlOW9iTDD
gpXBqF9s9dir76Nee9FHNOEKNGVXOzmAUifFYElhSfe/Mh/s52ulq1PDZMwhiLHJK6kJURM5R/Gu
Sl97ZNpewtzmBg0Vz2LG0FQiQfLKv7rdqGk+cjMJCPZczmHD9ZrXGVOnyixPkWjnX+mMYJ3bMdzp
skJ9oNr/XcMWOaxE7ktihWGnPFojZwIcx2dP5kEcDMSwfxHAyFfmsFqNv5HEz//was9P2C3Hl2Ot
JISG5Av78t25xbntgOEkh36QSbvN+dtxrMrXU698Wjk86GKTmrErEiX9m5J6X98TqMOH9PGVOnUY
ldkyWr5MhTLKtcJNGFBzvqP7M4MFEmflQc4k4hTg8UvCsb2wBdCkED2wEeOdoUTae+NuZI7Dm49k
RqkMPRvG1kkZCIo7oD+34ALJ7ef9OnjKYTQAsGGr8houCav6ETG+ohTL+dwCvY7Upa8RWUTUuJKR
5UPhbavDNrYRDnEe1FfsyG1MKKUop3cy1U17mTOes4Hxsk6igLw/Qg0Hqx0W2OnSp+1/y4yi2Y2p
6FoSLBkKFlEaHhKdL6+rIKtVlk0KTaZ3oz4PCq9U6aIyHy8eS124rZp36dxGU5XLduVV2jNTfPre
uZeMVDB72zesGgyjtiPxy9PkRcFc6U/F82bjH2hdM/PlabxIX4pFComVzc9m59eDrKycmqbg2NVY
qFjt9onh78+ytI6K3ExpQt3HHG6xENPf1h3Itk+TJEYifmFOHFgcfx8UNmTg2OkDwrxtWh1r9rwM
qLPdxyMbFgvtMW75vIxmo32njO8ZCirj/ZKLVssGhWdXU6ISamniwo4zo7f9Doqp6hXouB46aGRH
MaP0dHmVFsFLiXnPV/dRLqoiLg4LwhYlAZdwiwTaod4K48OEB4OvhX95kJXko24Mrk+hAVeZ9vdX
bhS0Fk2BOkiO1AIXILtDFIZpUXGY7VK/MTeMFqG3rOyaez8htfkjYJUohDVVa5LssPGWPWuACZ4J
G0I8ouaYnJQRsCjXhfzhLdnLBywkvejFXczfYxqxWbglnHxXuZepsLooVM6fSl22eeRlVAQKqCGa
c0QoSDSmTq9dtGOlKjzKSCAn8t+slm6WcLFML7oRnJjTunEtz1PqOaUPvp/t5cNTZqE+n+1V6T3/
+m2nbeW3GV8UmglM8OLVIvVZS3BJa+9bn8qcBn08um3/9w07LANt4XTG7CWBhokqtI3B0PrAcFNe
0jV3IVihbfXphaofdFWVCRGfm6pg1HfF2SczHhVCzwKRh5nCu9/d+ZDcyVyELXNU6TbxVMtpqTWT
X6cSwYd1Rm3Qx0Nu6i1WgUCmbtBdm9gJeiHIG4VVmWBweAcUYsWFF40O3eDKPTsgMucuC+tvUUjr
955ckzapJU+x4XP5IS0lYOw5QOr5LtTWhW6rr8+IRz+5uB935h2tfcPj5TxIfEQUH+e28JOn7g/M
0UvWay0QrsDj1l+H8FZfNfPVpUS3jU2+PYpqQoSrbwe9D+ybsBFraZd9S6DTI4XXlYWUWYdv5MYn
yzC/lgy/doCwzNLTnex9gOk+2ul2L7bbPtSQUxbMsDghZWn24/lKITgn/3GSlhdGiid2MIIGk160
ZDnE/k7cXXsNSXclrKu6eZ3/0Qqswnp5Dl+JdrcKAhlX70iXUptvP5F0ham6bsZVMtWsimhomQ73
jixdWi6LsL8T5JCf9c26+r8vXRfnlUWFdw9qHVq/1WJNHkOB8rHOrOotpn72JjFdkqy8TO6+MQN0
L4/UpyOvUOkRX49iMB46VMaJQXoXR4AaqgGt28BunOzIHrUwLqn3qAKDJkl1Zm9VjaqxmAxPJLqe
MudrKbkG+iCAGaBwHZqGIeMMgbTHSe02QxFp7mFjUrxKBgG3bSV6NSDPMMNOkjriVrej4bYc9lsC
9jD1/wTFccSR+9tBEcADwSXorn53+i9l8VD2mbg0j151VrZ0oKekZ/NQoNI+8w41zyqZgBBtjz6p
UTq8cIMfKV5RJn+XA6IAhx/yom7rqw0Cvh7kjoXAvoii9u0MYPSjSkMy1a1aSDuMOjC2uQzbVP+M
L3RJKcrw1NP+EOa5/sATmWIs0CBZv+nNgvkeHM+icmcgpFA9gmWitKb7d6U7iy+qZ9smAwBJgXES
wRX2OFKFbZeZ+Kpjp0riaX1xWSmaTlHlk2b1el7KKbV/tFHSrk8DJkfN4xPLQ4VVd/UnsopKWptd
MdYIKTf0ee8ZIc3HwnTfK0sdrjDWsScAcbzz0KAPw/RgnBkI4kQZiVmdr6/O456gbs4zhB2G15o4
PGu38VWAoFCk+zThndPtTx0n3b0jqHllD8C74rGrw6cIvMd5HAbMZwdGAT2CJaRddaLVnwAiCAo2
0BC1eOyyjGlRa5YsSUPALPUA7ba6DOqT5MY7qtoB2JnBKuslLAtatm1GcZSkXgF7mNNzNdNTRWaG
ZtB9fjw79QDzDg631ufY1JEPNsEtqtxbosKRjYG8oSXBHseevA7UXLTphyszjbOlSkJEhAA7Uq1r
oE6V4hriQHdw9AU9mtJ4qgMkF/IIgVC1cBzwNjxGYVxU5akVRI+yBys0KvUzooL8TOaFDbdicjaR
ETj8Z1l8rEttkcOkkhpXR5K3DFTz3DhP3XLlUXWOxZCCUVgVjDbUoIKqLmCs7yLcJ9fUaSDfmLbI
EjJCVCzA/oeeVnucFd5IFPvaAQP6rd5R7IC2WQDeK9S/lMoiKfWzt5VC4Z5hGrPOmGkq8Sdv7iqG
hXowKnwRQoTottct52NP5a2Gpv4PaGb/NWJxIed0i7tSimUyG+8wd3JFHs81W3lqFSHbxT6Oofun
B8ni1a/IE+F6vvw1WDpBjHbNiUZx44yNPc2t3EIbRVtBeJK+YVeBPxSUch5AvUzXqJQbRtDsMyy5
tRsW+A4v62vY9QTr3v1euGF4ibtGAzZ8PMTdUKD7psvo4bTiymk77srLJLVfIo2XL2phXkf9joP1
Y9mD+iQ3uS/M2MAYHiFyTTrxwIePXKshDEjVrCajyBeBn5R7M/NcsiNBhJhgbO6cbNtIdzHfFiO0
VDX6N8v6OCn438gtOqovYr+M9UeD8ii2vB2kTTY/HE3FhpImAgC/ZkwX1ARvijxO2snNvkjdXD2W
6Oh4Q2e1Us/0G+I7H9r3vREXM4n52sP8CEqrW+5PHPkC3NNRAr1pKUmkyBG3AG0jIyzRoFx1yPIX
Fcdan3eJJkxBKApzuF76bWki05wILGNF7/K8DQBVFz+94QQ0+2FsllCqjk3HE8+E1gsz7L9eEEh+
nemXLjSWaBGxdvhVFxsO2ndAeQIXbTujjCszlJD9e/8dYD9UIW5B9qAS5iHMC8ZDHt4fRGwfcgpM
msVFZ/iwJECvdayGLa8pHQ2EXmFLjaWao3NGBXAssaaKT++Cgg6qcFOY4h4KPEE6+f07thKyB2q/
Woj0jtpw4qwrPMfJRzDD38ukJyWMkRUOsJV7SnJY8FGrbK09ImwBWtPMrsiezH4A16rXk2kOCc/M
0JqrAXai4nu3+kUz9o7hO6PkdBTK3SgHRohL2+xzZ7ZN7w2VwB4SKpOM0SGYNShV7JDlDDZd8Z8j
oHFgyXz5D1OBBiggLPQzJtyPak5zLhxWsuTxL3X6hpopGSceuuKh29syNvb6Gyg2BXTqKpe9CIxX
oYegJD0KCRp6RIaph6Zy7Ef2tBdsX+HBTjZvDwA+o2FKmMIVLhn++YANCDypmf1SCkCJfx1rYLdu
IcVhBxo52xwMI0gXzDPmU11VQdppEjohjSyPOgijmi2DT7PoXVKDFNG9hUNEvSnIFBOxCK56ZdUJ
4Zu6bW/fuY31xyqP7bSm8jK/jCo6RW4+VBfVAeD+/ascBRC68cOaQmjAN44rzHwNMgqvGMC5UMDS
Y1yGibCeyAzh704l5BGOoX2NJZLdz1xZkuI9OeW9QvrdCQ/humdhZ1t5y/jlArEEmPMElkC1mtGd
IE1GXihI8upFvteGpSaAqlC1wjoNtFQocWm1yuyJSYjKm6ESZdFiADSkC0/KaKZJ3gOjOnHQHszq
nqTT/jqXBi+DUo/FhmN7lgtYLRuTXPtjpcNwnCSCps70a+rmRSCDwvQfnMGHJbeCaYYYymH7vEvO
gZ/d0hLxzwR160CtmlEjdtBOC2h8TsUlk4mwABJgFzvOJSEDd2WQ8Ke2+FoTWQtwfRtQ51frULdp
dixL5HwnedOiALeZwBY+rxmQ4GbOQVl3oVNVOsr9xNo0zk6+ineP/3WxS7PBeF3xKwzjahiffIB7
z/eIDyk90rtoXK9L3dysTa2GPI5c43qdjPgfR3cE9P71GSpMKkYBANcjOJCb8w7RgPhl6vgdLrdj
h+6iiFoPNB9FVQBywB+gcPgd4WUVWjttKM7HrxzXHO1q8PbWFBB0ZN3wm17ejTUPEKcYAVl+E5yA
Gy++bZYpdWKrW8gy0g51GgvXXZ4fVMW+omufkAJKiYWACL3CGsj9/1CDjG9r0ROKeBlU8cdlnhfq
SdfQmAhxVf/LYK0zFqofwaKGlY7K7RdMZhQ2RLP3IfBCziLSrtt1f05wBM7z8nfxexx0EzaIqfU8
fzaHn+OKzvYwYflwaGqV0e06vYjNH3J8WABS98tKm+7mVzDxwa3OspLo1/uZLYhaqgBocQT2kLbh
fvdrb1kRxssY4F88DlgB5XpI/g6MDRjfgSu3aZNp9YZGXxIHSe77FErn0+8JENe71Iv6xj17np66
iaj476cAKfz75wWyXS1oGgGqlt0zVk2jzw55OuxYG7LT+ga9XblOXSUURJ+IaPH6kIpLPrJkw9tP
XcWVDL/WivPvdCZkFdUKdZBm0piWYVUCuf6nzG1i/NI9HuQtE46XTIetsRRSEOqvkitfmNMSKtlI
Y3yIpu3PD+P5DxgRZIyo+fuq4KNYyFZWMkQucmZ7V7w+xACSTgKD0EutI5sGkk2g0OBK2U/Rygqp
nCNAq+0XXje/Qwbfddo+D8ibZ9yoRiJ2jM/7X1+w0Alfz9Nwf0vxrzWSDo/pI6Wu+5CHz+FPuqWV
JymV0zWbQzdO38HjgQdNLDlGR1PE4XakQeCh5/JD6eg9Y2pdPpre+oeN/b+Jb6rXQ+hpBXoWdN+6
Fo/lOKVHT7aWJZq2BEsTZcSpmsZT7JADO5X/BG4IDs55/vRkIfSysVrc4fdAhWIGy4tu3kxtAM+N
ftY/CN/tcDI0ixlZZVcUtRitBr8sZqQGB/u6O2lqQQsk+zEJ+Ee1FqmCo94tptpEdjRq7S42/gHz
xfShtB7ojyNv2CbbllUTInvS8cV4IqCE+SqsUZ05uxji6MSgloQ2KuKFa9j2XpmCrsiDalEHzghk
aGXimImv9g7FaYWYfP8EBEbi0XIdbzFBmgc6mx996xy+9TjBwZTvLpS+htfRdS+G4XRvTaE3s8hJ
3hJJuePNqG4RyYNMjVwWq2eVyglxoVp0LQgEsJxEzytCpYqG3aZ/qgkAUg0qTnNeb77wGdtEp7ST
PrityY56kj8keERVF2AM4SwxYRee+tOJOCZfaardXqKfGAcUBsCVouNpsT9qrAL44BvK8zFrRzYU
2iwLS8aq01HRu30NQjULXo1o70NMBjjaYjhqCiFM27LM61+TOhX9pkjBt/B6sV6/O89fk0cnTdFs
GNl03Ci7lsyjAKH/pChb49IwqyRZAc9iUimjkdZ7tZzgc7psbE4xKSxRySxKikFHhYbXcFk+AH4/
y3FQxjYXhoVlv8ho3EZ5ngeJpZKHgJX1IJbtlC6guxUxAEMiAIPs3cKC2IIlOZF6oq4IE4ArqDdX
6eBxZiOJFpO97bvq8iSoYE2JoWzbB40umqDGxP8O1kwpw6QbkSmMWiKa+98YMmAIogdyVGRI+v+L
khG5JqoYUK92vG6rnaMa/v4oBsqPuuSYTzQTDZWuh2blvRyUNKWiTTalCwg4i2rpoll9UZVK92DW
De+ubyrHKtET/jIyMThENuAfNb7/QNU/mPvs5IEhYSibDfs0VOJZufZxl45ruMgtSbIyNSQ08u1n
bAT6X2jl5AsnNGl+xjfXY7D/lXM4XvoJrArcszH5eWiiApkFxhq4Xj64PJ7n+0OLOgOHASF3j6M6
oSZk/Nk2ZKwtB+9bMzVN0qNfT8T9KqNUTASahZPG7o0HOwQld9u93HVOO9k0RZ4ZvN6Ddy2thY4K
z3MxMG9miff8XJB+f6U/rPisQ7pIC08650F7uZyFOc3hwzmTKnJsU1Xx94h+zgVkrhY7imwuw1hW
WMAlgmqLYNOWZ6WFwMbsZAzUfd+rXTzZY5786fLBO8y9DldrUegcp9C5zPMgGuFCmUfL5XUJl4OX
xBlYlYkDxtLfmQsX+iRtnVjTamKG13D4eamQkCR26zxAhTNP/01HmU6mlQpBri2OWBde+oQPvyJn
Zl7zK7yIwDA/Ol5MrkM+AZNrrxSR/LE0Zw+eTeN2CjaNEOuvjmt4B84PtpzEzrRuIIXBWx09lfqM
ARDrp/tJ86y2pZGY+pMXDpod+id0fyKMV5K/iIbXew1Kjh+RRZS+v1HE29XPCC5oDqd08b/JC6p6
Gr8CkAK1jVGBD/Vt9MPW7Cu2u1OyA0m0dSn4bae2iTx/rMWoQU/RUkdWMreTjnNmMPTdkZQmDMOB
MTM7xyH6mSZExZa4F5eoLwYPvABbhboaKftWu1xiCw7sxeofX/0zpF8lHawrnAfYRYjtzXZO7A+x
b8Y3cJGCau3YdDhEFFj2KtFZOlq4vNoW62Ou1XTJ3zL0NKqTSf1x0ifxZklgZKEK8qehhTz20mDJ
R4WRi+IVdCCwIFbVRCsYMM95so4QssddkYQkIHd7BQKaHQTgMT5kn1VFw2RlaSn8fBOcIDK5Kdea
N2s4pTYS6r0rwBPr25wApuLXyjryVnWnf2BIHEf9HeNUlgFELezbyyKhEoY3oMbzdQSqOIZbrBzk
A6KsjwBUfMNVDm8oiPR0ddbUyW2K82iLGDPVbeL42h1tVbKOEAx45qejav5vv86jakC+XFa/0zc5
Asnj0ENgJzsobIWooOdhKJePVPT0bpcrSu+H8MHidChHZRJUygoo/kwsInIPYPgMpm50412RiYov
es6eEXmPQaAaj4q1VL2OiMZPOp3GFtEIYOs+rRf/6Fqeer7PTeSqhm0ZLM+RrbFPDqqYEjKxws1x
Q6qgE2z2GC6+EETjUANZsTo6X0Wy/LGSOtInpX1LCPrD+3VaLReUm+Sue9IZJatawvdl2k0fM5Ui
ABUNEqlaVMrbolCdtbrSdslyL3TagXnmNWD6WlI2HSmtENQQDMuMDZ5SyBqh0P4v9+XgI6a1IPIk
8cEadjEMJyYjzDzms7hkkRxBJew3a3hxiMsfBVBY97VMAa/L7EkQ5ZaMOVOhpnbaYg7YzikavwXt
fO6VOV4lZV51wnrizZ2ZNcdI+qbga4AHlbE8wbCUV7yAAXbzMzWCQ9p6WDHEVRfJT4TWBUbMaeDn
lrt70NGuLsBl+uWJD4kiA08aSh5zXrsvAZp6uZa4H9PSb/LkvDSHt+ptkRSCvi88p57ClM5G/Zyb
eGhWLG9g5FsTA3vDCven5YBvXaQaEI9ESmD2Twe1/MM2YBDRpxRJbQe6hJG8N3zR9ztDdLJ0R+6m
AfOE9JBHU/Qk2ioT6lUkM//Nh186OBSx+deTWAfT8JA9/JW5dA9H69MOPmGaoPEekgtX2FrP4rsi
1NeNgT/Os3maQwGc7+vWOYoEsj8NB5N8PaS6Xhn2AbjFQgk7M+oKlJ3EX/QZNaO4NOZN9/m3mhJ0
KK74wDsk6IaUatAj739uPnEHzCtkTC/GLxpBZMGUMpXNQAjK9s2w2IA7VBNi96umwGrdC1wyIRZE
F73gReu0kdtgYjCD+KpLwIK44oBOxkN0/2i/QhgVWe9r/ctkyoCkn6Vt9befjAFRBt0USamn0b/9
Cq5qMinlA02jt2lQRMbXT8OBErsJkZeu64AFPjc+ZOc8bsVUljkyhprfd6DOwIyWDpmfHdc9NmQU
qrw/Pi9cw6D8HEYxVChmOqLCY67hxvT4le/OlY0R94dq7k1m2WnkHRsFFf+bPA8Z5o4e5zM81Lpo
7p5Gbm9I2fr5pA0moloCCiM9/q/4K6/44u2arXcc6OpJfCNyEckmbhB7znE4fbwfOpwA/MrJZFCM
7m5jddbVM6EdG5ZImVDN9T+jGXQZpgPge6ebGfxKCOuNFwSiqGz03J5gIPGDam904qPlmDvamWo/
lCrPrTKFb59YCRYfm67j/RIDDK2hmqlsprVTocUSsliw/6/bOSe4qC+I94O59380gaqjQopDjN7R
aEWtXM/0AMiFc/n8QjZ2MRfZ2WMeBcabQUnkDUteEXzfbP+p2y+cXGF/DNJA7xvMYP7zqI0sRDEY
wYEKrdjeT88Yz+yizWLSdA/c/xh6oOq6g2jchnH7skgoTRTJKdnaLhyK1Y9RDDgiAzjVDWFV8rD7
Y09a+h2sFmME1I9eNw5ZclHzL1wsJqZ9n9a7weRdcGzb3yKMC4HGnblrnwtPQKq+OG7cjuKisXnf
siS3UhnwU0vX5+fwLVe8rjxqFv1mWdiiA5OG8Ce6L87QmE+IZYrsdYLAVcAQtyGkPlG9WGBaSPwE
lZHZrS7dlNuBWaIRBGmHuvu06SEHMB4Y5EM3Ws4zG6Bs7i4ifZC4XbY1/JuyWZs+dKv3kin/vgCV
rzex294gTiuDK+FrVGiSQdZALajQGS4vNXL+ecaPtSS5oO4RbL378991206UMfj95MRLwULjPTkA
oKotxVJymAM1kfozPLGWWFPmQvwfSUQxwZFqjVWKOvaLfQj5fHhMk2o3YIhz9GgwaQ4yK/9KXeIQ
kH2GJowLbtzQsZi2KdSJFA5TXd/mRFpYFyKf2rR6CndMorzASj/Z6Kw3H8pC/e55Q3vyseeMagbc
fLIWkeuIXXkRrmO7FRF6+D26O1A1GeWr4wFYwrHQaKF6VJrXmbr0egHpokjWSZgVp2+U2c+PNoDA
kM/ekj/VkO9fcTQJmNALjmsr7u5VW3oYDs2QaLsWZR0StvJp1BuIyOgzdOUNgJ7RF/M97wxdP6gK
RpXSK6OjIn/szY9/vxbdJdoT8ZShh+3A/aEJyBTCR/5cTxE8Tw3zoCHCEVqMbcdOICAcj6ZUTJKz
9ksHfE7LVOShYRyAFMQrLGmPmzEd0eedaF6q4t6CwN0fmFd2gYy+9V5zAXzDUOkpc/ujqZzsfks8
OZN9D/wDRUVWtKGyB5oI9mlQaPVh9h9cglvY73wc26JsRKruirwmfB0FYbmOgti4O1iTWO+7LpEF
l+jDARnJYdkouPRz5zMI4Ta9yIKEy1rjQPB+cpVkGjlrMaVLWPYLWd5+OsFj0hZFU2+OkSSynxnY
3pY3s3CAri5psOzhegkUsUoD5atA2fKUNuTgzyWWJWF/HWG1Xc8H+KNChGYJMYGq2SdmJ6gegKtL
ejlRgE2GPiJPYrvNHZCPeKmoy4dKCIWkrljIHDknGJIPLggucFwqeTFedKPq6EK/6UEL3oNAJzZm
1LUn9zhzza6UuP5HEBZT9a1liGxoH1G6rlCmW7rrmOyG68gjh91IspT4/VSN5LPamgpHfSKV7XwR
wpoojpMyLlbjzAAzhl/LD5DzTdxHKopM68d8gpCxEde5NfRYMF/oX/qXNODcsMNxvW6Qk2oZLwED
hrKN+pkhyuKS5XO1zZ7McDSsLic28vXeesC9x+3lkEZhZr3l5Hr4z/0jvVarHtAf7cQV4rNt7PxH
6cfIRlzxbQAesJ9/7UcOPo2yG2zSmyCmgCASZgQJpeRqFEYhR0IMBzZT+TNbLUmyyiYYOXdzgZ+S
uTwRH5M/poZmpPsD+BmJghmyb3p1e9avxXIdFHUqm8Q1kBKGZNfvHezqTcMnXqTOnY1O4Dxx8Kra
MuXQs7wZPNDq4L9G02vVtG/mCLr5r7tUeW756LM9CKuVY7KPJselDNvGvTjqvSVuyr2+KSlzXyfI
j1H2r+wyz3N3dXSd+VWOV/cbBh0NqL7rtVaoE7qJwbuGHeFjRoTik3GwyOXK97NTmYiwOYbQLksc
dA9Ioum9h3vyTj3xzO2BHl2qGVCRc4I8mQNPQ8O/c5d1svz0vUOBFc9rCnlPbkzbjK/bG3hcnUfC
ez548h7ztRp/CP2PlTU+oDxvSMauG02A3UqKPdBCECEtcA2xoqjksMXo523kXGMYdZfJEX5AnGV0
4+OIPpSk07ZJ26qSrsA3y6yL4x66/F8nhV2/lPzXg37WaJ5Xd2qfd1QknAWwnyvxilG65VIQJS16
vDw4u1Nvh4T/qATs2j3pjK0GfKaO9Pvsa014RJ+3ySNstht3762Vp8Kp6XPpsPHWnmhxtE6qwv8T
h8bcSVKOgwB8g7MRLpKLRTnG7TwSMn/A26Nt3JKU3EvoxncBBdqbd3jRRgBxOXgWlmbtw8r0Gayv
HuQvJxSTSN8Au7A5gdl1CxXeT0YWUR5VftF9efyR30dNnXymCAyIhevo44DSAhAoL3iIeAGuS6gn
Xuv/KaExQG5ZI8KAGMUTJbXsG7R6g17wy83di1q2BtqFN4vZL73rOn7zTtlntgIhenBMbaRySpp0
jDH0x+6BGBIVOrCONqOohqKYNUXEry5R1KAD6Dp0JIfls8uSIwJYvd/cn1St4MGWK+HZeimuesEn
5rudCNTwWcJsuQBb+1V2O9oYdMJ4KWxm2A735RZB91NRmSYRkMEjFPEe2U6WtpeCy5de+/OIwKrt
xT04Za1M3bW96aQ1eEKOw1o+facglL/2MKk7YYKAYNru6DSXuzmv4UZ4041ENxlEpwg6EMnLGPg2
hytOIdtDKUgQT1OfGA/nx94LEHTpEKbhl1RaToDOwSbRLlLNAaPKlp6cigDDAmjBm/Bn6PkBCQzH
uuuPuxAr1+9dsO7U0KmKEhW21UhRwFtjSSVLeWBiM52isVq3ACzKPdqT7deik+6/ZwGb0gDhv8Q6
mNKafsMVT5Cvo2ShJ0saju7sBtMU67EIP7PbpJwxLBJy3108KTD/WtBXMpaVuMOwArZsgcZ8RZKw
06ihCnoVuM6DFYbCrNYrpcTsx54wMKDAFdXXIs0SYlWHS0KluFhj1kk8nVlAG2jKCiGRV15fw9Ou
MonKQAFxJn/7OXO8Sjw/V2UPUi+HE4NcQitGnZMQNiVF9y675T8lENxsDDd/oRD+mMrRNWihKVr4
2564mrkKxuF9HJEvOZ2bwNYcuoW+ey4jPRzJ2wRypT5Jd6gXZCZb/GDhKAicySU09VqmXgZBfAsR
wwH3g1FKffbsW0VPUIH4pRB6cWcndHvF+JwrwhDzM3u0wUxyN7aehvarAd9kd8eAqnTcuc+r/E1g
oxMdJlXlDtRiJkLdPTw+w6zCjBmuE70wCorl+GnOgcTLXZl4NmFXGw50lrV5Z+6pelHCc2r2tXGp
aevwYXz6aWpU9OU6o2uZ0GRjqxhs+nrT36e6cMyLORkW9izLiPis+w760zQUlk6p77HPkusVLkSf
dKL/ZbGkJTjL55VMuueFqK2UHmuGrxj/m3fF4biYzDnIkYbNth/FZpSWAsnAvEYkBpU+gMzU1D/8
3MqBTY9Kkah9DM4NYQe7Ih7XOSdFkb84bwhwNNQKQ0LmUyRLQMwrc1EbRz8ba7eE+/fwjCuUJx1o
seAAd3kdm0EMTWaBjTDGn6s211Ww3u/XZwKYr9rUP6ywh3jafUvMha+GXl94W264y6TtL4XHZTVG
4za4x62jhEuo4oaS+thj5CoxXdkyisdmJNEMRZW938VnTc7YDRMod2EwVYl+yf6B+TLeFuYCRll8
cplIMS/I1rZ1axBoqttPnc7JzajxnarmWzi9sf4/pSiNvNxCCzGslgJbZXoRXiI3IkszNDB6lvY9
Zw3vvKpkNEZsqrNgXZvVdBpx9+xx1v1rcG4FzWRckU/ux03Vb37bwbR3BCd5p7vt1gRfo0OQDDtD
vS7jw35iZTR1VkwPmo2MqsGinTomeaMkp9rNSdnMy2rIZaO+QP5Am3rYbJXMYioR2dXYbHJriGEg
+d+oS6SFyeTLZE6i1emkap2TNvxvLe6OYxUmVp+Slx+2hR+W6BdtH23ph1UEMjWg6C7F1TOHfpAp
Gj9sjNWH5DLoisYLJPiKieANQWlHQpEOcPYHjrd/SpRyvbGPKHtFfnnhXbjtFwzuDWX5Kif+KqEt
2uVheiT7dSyF/GfTjwoNuUwcRrsZLR1Mnz42FLAWycZQwzi24ce9xG+8LPUzTdZp2ZNbE+M1+Spc
20r12p/RFbNZabmXcuyvjsFRakn+h93x+i4gp+yxszqrT4U48s9PI3/ZuuR0kHO7sO9g5kLlgXjr
PEkcaKlcIMPIgBEV0PDHefP0eMsfD6RXKDAQoc02huhCzdp00SaTcHgCEa2Nr/1NettojTvB8vc0
yZooTTQA6ME9bsas6ee1c9HpSr/lC6eiB3aHG7O5XHs/kppGrmG5+FKLpzVDpp0On7gboJZTscBW
WRgZsfZbF2HbuLhQzUjO4OpMOrscRSa+tmtUXORfW9nFW7YxdxyxL/7cz036T2Fk8MAOWHlBYAWk
kcMY/acdIpp29bEKgTRZRfs7tOHwS1/ZMdA2TFMFbW4l8gH9a8Kez/OuwJYm95uUwtI1muFl9z/4
lxmIQf+YfCF+lwTh2wUz+KIVrOC5w3NfztpOR3Odeh31+KJGGhMN/MS1eKPtH5DlnwELWYnxt4rO
iv2B5ecxQpPPBspr5MPaWXVoApCEQ0T5Oro5fbbdC7uMukkr6nunOfRTl/0F1TBgP5BUNWKC+Vkf
o+wP2SmIvPqev6CO/2dI8m7KgdAkvxFOt8BkDFBTaUm/peN8qbRBzlIt/qEKyjUlqjGX5WzFx94L
ExWFBsR6J7RpZ6Xwaa1S9SWPUjUJu45OdTihiecc4A7ARv1LqYp7s/BTwYEJY534Ey7oU5SkAadt
y3z6NZe72DJFjav9NW9welryzhuqWtmA+VTzZXsLnxg/kC/WGBmfKS0RrcokbAZN7R8n2VQnj2GD
Ghmov+El8oN24K7bfhj1C117pxLsajn1lPQdZfI1etw8sAInFhBRdMx9PNiIwwKuP4lrr26l45nY
zdmop22qVkc9HcOiIj72jQWGF7s3cIOkjThgeP3Iwyw9e0H160RrNo6Bc8dMgqvcLvuQhCDV4M3Y
zQEt1UWc5AQ/OkwoKorowH/DO53A/Ql+sTLJMYbIKt4pfQvwqxNKAVRE2JVxZQJaG5hnNXQE0IDy
2di6uXLS9FvP3rGwVysWLsMMYxRHDVhKTkGJrC+O6U8WKhdzzVdwV0HTwMkPMJuQzXl5FXzGyz3a
Ofsmja3Ar4LnMV2vkECTmNHU3W7P8B16AHZruRD544Berf+Qu965/W68BDuWihnyA075Lm64Yqnl
t/QiFPjdnqTy5e6UIzB8VmMOr8WpJveBItQICf6wWyGuMj3x+zd6SJlr6StwrxzB0wxVYzllbt+S
osDYQK+/28F4IkERFbx6nv8SQtttNkX+AKlTmPv5JBlqv4W1CyFsXXylEPXaAptqOv/NCuaEMwEj
vMFN1fWa9m6pK+Lh22XlkqXewa2JPLqx9LREta0l7EyAs96ZtREkfdW6EabAHxT8tPyRF0cZ4e6G
AYGfJi9wi71C4a9wR6qO1a/NioR3i3MOmPGjjNR4Ou2R/Pc8c4DoJSumVQ6pUOEX1+ph/IwgVP2i
ydH1eyZ17HtEfO8NeHK4tGMBai+zF+N69sSqmw4BKdoTnDkzuVGc2znUet5yXQ+ydktXAH7TILRc
+p8xU2HGfpWDUCJVPQeljLwH87aEFr2bTeajoYjn7NbSVv24lz+31E1ERAqMLWvNuWF2iXW/myr5
LhhHWkR6u4XzX33tlMqZbrI0YvtrRYOQpCTJdZUtxoeWRTFfWv5rSel0TmzHPPWVomza1wb9YUdX
xVyqqB3XS/KMoOO+Dtkqv/fq1TdK2+jK/6yof0D6QO8ScLI85SZGpMORQL1OVA7I3UpqBZHM9WBR
TNntBTKpzaa+6TfhDI3BnzP9gG3lf0eL020x4fSPOWe5eWE6/Kve/SqbKWvI6bae23kKskzsjpHF
1/pmsGJAKhQENLawiahiPY+CXpMUA3x0SuTBYQy+LTaNvNYkRfJdhJeP0/4I1D7+AZU28HCjMJ5C
ty/svk9dn3sDD0ayN0LkWTNiuGuwzJ7y43LFwDq3F1FmbL43N/eNMq7wbkXqOYsG43AiItQtT/ws
8q4VY3ampw7HgjbFYybNK3To/bUzhuTJ5GOL51iOby92XGGSamrbWC1yrY1G4B04Fp/ZGLqp4/dx
OUW36q6309Q/sZAK1U5gFOh9ncyBcPW9xGBlVXgLx9kbizWkbN7/YajAR3873b2sBouDudMZJs9J
gk4JN3omYuos0KNvArfPddF6B0dUGci5IL4b9kKx0B6Z7wXAisM2izpfKbwbkqq2r+3tu/VAiuJS
2VRb5e13WK7kkB8SLgaOY/LkghR/xnPH8cgNe/BmDLYJZtoc33O65SehzHEjO7xOhsvh3W0fZw69
ID5LqTV25DI/OsRFBEPM8JuY0YeHOlmZ6ottQgRLp/6M5x+MsvPZeiFSur7jOWBXu10/nBj5BuOB
XBxXTEgYvvyjsg6qd2zwBQWSpoShk8/PzenWCWd7OMoHFn/rEFg7gnkGcqfxa0+2ZNNExTEqff5w
gjd6G6LekyeiW6+0/+TcJcCX0kS94sjd21PEamHIWBmXELg6WzWML2D2JUwfg5nWaNZsasCRJed8
aooyLhteWMbDhWvD1JbsGyhy0uoMdDvKLWdIhgcJG9O0HTpLZmUqhk8J/qZcHn5bicacwnCRKgSn
X7iJ8phtUgk2+h/n3ZXghfhU05HPfYcQxULfU7gbvipazVmKMmqk7JjBnXa22ohl13FcS/JQAyA1
+PHiRxHmDnwKh+ttnfPbcN1NyifJiedm/bKVI+GGmZsMDgvM5/qk0KotL26W3ie0UD2hJa2y4BOE
k2YgNOJ/477uFRUb5GxrM2KcDI+M3Oau+kXOZUd9Img8z2XbVyuoHVnHVYIDm/QktktZYMW3Dc3A
e8/VTt0OSzcGE6KjC5hrDNoDxOBRX5O92DeMAM8E+YpaTCC/o9TuQzxzMP2uIzwXX48U/3tNFQtM
qE07H3n/OiEjB17utvb0d45MyOj3MvXl9nCpAISQgd3fjf0D+xP7DhhKzJ1o1XyyJPeuqb4m+iEu
PulR9Xx6UgUDcYxZ+1MF3oHiYylBvG5GCwwVqr6o7bAchUa1WN6gEb7zyX322th+T8U1rsW95Qwj
JcV7yYjSO0e7SU4r1ZMzsl5+9iTRh+kDw553Lg7XBuW5VBQKzkWmBlGTX2OGbA/mCXsbVCF0gU3Z
uV4xNdapfuIluHfJ7shbSnulFk63uQBjClwGj/8xfc0wQKBLIKKDH9GEDzAgEZFfwLcSpEjegghS
dMP8nRVtOI3b0gnp5s+Q1oI0Psa0Gc5TMzPkeilZa748mFHz4qSIkl+/DgOGWZZ2EHBLcOMn3EMU
yZlLNfS7tESiF3+r55CjAdOgkIHvnKKgss5CFGEYuup2D+XzUDLT7neXkBJkUouPGefJhw6KjXMg
fGhcKLN9WZIOZQJyB1z5QOkXyVxeWjR8uHbFDGwasLFYOnFM1OzyV96JFkvqGWvaFfeGj60u5diS
utvTWqGNvirchEv3zrfaGdVS9OKzEzTiaO65rWw/fzn5YrCG7O31EQy+IWgv2JXSTdZ1NOZXocG+
9QvzM6FiiFZoBlIbKqWjsWl3wo0rWuldcAL51V/UXR8nE8Oxy5UI40mpmDuBWGYd3aBSfg/VbKCg
6+xFurnxvh990ERcRnKEhA+w2vrz2xEQ7WVUaZCasIiwt4j0a7KXHbYlaXW6QvdluwhZEdWCGRT2
lxA4/qTpJQuGiapBYC1DfqVbdN+gkJ9XjfAzIakrSLtay09UmANW1TNCHhEuM6sFEWlbB7DiJg68
tjhkd61iERqzeejovmm6fw8Ry5ip5pLDxTDq5jlaEWkwaZrTq9vEUthyOgAHqCR3GsyuUzJAdw/5
CFJuGIChf0S8jCA6qxIlyze0bs7SFUUVkFNMJ2AbOpv6mpbdfairS4UEFqmYrawI8289iARthlCE
uUBZ6kuVFEc8tjetOyjEbNPtSCggP/Z4zUPxuagiLP+9T8ihl94tWMpVsiJJahGWv0CWZdQ/uDrr
OARuhrX5OnES1QiP9asrARBgIys+BmrIX0Z8sq208BS8u357Utyd5bQaM6Bf5Uj3cVDsmZQTjdDl
9CPbeuWhARliWbHsNK0HXMClEb5sMVSoqRDmVq+XRv3h342/rBh63Mb07IroiXD4LwWsMMRX4y8y
y5/hDMjhsq9oY5rBKahf70uLHnvVW+EGOkI6/fKAUm+94de2DqjJM7uwBaGuu64ZgDTWnsv3Mt9R
NnDusaKlqVgKv8DekIha/oFIZxuWrefKn7nfQAqmjqAhvLT8bObbLAPsc2ys9QF8Oyu8jc9Ccm9f
qbDGT2AJiFamghzZ1BF3/2ErbMhuctsljrvgppJRZ+mf6A0kxVN7AgwvHWzeTEigDaDf/gLqp3uy
m7uGeVBrL6ro2GsG9jlkvW6GyqYWy9p+nkeZGklm4cPpDGHaGncHFONiuB68BP/I5Q0ZzrvHx1as
onJrOmKJaVsqfG1+1k8UJ3H+/gg6AikuI3cluXsoUMdfgaublwoxSgB4VByBr+Zk1Ya4suQ4U8qe
7IR6p0HrjpmFhvDZMkvVTiJvoHOKYgBtSNT68K8GR6vGELLsYDBcPk+jM7DqIFNyqnmyCUJ76TtO
NqiuErF/pzVRv17PT2pq2RYovzrRKmFoRyPvUVaRln2gK6GGr6H6qQxFHnjAAL9jMAkqXHfhplXo
1UEWXrqxbGIw9HxPr/v8whyMIhcaFrrVPSymlAb6IErzZt9ZPY1K1w2Y+aK8VkAQ+IXF6uthZwlv
qhQG/nEMulYLCDLLa3PMBOnvXWZ1axbXmAYtq5vEXF1t2QyVYe6FcSgeMy2TRiCoHDjC4mqgE0ot
RN4+idL6w3+70ye4GfghPWZv9aVJeu9Dsi65XR4ALKkcbpxBAUve0F/b4pRKfORKWxoulQgppGWI
9QNYiBwTWww2oA5GBR1/ABbjReWlSWvorQWhJrnDlz0V1HMDeyKadNRupwlsNN3MbYQwNEQSTjJa
8r+PX4MhLgULc84xwwhQFr6n5uTCK8w4df7mEx1gljWq+1jG+X1oHEX4s8QtQOgfPH4xyIlj1c3k
5LHzPcHsouW1sRBxTUBGwwrl0DjrNMzzmmDiSLvTk8uVc1y2Dy+rLgWm7pFIw5vYUC1v1ds7U5cP
ISDVAkE3/U/i2mw0U+RXtMx9Z0A0nZD8BmmIR42bB4WFHpIV3O2nlPY/4u1/WLdGbgWgfrgve1Wp
oLIO7JuXGq0Z1YbSiCjy9nm3rFAtCwYn/G3H/6cY2P7xVgs8BsbwHCN6rhan1SbVZyYzLA1ONA+f
xoDwwWJef0gMvFf0Rgub4FiTtvpyl4BPocV8A/cjlphr3TEV1VPt6fb9Ff1+/yhksmbEL1wBAbhy
4qBC429XGGb3ge0IN9qCn1nJc9Ob5Vh4uJYeX6QjjP4vvfGqziHxcT1m2+zKUyTPNhUMLG9BEXbY
v/cSfuJx9tn236Bady/z6WnovTqhgzEzueyE+Ff62fkY1CwqjFLcIilW1Oa1C8SmgygoAYa5bzQS
l7qLH3aeQzAE0Z68AAkAOtCpWZzLZKoGVegzWkXu8U+BKf9WNORCQWR0knznEVQNGkb+uI8fye3/
sJae8ZxxDT3Dw9QexLE87WrS2ufraMLjhT25/M6MaNlUanCokZBTOpxILsghLKGNK5xtgXjxXIqv
hup/zDgaROeFVqEajhTbMXVZ2lWbmmfBOROHXsR1HO14y+mxbGtkiiderqcjtK0BkbDLVcD5ziXB
uH9Ks468Nlhu97+YSiOpUmJDmPR4Sf8pPtNm5COYiNAUhBG45A/UNLivJKkfiPrrOFqm97LOSchv
jYXVSCBO7/0Vyf8K0iFXq5DJjnOFsliLNoHc2gWbhWZlteqgcKXy52x7MLm51LNE5uf4m9eK2O6Q
sglFKqyuFx2a/NQKv8ClxGT7NlHJLaezYR0ziKZUIrsr3vz6OCuoHvx4wj1v5QvH2YmyXV2tcOa9
0hdi1sQzgZnjyMTkqUvFdvlDVrNT3IjrLQPtDEsU9MHAI95Natg+osUs+421PqLsE6fdzVfuqUdp
126d6OMZVUaSkLzDUXm8FICirNH/jq6GdaHOmW4YAOeEzuNBc7GLQBSxJ8rpMJ/mCGAG7joO1Fg+
EJCHdgEAUDuofwPoL7JnUl902FL6wTTvd4eOZ0YnoWV2yivfOb8fSRB/R4461PrmMI59HnFyJFUY
VUCFMYfcAsNnJEZFXkxv2mqpIzzw8f2I/Sp/JxSF8S5flAaVS87KHzYEJq6Q3/smWBbGH0XT3DEQ
dUabXKawYP42C+rECyUdUkg7OsgIRAH/89BPwM0UA1vE05G9U2OD6EduBBaoMsboqi1/G0MzV9at
dUhkmNsUEaum43UbmzHnVbM3PEV97PT2JrW2gmxVgYMr+8cdebxHTcCDuqcN3uSqKr/PFvwd1gMg
wSkcWYxZvnE6D4pxAKDvTHGs+A6rHODoUpXSPdUo12y/uguUeECbVdWWWz7A/rBuiV9ZlQGkmTBN
nVoDYGhDVMU+6q9yWSZNSWFpmf3d6zCXM2x+U+eA+5g+orcdzIe19znjFkONr6HZtDIWaJb8qXJy
C0TIXAVQ/J2T0sT5AZIm2IEDxyOi9s9pZasMd15Zwuv9hh+w/7f2S7o1uYUgcZQo3iXmvnGP7d4m
2rCzVwCdmePXb94r3ogzJll5UueLtV0WvD1DY0skLA1Sfx/3hVoVS/zW7QUFn9OlVjqdJW2z8SLu
Ke+x7zlQTBS+/o+q3+givduG054tQbn2eaksysaSOWOu1TODtKYLxe7Shcp7yW7iDQ9X1YrGGjJH
EAcMtexQflbUUEbIPZGj6Zqckv739rS7u+SfYHoqaEYAorAVEdUbzF9bgQ0t5fJLbRORlNzWoGbJ
LKHlvkuAeWQY0HYBd0roBxCxPNXU+izcLYyfJmPNFagGTCbuCFA93Ur+qIkxrCG0a5T0nSDHk+XP
7ONj3NYy1aYn07mHt+kgbIQxAqKb1SzIec8mctYB8zte40l7jYMbYFYx0hVRYNh8NjXpn8pIzVcK
i0O9pi3hFueay3sHRQt3BOFpTODmArpLDRxeI4VSIwcKQHHlg3ICp7fLgpx85fD28dMwlwQxdhC3
s091WeOIPiNRImzfKpBzad5pE05iSlCu7jpekDZN8WYsmlZah8N+gtzNKLniV+QMBVUn+GVp1r1B
XvQjtVjMnxyzTez2qcHh5Jar2iklyyAX1OcJDuRXDroPCZ4GYWGIsd6R5GtJhGyzj+X+H6Z2QKNC
Nd+jy5EhYnh1yk2q8h6Sw4L5NOlAvT7VVS+yRgr5Nf/s9PpRNvyg82UBZUr4T/YzoMePAUZT+qek
cOGcU+XrFpoowIzWVczlQIgJKBX1W0Srux0roKYlBHykg4C1Wf95ivm4sl3nlclM5IJelnNW0iky
UvB9ai/Aqd2yeNiP0PQIf9dfdelBIU1Tens3CCiWUHBv2WRmXdCdHaJMcDrF5KQ4fH+v2zUFkHfI
vxXuatYpTYuZOXCTNvrCZo8mBC2icdauup2ApYeFKnNRueLdBCcKSBQqxhcRiAHP8quST1ihyWQa
qHomj6EWQeUBbI1K3nQsE/9Dak1zhY3M6x0YvkzZgzanMgruqxQPTQ2xPWiSJy9Va+LGgQlz6cEx
JApLHDE93CtmSRCK2N8zpwr/lN6B+kxL+2M9GdR4WITBKBatxxnEZVfcBG7A3dwn5Vtj9bBoseF0
NvQ8qLcUBWyW3ACWVlHJt2iPgdO7ne1HGZTTisIdvFblQYg5YMuEXzjSM4nxKsNAz4b3Ok/AYCSw
jY5NWBx+9vq9lryS02k4116WnsVhcNkx96bdiufYJU/its2ab4gVSs8zssrX/Y8FIgvLs74Um6d6
08F6JLaY7gL/mPT9N+FzfGfkDz7MNurZGWHrriPJoMLI8NyAG2dI0ZkzZouCRun6UH9YRtoX4ENq
kptarrUS1vnlBmL/yNrNwMsJZOjK+vnMTtqdvHX6V+VFP1YzIkkh4gYHOJ4atvWxLF18S02oY+NS
I9oiukpu9F5l4w8KVk4upCxwlTQ9sRGkz+KERH49D9bbKkO1uzKrGcbyD4wfgYUDSiV5+4b7R5zz
msQX2Tch51ro/WS/SZEFdsyTVcVhnaSRPylfYy9V/HF87SPzxoRC++9EicT2JgX1SHz8YTpft504
abU3FeHVLFnqeWw/pX3sKY3P68MG160Dx8Ebw0bycaeVD9ZxAl/eKbMys4jKjzozDe47IzWx0E+G
YLwg5/cHf1U/8DdwsdCe+iFAypEHZmZArWb+Zis9IRHW6Cctq8n6MTUVDqn1I7+WRwUWsdr0BPRj
G4oZpxy+1c0oniTVz4IP/m6QXNfjgUOVjbd7eJcD00wAe1+2eg3CMhYTnGiwciJcmurhGBrqwG0L
z1aW5YtpLI7wLRwWM5m6zMrbLfWmdnbywQ9FdYcN8XV7cxoMIL8t2GmuyuO3Ld/51D6BhqDddXPX
D4/Nh8NjSEpC+toCp1vF293CJbyoipH077q5uKT3G0Kasg/yt0vujxme7a21NV684Oxv+DN5XsJE
muKM0jlRn8lZbbDlpJvd4+BeoKfnkmYFSWHkt1zt2tZZrMjTulpRT2S7MFLuROuaQ5Ztmb9QqxCC
M6vdS1fQD8Czf7LYVHQBwzzGOTwm6knLi/YJnW9WYEEH0DfsxN06SBaB7TVWfoYmOQQVFSlC9gpK
+2W1jT3h1xEbJkf0AlwUuTp/kFUo/u0fJlTENixjP06iSBXMsaL+/sQNI4kLZWOdTc/CjGRHtkPR
VDugzG//ihrhFOGl68g3P43CBdrmoMgVhC1UU7B4SEAZVY3KD53qyilAKmJtBsGvnEhqRQ8vRmpj
NyGQepeQx/nbXZYMdMlLcANshLeBmR8wjAwF/tSDYL0qk8lfmRF0v2CMHWze/kpRBTdO6wvVnvmP
jSf5+WutvBr+L9oYkF8tzAD1tHOcUEwVEbcYrjJALWy5iitFBsF3af2zyl/6TD+QAJk+zjRIOwcU
v2J74xYZWlj1DSyLv5BCYB34bYfHDA59jJCNKyDL92pcUJKv27aVIpVtk6wWyMAFGrqbE+NSCxeg
yDRAME978pH9TUAIDFX9lQoyeSrQuDYdMmPk5c/ia4e90RmReREIirjF9W0vFhfxGGcf8diNUr64
/jBovAdLHMYg3wFWgPnMwsbWbtGMGV6gP3NxP5goBeYyF3E+2PcHzmGSl0z5xLTwx8yZ23HDlpLO
PuAaU95m2C2IS6443w/CSXsDZualLIqB0Xg+0ML/y2NQ+oIh/opXrHfRaCjbu3yrifwPZKfufdmG
4bQwj+M+Epvinf8BsIqFcntKZvRw03FL355TaJ4jdlHvBUZrDsvUcrQO3rilf5FKFD9AaM2gMMdo
xuTDgG67wjadqjgYvKYRASq4MGA58N1fs9IAON+hVm+g+JgvyrCUc4vq/1z0xzchVrnJ7HNuBl0k
I34GJXXSxV6PWGYOCWAxhbaR8fPby0OMAd73OyKbbDIhZzVSNzF5KPXtuE4fHKVLKTuQAgHm+PbW
c7F6Hrc2ZM75l1mtnHkBJaggq+ctDCFcERfOvImS9zzkvaMg9+cviK6hNmE4hneEeFGTFpBgQDFg
T4LUUa0W5Sri4k47n4gwh/0FolWEiPL/00fhbN3YrXipXiJEGmndGPG7TXdVEYIeXr4OvQKYcRdI
+ttURP3TWohivIexHUEiUsBGdO8cfDNwl66IXvbqQuWkg/wtIGnYsC1x//CGl87AtNWp5HyBYvw/
YSNKItI+wWrPr8stVkoZNfcdDYyn3fBq15BukESznFpVsJ3DWMpsePQcHtFlDwZcEHNUvYrlybt2
9x31IWF456u90Jig5+M5HmJILyyrK2FGIEUjzCisaNUWCFQ4iE6D545YCCVUyLpa5rOUG70inFCp
0Z2kteIYqj+Zg0f1gRn+de1elFKkyo0ofZGmYn+1xfeduVO2bsd4fE+oK2v8+MFgFWjb8rcU9mjO
Z/1WRqfwH1kAqAd3/z5ElG35NX2KHkboEes4Wilb4ApU3vXwrNCH98NReDYl6R9jRMRBJ/6k1PmO
bq/0yp5D40ewG+wD46j7CbdzawqIVRYG8u6HC3VV/NnSt9mYTQ2f3NRiyXJufdD/qvwX/m7fjmUb
vegM46IF+FwTfUBqwd+NIfZR8Hz0xEbaGIQUwyt+luEKoseohRVhjY+ETj4csdWwyYzR698vtvee
exCPs3+jWg24OKrwDJJH/9YJyaCZ6Askaf5WxEagdDC104zmPnYMn/m8Q6RKBRbVy4q9j9gGAMLa
3dZrEnrzEoLyGAbhbxgPprxb1IWnu6OiG1DC+MJHTJy69Gv2X3Eo0JRpKFtRY6LicWVeJ8HccnrH
EgOpCR71EmstDyRVpERjAfhESD4w388Nkds565RQtYHcpWpn4h2K1skTZXOuLotS8WN+ua1/Z0TO
q9DPXz51Ecm5E8yXCTFb5gtmEJnuscNUaWSJ5rAJoTQgYZQ5CiAq8x7cCMWOVVXdm6brr41yq6Mp
8yR6fgcskaaD7OLq6jdhITL3HdH4lK2mzUrqIjwT5q72Jjs9UChbC5R3QCQ09PZ3TYZvD9nqCcuZ
a+72a7XLYvmXqhMoFKjFi3OH/bEjSW/vvcIrWMJpEZYyU7C4Y55YiRyt5bmUM/hxhwPJvi4gaxkF
/2lMxhKTCE39lR0oezdS7AauDXLtUwubbvaLD0niclQ+xM4zGgAIiy7bEuHhK2ZnuIbqNr/DjFPj
bzvIEWwI7KrKGqfM6LmR/oE/d/JVHtoPI3CfFVa782j5cG7JmEHMxXf4wWJuLm3RM6cD1AVBAso5
UHIHYZJvuvw+8EHSGVF+6kstMkiHVbovTLZeVB5sEJXQSTanh8qsMXO2TKodJZQnHk6h+2CC8Y2p
EWVOLCfxZzeTvf6asE+CV0/fqirh9V/dxGIMHNWrE/ucekrBpYGsCqukM5fuNchPENG7K+IfGTPS
6mC6UyCLPnQMlfE30j86AOChfypzhdWheKaKbIBGM74YtKAB6nvWYbumbz/2yXZqw/dmI29nMD+w
FAXkq66KZUmtFCwCeFX9SbSOLr0pGslfPu2MtZkBYN7VoBDz4kcv3VUffS4G9u4bxMyULT2iwm+F
zq53cr7YhjJbNOarX8IAZ1g7Goqd7Q2pyXSTs+fSSUD+s2arW8wxkoEGAQIUMwYoj87r9LWcU8Mi
B8w89z5z8aCLLoQctVwEnEHeixMRyY04Rc+f+1Pkw/ZL7FBwPsi5rKq0e7nQscOo1MHWDXwUmEWc
eLjgvEmJurxPqXJIxFnMl8V61PNLBFIQsywZsAR84snwoFM10AkH+G9asip3w3OMitC5LPTxxzDF
eW0eCkVO70r3UEsKeR+krDDYGs9TYTZ98o+mZEaN1+f1X6//4ZD5s5bO23yeLZldFdaj/bgk2Fdc
wANM5yH1kH6k3hsvPgTAAmxsmv0A4ptXkwJctVr2AjlyNGqkKq7T/CoKwio1kcE4H4143nlZswR2
2bG/IyFe9+S69jdXI78pYmAWr+pqVvuxs1QCkwOH1H346TZVRGrLjsKjyKaN9tW6wjt+TfR831Jd
XlxgvZ761Gze20IOXLZk4mSnyO6Hq/oIWGG9st25xEXgkbhbRIW/AwcBVDlxCriok6w1HVMqkcXN
Q5mXfcNBUGOU1zCIopbdoepbcNe3zhWP2GxtO7FsBA1KRz2m5hL8XH4V+4SjtB+thP2nklKjrn/y
lALx/+5KBz22y36FOZNK2OBIKbsCvvKN8WwLcoyylWjHaW0Z5P68BfxkAyLAEEipOUWQVbnY7CNN
OKA0sUsMxxgkLWXATp0QhYiRtDoEY5ioYEhVs+EWKc3ptdMRvdoCsVk/W7+tvUfeLEfJ0jujqSwV
iBjIDQRHZj079ljyEcpHh0IYutI6hbAGH6vofozcYSepVyMQ4Sl2QWHPy4LaRPSaLdWGtRgW/ir0
UUp0AHWrpz/rIo10UyzzjpnfvHWg/VLwsYJlPQZB6wLRDccBjB/diWc2mPtQWqUT4k/Gfmq8gn27
I3MMBo1tD5+T+smTIXAJshLsmgrY6UxcoXOnIkeqxPWvkhgPBysHTOWw9mqAkZE+cF4lRiZmY0MT
GAkkMbTmI6tXWN8lNk3Nl7rUVphk7q+U1lK/lNrKDi2yXBousjJM+gduSL+De/amlJzAZ4jHT+1b
T8Kykmisns1g3Nqkd98xFancIMnqELU0l7mkrntdHpJ+/HzKk/We19kbc+2KL27kJIZ/s5HYLnoF
VXOMxCR9gUhqvkIrAzxGSr31tRuVtra7W6288Nytb4BJ/037qec8Wav8CmiiRye73NpkTjhiRj4w
GY9GaCBIZ2b4Be+ISPRNmjjJTpQFBPnkDITDF3yq+Ku/ByA+P1a5kmwV1wnmxw3g9a8nux3e+zh/
PJRGXxkgOqJpvBFnIN4kSGxrrEfIU33vtXlgBVlemuYTOY3/Tu0jh2W2rddWYy8lBh70pOfV+rMf
AYl3bImg6f1aW1zoP3PMRONdEY1Rr14XkypjCMdDvvAMF4hwrXSts5lS/jxyYW1PAY42xkV0Uc2m
EtRJo+RKEaDJjAEKzvpoQPNlQpqRRGHcobTGeKXUW14HG0FE7AatB9MhdydtOGsWjyRSfn04z4MO
dYFmpxqD2M0bIA3FE9mqBT9CrNpQS3p+JyCBRLFmTFgMfk7V/CS0O4IPH387/o6ilK/flkSNKOez
wMv/VQx9iEMZD9TRM5UQvVIeyOaBHX9bmxpBI/oe3gI0WfcZweyevIOmygMz+Zisqlu8KtXOjEgr
A9HvmdQXh65YwnX+8G+oCgItXd1OAzJVn54dRxQuVuf0alprc+Yxhvrzdn6kG1gcsESWaPbr2+DU
KY/k+Pmd+U67UBQwTQibZd7EKfeTzZ0Dese0xYvGhYnqnVACZmwil0yPkRMMfUfSMp9PHpmUd0tT
N4VsJ8YokpA4sm74NFyjiSPpWxLuamIRC163HTfurVOphjW8M5sFPgmr+uaTjKNUr4zp7a8+J+s4
L6PGjtGp5mNhbaYRqW6L7eKwNj5/CEUWhYuUhYprakplKQuSO3EM+bunRbIZBDHFPm7+JsuWkwWt
1SxqPaF4L7t2Ykrt9niaWCjxjlUKskE1um58h8LLrK1MxHloaT8V1sQEDiafBVgZXqaLrGE3o4DM
qRTcUyHHfaZpgJh4QbXHBZn1bmhvFrXeeesFvieOaWiGlBX4UjbB9J0dCMQjlasawBsFJLIgTqoR
Fj5eyR/PWN6GEyrniQixlg1sKdySvdT24KHjTq2nQ7Mq1j9oi6PIu9X9iU5IIrJ23PSNWaqjcJu+
hUwkUyw5BfCI/Cx5eimawnp3DkajkIv3evUrfiuLz+atAZjW/NPcoNm8EdbOPTqPnoFNPrksNaAj
ZvwM0lweoEhOFeWZ705U1zOFmIo3YKPuUpfGsdFL+yoFVI/btP0mWoNObuP0x8Mol3tG2LbPFO9S
/Dco1CKtAKuyEiYdKoIr0m/4zTIG2J4y/omZ3Mgeh520gpiPyKpTxXfVBQ1IsgoyAoLCAMQfQEv6
9ZIRz9KPoUepltnMmO2XnJvPXP6hpDbcXvIod/4ukLEBm43TAwXE5BUek/NxpJcD/WQ9RluPvXDL
ZrNZSoJ7MxRnhfbIiLrAu7w9pJaRETd0tODiZW5diM1xiAVe2+mJk9z+LjzidcoObl+U3tRUV8NZ
7ePkgxl7V1qiBbBb5eM6m4TwfiVGqGkDqY559Kab+Apb0Fwf1QzS9UcZm6FEaZGChuJp4rl9psNa
9vHMCItc6F5Cl5a97jmIYSl3BdL4TX0noJg1Jtqkogget4YSr5qZIv8l5POcbCkSwiqx4BUta8Zi
RshrkCnzRsPqQGK8ysV6ApWCg3rPTNQeMr3SJf6QtbNGLksBc0bQCOcNFs+gcr4Cjlhnc3ZsFoct
P9UoteBpE50gsptD0wuP/jgNBhLMdwb/WYyWbYNb9fqphnYixH/PvOmPi9nhdmpuRtwJ07fMy/O5
wX5EihkG5F+DFGXRKGtg5Y4d4pySWO3N4nZObCqffzRQTOkZhAJyEnyQUKJWcxRB8tD8+4ZC8CUA
yoCd9yzXp7ooppJQP27gM8549YldBme3xyqi9CqbbKgmRCw1XfSt4VSsfB1W9zKCni7PQOjSLxsp
su6WwDOsCVuYESEua72AIpmjNTjyhTZj7LsiU6G8S51BlJYErJtN3KqLMUXjhlBJm6amhM2ZNuSP
9iRWOF6+VSeeJyxHrYb6PkRzwgcsq4SChx0vORsfaW7J/EZiMQw4NlPpR3ts+w+En4h7X+X9CWrA
h0dJ8bWnxSmVzxji/sg4kYZhBDluCSNKNsz8yH7PHNclaqh61CikvpqXJk768HisCpU2ORnam/1c
22F1o6AyG8Z2q0a+Cb57rCyRxJILEoAHBqtwRTwLTsJeW2JxvhVlZlE5Pb88wzO1gc3GiM/xdu9d
db817X0L1ggewTYrP4a9Vm7LnezynaKljsJ9ogJV9B/gXr2JRE7PBSZU60GKFifiKUIZ0tZ5Qugn
C5LmM4cfflLJODV8wQpsZYJfto20wYniA3dkAnXPIfIiPEHcaNrnraA0B2/A/ItLM9APIGBFcHiT
cY9doJNBBfrHOo5nLeZ2CrXp4If/FtEeQGtwsSTFF/umcUQXNA3SgP5LScqJTgkrorwrp6PHvqE5
EkeMwmtc+chU4g4IDx1VaWz7uq4WCYCCDfR27BSPZX2D+a+f36aKocGt4Z6QTqeMIPgnFIwTsoAb
x7sAGOOhhtG0PGYlkIay6sSwOpENGCtn2N9p70DydTtk8S+LKdx2fhGa6B2onbV89n7HRqENtGYU
baNIBVPRElAxyFBfZC6YdA8SsYnZ/MWrKBPRpJKU3StMYWT0ENs5OroG5Qe3G8lSvxDVAR3jvhU8
1/EmSR7Mw5wzTkZw/Bpvvb32RVt4En18TrOmUULbS4Qcmvbwt8rZ5MbhR8e6Mj9XSNb4am1t9jeD
ZhWJawEIaKGUMUSGl+gBgXAiYde0UV6ZqKm89NYc0s0Z4PbBThPDozBYgg+42COtdfF1XjSbwPbq
1wnm3AYCtva1k2T/lfFgxTXkWWSo/t6dFuhiDhqZFM5W6BZVu6DfoULDhKxBWgI468WOd5SMJWLt
UxeVIfAlwi3AWxZ9fD92p8exy80htEsDC27BL3IPnYOqfW/gZQMbK2N5U6PaM5vZN/vAoBVxN+5v
yIcWt2vKhBH5JVKAWv3Qn0zv6I3kKG0lYQ75FXyCKo+RwqVZskMLx+oi9/hpJ7vKVkrCE9PSmKln
eguehBgbGnin013nduOQ6UsGw1d/CfuXGT31q3T2nbUJC77cIt2t1pYiV0TscDw/mMdnF4C/q2af
4ozT8PKgm59jvZ+4mlhTbP2PevCWVSTsIBOs+kEwd/ZUMxHxxnvUN6hnvHF8zioj3Bnp++qh2B6v
VFw9DqBvoE4kHBrjXrCzxn6CRYR0lBosKARSIoN2S8r4XVvMBEcd39ns3O7iSVQFF1Ed7lJqrq8v
8nJ9ocAiHua7DlptFmiliemne72aTkySC4i6811iV5zCp8KC3bRlGWl6SC1xujGtmFLTCSdHAk41
C82OiM2ypYliSVuALpS/hytRd2pyV6n0fvX1NgFeD0ZXf11rhbqOL3VtMHflQLu1Memv3bBKzuXp
jzpCvBmXbYkhOy/YOV5yKr+v7wWFXdjnwIHSxOOlrAXjIZ7NVMZ1ccTb2OBa7F8Tr6t5/tTsPEyW
BaUT3YxZtz10BVwojeaBPWfwbgL1bPOlzEPDYQx+jRgj/jn6Dm0ZiB1pI5nV9ZPWuiv3UHjPuNU0
mpCA3wDT17GbQqHuaCiyhf63riJzIudT+10pZPQ2LOU5a4IQkLhXlz3avZaNZZpNWHRgxF4LIY/p
YSbd8RWScMjaj4Ok/7u0e8kwN9zZAvDv6Iw2Y14r+YDDhSVwwzgqFbFnSWyev0Mas0FGOr5rL5fg
/VtH5aKOfEBnkOQJ1UbFBsMQ0yPFEImazipR5F2i7QYQafRWPmMzN0nBs74HAkyTLFVYtD5k7lw0
vbu4kXHW6gFLp4SqZrnoIRCtsCrE/kuqhL2pJ2kJRMhpkHHc9rRGHd7Haer7nCv/DgbF/8WP+kHo
bi1LXDFNEDwBrlQNP2y9q/494vnHPYzXLTwwJKKmBF5L9t8eGeyamyuSsfDeilHg8zw9QV1G0GMy
HLTd9GOjPRqQhvVAwVIPYtsyqnbJE9D8WqP82KPGgQkJ4zzcj7w9U3ayQlJA4oaQ4Q4roXPpf679
96dlpKLS094RnF8AXXHrcA1JtiTJuCPBEYZYoQF1nzxfv83oFKTatLbM1XpNiYPvIRN7ag2wG4ZM
p5EO/u6gpEiEiN5mKPPq1EPWxGprBZgLGjF8B2gzZBkvdPa9pIAuj6rBCAKh/G8xG5HsEO8yJaLA
AM6mqQOEer4zgUBo8msZVGtKLULwSkUOZieapKRgMtolD/Oi+f3nNVEES5JHyKx4aKSa2Lmb6VPS
tQvQwRXTxTx3BykBF9yGf78AL44RzEq5mea9BHmeShxzUvieij4g1Na1Qgou6u2VUMSnDB6YIkhB
6jaHcSq/7tiFP98e0gq62Vya1Xtdh9xRWENCaDph+aFUWwUAS8BI4W2NqHAzNJwAD9fXvoEv54PB
tfUlFVMR9e6YEI1OnXMaI+RoE2Qr5lDyC93PyE+syys9pPYjI+qNzq9IlaLYYJRbVvWmkZMwTBKy
5R8H5mbhZgDP1pvTMpszPshwpy6Ht6QYSjjpmPtv4EVwFmRFCLV+ZmudoapP8K3VwWQCjQKFkU3V
bBkZkvnDH1gjQOyHPRCpBgVpgAQu/ATniRB9lCzAopSFq6gtXOrF73fVkPCeWuYJ02WJt0zIB0B8
Gxf4dGgZWCk7Wfs+FgEYtEbqzRqdxVwhySMNJJkgMi/0DtSSSM6S2IrpUVbxsyvjcbqVNjvN42V0
gCCkVKKbcSL0WW5mJSUNq83lLhWSXiN5N+fxInAmgoCHMtFoCCjmKs9S7eyhxyVre36ztzlwSI77
WYQfxK1xspvLbct9OVKHNKh+BGUQbXXiJhWw33ExwmvwN3V8dOwmzzpShilD+wgLG9ZYObX+H1D5
A9tkIG3xHOT/w8tp+kgJbirorQOdSEe9Szp1fuzDCky2vXgUVVbvolTjofqC2kf/vkKHeMG+wu0L
rwslBP9aHpO+CeIHAEhNiQsTUMex2qZdyzUyKdG21h5c0XlZZAIUHTK5L4xXyE6susW+HI2Z4L7Q
demnFZxR7kWAKy348xyKjy0fOX2W0YDbD0tEkxRYENEOZm4MLIhNgZqdvf7uz6VRIkq5IPmXRnX8
85JqIgFaV+eJvS57tZFFo8J8V3Y1XsIdERAZAgDPcG8VNNEUY3TCtkwHjCCR1UOnj57F3w4Ayhxi
b781SL0XOCTspDd2KMnPe7JOwZG+7O1ZdC10VaU9wjg2wdZGvKZP120ciTTa3qWr5/4G2rfKPh1o
+0lYGKzPu4lY/elHHriIzbov6UWKqUNMk/Zu9f8oba6x+Pb+VqCR+7EvR3yKhO4din8pDsuRandh
cMrNHAMZwM5QW4AgP2HXjZLSEdWOdLWw2BH+UOX8Umhuq1UoK+EAws4ETecxbk8xktrhjc5Izes7
S078fvQs/a5DmzhQfWkbjNU3v9AtrtQCdJNi6HjE9+yj+42I3td6Kox8Ulsnd65VX5pBm8TT0JDk
buYXTBRkHJoxykXhpC3ui3Og4JiQtBukdWSu2VY1C7MgfoF75TuYLkej5dH/FBFhuIz8Dd9jY947
pH/1qiQWEVrUiOZiQSKZIVZJbP/lG3PDbGJFCo3uciFiGGe8eZmZRT3UNEKqHfGJRhq3P/B97D8O
jwpHUYnUJ5fHf3i9xUwkDpK7NG7Q3eoaKMdbHxxD1q1DvtrSE4gp5YJExZaCyaTMeaA5rHojBQYO
QgSrmcC5dlJITp9sH1bmJFPiU7B/wTSw+Nd080cSGAH4T7eh7hBxhP89V4GLg9rAbHT9E/XABkC7
ucfgImhPQ33IYeT/qQ3SnJWA/s8+fUFTEPOLodIb1rS/XaJCIwxnqxxLwkfecEGDlz1Cw4K8Yz1c
2mQxuArxtaAXlweSw5XN6VvZjR9UqZbrLAJE79qjQuA6+M6/GtNWtiL5dqKckzBtwCkC/86oKmTk
4Ex93QlZJwlY/EGCZYZPi+6xhomnatN44qptj2Y1mp99uMIGcMkeZ0PEiR58rvY8XlcyUOolTYM/
VHuo3lRpD14bJAiKK7nwreP3dciheCzAclzuLKmsMUoZH50+crpl4UIy5jbgIj88hfG+6CpBZZWg
+DTzAJbnb/AEDRRS6ua0Q2t6v0WaxUgS3JNAc6tHIqIPebxbNIcDSXQIca4RoZQdW6sMrdg6i2hB
ig6LvrqErwGOP+Nk8AZvcD0XzagAiBp73HwHb5+8FURPkoPxxEAyxHyC2NmhN+ZireD7bf1WImkh
io7xZPSufK/pR0UMYArEv9bg/93G7od95kwLd8s1f35XFDF3U6eaX9uI7K0ocEeGWXYFQsnnTZaV
3tEYEhAjzJn4y+v4YeIgDCGqn17e7w94PcoeOP9CV9zWJn7Z1SqFjSi5lVaWZMi86A3MhEDHIk1R
M9OLdfz3q3HpuVG3RYLrT47n+pXJ36pHaSOD06Bfoyo+wh9PrB/zqHBd4KOxpGSwnJybKWtthQqk
4QrNP+qxccmZYAPj+ZHcqbDAs3+QKRR619oZeQCx5XAl0GiycgohhDpn7SnDZ4epUcD8thXAP3jd
VmXu6v0/HQz/kqwPBBY98B/wb1/Yd1fXWxMAQtdPasLNh+pk3tSLZpvuNm1WeVEvqozUN5w/9EMZ
GHQbEfkLSXpcN5L6Vf1fya4UmoSOi0ZGsiF8oqOAEnohFRDx1UBGiDc7shPWF2QwaZp5ptAbiEMP
mCyz3OcgOSGytPpp/chcTA7qITDs+DlAet0fK5PzxkmhtfF27OyoN043usFexaxs22bwYH3I1KWR
lNNfJ4/Y1IA82iI5Bg4rFvAQ1WVCL8QrX/r/+yyjnmdL1104VDxN78gyqH01/V0NsVAyX6Wi8yUl
6fedreAa7Yp7gOt9x3rmIIl4xW7+LIbGYVWIt1vg3XnwkJD/vZCfac/la7b+GAp9VncdpCCf8xka
uYRKvdrpwVMXMAsBimRvFSHl3MHki2Cw2jXcv+dsrybPI4uHK2m1OP1sJLVRxBGTg8BrfRyHjqPs
6XauC9UVLnmXZn63B4FMBVllJW5w5iPwEVMjDu8aur6b7Z7fvTOOR7VTYWQa8sSbSJr3aTGLaU7E
51kG6OKyzB57gNbRtofPvDvbmA+8GbFcpqnO87dU3O9r9kkzNCASDXgN+Dijpe2U8PnfeGr1/V0S
WF59yh//D5vlqR5YjFDd492le8sJVWhEPCIaE5Y/jRiL16p2QXwU2drbCd+Wd+HwxC1Nj7YOGtx8
Tbwop6sWMV7JkgTCSHpLKAq/9Mx+fuEYFdpfykWK+wW06DNgLatSAGKZYcCwywjyblqKwW+sbPZG
4meIqp1P+a3q3frHr76rrhJ5xxQWtAGSIdw8DhojvbZzR04yURW21MSacBNZ5+hAsnsK3y4vSWXD
tNWmutlLwMrc8Zjnb5a5dNpy75h+jaTPgs/q+/fG0ozse6moIJXwO04fgjEkXPmffjgfDR9CJztN
hgR1lW47mSTmoV/O7EVEsH3SGHGzHuDGj09eA8O3TeVLpmidRtfEshCshsde52iTWGUOww4cSZ9m
24qbYQE2BZ1Aj0H/82+w7OyWLLfNIQG6mvzAvOxuWdLgELE3tgjTocS8ExSIHuSI00OUVmWOP708
I1JjoUG5aVjTE+VdqeTLp6FaduoivnfZeJ4lnpxNFZU5tXPOQPwK/11CyFjgfnW6fh+9K29g2nk5
xNynaxsNj9YBYSR2cujYNYaYWInf4GfUR1Iox8YxqUUrM6+m195BZ6AXuUUvW67gF3SFQzqEMJfi
hQKiftUPTpkbO1RFATHwfvXZINQBsyUnOxIKQjgmqDDJtWMzxXuKJPI72D1BDY52hxMGr4FWDmUs
6oSFTqHaBLgJEe7f/C2n3aCbDRf7IS05o4BkV6n0KEkmBpzNCR66asOylhyHSMIkxivVpRVIQ2Dg
UvQFihever0C6DUWXAarnkd8VCMZA6bq89KsLfwgDBfqPamSzbcxP/a3x1ryu2XAMJvga14p0tiS
0sGSDveSUpgknqy1O5c4HkZWrHjz0xfL89ZCZeQttSXe62dFicvXsLZ5JZUqku2RiC/XbIOF1WYu
P0ANwYaiUjSZBAFD36FaKFarzs4O2Chz46rTcVIs9vPt0UYdMcLBDEhx+Pr+ql9FE3KW8K4ChgX7
JdJERaUvTZZjAcI2kJy1T0CMmNQo1u2+xwQfiUJNJljh8/oX2Pco8ttmhwpTOPToRjFUGsoXHLBv
MsyF93hiIRqWCMQJby7p/b7yZ72+rRfNve+5kWwm0+BwoTA3cDM9xokVrYAOYjObdSIzqhNvh7uj
5rAYgEHt/HGEvM65XjxsXwOVylUcOwulXSH7bMVIMxul8zKshzqvPL9/d4IO04SeNXhNWYDMufaJ
uhKlDYGq2l2GVWpZQEFYyBhIn9qwqpPb5/KRMQPv7vPvo6e4rnNHTrOc1Q5H/Sqxjw/XPfDxQ2yf
+ChgJI3FCTBZX5Zv7DqwP16aUzckiENOd8HWS9NymPIAWjIerrOIKqyC7BjhBBTtWngzRw/35F+i
Vf3gglJi5Hj9eUV46SeEqk9SpRZv1Geyfw7qomfKmBWrhQcDzoWMIVIH/D7mckEA4v7qeNUJt6gb
LKkbPzkrMbWXSxVfwvcc9qdNisDOHaoPJaVoV6EYT6H83i4NUybtqLcMwV6l+K0sYU4Q/4HZs3p1
YFZiCCQdeUNzygdkmfLfct7Mjp4wERoYACWZID/cRUPTt5hEuw21G50wh2b/EOPwky9vLTCdwWG2
iu1gpR5Owl28uAaDfGlrSsUT5TqvMXsfu+clvKP88eSBlRHo8SCaqypABxwPX/PDl6AlozVCNvMA
CbpJ+P4u2MyK7r8ZMkTmoX9/CYbwSHXu2sUSnnxQIloq22M50ICq3nNVtUmQ6sL+RvIlY9NRgXcP
b4ZrfLWUrGZo3m8O+/DoAotzcyzc5rj/paBBcYRrDPbJctX8Ovetc6J5V4+2wathexBWecgPMPXq
l+1U6OB8bXVff6NZqK9F+f5SzA4hIB8wA7Q4G4WwwYzuxEUDqBuI3qv1okWjhCwM09UMXgXDRiiv
hG2fmgGvo85JFwBiWe2Eur5FtUPtW5b6+nQ1mmltrIRm5AZ9bJadG5CDQqC/rUpBdJoGDvH3K8gW
lFFvDJU25v2F8gcFNnUNctkb4Gad12o55/fDfhFh7uimWgmr1DNMHdFGceOMh9KFSMc8nYjaFZ60
lks4mXMdgfXkjXlrFxQqBphzfxyUPPyR4PHL04ShYiR59p29pMZfWjT334EbF+LGGoKMEM94/mEQ
nP32Jld2AJy1DrfTbWEzaV+cWvHU/eNz5NzQkdqXP2wqL1ZVNNAG4uwaEgAUFPMwpyMyxoy2KeMy
yyWe08Tt1GkysKaJ1FfVZOS4qxqkH45lBl0BsMQ9gBYDvw3a6eGUUT4BIYQeA9/4/5bWFVYHvX9W
jkQ5tFbkKVN+vbyyFXLmpBLNlTvwgAmRWnYYrmcZNm+0ulG9CqNQXp6ucFACjD0K6Y9PCDvAfdgs
Cppv7q4Gl5DMsUv2lOp+E1FCO+8RFUL5t1dumQITTn3fkIbFIxzrFY3OKekHzZr8GOapd2QNkuS4
AYyZ1NgzUfGm/pis7dxZFdLtPgc8YN/4PWbB98Kag5tlNssOVclMeKCAtbJfy8VM8nlpT6gPeZ1Y
X7q9odFsuydBbx/e2pT02y3qmk+OeG0ZsfBwgdSJAwDe/tNrgFPpHZMyf3a/EIqFv5l4HZzp2vty
vlJDpFdh6uDarkXlSAPZ42XxUqY37dIUETRUa0wHMX26MwredenhFFzMzidxKLz7HDLBsZHlAo4A
u3/oFCqEPCD+l84hTgMkdZWl6R16+SUt4XViTxCc7WHp9usMVIFqx/B0kRxxz7kaYqwUbszBvbNU
MVV/2yU7iJ0HkfozCg3I47qndawz7mJ5kzENPErIjb0ZLjTCYRzziIVv6l6ixz3joYAzYf9a831t
M0uGpLQ9cmkGaIa3NLFg8H3DQKEvJAqmyHVlYeIaDalqgKHR5P3e5S63mihV8OD4qAG+L0LXb/pG
/R6evHxAXEfEF0iOdBR2UR4VOUbI+FApNqIPsZ6o3PxCh3SsdULrcAjsa38TqNqYMySDV02Es7BR
mo1qYboRV9PIPa2MCjepgKhuS5UVHk34DI5eCV3WtNcC2vXxNUi12EheMMcxS5sd49TpyUK94pLS
oWIZOMhBI8OPN3fkrFESCuNlJWwQ5rbaVRwhnAEb9kbh6ygLM9KLUsTr+4kKncIH8Z92H5hj/Trm
ZUUWbwkJlQ/v+WBWeEBPQJoueScyvhhxc12T3MhEXiCJUMDdL3Z2XDyHWq1U2XaAcZW1y/rI63yR
7rO7k+QdJOESYVwbDZOLA2x0wrGmlxzotVlFunbfT6Tm9rKeS96yXqeq15Dx9K0eIsMpZKVYyT7p
n8oCCzD1j4aFrhI/IkRGmzTOwyI/iCzc+5cxtOtcC6avMHoV7IA0yTpe1SNb5NSO+ITTg7ZUSeFZ
SCtv+XB9eACp7DKZY3WXtHVoYG81xU57/JeNRZAznFlyMLpRq8YBrAw8lGfeYbniaK8B913FkQsj
3Qwkf3v7QJC8u+wkB82RElWa0CzwcTQ+l4pOFNM97ODKGBL918ghxfNjoTKiurwIDWnGG+v9ZRnZ
ZxN9n76gdQ33J7lgWgSi9mtmVjbe5y8uUohispAFQ+aA67+x78g2bvX5kB7IzfU5E2HjThb3T3XN
0ogxh16mypvCCyTCTWt/XZ4REFsEwP9kIp75uanSQ2oc6kQA5Ve2ejD7QiZudJEObWOx12GP+0cn
ictFajccn1Dub91OY/yApqyiiVtM6BaQCvnMi9gFv9ncuZ1udnfdbbvD9amNl7g+cZww2iJCzncx
WZ3k+6f2v8UqGHDTGNBHlJbg1B6JInLXEghN9j5lx65JB1LWsCnJfO6bxJLBkMR/D3etY4iF1C9Q
lUobJwrmTpdK8JdgMxft9kptC7FmOBMZM1kTKeJXVkhkQJbGncAuFZKxUQMw6ZorR7QKk3DT91oI
l6XivlLYMkRa3/jTf/IKqbS92taV4r/8vwX8q6VPboeMgvZFP88MPZ5jvELdeoPCs5fvV6QdysAm
j1OOWsg35HkwrMyl45jwU6tRqfVbzCCjo3luJ1vXfqQGtW28pcieE2qC78+iXWa4W7DIcoE4FW81
NZlvlrWS6q0gH4eGZEKKDqvyX0bPtcDa8oVMEHfBZIw5+c1XritbJkATVC60SVtMSDxJTCFbpnrv
abGE4wSbnsXf+SBzJAnQBn7tj23DXrAM+1o/yoJLWXkhuGmDUDmm5ev9l0/AzH5GknEzVmFAgCLh
XWfphEBScM+3xd+svGcYEERnQpWYHxagM5X+aS9AxZ5ieqnuhnTZPwR6bMx26ff6BZh3KMo0X7hF
q9o9Npitnf6fE8r5UtNKDo+hhEZG0ZIXL2JWJ53m3kAgd/nSd9SP1vX/roe0VHJelpHcEpe4BKvJ
12BbUFHxy1/vGVT5fZATfYOlJpNBElmNd3dSjeSjcI9pGU2sNEaEC50aCiko9AiunzAs47vWuMz5
Pd6LUeyS812URnYQFhI9PcAFhHUdRbXAc0jmz9hjvL7zu/juqV6uMQVRCUxVAxRm0UEZGhi0JniJ
/njNTOxkL+IsSZhnaeK2Uik9DkQGbxJQTt2WEDJi4Aycns5fBf0OMRE6yAwjBwOPfb9ToVd/1f1/
fJn8UEE11fr0vboWD1WcWB2ZAhD/cou7ushPc6SULa5AYEBx/6RK+YWIhuWSnEetBlUrzOkgyX7Y
3ZPNb9iEzsEjDoAaNlAP1X9fmFwgNi3xahWovLnoyEM3ERZFlx7QaRShAl5ygXKcW14W8hos6RIX
whLTe2doj7jdpItFjg4talr5XfkNm/XZSifpcOHZnjcqVJTWCfvASrjSP9rE+FoNqudhibJBkcoJ
udGZGPtWp+03ubuny0BL2rv+RkCOtBhOvAlIXWCXNGaC+kdxpScQlnFoHfKWKweYsKhszDu8nBxY
FjpjRqCN+XXr+YP4bn38t+QTm/wC6rdhsjjDNr33DzgeGgmYjhPeWfprxWst7qR2S6k81ImhHQvk
yVdN3H90PJWmn7jQwWvW0etTzQkbLK7EAmERQ7rn+sFmQHqHFgAHfETsXNU5e71G3MgM9yK+33ml
cj+WuN+qs/yzVWnYeUqyYG841WxiD+Cf2YMZ7KnWkYhSXGPh3QBtUWVEPHfJDr1yVMAjva+3BUj4
X2FwvRXPWYgUcu0KmwUHxsUms15cjdYj14bKtLJ43zld/0XhhwGlwGF24FXYauvBfby4Zf8qTbTG
KaMtebgt5G0JZ1634wOIuSRaLkwB/aGdQ0nUVQKsq2KPC3xBv3p76jPao1ftQTIIQR7a4cDBKDXC
3Eox9meDJ2SNwbz2A40wl1EBYPj7+Iq/JEcZpmGwo2JmZGwBJe2NU4OkFn7iBuJ7RmbSf/K1SEMP
cmS0GfeutQJp+rLmOEKWHSPMc9AuSz5jSBt/VRQgEPTRwFnhrEzVdDHxrrKjPuCKMCALiVsBAAxo
IcCCQD6FbcW1yeZ1xlU/9vCYG+7vu68bqBV1eTUcb/siAca/yibKqPSEg65rfeTARRRTp6+JvKUD
8686cr2Xsy2dQfTaxVbIWk2vLsop0DL23T6wioGLVyg+1IrbDCW+ICtwYYVIKgiuTRvQtc1xH0aI
8KtR+P/IsPtSZaku4RW5lqzYJVMrPyfHWvJgDCWHlhlkW2KfkcSTfSHw4YeeaaZrQ33QpnOHQ6RE
IYxv7WguNQwJ6T/gdF140oXjK+BgAPx0DdiRwVaXoPQcF6xQBOOe8gXF+kR1L0AXRbrnBKBI3F2X
tKpzVqHGmCeDiFYNpZrFOLrhY4NyMojWlTCa9AhoN1owYCVeIeNZWiFnUoH2OaOdhv5Emgjm7/AY
QnMmXH9vDIT4yXVMqNQ2Tnhq9vlhEWyE5lNhTtJfDBFmAiciZ1U7iJ1Ns3btJgJz1HVe3RxK9/lN
aFHOfVLrnSZPaOwST+iDxlYqufPJOmRuhxwqEHAdX8bjNjMNxdmr5hsveTUqfp1+dYgytnq7ySiS
/kOrlDa7GhAAgRYCuX8ZWyN7AebJMqDjPdnXPU7tFE8tDhBA8aPqhxNWtMrx125ycnu2QsGIKq3n
usv19NFePR2K108/n/mL3+7JYco4ULx0Zk0kYHbGOw/qvoSJF+L2CGa1WDF/WeySsU6AtJYGLiM/
xmfGy9EC9ZwvoCgkWBUyqAG2JI07tTOzf/ADmbn6kY0B8yftRnz3Yzze38CeR4nrIUTYDLaYqU3M
cQ5sw8E0+pvrQ+r5KEmgeP18UDB2dL9FqaLgElKpC6VWDJbznLyr0U2+8+Gv7KXVBZ6TT2lnWYpp
ngN3lHp7GvIjI/17CrkrIXTVqClYa77rCa+spne34/do/BgEWg8M1Yjh+V9JxyuHVvEdzHE/IHwA
J8c/gog9pd9OD6gpbo7rfI4LtctCL6RM+JwYtGd1rxW5wCG/FNuIB21wXBDkEhF1RcuKUTr/AMxn
2hom5s0iYIJ28y7nv6V82Clzi5GmbqW8iYcQSlOI0SQezmwPPaAg8lybKXO3PxQIWuCq3JkjnCBZ
rF4z1HFESAG78xB4Vk+wNEIemuFecvlGcZ5laQU1Z/XuKMCtuJBdIR/f2BNbl6fis/XYTh7j7rqv
Z73hv9MHF/39KkhhsnIXZdQtWQRva8uz2Ye0EV9/vIzQx9eXxlvGfgcAdYJzuq5/h5BaJRRpciYo
eAu1/0MFW4obLPK8unEu7m+NOtBlNM2OoQxcunBufVS/gcBIbjlGzZRcEaz34x99eWb3u2hULFt5
zbuT9szxma1NBsacYw+8bQCoa/k4sXAzvOY77AyDovRul74MgxOD5AZRmfXO6oM6VTi2ZnhKkvIz
EBuL/7HZ1Lzi4Lwy52K/OzCl4dANDRN7sL2t+MggUUSYp4Qk1AbfOIJXILccNrUr/Gt4QF5AB1i7
M9yLC4T4ClmGGYQEX/HRqb0wEN7OUY3oF3113o3LbnN70JZr+zSc5iKDrMpQdzTJfCIzPO1cgYQt
ciPw/lS7v6xvjOtJXmJ0Q+k7VNNdoNy3jW+AyW/hs9ri52I6K+RJSPqSM5hS5dc2WcSg6BNHX+oR
5VDrRFbWPfTtY5hIPBszZmuKQQWNSsT/WlzjGl0J8IQXDi879B/24MEoq00+pSDwe7M2lpmGOvEF
KFmRrrv3m3cMN4GKzsPro2g+f8aVS5cin7suFwQgM1N+1sSFL99RApsRKxjzE6gFyhcvysv4p4+A
S2LG4AQDb3/zcijHYjHcUS0eqZhj0vmcdp3OC9KFhO16nI/pkC5NEExuKsza2x7RaGgDbsNGLbVK
QSbJlNNQ+ueK1mmeJRBFiWKCgtv34y7cxesWysfbG7P8nVVAtLMmmDdJ0Al/jvLLROrAW1VOu/4/
Y1DmjLgTIfQqqtuCt1wepuffmXv7vQb5bz3BgeiCw6MSzE+zgKOZuSXvj+FpN5kI0NGzW4s9n9vx
DrQt0Cb04mL/3ozmsE09PMO8c8I0ZkE3y24Kn0xxt31mkfcpyLAlgD3Qdr5gF1SVn9A6QgLmzgbN
Cp1jNTYfW93cYYARGywIrYzu1UPJ3jiTna4p1dKoL/dfYQViWO00EgsKIcd2pPsNWcjEoL9UqKoO
mA71uvXt5xnn7TQTB+oils35j7Fm7Fd7X72Dif43t3xsIu6WXAwSMOLxbhuSHEqb0PkX32scsHwk
FR6mo+0qH13vDEoiTh9nMGtSe7TZZSoijhkJvK1ebDcpBV+AKbwjm5NEPRV3p1KiFUbgJjpzRDiW
2HnuJ7hRLjK5Fx5IZP7I2pLrflIqNyWahGyfzsp9X2mJnMcaCTLYrqfeiHo6EAymtdnrCalAd0LR
v3F1ZP7V5K3AUR5rt8bjHueBTm2bjSzcHdVuanzrD0yvcz96nRM6o8LyuVHrEq9gpzH+XlQVIxg9
iEJIopLHpwtP4XDBZ+BXQGKsu+NR1RDZvg83TqlVYi5ls6gRWQ0W5juzDEAjPiYVwlYzm5Ez7N1p
PKeb/8J0PKxKeFEyUCNBbKi/QFKBQEUh4BafY1LlPn31DvJRNugICfPQXNSLMjmKybDy9Mc9vSDa
vI9fRh6i6jceOdavEy0lhn2dVAcR2XPTy2j9ZuZ+/sgxDj5TOofI1Fd1/gTtQACLKkiunb0G/b7j
o6J3ESx1Rraas3eYouBhmkpBugmtJNeqWz7zpy1gTxyiVkHNC72F3E8yKhwgt7Hdqjy61uvyrKN0
MNh4PbXLBGyPq8fWtpYl9or5yzlko/CF5agZp7gdfH0zwSvGsZG3rDGxHdPrq6QnF2zI/3J9BzaE
EXSTTCXfF9vFzFEkEnZuf68yEXC14Cs+jcvQ+tzpmCSmJPt/JALyFP03PU5aOUUKBxyd+60Q7/Ur
yBTtlJYdPpraGhEKVQazH4bFsxyLowAB2yaxPMyCoHpIWEXvoOt7E8bhM6ECnBBGPXpMsR6jozKX
i5ZYf4w5jggN6rUxfwPXm4zr0Lpaw8G8A3c0phqKKh8JOgtRLhHlcHMbDpEPVXR26FdEPpaFAX/b
ks31a6KRsjhNXntJgordysOk3LvV0RkdltV72/ZU7w154Gzc/aZkIY61wTBqfZ5F4piHBjGEcqPF
vvhwzCMPeqokIUnWW7vHueSrKLIf5MRaYflf3rDwh7I813bo4y45O+vAYTmLI/5i2f7MAWWqwEOr
fr8t9tXIDATAhDaFVem8PLPD/9/+WIMuT9wMStUbonUBQN0ihV8Q8LQfZsKonjSJMX2DFjXcfTmi
zIixA9Aiv3HW2ITygGYnRvSVXa1P74SuufZ6Sfv3VY5gTc6EVHDO3px8lgXd1ktFur5mbQTaCuqn
2BWARO0yLGC0RUVe4UvLeSg6448k4Cn7PxYtitMo1BZJ0Ru+oB1n+e6Oip3y8FMzdRA4KeIBAQs+
05UQTugYrsFRswWe6vgTvUB9nIcBJXMbvIIM+NAqrkw+n1Ben2n8BEkOcZjwTy0y4P120qFwBuPY
yc+HC1z0HoR2cfUzj+wZBVjGMj+/UrpJPGVDuN7Uh4+QqY2/fcptB5tPPikzFRYpq7jS1+TvSLKR
3tX9sous8bAR6SsWAvFO8OMgesDwZTpESd+cjCqcGBbcz+Hh/MmfkGFkebaZRdvk2UJkbFlV9wna
IPob7YFgrLG+dmuOOwl4FCioTgRsoYtSLjBToxangUU3LTEMSBRkW/6IyPCi/oQR7oDlrLqeO7Hp
mgCFeACGvmP9Pn4BF4cxVZCSBLI+8GgEccMYIQkhW6Sx+sUcrX8OvzsiaIT/tGShV2t3NtHvsooM
kdlT7HVYpgEj+lJZslPb3UDcVBHbWa1n0TnJxzcXmlCI2Oe8Lky05D41J37hOaxsq/P5bWPz6k7S
KC27fo5JLnPWPumBQ5K8QUa9dwRWWuqwpol9ScK5RPPZZ4c5DHr5VKFViDuhmTgtxOae/CeYxSx6
GUb6BUxrMeT3MXPgvHsvVYutLTrXRYH4+R7hYkWRQP/VPAVyQ6jSRcg1VowiGTRJeItU2qpTcJQp
2qcFbJpiTgj4IDz1s0TcHDRR/pNnKfnp0n+jO55BIxs/ZimO/0P5yEMbn6KHm8UOkMyYb+yH0ib9
grvw3e1GOEZ6dhmrmFWGoAlnzczPcXmzU9Kl94qgDJCquCrVPecD2+QBUzlLpw3B6tpNht6jRe8u
jPj9TDUjAUk46EsKr82cTP0H5vPs7CZA1s6ovGWAOQBZSj5iPj9t4k1vACqIZZsFa6kK0akehrr3
po0Ews4mp+9EnB/Hzu/ipr8b6c++gnE8NrrjGPDfwlbnHklQBHGTl5uTvpSyRpfXPffnhjGT/fk+
fzqonxkyF+HQ72Ss3SBjfcBnboEDusMswIcmHPSheXJH1zdgBchL0lBZ9tfYe0+gasLTEQB/p/7S
MUdDx8QetYbcjVbzf3c/cQo0BZASuN6HN6ELxU+x+l3kVnCZKW8phmUXGjblYf12MCi69KPIS/Nf
zdf1SfA8rz/FEMKdCclBB37R4aiu0AlmS2HtVzz+IUWCupz3mTvcRAvQjuwPANxLf+MBt/BdBdWV
h8rGS/YmVM26bzRBHQn42hMBdaD7ulCnZFqrRvllrfPu9f5OkbJBiWUvhTMiu0sKVWOUqNBKao++
h9oFmq19Neb4QTbppMc2R6l5i9n44dRYC1y1/QrXP/8V8vdGEIYbmm1xPu5uMZ8FkTvx36yh3Qj3
smZ/WEqzR54pQTdXSgKQu088Z0nW7pA/1SstihRqwjMfeMofPJVK9F8dVRGAqiSmYrQX3MGMk3VM
GfSlys1d2XKfoRy5+4XfVBT77xO8ooAQJaQqL2JObR/7BiZ/TVXkYEhYMuxdJIJ/oEvYL2Chpn12
mcCZBQ4T1bpcy4bD6rG2rhZ5jm108VTN7IvcRbM2yxXLJrn5xZX0U4f9GgYdEWMgwaozcCdfzbJd
gQdCl6FJREkXWq21FImQxnr17ecy2RBkawxr6sjKQpkDTZcH7+ESSKgJKBzec/BrXC3fO5MeIFlZ
f4aDF31c5NtQHhAsUuK7ygfI/7V246WpiaesAfnY+K3+sggqkxpkFVjBQ1VvzHEapCuFDq+TGzTW
7zahAUd+Jff/bOIEG51lU6c0jJbQH+2gjhJdXLRRX0+knCi3T8/XDiOhuw+em8/skDGLxFnYYyp5
IgRMiQPzrOmBu1WTIZC1d9RmYwim/g8eCwvKSdsV/5oK8AhO8PUceHX+GZv9PTxtNwOJHLP6mpvc
iXPixZV+89QsSBUVg12sEdA08XIbLS4nL26KGzofvecMZXPIZcd3SS/ZFyXu3/LUruxZy5JdBgfW
K7Iw+IHMySOgLFg+rL59TQxBgqkjkgzSKcHYEoj1WhE/NpQjULjtZfLpvjtZCQ7itwkugRij/JfM
31sp7PfVrxMRdT7GkIXJXY+1FVHP/iRydeL0MGBDgkV4JEPgeSVTfW00nT7hFf/Xhu6757z+WGSi
2C20x6x1AgZWOTr+oLm8nP+d8O+7kcZu0kCxcugqxDQAq0Jx/OuBBFmsM8osTYYZXzQ3EceAtmdh
pRx2aZhyRLJZVnfA7cA/6XGM1q8HTL7rdMSAF9SagvyQyTTf5DsiiPJ7oSfjAfusRD1FeZU6xzC2
M6PDgEi2Zwx9BcY90U4HWR8QCTGaGmyf4EzFXz8dql3SpUMC4D/UAS6VAaWrCH+xi5oEBg2NBIGT
qnuHkRONQl8jQn8rsPr0Wk3fatVZ7PiQw4X5ei8lryG2g6OQnROMd2ve1PybtlENglRQY8A7Z16m
wJqSRW7RFX5u/m+EUlWzO/uedah46tsoLe4pf7BIOI1W213daBNeG7JHCcGzikdRgIFO/tyAXpWa
Zj0P7UIB6gWPdK6bWdjhwhPKSGjggTQsMoN5lqXOH24OKFeLYaGWgPmtjLFvtPa5W96uG5iNDg70
PXcBimMo/n0gksc0cLDhzxVoOXqDGsiLTvHM3CjL1MyzhB/rLBTzNpOGJxx929F6gvQuMsek8P8T
pndtUmXtst7itNzaqAFBxhy9hcrIjKu/ltPYEVJADMh+UsGbmYwjpRCcUxsPgW9XflFTmqYnNkPE
973Wv5o/ZlRdwtwT5fDvIFcC8NtvvS8iXGpnPx816KorDDtluSbm+HwCoxKUQzvekya9Me3RMh3P
W+DRZnEFMdNbdl5etQcvlthegQyfJQTlS9ueVSfHcAye54NC4E3QybI65qaOeQxzAyAHe3ZsoLE4
xPbBdJo/ml3iEIT3kdxGYwDclp/sPZ/axCNcY4SDIf7UvWmAV+9t+yME1sf//yrmIoRgEOI9ns2P
k3/aS94jKYdpERidClNRQ+QG2K5vX3MuF8Mc868jbT4CEOFjMJI+X1NfnBZ6VgA1U55RmuzygI6t
ruqolPT4Glt0aL71o5QdEb7IVTK3oh3L1j3TSWuQSsaO9wEc+L174LLogI8jH6knCj9MMInHHPQy
z6E8AdrFZoVhKzpk4EaIg1yXjSWj19JCpYaqc6SyRe8E4sBjrToDHgIPjkvBotfig84Z+4Tal8Ow
XCGIj0NHIRl9FXUNv1kGi5Tn4SJjxePtuVLaGzbZtkPvLlnSREs6ol9/vhlenjsGi8YPwPStRl21
iLEZPo9RBI9ZhZQdffg4Ehhb7xlVnmkb5j4YDSo00tCnxUvm6pfXoEi6cozyQXIJhny2FqW9dROK
Z37UTG6fccYPJXsvSPxmfigBlP6Fm5MT4rWqInmJ3izhVDRKOqW6am1lFFWc4YbzUXsJOLj+/y6q
LRrwaoTXuZGA6e3nVyGTi+JrHtaGHwp9i9Bc0qqlu3bKLtGNdO3PFG96XNUiL7wxws4VtmERIhc5
5urxPhLHwLLX2/n5NyoeRJYxFBNMra5uUyhRmY6NmUZlGCfQImaKJqzVZdsoSNg5gbDyZI0kFq5w
ripbg5vkMKt0DoL0tTikKWnazQllVLBl+Bo15LvcwG7kFnm76DVhmeC5suNbTGe9Tw3u7rI9QFd1
YbiZ/tkJrbzy4UXwjNom5SO/zPNyxyHAag3/K/igrUQVVn7i44kodEOxQK7KZ1ytaXItQbm/KWgL
cab0s2UKADw1KJMCaLfVy2O6WuOOGULoCOJEMF5chPsLP4laSBuRii7jha1xJHn0tKOvQyTfs3tn
A6Mbhcug+j73/0j9N8tO4M/54JYEeUxmY3JnyNEZms+yn5Pb0ZMIGBe3CEE4U5k/LccS9AZJuJO6
OvkPFTwIllnWwXqKEOfcKEMzaefrMNyvthbehkEHoI9UBCs9N/5FP+vKCp1F3sv8XYAv2I19nfip
O1Lgmg3k/JZWrkGfeW8qBNgu1j3Ke+o2lmSwi6vDvvT4B6FJM8eOPwMGXWbGtorzbQTZetSIZZsn
J4s1b28GRTh0J8HMc7xWxsEFW2QhqMB8+F0C7jUo/jsJcd+6Cye6ti/I/oUU1Yx5FjehhS4R05i7
MHgFOg5LxH7ve7AOTZB6lIgkAEqfRwb2LT+QiAk28rjXu/QZurRKV34LuiN5H9TubJYF5wNewMBz
8Zc6LbT6MH4P5UPZpvm82HhNrMfERF7stLPZZjg2N6baG5lXeZGKO0IQmjC2De3iRa/qQb2QIC8l
3HXh8D3X1d/iXV0NerX9+6WdDM1fNY/wAiKmeugYwvtitTWGXUMaDSSYnhLdJTa5J5Rec+8DipdZ
lOPc1Ce69xtm25Buz5UTkztUyzbSQtvUGhS0AASn4bhdTbfBPFSqyyrOPWfN1HkoovEr+RRRiBTM
V5x+Qk8zPSud+y/ixsUrGVRdJYABBaiTUnCJlKlzOlanUMCqj4Fazut5pyi0YDgIzi4B/OeI58Qc
e4tBp6uQyhZlrYS0bfQHy2+hmFwCNw4NU25VpzdiCB1UAROMb5RWXomJ3f7V/MA9xqIWWoZDBwAV
ID4sUkgMcfom/roC10gPA47xOW+99T/ErtmeYU/RZiw+x4sSWU4twlyuNrHFQ9oBtzM3+1uqM44E
LhW1Yzjy1WXPth+Pj9qUUGr+rBNukho0VqssnjQAGiO7M0HkW0Ing1TNAhOPAY8S2ZvG3kcd5ocg
HlQf0oCZRtLeDAIK+tTlqp1wiH+thqQSLfKCoJGVVlUkEozujMOejAK0p7y/ECauVfYSm5OAzN5C
419YOkXZtkfB94WhyOZgAL9SEWfLAYSIaftpiBuoJxQVPD2y2z5ZDjmoaBgud13vWrEvu+KXw5I4
do413pXszLk0/vM8ww+KDvsc+R6BwvraNdOedle2KI3H12OhWNIiiiQxvB6w9Vaqp5pTHOiNyPnt
WIKoLbXrAVRMIg3TYpVIgjOCkCsnAsJMWwezfeMp1yRvJFayqJPPpBwv/9mNxnn/qdtxeSTmraZU
5te2QGEo07oYDcJI6Lj5SrPDktH7i6QCxwUVDq0g0yN5Fj/sO+dBddLRs30mIf4H/IF0qiOPcL5X
IKELkv6dF0cS7bz01CkT7S5UVYretoQemPn/jCr2pzi0okYHbUC5Qa28txXxhxYnTS//63iryfAP
OIEpLEaFebRYdaWGMKO4MIb/1nqlR0Y9wMGY/IYxHp0QxU0fFGVOr3+8TFG73d7YoXDem6Tr5lqR
zBvSfFVcil4ECEVMczFjdYLJdPPeWDuxaR+hjBkjd2MW9k8FlLZspH6DCqEfqfpjjkSf8SKr3PpM
pwElEXXvSqjyw/cpzsnAz4g7jJCy4ERRH3L7yQDBJ078mLtm8TwNLz9dhkm7mnWruI7zdE5DXn8c
Y7Ww2SoDlNLfRs/Wh4QXn27Bq+4SgRWoXe6k6Rb7tkir0SF21pnoHiiSZo62UkuWCAy0gyr1eIiz
TAJq4XM3pEg8QM+dQzQUC63ZUAeQ99mspmIZgJqeKjq3KtXc69Adp1QnEaWIRCnALdP4Gl/e/BaP
cx0eL+6+6KLlz3viej/z80QGnfiRLqjsqx58Q9w6tyLB2853VYqUuxYh8/mQ3YKeFXQ9abSmqXIO
ztuYYgLAVXnfZ3106v03k38PuEO+QdJJFgS1bHjahAIYKjbD9Dqf0Kf+kexjADqYJK2ofYdDoTRF
VWunMKscWnX64ivr8pTIjR3HU21Jugt5MU3XKt0WzYbVAtS3eKNtwxNh0KP+rixOXlu3ixoUceXu
pi4nD73F8xlQF/yXAw0ABs4ToFQSXhJ0QASMeKhiwR+2AZ6tUyTK8etymiEAiQib6cUHkTI0HjKC
7ui+G98gClW8wrtCdte5PcDX5QFfB3htRSHHwbNj57JOOgJePoLi6v9S/3kSrfdDDL8w/CRxE5vs
miunc1UCgH6i37U/YRax13JBpixA7sPxODTANQQkoCqgf5nXn014hOCmBW37ByvXN5UNa2P8rKnZ
ErODmpq0R78WgLJXOLEHg0HwkigsOi1Blkf6B6B1+/tyH1wB/P9dwX7C6yHLyWQ69kAf83vyOBEg
O9+QwlL3Lzw2UND1x8t4nrhvg4xUR7S8hNPWsoT/EMA3IPkx4sycs1ZQrEGbzbowmd41ZaFghqVT
/i/sVY4thGrJldQhrVN5epq5ID3OnT30qpaNsExOIkri+fOaMBtAjwJrElQJRSTGQMSzqpeZMdgX
SSDR3g/z0KZ59ueZFhq+7y8JlnOH6rGv2KFni5KWR7Ei+Qdw8sJkY781Yn1WyRQO2YV8JcloI877
bfuRIm8xrb61atjpWbfNl84FTLmP051rBUCpMK/nxjrSJFWrCg58mJqDybCA8UzU2hM7JKNGD0aS
qBsRzRdVI5V/dTeLhVyYBnt5c8pG6bpabAXxnYbbl28Up9kTj+z6VFE2TRV7nh7sMolRlStYwmrc
BAkHWE/kPeLKk4cIzj7TaTXs6ALllTmDEVxq9pBYQTzfv5BCi9JJ3VIYhkJjlKO/g9TVM0BJm3Sn
afOIpEueILJgOZk2xy3CPtL0i5FbuQXUEtCsGwbXMF9fYmWVxPWE/1cCrf/jF+n6LdQjmU61ZRmF
nJvCORDGcvhdL+W2KD+RqAP6KWF+rclJEQbmhkPQwV2jAGYcpUIjbn4qYgZsNdn9vxFlo2rfghEi
JBwcysVd9ondJVDazqBzPZYdh14UyA7UI3ZXwO+4q2hH2aO9hZ5iG3qdvB+Pj4KgWosIlxqS7Zp+
kWXvBR4oz+mGI/XKGHVvug/44m/DltzhotDv7MZwyPXDdibop+7cfpggh2y0UUXkAgnfuA9iYyPq
8V/fSyGeOOrLbBWHqjkBMAcH6EqAfQc1P7rKzrhZQHWSh/rGKwHFVMW9e7N8lAFW8CrncizrvVJO
2EDFUM/DZypAF6mLrkgM/KhDggwqRWdcgOrfWnenubyuxILwFdMNoszJTBfqS5vcQzFpXA6fYXib
R+sGkgQlcwpUzzUfgLNbV9PmXjs/7IVTG9n0cJgGSwpgIAX4JZU6pBmcXrwJb6Q+sT8F0OOg4ESS
QRqu9ti/scGzL52PdTCh5HzZuno8hGg1QUzqNV7CuJ4XmKq6pxOXKxOHpT19kVgVAjGuE4i9wBGI
hBu/OgsjzQiAFS7rtid8upTnX0Dt+RHJXdOQmrHTtar+eY3eo5YUJY4z9WCn+GgTO4cC/htXx9Xl
Fpml6twp5RLXj1VtcjIdp7HB2DoG3SLli7TGciI8Rbz/iSolpp0pIHNMNOGultcfcXbuPijnXtDo
SSqnFyhlloiivMOMkNowIV9O7Rhot2HhC4JoESu8r9HSR4tqQ28ZchvSb11+fHA3LvwteCDhfl6j
QJ6NbjrC3Sa/qPqhtprhMON55laJV/jOWUl1ANgOnelhanDSsXa5aKrxAuaQkEc0386qBshL2aE5
v9rg5hR7paeqZQr/pXEZxGiDQ6LRyZscunSv+j7SK/BP/pekSWeWntTqUVn7ABrV/hFogQc3YqDj
YffkwqB49gbh8NEqFZjevSBLt4pYSgD5KPgwW26ZFN+O2fNdsqeFbop1+4u4BAAViMmCxZvRRux5
pxRPISo8Q7ljgApppz4iVBYM9Si+kLZgv751w3vYPp1a8tCytpE1jQ7b5L4/Qodc479UzkUNzKVD
ytpgCjYuEstLUJrS22ZsXobuFbo//c4LdvUT2k2JMAJwPzu4AWG6FT3wl7Rk4Gq+a7KczO0GsZJL
FWoXr2J/7JvzOcx32uO0O2w3RK3rLzMx87PamfezZE5njm149aVVyl7/mXWXc9nv4VVovCGevoed
5DnzzBxHzHqrEvlIrQ+Yf45wfjJUCPC+Mm6Es1foiZDTdJOrJs9rGX3rOXMe47rec6ZyORHNNO9d
or/X1Cl7xoT+tpCl06azI7dujMpo8vRygoy49XX6AIL8mdqDNqiFAVs/3jASu6FJBARiDHJfpO+B
okvaPgja3bCWKPQ8gmE9RjWkevO8KA1uEY6u+dFXfQywKQewWnyEipGZ8XEJjvo2uge2NyfhkQk9
poMikGs/fKhFSt7Ic9QK6BQqo2n1AouUoDDWRObkCmj9WcyGwFzAY67fGYm0i9paV6rDCWoYWs9w
Hw248Yu1Tzx4tdH8nB3wy3KUpyCLlu7M4ADNT3P7uy05HanfW+BcCmsCw7OYDIFy8+JznriVM5b3
Zpjt15VjIun9zb7kVXhJe1joeYysswRFU3Hhnh1wYO0PjUirZ070O2ClRSVnyUZK4Mk3sUdLCbO1
iKAMOEWJ6kdIyzCo1aoW39HttqJ39t2Fdag+Ed3niLq+juUDygQRBn0l/YYQETSuSy/eiOMuUJVT
nu1QB3ZNAQMA4ei287NzI9HQ6BrI+1We0KKQBelYhUpgud3fW2CpqrnhvR4bKSjVPxzZ7PbGdy2L
7+G9QTm7byM07JAFz+kbl4ySQmGoOONLxXDrkCl3iRVyRb3SeksuKNbT/LRybdth761xkp/8mPfJ
tM/rszishyXvYC6zAEmnCq4MuNqC5bU/9nhxxHd/nBnnMsST5bXPAqlh6uyFLDANcFOUMhNg9IK5
blg+vVLQu9NOv1JhsH3m+7p99A4wAe/9DOfrVgo+0ykXIBbe7vxcFsch6vlLM18RICITgjSbpIv4
2VrmFHwqg2bueYfC3/QfmRiGxsiTcJXb8sZeIKr3hgOyYrcuYCfPnpEqv1pdbpZw2WvG7n4Sbq4k
LsY8vgJ4UWCXqSHC9rDJHNQqJkv9CTOfj/gbxF54BaMRQChJpho5jbpME0wm6lOgO8CM3b0tvlUE
m6+inhnE+ApOBsasDXR10NKHRzIA0c6ScFtWu9Q+qwAqQzQFRMx3Ii4a4/pL/rF6YxEmkmqN3oJx
bvm/mYixNCHLjtL1VKLdli0wCsa0gdK6EX8b37oLiGG1ECiy/CJblPDXHgXeUMRNbTY4s0xERm1A
sii3nQigpSTalYBFCOyPRkCVS9nPb+RtjekBJyfpAELeirnDjW9uRHGwJLKFKZYHzsQOLuuVsjrY
5Ye5dB+vMI35tDdAQihECSosKTpWBijsqBEsgCsh+t7hasL3UucbIvrvdkF+EP5vZR8AfH5DPG30
1r2DyCPXWmL/ER7wkbi8KtR5jdpc24NaxPiAiB6S4o/1cPmDoCEbjKdYYDOwuns4BN6p7GnRW5Tf
9MwGzIZ38Ct2R2k3JMTPp067veEdiW+3GHLwJN635mP41zrfVJvVx0x7gibmb/UM0ZlmWA6PdzBM
FdOSBJHokp5wniiB4uJlgwcnoU+LO6Ko3qaBJMTUwIoCQHJVQ+eArm8cCAALWU4BfWrq3o+mSY8L
9vjhgaLMGWfS6uvpKuIX6ybXsQpB4k9tlHV0YXDJMxVXkgseDMHqJgb7i891+M4FXx40yXKJQQ62
s6Gs1yMXnKeW2pqUMaYXQN+AyDQ0VrMSogUP0PhEkhj5EXQwUWuNZvsX5Vf7oJGuwaO7CNkDpLNH
63AsGsgjVO0dWvcwK2Ihn9GiLO+a6tVK1OXFZ37B9JmZbzQH38Cd7EPTAZGbvFnQx+08Eyft2yrN
QDp7CsNLEEea9GQlEej+9COlQJHZmkYarSQ+buCXtT0YEM/a/XkEJlaGxvg0f7y7/NH/3sTh7d6P
sUahfJ7BMyPoyAbn8+4SROFkh8z+rnLV5LVrNKt35F3KrN95CbQfgfAGe7qsehPvVqQva30rKJvF
eWxeTuuEXn0/kj1f1rpIdF6g4e5f+KjgcIDiJ4XUH7+7jiWvqLm6cv6BwozvkYnouWKbpB+G7Mtb
/WyzuO2m4RKzju7MtzT/ieIVdhI1AmECxxm5s75omjlW6KEzAZUBl3WB1NeH6eWr1VL4wkz+AEF2
Nb8d6GqPULEz7A0uCUebq2PK/gU2JET3We6feF3TR7DhQ+nIyu8lR5QWQP6s4hv/fwmWGiAFpZkU
ZlnxDNNeoEMr00hSO9qHikHZ66vjMZI6/eD3zPREr3xbH9X1g5fiUDljftP8zdQCbtkIQiqdBtcK
xDb4F1ZXmvw/xSVZh4x2LW+J+Re9Ii7mQ3P5OwOb5XQa+YBH13aDzWQhkWqJvZLEtMLvcDGHTxQs
TPh7Q4d1YehSwAPsNZ/eDrG24Wg/CK14My5CCWsdNkbawpi79pgkl+WoRk0Ij9AOjMfX7cP6S8P4
dELXDGvcW6xVdh5bpQ8ZXQGI5a0qGJ7v1nLIyeHRGhStvEI4myFV7EN0+QhryYSS+so+G64gzv7y
fehMGZkSLyx/Tb2nwM+hBTDp1NMaTTygKBRhGlWylSjVr+FCoCxgSN0L89LKIfoeoMydSWhQ4FFP
Dpo7WLR6sSf6D1a6j9gnDzkKA/9vhQB6c/hE7eH2Y9rxphxdMSITm7p83dJhp+NAxLe0nrCQ+XMM
Z37wgQqysqjroTK+beNSLMUhMJkJSbO6M+wgQkybsP9newP3U68Nk62o28igLl2i3XrxUp71aFV0
+FOPFax8kBeWyKBYTDIS8eruQw0aXcLsoTtzICjEz+dXTe5xXWEbMVjO/W5IJV0lzQYQ7YAPo+kT
MBDnCRfjwWE4gL2fh2Q7o8khyXVvE8uHUxm073xErkfniB06tNn14YkJE/2f8JIIbhEFO0ByBFOu
3iVELaUbl4vhIvLSVFmLQRk1ua4YpSZA3snqcxdDe4jlVhFNScOYko0WrpDTQDMNtjdU6oWNHk/0
crKw61pn6x+Bi9eSS/JUx8+fR/Plq/oS+eCI3SNeoC4IXz/dhm1gbYp3c9Lh7A4pAL3uGdgR45P1
9iP7sCbxyN9jzc/+rNOSbP2gEvQDK78VUDyQYU2yWyl0P+PaEItWTGGpMihqZsZbAOetKP2vkfaS
nATbtejXmDjTE8BRw9YheuxcXFGwElKH3v/IFeJ5fx40sw1HxSRJCNa2sQRAADkTPs74fbrmtX8Q
Jc50VR83slfaG2Q70nVW9UwYNVWho/oX+DYCA5i6hdqwxvbreRhrpNm9fulz9hvaiLAaaC9VtqOw
aJpi8usjzbGYsxze7OBuKofM+BXKlwzhU0GYYa0EjxgrL9ySGj2nDcUNwDWQ2F8gHcxRKlgegake
XnaGLlF0OnOjsijtjdlKwMXDO+yf0BYeRPmWn0uDYi0R69GSnP2bB3IZvYY0fQ+zI/p2Kla4k/sO
sDYlxLuMT8En45mxoGWebHIBjfIEdlaLN7ICWYtQ6cIPNBWMB8FdDt6jBz8Ro520465s92m0rUfK
x6HI6mCFPgD9MoxGk9whM9nAZEjjjJ/ZNA92cXP7fg+/GHqbQimQKgQP+ReAj8UpWIrMKkXhEcG6
qVICO5QULGKwNPcmOBh8qWLU5c2ZQWiXA2LLVRf1sFiAyNAe2nJ2lOZwgl00rog4+y4VfnrQAhXu
EEs0yLakjWCkYlf6wC+6TL2Axj4gCriczPC6exeZNS7caZdgx2kQQMTXAcb2RFwI665k3wqSFlnP
4JL3bF1++XJ9GUi32M67FiGdEJlh/a6AChlFQcuvaMe5ik71p7LNUuF9MWVKtlQbmr57CgNCoRzu
KHHx1RmpBb4q6VR/9DEyKCc+rYpeCIo5RJJ3RkT2UeukvsFaWQVol7zkT2tfzLp4H6XeqgSTTNcU
J0wj8jTIFTDtJ7hHKJYnFMIRZyXb87F/AlZeGYvnPXOlygImtt2DmJZZrLS0urK29aA8ahZ1T0r3
0dg+fpCtxdKSrem4gz7kD6ujZ3ovzp0ON6WZLjcUY9J0W4wtwjrPbivPzIGi8EoiYmkRzUssfzzO
7y/QfmXqSfilh6RT4wYfWNzXvZ2iL1JNu4xUftyNH/1slyVNqbQVt9ZQpuU+3tHgpZqJQJkRhXf5
qlhef8EqmCS2MakbZCb+9Zdl6LYhxGTHI7AVHnyZ69wMo9mp7uwm77cKRvB3P+flQfw9D/yfwR59
kbaX8Atrphp4D1A3jH+QlJjHQXgOZAEUH4wQn4YGCTB9qBcjbS1/WZpq7iX7cTlZG17ta/2B+0Ef
LvLnW5TMmHS9V8yz4A9PApK+e/hbjOXGFez1OJT5Q6ZMG6TdnBIRU+UFKUbDxd7jG0XIQS9tTMoT
9GZhUcm4al7LWPAzh4U/bUtOQWwHYlaJZeEvkEIk/KORHe0Hh6HS9IprbUVfxYnCjBIJUvnCcxBv
jKun3lB8NRZDt4jfrnkqiPIenFeCi7FTzUwWWEBgfBYx1KjkRs1JsF07S3+vY6Pd5cGpB9QXjpgb
dgM+I+pMf96o7OgLCF1hf4mOTcq/1NYuAz5NufCp9AMdUk582nGeIqeebRLgo19D7UwTUg+z6Xcn
yA4sz2GT3MkthzzKkefuOxAZ7l8bWoSeFHomulUirePd8N1IftPEw6eP4KknWmB6w63mrMOQKOfk
HBusRm1kl3GHQCb3GJq9CyBaW8GTSlTiUxLHVaxhL9PHhsjZymjhSydlXe+7Kov7lJ/Q5aZD8G0W
ON+5F1A37ZhlMRpvBCw5zGIpbWWxlDdg0tY9kq/FkBKtcj0Xk7DUgW1sv94Wow13ELNc0loSczKt
RJKQXXcykzQ6Ogq4yuS5xB12IknuHov8l7bbnyC5dwF3qGryo0rxsrX4OllGJo3w1Zjuo/WpGTUi
6qdrqIG8fcxmbQRgPTv8FV+PnmaXFhjNA+Fpksc8RE3vWwj0jm+MzX6ns4A8obuqdJQKPY1jeuFV
qcInst1U0iD56+swlwS05mxqjkk7Ica2SlWVexDDp1zzgb781AjNBU5mLAa39wHXX/SEzDw93r/A
71USwQ5HfFh4tFtp2PJpwQtxXfZ1j95VGbMICtepQCS0bS8S8kwIQr2VwRKGsXJY0qzgRlH0FIvb
mM3/QYI5jgJbte7KNCVfqSru2D1bQIkbBfDrywiYuTaN+H6YzHLvp//qVm1uYISOJblcXewRMFOc
z4QhnnXrkm2EIMiCfmTcT5GN0GJG4p1TKO/fL9t4BJDELqOGT4S6KgpiRwJrzqVvsOJAwZtfD7vQ
6HqMt7lrjCUMsZ6TngbnsNPsj5/92afsCeIDK1ivwJa1Z1iFW/VaDwrGgBRpsQ5N9UKR3oa8N1Mh
e6heztmwraC/PzJl3FlRJTcQACUIOsIJknjyTVXcVtmwLVB/CWs/WNZ3Gu05uwLUmppvoGr+vtXU
3JguLunqyesdSQ2Tl1ZRi9zJysUhp7Pcs7bVA02ujOHiz7kNqQdme18YhMIEkj2j67h6TD7cSc36
ZgY3YiJnd6LNOGNvwqm+WKQf9CX0o4PKx7iYgKZfh2SD7cQKZhYI3EeDUBr/HtgdwwFcKoPQEo0i
Uqa6+pvkAhOXlIdXVkwTuBjxNUzqF5OZJ3GQzw3K6vZZkjciogN/tR5BBnyJFPDzUKh9oazqKfgl
swtjLU5hbffrnuq0DEyNbmbgY34R10PQB7wqmBg2l4LVSlLVwqoRXDE6wL7RF/vXBPCH5Dkaw+K2
YPIO0EANEemgwpUpYQRv6oqO8gDIuE1K9FDEqE7CXaWYdviYvp3Ob+9ZYpsYB+QaQkYGqc1uGjaB
/kEdQAi1awR8IU3PeBJ+qtrwJKHuPawL7E+Jx8XSv+ezHK7ibEXnTJieYjwS8tZQ36O5eYLxZsJ9
zaVH49ZiIWXNCiqxGxwwhppWuHlfU1pNSYqBQKJuIvLHtzwDaZC0InyhiMd6ot7q4HaqTo+sKZSz
mqhV6nCMQV+GaCxVfvKL7DgEBgcsSmWwKx6EPNpNugcfq83/LtVfF6IWhCPJkJlGtyxH5/U5DhUF
9X+MBAZOR/I5VUi6AOdMePi361SVfFmpkx/d+YN+VMy7n7aNv8LKu+Jg0bJwKnH+0w+5I3y1ekoi
c2ZRshgIU6Bn+O6JiS0k44rpSmM+WczIkmFTH8YhYzF1UcgohQRFzzmQuT4B9EfAFMfr902UA2C1
xAEl+ker4+brHeOr07wpBISUH1Zip4AwMoIf5O9fiaVQM5/8Kz4r871xDBCTa595DC9IX0O1LHVc
5sWoqKaIt/qY7xNPX+/E8zxUlXbCXdUPib0oYcJvkHKR0sdxeudwrqgxsLR5OTqRxqHOM2Ck2Ukd
j7Bo7a1obUvQunNp4Qy1wZYd/+FhnvsZjj4BN2PV4+2CuD/yg02P0G/c/aDbIm4JDi8jJHn8vHGm
LhwSjWksr7kIbePJAV6aCWWbr1kyF7D7XC2jVop9K6HOZ1bVv7D3EM6o0FGEObw3NVdomqEN+Zfx
gz9C3JLVkhWQfUTvX5bzfYudFsdJRtz+XpcsarThkVMJ+Ju0jv0QATTeCrxAmPRlrZYsFeAkEyYe
VS9i+aIaRr83QZTOH4wRpW6mxM6RxUZwtaCQjmisOOTIWfyXL5E1AgiuKv8fKoWmkKqRZ5ZUZjbl
Kbz+RRPO4zM7LAS1tcTeVqNaPP3+kAlNo4WLcGymVkuZeMeE1kGjo8BsjnpBvU7q2Mc+SZz/lRQo
8Eqt62ML6G6tzNkjayhnYV1igeiwde9Hv/YKKXo++LOghr9bwdJDVHpQATq5eu/rQgWZf+x0aaP2
Tr2WdjwLEHbtOvIRSU/OuP1jC+Z1dYKrQLOVc1I7HKXsE8YLMV8O7geL/CrhWeDouQWYRemtSRF9
bjjLdtjRVq61+U/anvUK3fCb6GBpSjNEXP/6l7frxJUE8UuAZGqmS96tQeoiU/oEub9WJw6NZhNL
3B2+tdSVBHdRmUA4eDxla3oRE93oGhRYHukLDP+oFVLsMPl/FPaa70ZCD1sb+04UGd6ae92Gjyhj
un5fCq5SF3AQlVTp7I/0Qo+JiX9OwQLdx1Q98tpL9G9Ttv22jzVIWLhj5/2HiH0MMT393kN2huxC
8JlCaivdSKoxPRZuhxUn1gQ111+I3eRLUcPyqnwVt9egTzi/F+upyv8EWgGYS4vrhhgwQe547xDi
KL4IumK+LT0r45V9dDJ/QiM15UPovpKc54O4ZdrnoEWnBBt+gGYzgHMDVoL3FaKEovhQm75JOmPg
uj5MU56o5PvZCp9LfCuePLeUPxJQa+wIqK8sp9KB36FTUI+Rr1sfD339lz21Ye1EpoGbTd+NtlFL
CMNks9iHm51fnAH9+7jJ7DMWpmQMWJWBdUCVPkhILLjIVxaeoNzIwnv+F4mqGC1dLy77FOBbYM+Z
X4nQauN9IeiK9nivrays2FF+pd8NSNPzNQUDvBGqGZ4KJRieCd4zjSLMWqNNELcekQdB5wBk2apk
KcDFhwmbjFS5zeL9f/nUZgP2T+/GcXwibrAoKzweUuTLCQOe8/T3g0V+9N9Nngt5qpZUqfByKKwE
7IQFlTn8Qhx1UBIY8y1nq4PD2cNZ6yEQ1UE4HL/DHxhm2RLQMHMnXyHw+eWDf+Ou1DpTr7eS6idN
riBPSCX39g2ncbvL38SVNgsEiry1tkFdCbEXHrgVZG6DTbtvjZ2hZDho10zoDaEqIvpiKmSgwuxN
Ur3Kh6eR2W0I+CaRSnj34WES6t4WV8irW1O54ngTsDE0bow1OiHmXjGsf/bNamar2xeZxfykBJ89
vnBGmPBLBGLjks1LjB04NLJVUslE3iW2Wb9ji8II7aKM17LAZAJmshfgZryP2pIN+BX5qQD0bdmK
YvMN9BrLTdMZLbYa+HvW0IhLKR23dM+zyF/QO30hdMtDth9hTXEABYr4GAFS153cMTntd1tMFNHM
3oj+DauCTW5YbHc/PGtDZA72S0jjXs62upe9VutSpBXyeBxEf1lOXSoKzuhzw7fl/8HJ327UKmtR
HH3vLS7kJryTahrKWq3ZJNzK9hlCJNlDBio5jBdcWUNKFqhJ7Xt1wpyB2IQtMZl9kmBqwVGQLEqf
mogwtSOrTaDYgBW7X+rxkgx5hGtxHdXvMd8vb+j91YkpCAQP1V4GyoYcSjRjWqQ788jeM9IIW2dR
ntfPrmQ8/8zYMxD77P+QdADrngPMJuIDS6nVAKlQRxL+GHCswN08ufpab8m/lt4IJNnC2owgH69E
uQ2Jf1Ntnh+HLaXkeSeE7Bd99uZjaI7QHR7AGQC7VUWmxGljkWYdgGPxAT2I/EerrlfG9L2FZCGl
bf8f5EA2eIoAbV6XvUx2Pjpj5NzmObJz5yXyNbLNRulpApeb4AnwUxDMCB6YBgGIqBNnoJkgKFdC
ceFM8EY65VL3MeYt/bZQfDEd8bN7Az1tho5zJhk6Nxrlm5SeyQlFR8RFZPBmwyCPI8l+63vi1s6V
m8RoMLl90N5D1SOgpalXIqf7ok8U3De0EM+tLYzbax/8hKJnP9qpk2jS9QkzRGuDB2bxnNn2F7KV
/B2zz1MS0elxpT7kmlogQY4+9/RXD1wUGTR6T11CqL/Z3Cwy8wqXTbEBp2Ifq62Qs7Mpr7ss62FX
LGLhkyfPaqnwmsoPdtkqihMDpau1bVzfWIjfTOa7T7DxueOC/i/NJjW8gcOet/JH36r8vafKjjvI
/PpBQn/X+LMXZ3mgJlMpkprer4Zx5S+9AHgcnTg12TymevJhFNAyrSEQzmN9ivD6h2qFcJ0+2SeS
ebtqgwaFz2o9qsX8GnLwsNqg4Y7p6OHI3pIgM76aA2BHydp17byEJYiNJZPw3bPLWrEsLerptyoC
T2YihHbxx108WQW+x99WhucdsCoznwB+q6XWQsh80cRP3zLSN2Dxoufnp3o3oZLG3NHEb2tlqTyV
tYhI5uCJwRt9G2I6d1CC6tThQK+PFpBK0MxoQI+ByZshtmltPoi+I+5h+Gh3Hg9i3nnmmxXWpTT4
hk2Iz74ryCEiZUf0lFmJrJjEOfDyk/FIlhkj6GbuUya8xvjkaJAWuPvo+xdNJ6EuhMYTzcaU47kt
76sPfX/QZVovBoJlOb/SqSItT/t1NswMC3a+RGbt/qmsvWvE3kWdu90K17cdxq69rNYoUvfeOeBp
OdoRTt4EXs5eIcq2K9Tv3ryEdexyJeyNsHpk08i1UTDlRoUyx6MN3wk0lR6PsjZoTHtOTjtMSkjj
aXTga5j0XlPh1l5Mq0zYo2Z9GCXF0q6c2hZNN/1ZtFOLYkWRCykrcMnV9VdfTsexz+gHoDk5LhiG
MnJYOT4zAjvwm2+/E6WqEavBrCQsJRSpNC7kahI73pDDieGKY2cWl3OKnrKEIRd+z65WbLOa3Q8e
8YR5zlPkygBbhnruh3VClxtok7NSaw/+DGjMbwx5l385+0XBuHj/pvEy1fTGCLVi1adi6DB114pA
8KcTFNMTu65W7aotnGfUzMEGobmFBGS55PKbxIdsBlA86uJp1iygqXZF5Q8OoyLi4V0xnN9//OFw
wDirXaljI154KzWFVs/i4hqiq0UR9XKQQ3ojOdERNXUXrZkea02aZGJbdIB+sywpSuZvu+/1pMVJ
LBZLBWk1PkXDEsEjlOKYbJXYoFKHdcFqVME2gm1zhZh2KkejC4B3peam6W96ZyHoD8Xb3SbfJ75X
AWb4qnpna9J1Q9fre/alglUENzmz4LNfxJtGGuCv4wlx6cOrLqfHcP/ro4bTrVtHwI6/YN4i+1W9
mSB216eoF4oFAlGk7KCykxHNjx0e2TkVxznQXzrHaI/W4RAgjr7+EgbBz/Un8iv3wZZVPzsUKvfN
gaa5lbXFq6ji+t6RfqXrVJLAmDaa0f5d5MJQSgrqHZYVr9zkVFCNuPMOnunNRkad/3qA2zkcC9uV
uZfMea2l177J9NTTa5ZsuRZt/Njd2xA8jjPIhDdyfkOOxBePGG/QE1NlLgPmfH0XPcX3XAmZpboJ
c4SQz9ni6DzqEUQ93vWF3sTQEkFLNy1zx3aNl3CCIH/sF34l3KkurBEBFBjm9iNVYpTDpu2sIj0K
raJQeKfcm7Nw1p9vPJ6P+gkK8lj98vhiTi2ZVFc1AGn8Je0Ri6OxKd56rmzR/5i686zebYVDmnh/
lIdABTeapgQI3L69AsMw74PxX1TRWbKWIgGR3eLwHk7Ulfnh2GBxNFdrNjHDHkW/I31Oe3KPXbcg
wcnXeeoO6i6ckwFMnrlJj0HnFCkDVo9Pr6zauc8YH+YxZMdMlc3dYCpJnLMrjVz+UFr+oiONMgxn
d/YW0iLGJbUMIriNLPd3NXOhQAsNGKuYhfpzKhSyJkx9FIsWprDunF1aRFbc8h3ERrPua2ZbNziU
c28VhJJjpa9PYZ2f7c72Wfdd6WxlO08hmLPbjnXbOnA3N0pk27gCfuvVruromyGuT4CHE7TNxrNN
AZskulSjyfjySH54sr3drqe5T4bwDlIQrwKvfQK/aD1x4eW1vn5A91BilFLDGd4R4gjftOYePiwx
Tcyqa/D1lTfjr7WzPzjGtFGKFuddEZNtA9Wz4pAF3mSGrHQLn1Z3pS+EmUOHDAczTYjQLEPqMMpQ
P/ILN0fY1sfEBswkI4jR40R9Is515zYpZpvemiOBoPe7Xm1YFcc/Plb6r7Kooz54/9MSmoSaC0gu
I+76nCtV9/g0LEBkGNGcQtlf4mTTOWb5t9FO/nGiTPGZQtRUrwF8T6Dpr+RWpP5xu/4mVC90NOkp
W/u47VuY3u/JZrhNtzQV5K94yVqaqRiT2+0Rj8j9oLvi2R18Hpk3agLyrxCRdovRXiM0scA3Js1U
oOIJiKJfyBpyTPDCxAlm36T49dhWv3A+zLXO3EmztWFnv/04E8e+WSPHVyLSBLqZ1oDGTQsuGw/k
1XJh7bFqasfebjKwjFPhrjQf4j5q+ZMGGAPFxQgkkllVREjU7UpYJMwZEtvaOa47Wesp9uAb9ZG5
8OrBsBWk5oGbGHXAgJJHtf6qPPdDrs/ryRf4xa3fl/r019VayCcK8DjMQn6yjKEy0fh1neih7J6q
meXAVRLxZaUlc5i5Xw2Yg5Hrca3ONkijm1CyVaeuVbYKY51ojIudnDnYzlpmtDgvh0hKiBaf0aUy
GfrKWb4VOKLYAHEIrpRKNKRxkzmGApDKZUguz2oQCtvZeAEomptLlJ4mgcjE1fWeuQg3Hr8k53IS
k0xrVrMD8JGA57Fh8ozA04DfJAIzdg+UWBgA3/u5YQ4obK1z8dXUTA8za1I13FhOaF9+inJaTQ/w
/93W2KUtUMOhr2y+eZC+Yox1ywiEg91XggkRP1T9gbaVEHVrvFuehf354/vl8qELTwgks2zIECkt
PZk40OGtF0WSKTBcDU5H1pk0UnlJvL1HnvW3w4lLp7okSPM3dwEPFNSrj0CZ6WPhivuBYqoDliuA
tdkNihQBoIF51DHo3UcjICOHyIxolDU6fRHT+BK3i5rUwMFBD40afOhEvd138bdZisIjtbR5YAYa
zV9R2dv4aynt79z6gb6VDNqOYPGKzOKt5MxfsIQeSZ7fVCLnlzVUi+Bh4O7ZVdODZhuANYwOUu5z
cKXVyyVYtEgCBzQonSVkg/Xbd5hKJI991bZ2qI7Qk9zTR4EOLa/t3ApTdtnNV78y/FGkqRupE5qE
DbZEvp67q51vR3wgFEdRAQ7XO1RqwWZsxoSVF0wUhIcI9lIpNEGLBrxL8lUM2S00wIZCzR2cebYs
lg5r5LUYoaPam7fyZCFjevMGaPR3934BIE+i+zpHoS/ziuNc1fPsAc9BJDvP2j1Y5Dcqtb4ANJpx
uxNn5zPsyXK0R5dRvLzpuTFtOq9MAs5ErvPj1CytBYKKASBHmSgkSxmb2OPDK/zR0rHP89GpILMF
FiLhAck+EpDbg68ssZBjR5GzSuCfhfKG7VbXQ/0cADXpp9qZPfJgWT9cXODY6PzE/xU+IpMDhqpJ
9yVQqalWuWKMHDGlk6/5tiiWLMh/RGU+yPEo458T12Cz55vhiECBFYXKpQecT0hdk8ZWPWwri2+d
xO09lxSw0cBo/ZvLSxdsjES07M1aL1koTNbxuyB58mlFj8dXKtAhNH6lHJwUBxlunpo7R/kds9uf
GUMr6rV+WCreiXVR0s5h1sw8F1YeMwr+glnG+1apuwkmjQ4Thzrq2OvQJ7lDjY+FqxPlDz2FzXYX
nOjhoR73cVvOF+wvxsBAYptd4KyCR3IL9oNf6VVI7lXkMrsjgnWTTCWzrV8lctNgrOodCcqPJUQw
iK3wuD6Cctk8JlTVEHDfxb463lVSDVKHW0M7kFu2dKJ5KcdCc/O1XqJ5ewK3zo9bUni8X+u8Lvlj
M0P7vG+44sn15HNiLfrGe9+fc1/B5AOolO4LOtYpALt6ALm3fygVaBhTxZkX/Ii4l4PnX4j+avB4
eDsAeml1DJLckNV0IE1kqk7FAyaBu6HWtsET++B3Mr2eTs8szDbboopvMcseanCxGJsA/u3GvVya
3416Fo3pGrK4H+GGvOGCL2nFa3NR5GneKWTfSYdbIpkIfiPI9eVuxwKZIArmtGNSeUQ3A9KiSFnP
Yu7u6bS0maSrQyShSLxJOnc+rX/4pM1oCdUvlY0CLS4leW83HZK7c9v7YXnFbC0yy57HoL8lH5+E
ECrLfhiDyWRNqRSM3zfYaLXg/TQNZIOuX2bskJ8G6onfiEJDXSyY9HIJ5oMvdXSdl3HEV3PfU4qg
3G0XHzYPUKvu6WpA4b51g6bwjyvC1Gsq5eWLqxXEX1n1RIdjN9y8OWAADdjzuxYisaVDMmfgXiDF
xmuHSszjHOmjHj15xxUDqIuKF10garCKSxBAPolYOI2dJmPaBS8KpY0Mw9gXMJnhS3fNdJRVk0y2
Fcq+HDMk5FsYBDg08/WfJmg7mQsl1DNHKAmsD5ngW6xwQ8zLvtoKU2Ya3m/kSeIJC1ltqg8o8oUo
bfiQdmCzQwlWqjmoFoEk/8NZXqr61nN8bmyUA0DpteNsMGg1knC+Elty4DldkfXBfMRgLeN9WDTs
K0TWd+a418AuSTZ0pPLtKBhDmjbGVuR7NX0FPSLKuliUzPO5Fi3pqtUlhKJJdHaJ8HDuER/eMhvj
dn4+XbjxrNO4kPRcACxCDLiLKeBNEktRD/7v29WK43nXWDYcgb1aKDg+oNHTeYawr2AIeOGMslO0
f1+z3ujLqu2oCG4TcwFB9TKWZ66wzjRWd7+1Kp7i4k5aUhZ2TxfuGlyITOrk0zPoZsr+CUFqPIds
m1f88mTAeA8Cf/MqjTjMgoSSX/DT8Cyhzxzwa1UzROppj+u/qgJfNXtJYLXfwUakjaNH6EQJ6Pzg
iFa5wjaWRMYkFWBxBRIGO6cmS8Scx8vfhkvvoFjX2oFhjXP910qhuCm33mSZ+T6OrGcLzpIFonbE
GkeJIUtYXs8xi678dRM/trU4DZKaJrBX/e+90Unpy0tyjApdOSp0sjwdtg5kuptHPE4EtuAZYlq9
3I8SBTqBzU6jYT69dHWIjQXhdxU7DvTeYVehf9El5Q85aTu7Pic3uF30HW+O4MAE0YgD4mCJaJgq
PRzPZgyJzK/r4OWBVtwcgjipzJ65HFtTvaN7teEs0S2UdEy7vigQnC+rGHy5N2stHCcLI1d0+2rE
p7NSSHzs8a3VuqNI3KyW/CyAQFKGGoV3zYkHlFVj4WgcLgPDmG2mwYmo1I/Rv+lrLpNZhs1jue0W
89zV/0qqRwyf2NguGiTMpJXlkOnhZNxs31avKfdLhmxA4Rkr+pjY1Q5QP353REOhA58dPsjsVuTQ
k11DCrjPrceYsP9E3Pz6uhuH8X6echR/itGi93e/TXz6AHx7AULsIEV6OmambzPSrF8ltmyXk7e6
Q5YNSSUJo2JuGgM/VJ0W80wyAwULwD8aE4KMkzvYGSczd5i5BeSbaeton5ryxgRemfprfcaVW+NC
i53lb+3lXaMuzBBlnBflk2sVwubHb3Lg1nsv6XiIcWysOA54uhTROyO36kBNvtQu6X31hZlxYI3c
WrCC1uIIRSlB6hIGVS0WtIhXKxQB7Rkw8Zd7+Hg/tKs08Do3v576RfqFf7JZDn9zVq+ExwuqAZmv
Fr96lLMJIo06ahe3vMqpCLbsM8SOCWRLjuoWhUDl37gokJwTqDIMSuZVf2RFieXdduzOIRsH+4C0
q+SYG/NAi0N5NBPIbuIOnQWuqaFYgWF9k+Vkp1PSTCcLNpFtV/X7tHwAY8ygCPMekyBsH935Xrfv
RR3SySc44dCEuh+/PbvBTxQPe2IoqtGR4WPUsZ355FuOQwC53xtRmDc8wjFG6uOfBHlHP0LM/1O9
ZcMcSM0Tb1+UlECav/WzRfp5AvroIqT8zYcVadyETtAxv/ZMMvuC6rtEk2oK9VkXvssV4CS0EIjM
YuxokuT678EUwkAvPR501kkUxKKqvIW7JTkSzxrgexguJQd8uAT21pF1XNWeK6PjANWw7R9QbFZz
sLyQPclx0o0VRd+269J85oPYgYRpNUiOezJn4vbgfaX9mDfTUmR7Vq+mwPGOcr5QRxNazh6rgU+R
K6EfjRHa8nQyDvDQDg5EWjR4KDVAuEjNiTKUPKjDARpfwBhlQp69ea82FqKuLOQ8GPJnO/ExrNHo
fMHunPPkb9Ui/hhfpHZloWciE6Jomh2aqsZmkCM0wQr3B19leiB983iwGxf8hyeax2KvpnsZEDDX
MJeyZgqdEUvjSvcCkKhV8FDB6gcseOEHZOkQwL+387Qujc8ILdXV5nb53EEhVRBHn6uA2POcAYAt
ZtoTbN64W2IfOvbMXdEOwQsHqw4J6yEVJ0aOGsdbCdPL4hzlb8KYkOIrQVws8Ql5AabkYaWseohV
ATO9s4YT6VWc7aUSs8h0/KuKjXZHwnnVJtQ0rBM0Lh23a/dbffJNwu7l/MnB6c33Xmd4wM8r1bGZ
nqxRIqq2Ph8nk93SW5/PTYE+stXZiUZjKDGKL8TGpdC/WVWOcPNj10BHghuDX7iwDuMuOlE7v1aV
YQ4SoMvGr8kxN65W8iaq7KNffEYNGImmOkWsqUfrCrGbuYTcQ0JMWCeSMuJueMleNMFVJaGpk0io
QeU3p22iyzNC7dpsJSm909QZyTYJKg9jSGh+RcxvHmk14u+hGLNKDkMZvA29Ki98b6aiV490oTzJ
nhK3bs5Mhn/HE0wulXmGD0T32AS3HfZYRPZF2Q7ZRfP3S61mIJJZ4Pw+QlXeeQUmm+jYxYGiV8VB
7F/h01hVbj1aFKhGqEZR83xXhMNhuwjNJnt8bTHBb/YY0xIca+wye255yBShBi0HusFEUryszUxK
dLom7HUgCBm6Ch2ZjwGdHgc84b7sNS+1l6PaO+fcVRoQXiOjsVoJjWfbVtmsCDWkKREUGukdR8DZ
lGRxqJeolTDQ5YsTiM+bi3VeMZW9+ZJ9T8mIqc4LEhENS/ifERhMj5QDonh7/26RyapNdmJ/IFd0
84xoxXohJV6DSIalQkDWQd4BnhVEDMP1Na/mg3OTMWSxR1HbGMGOgG7lDv1khfJMSjsPlqfNHGw4
gjAJDFubOxlQL49BVydS2r0Td87N0DhGaU+zSrTg7psFUtgE694NNzG0CmBGBqETf7inZr3jg0pI
IhPV17ue1jtxbpt5v3BLpFN93/aRPnKb2f7h+02ufv0MrgKWNA0CO92GHc/papyg1AgVj9pV+8cL
eZY67rPPyfBF9PImI6UvepNE2HA/6nxvX5NvNJMIjRGk6QzhOq1+/Nl6ZETM3tXcQu7fidnlnSUr
HwtP8N7VDIgPxmENahGlxYU0yAlam12TgQgUzl5ygWBHFaLHdClyNX3wbBPd9jv3jqq9QKSopr/J
Zaz+bk2e4jhaVZlpi0SJQmUoociazVmP1uHhsPILJF4yK/1bdG4XRdwooAk70x/Pj9CFQDhipdwE
PnNZvvfiZACbG44Sti2mDu2qt0JvW2qI8cbYXW4TytohfRrk7Pr8XYJU0cIxkJ+15fNxT3CZbIGK
oRM9wXsDOZlXUCu1pdrVXl3OtANEimXT3PLN9SETbBmzXqcdNQ++ScVeYpMjtbHNwHeOypm5O3xu
FHg6b3eibR+G1KP3sLUWxBX58On1dXmJU+fLt9tZyF1LxVmpQjHmndVyypqNWbYnhtyeiJHcNk4A
wBaPzVcVPJQNTLYUQz4vOZ153XIr2Tvh0I77FpLKuGwNEgMVa0rUV1cbe4P475OLn2X4JGJZBKe1
Yvj1twwCSStQcofWN2xakL2TCrkIWbKFY2NzjZSCJd9ZG6+GaqWcXguYu9J7cOWykkh7SUm8spz5
/htb/oNifhlXsDFKR+qZrqF89ka61Hk5Fg07RC6b+y3+L3b0mmNWLCU1tGsnOlw/34pPQWRIxQJZ
JG+e+SjVKwJuO1s308W3uJqicZ8pu1pEpOZO4g4N6/QM8mZIe4kjbxi8hf4zIEjdL6D55UqOpJ6c
Eb/Sy894MrZxrJrIWc2K4QF2iSZZnxUOwBnYXgmEeF0YPzd2bzfKUsfj589ADPg0r0c7Hax9F2fZ
pvrbJKYv1iKBxQqHuf7ugfRLQ8f1pb6Mv/5Z+xFVWp38b6JdYgrInWWNrPOMHcB7yKxeDFaweDD0
TiNZ2HBY5wlHDr3GZA7CIepuZSuHwR1vyA72CRq2f//8D14YIHr6CG3mdwmgBb00S/3fkvA/lslf
X0DB1Arm8zwcud1qIMCCHFAuKx/PWDhDVEqkrA938SQA1ZQRohN3SFRk/MfPmX/PCTJVWOM/ii1+
LF3+JHFFzSZDLdUNH906vitv6nD03IZQW+ItflRcKbf1UBHjaCS8ic1y9NH7vAL4wbDD5nYt3ZQr
Em2bbSld+qHaHMmlnBCmI5aX4SvCt4fd3eIs+va1Bg6l7tBOTuy8izEdWE8h3E5XsJ7oblkhtoed
6xU/9dI1OB8lNEQGcnOwsdG2hGYQOD11+/WAHwpGL+28ETjPR9/+1dz8jIVA/J8DeFuzUbPWl+IQ
7pJ1OuUKE4FgsbVF1GHuYOs1t/xRZukphLfgbL/GA2kH1zc8WBk6VKaX/jVo/alqCu3B/uO9/qLn
DhSbkxEpG+UKoQ1O3cXn9v1R19K1U5i1dzF/a/aHiAAatXKrr7SqXLB3HitGH7Az0IZq/Ymkyj/B
PwxULVmBVEifX50UOkHZaqY89YYP5miVskpDi9ZMr8YEMvIwXM+wYpmCALSoeDOQ1x1tAHDjWbWg
GibOh3SRtMtL/896mV8aT5KoszsWqu16VjnkqwkB7yqEhqc0G6ubOZv8YZ5RXm6aDVwLzMcaLjF6
aF6VXZ4iZbO68Js/7pqiLRhTS5ZRpWQD0JuBsq7uQN0vp6CKBb94t9cLiJbVeve5B+LIyDuMsvY2
MkiNrlREvG/UgX0YPTKjIuYAUwRQu8mw4F+2YdzIuQG037LdiL2S7w7RA9aZlyw5bDgcLihu7abd
jQzVng7OvtZ8uyubRCN7GUS46Xc7JtITb44pN4yFG1roRkTHu0BMzm5ihQkZYayAIkoCRMW40aGD
zdn/nV8GYePZB8tqKEJREWkmRs+JfLFPYq2RrOk5/Ui5sg8YKPzygWdfYQNMSq5bDMiW0TIS8tZ+
tgNvWwdPSPTplQaedPHn3ZjB7pXY8ht2cKnN4RQhjqzNIj9RL/kPWSrcXfWx/R8oERUoA7rFRpwH
axESVJxJiE/Yu79v7FC1LJ1nyMJojnXTGF5M8F4TKoXEruLJpmytLOYSntFLIzwCGx++62vhzBWR
B8jV9mYOMPPLZZDe/lVTgCr6Zyfrtn6JUmunyacKkvRhpyzoWiormCYrvPKHkaK0ntzncgWVlEPk
WNdg822TwegJ1PtloVaNp+F/6LUctXICW0xjyH4J4t7S+XZXLxsU/2ZjnIgKH1Z/aJIdVk5/kk6H
x8ia4VP0m9sanweWTr+u2XlAkq25xOPVDDgFsaac314ZoXawpjtGd7rogeq+480cGzneB9YMgFvG
RsNzxhsrjpH27nTo0LllqPlZmgFRYCvr3kVV6yig0sxtf5IHFrHn3TshUmKGToqSwylKx7F3rkHz
1LU4IhqUMVEeI/noLgCutAB8Mk373b/7QR6VIrXmu+ej4mRGxEbVhmoOFZddER+x30vYvlNfvp0Z
YyqJJY2EVVlXCdqJ6MvYt0VKKZjyjG2D+4BV0enljAysdVY0tl2pAaJkm+/1RVyx1vE6jUE8jVDy
4QDukEGm/OWOGiCToPMlsy+C1f/IxhWRdaoBUAwA3rYfCrteOSib1o4d5WYAJv9OHq+6qTpaTBoa
gYO9XrfLeg8Mu/yVbYTbMFO4MErDC4QtT3P572Skhx/oKGFUOdcy5/FqG028oi4SIF5t1MvzJMH4
uQLIeQDStpi36OFtt6NIKvZJvaWTT4v+mlw0MsAITfnM4oOnoQuUjMHS6KHVwxrRKcBJjIg/uEux
pWvfcKYcodVFWZDnRaRYcC0hir6vORyi2ewL8v/XpclyeO/8AeqKEQdECtmHm9FLmBfQ8nWp9Xpq
xfOt0vH90ScX1UI47Qo7l8grFKh1fHvXd+DcAbwDuhJU2wRCfDJXbFExtABoRBF4irLA/1KY4YDC
vYLzwIbqYRhIMTsqtav0qNMT4b8HHIuFxp/wtsn1pT72J5uq5fVMCx8UE3D6u7Kz3SeQSfzR9O7c
tnm3M8KFshoIRh7sxN3q4BGn5aw5qaMvtHdN+ct3k0lagAV4c/pu6okr6CfCLhCpKyv7PIEhGbur
8t2pNmgNoH1Y9hT6YHZI5r5GIKhWgJPLOo6wCql0j0j+JN10uJpKBGyz9sPAclMP7Y8cwr/uZlz8
YVNAVL3Sbt+mCUHC+yHwzuCzRnUiTlu7OqqQ7qKyz3AwXe63x48JA36KvKQ/ewzWTX5TZBlR2Xqu
08HoCI5yMqwhbLD9DWkCNEm6TmaLqrd/FHs6NQK8JhDBiwVwnpRKgEBhBzAPn7wej70qMEP09ibb
UMX8JNF3Q6LQPzkr4qH9ND7SIvBEc5ispEP23b9FSYVxGZkFijU5ihigpUrGCi+zZuEslDsmbjJr
FNOU37mchnigqBFwo6IBbb6N+n1wNj5ZkVpezdfYWyYIM1G+DOzuSsHV5/aREHZ/qkXv8hdmj9Xi
1OdnOPP6oTAvnzwQC/8Q65+ahrYcQxErygxlrce6WYqPswfUYMqaxD+hZF+bLHAaOWHfQTRfVj/l
hvyJktbMV/bW5X09xeTJ5GUIThd73KRNn7l9YldK3v67Bh1MVrIGjtM7I/32fyf/LtVgp2VdF2BS
RVcrfypoqnMiWE8dYurkAvebGwIvpd+nleOgOr6ohgGAndyYq6TtEzftpoqS4UqjD7MA158602OU
p8uoP9HC5Qo03bL8Ifqq/O/UaJSlMYwvjLpO65Hp+Q+G6WxH+eIOIdsCBvExpo1e16tsSIaWq6WG
3SN14M4bjWYV+0wD0Mpi1QrlIRrPjCDXs5TjctvwuRWK/e8Fxf+RXEQ9IRhNcG+LJGTbvuPYNtCv
gygIbXnnmmedMXaQ+QbYvVNdeb7KB4vP1lkkCBY86aXhaF4EVHwEr/WkRZhocpxmF+zvsnmozfrH
9VSK1KQvkcvVlroqaV9HMu8+tDR2a7uPlZHeRxBhC1g7zIqS15HMTDY/ZfcAxKlTz8ElYj82Yz8J
PyryI/0T2DlcbzCtPXmzSrvyWAuzeRABih5bGatkUeE07r8BHKsciI1oU2HiQMbjBI9tpoxCKsLL
xLI4v2EwFYDtOoCOzXh+XAdnKvVFt67UXOn42Ph3qeL23/m/BcYCF28FQEy3MXNDZ4jg30oYhnwv
3jal7P/D6EHyLpAg/iDpAdpbwFMzfGcQV4p3t5ukxjBF/FXLgsD7ta/cu04mptaeU8jOoQJ0nXL2
icbmed/F5LN5HdKtMxb6lmChTV8pc1Muh3xSWvv53jqxY51hYOQl7VXSM96wLR+fPMzKztErIlLZ
fH/dfQ5wkO6zLyATT6TGHA2CUV67VX9vGo3S4SVyii7X9r6tEd/rS1Pm8LFkL6bJtnb/NJ/72xL4
fyf4xlCaBH97C2QMicjkWBNMrCoOi9kz5umzIDXy97vPy1QWgo5L/75tzBNR3hq6dfHgqdx4fytd
6jT6uNC6YKPxEZujIbTXukJUHaYkhsEifZRPiefhGYBByKLz4jaL0AlB+ftuW3d/mV1EqA6ckELc
WvGbmsv3czhBrJWGah/wicW5EHvMppmNNEcZK00zo2l8DWAfzBwEjYDwxrHHuuJ8DBCWJNUx+nN4
PLkhkE2D9BIbqr4bh60N3ssAYZzCdNz+Ffl41zSDffzyvOEdJjQpA/rurTFr3p/L3RNBDrbQS/Cr
1wSqGrSGsGzD48qwC7gbtQJR7w9gTJ41+sdr1J3K4Ijmq82hxq5trV/0h/8ym+cuATEsGPWK1zwh
Igds52/OmsrLi8YNFLumHYBxqZwusBKlQjRKZNAVGg8sKWjTkJfa3zjEXiX7DpD4ByOiTYA10FZz
6j81jUAJXumHziu7WREOWxFcxAJY2ziTZNAWnFuH6uyK2S+6+yEdDgZw1cBDkggcX8sOf/wmm9SG
cqy4kBvIefZon/tqvblqobiN2KKP4s4hZQnZSoxlSS0M4zdBKEFa7XgacH7FW7wXNvLzZYnXjpFG
ic+DV44I534HtTrNwNOz5ILdVX+wd6EJE/QvGfRC7NOf1RqVFSaI/J03z4M2+a3pDJtxqTX1DCdJ
bWea3nO447kcqXWAcGZ+c267372FpWYKE1so0gV9reuiUQF+ZMpROIIoOwnu9ZUrcap+Z4GrH1nh
eW22c75KvwkKBr30z9a5DTOQqRFBmUhsdrNJCsNVVRNbM+iEv2H0+WfEyHLjJ5UFVZL6PFNnkyfb
j7Oo+H4uwcUAX0EyWnqVl40kIkXeTL2kgbooz6gF+mhq5I3lDiAhPqgRTXp5aeuC+vBLF3OkeBNZ
zulu2+xNCa4xm+tlP5+B6DPKw759W+UvL13VPKy/8PM6fiDYRudl/bApKku8mcMpCuqodL06KGvL
qAz8DviVsZw14ZXMZxBl4FD9yq5vTzEMUWPdrqbu9KFPZeDGkNz5dVwDWDjnsSM1O1S8nHoxvcbE
XO8T8gQT4a+G6OgVzbuHEfuhbABeWV1fFUvlSw/nA6VSORTfcMPiLRM31wvOqplJwLHSXUcLeELh
9fPnbXHmcnwHZWOXNTlaURLS/TtEQwiWA+ofZzeu3JVaP4ykrSa2u9gJXRh/VP2IQvWLlEI4NOTc
vqwVFOMIoK7xuVRcbjCKkQtlWMNvcOq79ac4xlGh+PqJdabQUwWn62aFRgDsTq5IRtYej29hd5Ez
DOsxAdTKtX0m3uQhcj63Owp+ZD9zhBvCtcQYA2VtO9hVcgMK5aThJkvRj3NiQvIbM+Hjv2ri/1Nd
LR6nGAK3Gs9lM8Tq1sSRxZyAP8t95OQyMGKqremE0+8xcaDb14T4cQdPHOHSxQHygylg0KMNvdOu
G74ZpBUUolurzeyokeT+onLrbIdnu7W4PPHlXXSkbJFYkPE91L6HLnMd2dyCVVhLtf+3/6ueXoCx
RZMPbGQ8zWGsQMnP/AZgwxTZfsx+OdfyJZtk+JegfnL/eS97gOtBOniynxHdEW3dN0l9LO9jOcfc
UABBFfAjiX6pf4Cfi9TEVyJuJBxPKzNgUyKH2ivXRBX8JvuvZgG2EZdZsgX8bBjNdmmRcS3pbkVY
RwZQS0XJ8lI76TZZic2cuJXJd4OljNg9YU5X7JsswFtfcotyLuPY9d0oQvDwOjZA7NkbiPbtatb2
Nczi/1Vhexh2w9rfZ0u4cbHuV8fZHNRspYUnQxU/v6mOe2ifYlx54sCAHIg1X7nlrydY+h5XA5cG
K9Wp/ItM+bbG3yLoKNPUZgd5+88m/scKKwTQ1dIA8YYK96GIFkFMU5QNQdxulOn5Nr6L8kXdh7TN
/jIvML/LKr2lcGkqjkfeYJkdZLpfEBOcRYTUBYNOUXOWHZ0Da/W+CIULqBRe3ihNczRSVxsWE03d
QOt3100CrBp4BtS2cu9Fs71Z26XOfcAR7/a84WDWX+Gl9abo79H2ToQVz7yF7WXHyoK+jZ3Idf9q
b5D/dtll8YAGs0fXtfYKDbnZt8sdRAxkHs4dy3FZIeeTOQ8LzWFOavISP8KAE7kKyRjtWqiqgLIi
Tqm95lA79nPXSV00XkRvp/GR0WR/r4ELcrPUCLZc4E8ghmSXPxH+pjMd7poqtv5Oa1CHtqq0YIyH
jklG4R8CGQtu0tsEYqW2p4dfZlqHkqumAi02sljKKUW3DpljhoRFJv5s+ox/ywMCxb+tjZbX1Cvc
WfimJyYcuWJFwMDkDGo87y459PR9XzO8FPlJ7qvliTDUTxTD96T1+PWhvCqPvHl6IEksYVYzrfvS
yuX7Qdimap2PWC9FLFviRErqB/9VlQQlkrO9SpM2bI747abDoVf5azUccEKunWw1HviFjTZ8TSrn
uI7rOtpnFKt586cp4DxlmluAp/GTH9tvLo48vL4E7ubEBtWS4njEF6Q4B7IxWK6Z4KkAWaqnvl2d
KsEtwj9u/DvYj3pdbkoTAPKklXvKti0PB2sFGgcnZs8tm0XmD3Huv8ijLjQK+7qz0k3Wa1BImkAC
IV4snryI2bLYSPEAAz4HSaqJhXcegCtdaq5Z0T28Wvrq/b++VMcHC+BOuiDMac1m6KVZolv1FeSs
EFK+GHTkw9lA5n/8GJWjvHlmQ4eT0Hf8deycJ0NzAMZsJCky5dGspfaGzKHyNhAAZ9C6WEhpLL4s
Ms+3OmZr0creCDUh4rQaOrv4Ffg5KfQp3DrXNEHRoeEuGYZeJ1sfNr2rX4C3lKQrZEDx8vRNAHoO
DSSz0VjaF/h2N3K//2S7Sdl+HP25wYUlJTOg0VBzAF8d1jgxpkL/qf06/5Ehd1tQa+huGhGe3Spf
+5u0pHpMiLhaXbHMyZ9UaQ8I7tpAUwCt1QCJKfoYkaOB84AM8xyaTrkuzInR/Ph0K9Abj35iH9Lf
z6jS7NcQWFj9qF8p9Qaf5q6V77T/s+nWGKOHgQVobJJGWKr1ZdBY+kAasHAgSxK8QPajQcghsFzO
BNmZpG9yKZgjmEM8iNqag3pz6NMuWQ45qC9YCz+5g18VzXcsZqK1E9Kt4VgUL8FoLDdw9Rv4KYHu
rOlDCFQpoRpGBaDLeO35WHVvt/nel5Y5BIKc0ePlaAIsk+s0Xwset2EN9RXX87O7a5EhnGvae+Oj
9DTWJQ6LiX+c/dEYj9JAsoJU7tEG6AvCdJoHH63ShURwn9KmuD9dFzSCSn0eCsPA3PAylutMtNXr
5aOxw6kUk5RYwZNjm0+iSsR5O3Xr539CXONhGYo4eA+e+sHKM9B27bYAzUF0QLS/QZB8nNJOfTbL
RhiKYK5b3gokOACYotJ8NT+/nzTeNfauAGlRiNKes4kkpQILHGrf/GoLd4x0J92sdVnCfVmoD8Uh
wSXPNpM3DsM4H/Q2DLLpEAB/dD4zrGZuBDN+geajdJZLPxe6VIvbmVvsH4Uh9SXgeBObj4wj9cEa
OARb/qW8tPFRtBZXsmlibgcEZzxtbIXGswOEbnZdvg9rq5PjaeRNW5MdkhSxLTShwIeJi6Yzf8Tp
RPDX9ThjszISBbVvc+YPznfUSpAiQoMTi5yphBumeuE+hbamf3UCKf/rgz+I4RBchGm6fqyaUv2c
SiHACehAJylgJquy6ArYx7wkxqYlHq4PsJAvFqNe6KJej3+yNUrUu/aywUANDW/8jyL5xJJff4l0
4BHVYL1udz8rhoOTLmlsaVOOBwbwvsAxmD7NtTidKZtT67rYqsfiXBa+AvM5d8zH7VogOyhIYoyS
xvs87ZPGyMZdVnSzl29RANpH2vQcY+F1jDOxIw/KtMQV4fHJk4x8wRzxCB5F4aKLPQwvvut/tTyb
fDOCUP+/VhQSidBfr1HEXXtE58xQ6jds5uXmuSplCOsadpp3MttelkRqLha+oPNCo5FCi8qL9dK3
UBkuvGohIimUhsvxCCYRGv+MzkXJjGBfFIq08U4sU3ei3KuIZgwxvap/QsRxtPNGor0V1HUq1xX2
nLh8ObPrLM4rPaNJUJ/qseydeDmjLm6bCCc83oYLRWuC0KDAjyJzTenOEe2uF5fNxWwd/MnePpmM
lgsjs3Kbhv6q9LsYxI9ENO42yeUKiDZC1v0XcF20vmZwiJ6uE82HNBpfODgn6s9Z9vYMLcXo5+S2
NQ+CtpW307IRPU51KdrkNkRJ9JbO+LloPqcaWElMDNCNOOSwzSwBsTYYh0uv71lm4wkeN3BMq/Ip
A7bodTyk4sBtN3GX91feWqH5TdjYALOz4db8LjDTsZWJWWv6u/ItugNau1QCfxvmjZTCYa4KVZfs
OSNYou47ZdEXSlY5MH/WqqXtqYzcVSJTTCLf/M6TEFotw8lgRDhKXc9KgruZVmYifaf/m2HeZWA7
BDHyPAQb5cfuLKM47oiQ3/A48fCi5d+Xxas38celWIoO100m4sjCbpwjB2CZ//vc5ZcUdjRmLq4g
osTURM9tzsNVZbsTS1jxZ5veD/jbzbCb8m5fPSSY9as9D6paOQCViyFu8zhnbCvKKFstGUc5Vkwj
JTmWJpkz1ouEWK36c1XF5IAYloQFe7XTxtHjS4VThPHPuVCn0VO71qCtruSiolguXVI1kdEFR36M
lxB/uSrli7+s+9mXf+Rfsw3fOsTx88yjbLck/cSKhJ7pyftU3ue3GnHbfQ8DCNUATDZXVIEdafoi
hkNqfObHQ4eXHLKCiFjjQy7VE6MTxHAbl4q/NuF7eKsW/CnZh+02e/NJh1fBuYqlz7SWFXzSi+3K
+o6inS5OLF6RJdrB79mV4nkOcIACY4204Lpbt5kVIQCMK22tvfsR/ysaiJ/rWYCVZ6OVOgkHxJbq
nFC4K6T+W0U3AjVdyfgZuzP5svNnJgz0MCf1AH6q1aMeGDsOrJsZBfbq/b+XNNJJ560houB60bOF
5+JmJ3+Q0VoXaS5JXwobaDYIYqd/Rnb7VR2DH4m0z74tueMLz04QONQOsCYQe6EVjQ1IslAMX0Zs
nuKSLcaix97IYvbGYBZda4jgG+kjBpjnmgp7tVSRufPMOOyPmGmdxG4hVgKuO1xalMu+BwyeEFoW
d9TNKK7G1elCQartV/CfY1D8MREn0Za43syMUtBEBMPgmJo68fsN6/vXADnk499stZT1c9lsllw0
9CPc+8HQRk7OG466JLteqshc72dcwa+6vQUsLYykiiuooSIoaFTE7wjop7bS2SioJILrqwtFZSPS
2GZlsd5ffpN6WHNuwHK7JGjWMccD/0dlNL2DK4HqREKZwBuV1j43ubqmQfEgtMaczSmx1SvyBdc/
gmjmX6mixJ4IrdvDytwHy5pcap+huV1Lk9Cu60ycu29/1LkqWqWOPdiUDukt/8s1BB8XAkMOI46y
ULHROrfQ4pmD2R7PaXMRzn1wNw58ud4kGeEMn7J41KQkLHBU7xi5OUtFr+vWIIUQ1cgHLB5e2Pmc
i8p4i0osVFwT+gDzFk/N9yxmtJ4+fr1IjtN1HzeuamgwsQdWGjUpIRjK80WBaDCx/eyM05K17PlP
LopNy5xv/ts7nLehyuWyJLkDXaswoFaCa10/XXtQvDhEgCAzBdlBVYo/OaZ95NwpC5KqnPw00LGr
5Nqn5dQtmyj9M+yKFWGujm5Honhr++vF26sGxcP2intZi5tAIyA8otYYi5IuSMMxLAV/kDbCNwfj
r2/DHnGyUMFriIkGULHp56+NP9g29YZ42StiMMpHN/b7PdpIcKY0ZKoDvxipoh5eat5LJk8WcI0X
2fIposyoe5G+GPT4buQEJghV/uWXGwDI3uqrHrjs0VINsw89/3TtBNrFiBLCP31gGIeTcQNlDB4x
FRWsg468YacSUz69+dmZvX5bS6ioaHzREtEnBPrCCMis/qx63styWy+WYFdHGM2C0qvDrxfBAj2r
8R/lDJ9ZOZuiOR4pJQ/rPPadCc2bUMiKHkDLNK55IWFw7PpThIDnVYpqw4Wm4RfD12bG4TR+OLop
5S2eoCVLZfhQGvciJ6lbkDXhjGnMAU5T83RJoyIt9e7SbT370Vo/TMb0SOw7Fjv6zZsaZXP27gQV
m6Q5GcZpSXM0SWXuI7+fJlpK9uoyWgjnOx1dHBj7i2tNM4M9FvZqWKWFVvP5ln699laEdVmNDBpm
v6ydSkj9qWRVxoQzOep642LxCC/E1XhCA9KLNhKKEbDkVlbszi5RaKrnGfDDvcaB9q9BKXU+GTAI
yqVrLOC1EensYJskuhzQG5esi4P3DiATBHOz1obm7Yq2kKBHBWYn9t9VJ3tVbj2bm6u8p3NUU4HM
fOjlaCfr9672uSO4b3/H5RRw0VjhLJ79YvPEVKHP2P23QfS0VLPP/WTtzHStmwQL5emUFWx09PTN
AFh26HLnRqKou/Kx2B+IetPPoTEbGZXVEcC6CxJgcNbCDpIrTc9LLNKKqmtbb0yqro+qXmcHC2Ld
6Nqi4LRkIn5CBl1dr0K5mzH3BiZIs94r2TQNkmRka64W45pc/im+TaEMtrP9n3jfG0OFMisBf5Iu
+y3uPvQiSJi6Cbd+g54u1w6Kx5PvmLoGgx9ulhm96TXYJKMl1B6YQj/xGcT62Hh/NrxKiUCkl/j6
g72esImyYu2Txf5UdJW34tLC0gc+SdHSM5RsRBOaRCe5JC0bJK3cJCMxQ9TDWPid1KCjexLNoiQi
W0vUNsdWOkzPJjagrxibz43BkS/FByG8J1/198SbcJFvIFNuxPsggvzck978KJdhve3wrFdcn6kP
00Oa0JWVXvKsxQNU8BbuARXFz2Li2KDEdKiQY7ViwzNwwpI3wYgOGf7oV5nWURpOT6qu9TTq9gIY
2UwX0Z6wueuYXW7DylYDdaqNZYbEg4KA3Nbcwtecap9WH7Xss8NYpqe3ytEqgIYW6/upVuYSZlN/
IIa+EcWSXgP/LMYjmDak6vE9nDfJwKLthfOBQ3exVCeHlMbNsP9VqDTyGYpUNaoLZ2l0P+XCZHFd
vfff+j3QXZclKVivjtyDXhbwGYxkZDYNR8F5L/sGL0X4Yw7o/sfFrHa+sTahoiWJUtTWgpfLOL9u
5xZvNdDiI/YzBZWhaWtM3sL9VaQbvjhpkIc3DLUum/lGWjW5R3+MDi1qNXI3ap3vFLJjD13wBeV3
5b4Q3aEUR8iXTobqedm5Q5WPQa3ix/9cmlZp5DWZxPe3xSPyX0rgXugKx51ibgj3WRqUjpTH1HD9
O/oT4LNXPHQ0YN2/mHm6lFpenFlrtB6JUV0jsi/50SXaQt9OmM9ADR/HlI9f9j/tEVt57Of/ub42
Cka8Wr9OWH2Bs+rX1iz4H7KivHaMeRdb81eKzhQdvKxcvOqX2aUqkPI53BSBFvU10mFDshy6RswG
ytDUFm63Vj4s5Z89luMsh3cBffcXZk9cjgPWygT+PM5OPALzOkRAhvRX/ZPmNr6Y9soa/pRe7f7n
7iESMwTeS9Wo0kahPrkgMe6+A+tUuGlox6OYE1PGt0Cev74F74GugJbV1LN/FWf/kKJMpBhhROOT
HcTwqk6lw3tfEtxYNwtyVNFVi/BPZsGBSD2cFhNGOfD6f3Byhag/wwCxd8YsKaSo1ILb2AKMMUz/
HwswKbLavnbaqtgRrVzim2H/pEqSUvnGOnzH5Ci/vgV88wTjAmBzTCMrshpkPYi8fWEL5oLprksl
ebAmsAUjlRsIHlmG/FEoXkchL/kv1thPvcRhwNdIfDs1Fi2fX9zaFowsOph5wnKNMjJfZy5h/NmE
XpwgwE15L/GLHQUImpZzGETkmpZmSkr8VSyfuVRvRqfwqNJMskpp1myt/hvcFnVVS3P4kaQSRWxR
CMM8kuX1Rfhjec0LEqUd7hSW3jJfM56Z5rZEtGYW5E0IzJkfEc/a2aV2jFIxAccdI9liMVU3AdYd
Qh7N5QxBVAbWwOcWyFxFYKiMCpyO0pkaNVtbauh1mFqJtlIQKc1fGas3timyocII16JnZWH1FKk5
8HL1Q9MrFjF2fDkHkhLkiPXdaoxBivI5kwhVHAwyjMCQI335eRLhUd76AqxI3AfTb89WqHjXKxpn
emPprbx5L/dPaYHBmf22WH/PsDJIF7e6/x46I7kc8JbzSIvn/ytAu54wMRKERDqpnfX9KMZRfY4v
f1W9tjjgVI+zJFXDDPg2aCamDhe4+6OVEtVpNEKr158SIjjeYi0jWiMSf9Be/jM2vEXOI6T3CmNv
Eb3Q2aQ+QEPUYLYb7ST3mCXi9MLLzP8fEJLHkWb49USCr27u0kCKjrbzIQlF5ft0DzBRAu9EFc9C
/grMca8VnixlJdmV7UfhzRpJU9v7l2Bm3Ve48h8Qb0TP70ngS12zLlkXTLQFYi0YuJTXSIU9QR3x
o8eTw2Ho8LYaccQxb48GClp4oTNCXYZTOl4c8b7+PBDExHZMEUVN0mPjNNA5as8Js05r07NpCoSg
sfIJNKt2Dwd6JX14wZi3Wk5MkeiH8SjEiNzYCbOMyKBjihP2U3TBM9gH4g04h20MVppqdG0h0W0J
rUalgo00ddrKUR61BqQmnMbfukgy3zranqBgct7nYQy3ZJ+n3HoR3qPyKnGkEn/afFnwjDlgzqs9
sHCeFSh9kQgkbfcvaML7zxGiBeTd4q3IKa58xDafTs0v1EC9d/+Lwun4cBwporOZVb+ZFFMToKO9
LMxiki2NwpgsX4lb/Yv96cbumJx4kEnk7oi5KTWeMZ3iYZgt1iGWwzsBLBN+L5ZYRlhJfnUos7ZL
NQT6uhgPZSBkKu5uyYxnryAyj1Cs0FBHvz6gzsmwMzNV5nVaKUbww8SSKWFbwtpkBPAl/r6Pp2M1
HbU4BTzMev4yybQMc+tibP5mI4s/mqgi6qwJ/Sb9N8azxlWHzuWecP/WvUdpQ5tC5LisD3FmvPut
CC3vQ3xzIBdgpcSapuUT3OPc9eo0SWAO6RP+56XoEPWdFRiw+GovxPBByG/vq5gdHENxxuA4zmDL
t+CzvJT+kssG/eyWDmFiFHApOXxayJx4jOTnzuIRzW4n8GzA+fpGdA1eU8F2YuCi46BXvF8WhjmT
ZIF7lfRGMai2owuD25iaDtqChfxyo5A43Nx0cNWo7S8v6g9WeuvCFbEeLVSPMiLG2sF2LS+fG/YY
nzwbwI74OWSepdYWOnhwASQFxx8vcmlyGgZZ9V/Y5RpBrY1L9x+4spFP2Je9QQ5UqgLStdRZjzhf
oI1zzkV59GqAAh9R8AeA9Btyzye+uf6oNo7AEoYbs6lhtGOTosw3ZXUAk9cgdzT3eWlsGP6kaDJA
2g7RLQliOLDFRlIhI7P3ELD9xwV/HNflGZFtPd7KS2ObuwSWdLLNcO4mUXFXYxuvoZz0YZpBx+bH
c2TpyXxi15pmzyrMyGm55vIJFxGJNwu8Z7eUlNYx9kcIAjwt/pt1NEnxH2T9nbCDR6x3m/TOJVFE
N3aV6uSeo2BTTt8BIOg9vkVrLX739ZVusUt8XZXdZxS1fr0VOHpFpc/szR2uuYKAXGYJpdrL0mkL
v2zQuvUFp/CmTqGLbXyJuLGaVwTRJ+lMm1oUB1gca02N/d69jTO3/zas9hqqB+cOWjUbz4IP3W0J
zEvhxlDOvItvURBzUPDlbfc22ZqsYGykmZsISBZ/QfJ522Iv+SCfMrff7NdFGfqEPxjl1OElg4J4
rSoyjt+WPLwa3UeyvC6IbHyHSxgKLVoBY6/D6uD5LqMwC4UKe1/QuGVU/nd8DNRcZcnkazu26NpN
twiWvKgkXRPzxUjURBLOxE2Vec3GcI8j8iOBVcTOTwVha+eBeJvZTjhg++oYM3JAqZ9dRgjrXwuX
v6xE5u/Fwg3wsEaudc7HWKGXJtRQFUoSf/78rVRUbsNM5qoACzk1tzOB9vT0c6JuYFE2IXpkrnXD
dPbhZOrrWRyp77GtRq/ajULg8XdMgMCi3Ncil/jtHToyjplLk0RT1rqd5o+KPCryGvi2YI6EUgwv
RQX2WmoqhSW2Ru1QpqX6YiL3dMDpXwbLQZduaRvwfVALE/SLSmZfsDgsUDQCWjAazNDIJkk/Tp5W
TAHMKpHm3FJH7NX+zfpurvMuy5xdA7unE2EVxB9AUBCEf37JVsb37/6MMWLGlLpYjo6TlvgkTrQX
bztsAKLemkJ+5bhNG1t2rUl3duVk82I9/i6J68JK91p8QbEk3C3oFKfhdxwiIA5ApxdJz8jMNBA6
ojTPEPYnEKKTXp3PfWtIYGWHFpXYCCX0rzQbxuRf0I3PBaF6IZEVzz8sn3LDf5g/cvedLXFUNiFH
/RbzubayY5qRiBB0LzMnfYJOn7zy5SiX19YjFzOc5vpHO33MecF50q/ounc1HnV3dxRf3khSS7YW
Vp4We3SVtzQgYS9actfljuhzC87FdTrGOawJGjYO1kug2OyiJCGMTammLk04p3D2q/cbrcFUcWwN
2NUhc67NBJsldYUdL4Bd5SRQgn7Wmb492JLWGhI7CHrokoqNGX0pC+zlwj0yGCYOOFY11gua3zlN
fyKdfDYt8ro3qgN5GlcwjjZOannI3q6dp12R2ul7fiEiJ1nS8RnWDXn208b409iLhFPjY4mPhqFs
jlniHiG9JFyQMuJEIh0zTqKeKKudbhK8/Sd07HE7l8G2WJS/QL3h0gR0MFI285pKlqED6WV0ImZP
3rNJdV36DAINhlWq4LklkptaGDw209DQAcFSHHLxbH8O9bg9p6ow2MUPjw23yVoShwh/4sZVsWZg
I0j0nSvMftN8/zojOUXl5k9qLbr7VQ3tyLeMexqmuRJpm9fyxFLwTWvmIsz+tu9KrftDPe7UznTF
rJflmioZoDFoaDiKqZ8sShzPvMcQgNNWbBG1sm0aybzCwj/5udJx7Eezz7rgQCdODMo46EeXXNvC
6OdSTDRvL4KE53K3nVcvjAK7F76RQobodECKNZqbGH7EVEjTFvrplhB0qQKsiz5X0WFQkM2bEuk8
4mIPnebLeRXroTpw/fXqbEvYcYlSV1c1CP9L1iB3EsVTwpdm52gqiuwODD6d/7dsnUUowQDdP8sC
mjRAjMMcYk4MMDok2UuNsM9/2glYYnxHTdJ6wsbprN7pEY7ErxdY8kMvbye//heX4q2XP62yW/pD
bNXxQLeuUke/93EazOpYJ70R8CFC9kq7qR1wTWJuEIwCFpwpk8P48PQZRMcT9p5E77ASsa6bpJ9w
KhQE58iCYFuC8/th3UvLWpd1VmHYXFRM4PwDFcPFPvyy5DSJ4niyqMS4EeMQ4HOGxleuk6E1jKF+
HvgRAL8Ue5NbOQdDOQ0tYknj0ai9XcM+fXtlU4WhtO7Z/ijg0phMEOFCnQMylt05qRdP/GXUX5SH
WhQJBiewn9ed1bE2mZULyvzdar6mTKiyZWQyf49JUpu1g7ZEyPxCABuy6LYXGN0Am2ZOMFzRjjA2
Wm/kDBxSZmLuT+SCu9fOsmwULXgJXH4Ody5Y7WX9fgsqTl38vNn5r8vSQjj8vpPgO+r2DnVQxnlS
5hLd1PuGGLDbepA18YaBZmUc/QTj4iU0EP34tl1yuGwbW3OpusOfV6BDjYLQYuiLd90wSKXqYHyK
CqV3o9Ibfn32wNs0oUSSKWWOSvWIYkMPzwqzmlXjAONWHhVdedQHCNSsbMZbmyLaLxnt9lUvJK/D
SGdI+wd7VGBKXI0d1PPNXsz1lxLcjsDMjzWUcjS0786nXNoiUcKubzOLFRT5AOoTK9n8vzSNuGNV
r9oOBncaN2IQemgXjvMZlodl/p2yChbn/5J6rh2BipWY73Yz+yzFmC/uHAkbU4YU+edUT2bW+bBT
7dHeqiN3eEqnMYCIdUfdF81jJEWammpA68nywth2QOn3Ga+hahQ9++vw0l8jWNsMROsZdKkAwo7Z
00L0TY0Ff+5L1HIo/lT5mrbINSolgsx0WnodaKHgr9PgpHip8A86N9M25k6mmeLldlL76KxsrGdJ
HDVmTuCHoOGRYHgvsvfGi+HBMmaEsTcQgfxicmTVll7bK4LTm9XaAUNcatQQrW1roV/eC790QuUd
o/redu11TIKCMRaBFITEv+l5gNLYkzaOz0W0qU5YCOYW7ZaXAvN7HLfsQGA7ZWfJJLbEnKwa7c0h
5KzZ1TB6i9lULNkdXvkcjpTrIcB3E201mklvVvBpePR+baGgXbo2dVutA3FuXwwJ4AHcCBMQmIwS
CouHQFUcmJDMvrml7JEih9IiyzdnLN0geX5eVr+nST2G8+pnMduC+XR/vjbSGAk5/jTY63d7djTp
P+/X1++NvyejYM2DSZkVR7ChW27rBgBXoWqLu4Dnd0HPigUrrQQj2SyZfEOFWe6/1ctM2QQlUMuM
755DoCgW+uUn5+D/U+7Hl4E2BkCIjkkfk0SKTIL+weAkONpsbAOaAxWKNMLLaS4nLjQUCQufaLIa
jsVRLTeL5gFMl/8tj3Gyhk10TSKV1UGBmzs1L5czuDbC2VbnezQOB+qUHYWJZ7sVKzcWa1NH3XXa
p+G73tYTCnypAIfzdCYTS/jwjum0GG1+lPUx1HBLw0TrGmBrNVlx4IHjif49vA+w2cnduTU+S2A0
Q8slKm5vv5LCCpB4Cf+36vr6L5tav+QQt3pog0Z+uWXqiF2LKx5ktxchTazhHuzjpNvXEWT2NF2L
kNs8wCMmgtlyyAMSNqiB/Vzhy/C9xVM9a/eP7ybsrUzhn6YR8d8vLYE4HlarR6m91w9L9YyVMh+z
d3wKEs8gqpA7LM8d0XoCpRP0w/8iyO6qYDOOnP7rMbasXrGgq5AF3L6cl5xp6dDJR0f8Xn6MV5VL
YkDrsKYe/yzJTZFA4xvPfFA/r5rsbMm/TxOHdg7dW5DQIL+R1Lz+G6f1OBjdSPFyoZnQQTTjBmOz
8mGJY0a7KIlngR0GXKmI/G0BQbgMeuVPDIPvkCwMlkyTbptLLbwy9LXXukhsvop9hzOHDKsK6RO1
/EAhh9Lt+Y9rzBubQMwIHHdZfAtQ/T/oJEcsfcuflWJaQdnX+Q3scd3BZQM4QHp4uRgtra2eQ3JH
/sxL+i+CV0hLOe968b03VZgQbEc+0gdooTEKtFwtA84Mq6z7DBjeL3/hmNvFAmccekcviVQZs3+2
due1MQdYr0KNn3iIO2htnY7B6XmsHkLORwLZKi72qdbe8+u0GN7+m8tN8jcpnVendJq9nr4cglKi
dY0KyW7SiukYBAeRdUR4CgeQPU5ZVlcNUUscUXKUMGroL1lnxIsSu47hGzE6d72rvtyHIzwteoa3
WyTwENbYScGfWU9IWyoQ/FmxK+IwOxQUyuKvBy5Ros0ZcnKNl/DG5gLu2YVnS2qHveDf5+/NL9uR
dOTDhB8Mkws5stQcZ6VQy430rNei1hZQuKiPlXom1jOsSLT3yW0sLc0qH1lSSR2/b78ZR1vNMjT0
kl0n9lovMEjOih991qWxSPST6hfDy7b2KT3nJ1Ep3hg1qiacoXyOhgoqLvAqsSwkiZJ6vAoXBm7z
kGBvGh24WNFbaKwz96MQnG3OB6R/WFKQir8WfZASKSw4FPmSDLpXhVKX6mFicVRaGbgzE3J8ygcN
/RTXSUDOgC38iIlJInp13d5A/mnMsDTkW21Dnj1Rwvkc0T0VJ6f8jqKtCo9nxCVC30tJQPdJtGC/
jNPO9DKTW7KCQXmDyHwamcnpjzh//asEEGDpdfxfrko5g4LxiYPIBaINKd93oslw1teE5HckuDLG
jagKWHnHNX18lkYDBXds6R3tYFyqVxu5pLJ1GiT4WH6RJp6QHLPCaHwhMAeVPWyJU843RPeTITE1
oBDbU96li6mOw2tQyuHaeDSRsF7v3OkAjEY0Jy+cIBqN30eDYEnvXoOKfuhW6rbaXbB6F3m5Ua1k
rV3rhnBsAdO2KufWQxE2m0aer04T9ejBp0Fej+V+W6z3UqOjNEwMwk+tWhyWAnfxTzCttY6IjvlQ
AFz5SIPdwkrw4hPKqhmk9ymOZMrQHfxJeHU7IvSvATVL9cS4XEfrBGIe/nG7OpkSlitkE/OYMwpj
YVt6zJwwR7A+ETmiFLYISVUh0cCA+7F0h0AF32ymlXtWCFUQoVqDcXV//wj351dQOV3m/zZvbilJ
x+JNAo97k9cYmd7ngElG5Y1ZpVAkU7ssf1kGPUEWHQfCdqzg3LORihPgDJW7DRbg2+A9PzZI/845
ikjlFhUoSAsXQJ4wXK/yZWf96TrzvQxTezeVBbK3WXc0j8/ATSSSVSRvVqhOjH0tPtDY6YZaDs+e
crKN7wzMf7kLfc/RJa/Evkx5vW6jArEnahOQryp1LxSLYL47BGSCtM1lSt7vH4ze6CbEbeeOelvX
rf6R51tj1EeIMB4uSj4lcnaj3KS2UH03O7+SaxHHx7jQTMhcGsQSyiBVQCM6zvBsyHGeuyV6oiHc
UVYNJuCa3dP5XhHbSYfFG6fUws9CyQbtwa6hAnuv5OGMNudRto+jdeZ5G2AItQqu/CwI0Kgy3Hlr
/CcxO8Mj00ZyqLDx+qJa8zeAzTPPGie0MQGRvMWFAY33Y7bCys6xS8RI05MeqR+fn9ddUBT7Jcbo
JVIUHET+53wPCrcJug4T2V8tv0q+4TGYT5wVWLBJHndkbWhL6+7ST75rg4hHOOjldaCodshb+wCa
IE5+2Pt4mOUzsm9GTqQaUIy21QJxeNNQeLYnDWMjyq+cWtrwYAYn2+/w39ersWbVYJt1qgCliixy
NVuDId4/6YUEO8t41gSee5qotPeDKhDS3gQLuHQMHHmekMXmof374v9hkQWtY04z5bh168EWYGqM
QrdMBkHgWnAL9EPOjR793ppS83ajDsbchLx8QXPL0UbuP0Wl4hKH/lXxddrJlo1WqCww/HWfKSwK
zfGLvb84z1AOuLv94zBGaWHeQKzrG25sM5xO3ONtDJoJjDwWPaygJEdVIcCdVomnyidCZInivXD+
xrX1Zg+QJES1/wjukPIZmbovQVQWeIY8w+hDFLcaoYtHR5LDOzAfxFUz3APsy3xwda1lXu/j4p1w
+WvETVPAnmHrAOUij4iiY5pnccFIStRCpuJdn1bQ6AuBVsgdq0gaSk7H0KKZj1oIYL89bkayUbcO
KnP0TQzaTWwJ+1lN0+0/WqiFUFFKXL+l2hW01svjzjV8aQG/WaTUfLl0ojPM+NqL97Y2lKIIyoXh
eZEnNiMxDBUYgwkNQLG5ccr10Kp/xThPuBWbXf4abBnIrNEGj7zh3iUXouTA5szEs/9VVcvyHzW6
Bczc8pwpLQqHzEicB9K9QHc9QJYZ8qaTRxx3fdbl1Qo6jNAIxbp69gfIQJvsNjZyawT0Bpbi4TdW
CQVvfx2bBhuoI4DM/k+jrzetTqXPE7vVEza2h61OcwM3h+C5U+MUuHDmmrYwpXODEh3NcDWn0Bvx
e4pAoocaqQnVH50MfpxIzGjHe401II8B+Jfhpi99KH7Kpr7o0LyqmYfviCyxsyNncicyq3u4aIdt
e7srx3nVDjygehvQ5I6YpF63xLIer5cPT66bpqygD3uGyKngyoAPwVSULTJ7srmT4ret+YAj01Iz
Kv6KabqLjR3hpy8lo3XAVniGL1QQ5qQvPEu/kl2M9DOUYILltZeUUnpKsitMRLb4f6ih4nUzkPBG
K5wfdL+Gkj6xzSc2mMOt+8LRP8pSlFede4Arg8zNtgU+6QPGTxcHeWnUb3ySoddgyQPtMB2E5gE2
hfb4gsSIVb+54ZzygX5IHbuOOgPAS9IAn7MlP7goDAKF8XDqzWbc6RMt+I3sDBx2hgu2aM47WDtK
9mMQnLlkFe+d3a+1t48ZjEvsqk9QqrPud8wWqq5fJ2l6oxJyBNsXqMRSuSt/A0j+yKmGOJ5lEvDN
TqxPuOs4fe7ucdZSKCqu5i753P+i0VS0dbC8lbSQ+u+u+BfIBftLz3IRYpLdDxpfRNBOxqpXky/t
mxKLLjATPxOKvqZ7UWr6IwGoD+SLugz5HoIP3pSNyr4MX7iQ9fufj2pP3FH441RwtC1vWQobz+Hj
MvkBpDUyeLEUJhILwyKZgkJopqxJtzw1lcWBBEBST6VkTCOlslCUlTq4Ttd3VejObHIrl+GCV+90
kWJGfwsi5D9xMOjv5TRQhxjhFhIXrSwUEQPAEGYDO7azhnkZTUqcpuNdvnsSbcZldNx/UheKcIhn
scMJMYUd524KxLhT5Nq6wvwtruXui1hUWQBDHN7Y/k0w1RQrS+l22PY7wjB5w5iLms5OO2DICFSa
9y4+rIL/9gYqVB1ngWyJom4TIWMET8hmMLLd98oPerC2Bj8vXWZRm/LUZXrYVyU0BLkTySicXIyc
Ce9olY3FynZ3F5TLLmRM/MHzke6hUda5/IFKNhOnfXXe4/54HyULzhOPv1HeffJDIc+k5uR/RpCa
ADp83IFLZxPHqFYR2+ja11ZR5ptEIw6cdFVd0qoK6yW0fO8L7xZY1nNfCDcrKOy+B3OiGPhvVpTm
KtBJA22mE6MyvoMUlnNBoj9skPtphTmQvF4g/FVw+lv9bq0+cjjEjE63Q3Euf6hjluwaYEFuYiDk
WiRrQF8C8aqN7yhB/STALcgQr33VwHtKAy9lliYi1o8jqtfBVi9Chh5gm3SBj4uo3h04eZciAkfp
a/Rq7ECD53XO1wmgQlxd+scVI3U4gR4QTHSgo1Ok5KaqXCXdUZIPTuDK6mF+8i/YHnMelftL0UUI
h1EhJRl0YUaQixAZZgYkxOPWztsrwarPucSQe0BCMmo93/BOwONi6Z/mvIW3fOPwzsWx5/v6XtqZ
+g4wTVjIlXXENFJk1JEgwtnB1FnZJQauIdEd2PNADxM02P4lum90DEs4D+Tsj5aXbq+pHWxl+fHq
kSgnLTg1w2yHopAGCF2bjgSCRJM3jvdT6fCUjhAFvcgyhR50qEIGzcUEEct4OZGGV+9QNa2mWbDw
3q43TUGxPwKKWzZ5TyZ6mxgtrVmgh7C5snq6cKd5Pj2ETREQoC7Aax5R63gLrWotMprbyyNUuBNZ
KhtKcPEQHHfV34sTtmdVYByBrSirL81lceXZ5sxfDEVANbO7cUuxpTNO2jWOplMFRhwjsu5gBVV7
O2sk4Bsj7Yo8tiYTEo8c+sh1IV8ImihphgeWekhON6KkH+54VgCPG6LF5CXdlkbehuhxGB/YXVOV
aXUMY8QR2P1CwFCYOft0Gi7Wmp2qACXwShxdSzIKgfmrsPEBaPTCz+VjIeUCKBl18ExofWYPdkw7
pTV+WOduzzZCaw0UGiUskvyB+ld4NwJJmVYsJ3+Bkoi1m32Sevciow2HHl81uZ55FLmUK0prSBQe
rBxw8qV8QG1SKPLUiHoZjyB23vqp5MfqTSgQK65+yWWX1VnCuhP7g05DbigPwhx9MBQyBrsbhJSt
LbJ+JJCkI+dSsyfajbJ3ZWTD/+T+YJ2nkKEBg/9qe07nvk4tmyvhloKMLXcOGu5IkAqaT1jpUYd9
hVwbZzkjqNhmUYh3rLRO4gvVNM/9JfA1NYF4bOUSDLZTRCqVjQk2f1fa4yMRhb2JfbBFMhiE+aOr
T3xgMO971MFKHYyeFfR6vIWNsyZTNyXy6t9ba2z9W3iZOtLSSm4A4EgZj13PI4WA4y1qnfhV3adr
afGPYbKp8w3AJdrLle+fApIWcAS/gGhmQBD9EOHe0ZXsJqPs+M4QZ4O4xCkagSJ0gG1rlM8kVAfR
Piyz/uWV0BSPadk807cLBBnSGM8ysrPZ/MbIjsvEXzUW/HrIQs5UCuLbAnys9noKZeyzdzKxTGqv
ZbDb4PvzT/H/OyL9jtV1Gkyp+AQsnRNpsO1sP+9EQxgYCNXsaJO4TMwAFQkZroI32teguFqhpaRb
9NMdSLodAsfQMVZa7DFtA2sbIgi91EpMc/WpU/YI33LZHPovLjaXv4h38izPnw0eRiqQPsAcYvuT
cbbdfFwSeUUYutrIbJs/KCnPAwWJgGgjMZiwNuh6wWjUcvKmnvOaird0Y7wR3916+ROdV6Rj8Cgd
+Jc3sbs5kRqbsSyhFuKs5DK+h02Tue4tnDGl9koEQroE8kTMRHR5IfSBdqfw+WsIOh/qq8G7epKL
ayKELdSiWLwTySkFeX1q3N1bBtMpZtfgHJxv6rjqI1S1Z2y/T2NCUcwNz8lSAPbhmwl1nSHmEe5z
5uMMOlu8c/IbekPXbYA4wzbO6G1uVUhyVkjTfCxLNv+tqH93RNyN0IEg2vEvEfmgpNAj21EZB0MS
91hSn8AcV+CZlKLDTb1b1o60F9lp1KLHo4T9EdTs6miOwUUxkNK541MoC+OxUMv+LbN93RWBvKNM
QPUV9idrbSzNu4IobLLfdzJz0DNEf3XL62j2R3jDMqHdKPza9OKmqo0i72fVK5hxXAqS6NTMQR+a
jHHT9ORnIrQqiNPsjiqZqOegGPyhLQ1r5+pwUq+VJquzBUTXe1l18H+zqAm2qf9ZXC/M2MuQle9K
832xUVTGaysh8UozExtxus5UKrmc74NKo9OiNJqfboA/PbvT8fh5t0M/JdG4OxUTs7+c00D4C3uP
Elc00i+Et7GO6J8Umh13NzbjjRqdvRwGbMovdx3gnhqjK8v55Nfzf/OQiaZWBHjoAP05OVrWdYPR
oLyzaAhLLDbbaSykgpcKP67ebH1AMCjpTB4yxqFksBzgkOvvfEk0TlCyF6RmPBIPesO4OFDXidy1
OJtTv9vg193VnFo43DhfCB2yISK+bWEkjgCuRjc27mvI7fvwm9em/NO0IdygiTfs8QJ6E1xQXD+C
0Zv2j+HGFgOlC4/ueBj1Zw97UGRHlN0LNzsTcoAxgs5OUzDIUt7/V/QU9Gc5ccTj7b2YawEr5l5y
R+bWg8dT4Epl7Snt6vlLld0mZQXUqTczoygQpfLQs71Kimwm6PDip/Esbc1i677wDFThu5D5MWuT
robS+DSCaNaDL1dzyQpCc5R5lqzGc3QdYYixOPC+ja/y7rJ3IdGnmmmrhWVAB11nAgLlukyyZz1i
zGUjhzQd90Z+n1UGzA53SedJ7QXTCS5Fkmf5o4JUL4Z6qKRTkaDXlTrIHbGJcWkyjMYEB1l3aZmM
K5kArAhPBU7Gfz9stIySugSOJaNPdKIS/f7Za2sKUrr+0BoiQYSjeTG5ooIhYif0rs7vbrTdEXXG
EBS3o7TrD5Asv4flaAU87sN7W8lfL9neNhErPRJM0Mc0FGDaPJtMEUFTr+znBSp1LE0eSO72FT6q
at7QSfgIls1ogdfbItWO0VV70oWUFXM64erbdYBT61+LT34IUkykdrHVsVf+rxwYNED0aTq4p47o
OS8DHXm1DolOmmoGQVDT9nLhwJS4J+Tso4SHb95qoH9MnpgpAoA4WBeIy6xYCh3A+DGFz3lfzt3H
pzrEp82hzild1FZBNykx+skAGSnV1JP5XYMjH0y5UFoMit4yqQ0KFkKHlApEjukBjAEl6CDiM++f
PoZfhVkDdxz3ERFmQa69F2MkWFdzU+CSid7YVOd8C4UtYDOujsXMaTYs39v+uhbabqJCj2ZuMSAR
4b9WFSQ3tq5wN7Eb7J3nsUWnmH4QdS1VXRmy21T7ZVFXKZUWCvcT2BSTkauKkHxkTcHip3J53zow
a4ceOi/h26qrB5bl5KrmC5DrucM4n1hHLiAl5lI1HjKyWy6rlDJV8fYyPq8hAtY+2n6O7XKCNWg1
d7Lmjq8KICDJTeuMBhq9JeJ+jVWyRtjaZJsZ60yJebirgtobT/eF2DoZbt3yVM21JroK3/4zmrlN
/D2hlnDgPKx6+3V+yuNHAai/UUQwB+aymdHrZyWpmFCRa2GZuSNz+qm13c8YEZCwCp48ySEW/z3J
gi6ptMChv+1ODRv9vnJHMStFbjBdZKXu709DE59MGRGGLQuixMmmeo9o67a8uEcwoXuHZu09q+0U
Yt6X1Fm10nzOFqZjJ+rhLrR/Y/We2Q+FmkldxGKKXwfdBbxwahN6mq3CCHdx6BSv29pCFnDLk5uc
mgvAOTGfzJ939OmBrYN3GKPmuOkZBdfM3F1LKK+UGkwajQXNLLheqaVzbzcit2Npar+Ood3f2kDa
ej/pvt5AekzySRFmuGfBV17uHBxVxsFQKJ3E0sEQ25sE7EZXcNkqwotB4L9jpyRNZR3CMK9M2ibU
9rqk69RkjQ9hmKFUU1dyybM0S56BCNqtiwMbgTvNEvHgmcaQs/G8ThSqSVikR6nwtt489Zn3IgG1
1mOrct0V/6wKdIOoX+/CjHcpVan/kx2jSgaAXDZNX2zn8cfKQnWPzfaGGGP0Pwgo+JsRu9BSUzVz
3UollchTUM5T22AATCKopveSnSE6l2qRu9aCs/bg79qRwSV23waxYUDUzuLbangW0OlNgjh43ZtZ
ZdZeanMsHL5rXMYv7Cu+7fPEH5dso3fqTj2zYGUUBTq/S6xmeO7Z7X82tbsfgC8pNkn3vZECxCvA
MXUjTn49EUAp4PLvVR1NLyt5GGjTVcDRWRCEpvEMJq10gmBjx3LGgpc1E6ENX6kXKf343sVfumiE
hKOUa1kgEcwoz2cAbRTCpcqinmf37UcOsazkET/XkF3YHPNqQYXxRJPRJSU++5T+yN7x9jgj7oNv
qtQm0tnYilMmTm08hskICTbQ5WjZZGLCKsA9xfsxinK23W7UArXb5oqECpwr8kKwGHyPn+BSi4tA
MHqybVXZMDjFswsrgsACDoWC9HjGcJ7lFz21AEjZlEA963u7kSpNThKZSra9Ft7mYMaYro3CzGaX
xz57EUVJ/g3awmoiIC1IUztxvKu8WlkajZvGo52OBTilkrvK4nZFDxr4lBW5Ma4ut8dxJje5Xcep
zkKafT4c2D+p1o5TaShe3VY53BeWvSM7bAFS19WotWGKHFW+8QYc5TD0CC4mC6RudS8+OPWks3XM
zIXGhtV//U9OfgH8JKYSwBuTkhp1c0h0HPgpNK6OyLVFRcFkGE+exDC/s194Mw7NRFlEgX0v9Qlz
Bc6eijRyWfEETwJv8takEmLUqjnn+wT7YvQ2J3TcsS1QPit8fr3WTCUdbv452F41aM2cMgMdFrRg
CxBUYQBgtn0yVodXbLyRUXLBZfS8mqiXaUu04+9+PYkU2/l6hNC53Yj829du12wm8g94c0K9j9T2
S15UDXtUdzofwkN6GNJ2oCxrNHZRaHY73ysvJA8GUfTlB80o7iiitc7Uoq+A0vBj5fXNktvl51lB
654w37Tw8ugBRfYqDGSlH5dovkWtoTjVmtNQ4nvHvgjFZbGbOEdGMtkZt2TIfi/1dZpSRVPTAQRi
xzdewY0Pr4d296eWHHwbURXdoDu0LNd9Vh7F+nxvkdGb9BeMrnIs1Il8txooArK4mZa8gdVkYmEf
RXwwkj0t/15J2ibNX2Z/Kx19qeF/v9ubXEt0742xuWP+anpgPOI2l2A2oNiPXTQS0TYPem3YNSN2
hteGkW+UsbJq2nXrKz8MaTDceYnChbGGNU+2/JAqmbYQs9bOTyhyopfWCQ10vDEw2pGy8l6QWVK+
TsSYjXtUpHEYo6K9FneePsyPbH4sqKwFKNeN5PaHyiApz4ARRpeDAzYUUGtfWX8ISDQSw1aPf00S
RHhT66nJvPK3SA/7AkFuV358Fxrav2j62Q+F0swHikNwNQr39+s2eJ3Uj7vxaQgKF05onTFL+81v
9P3nGvuoDebYXqOtLcuZujdl/4Gnetjs+ciS3zpsHnfOgRERQ9vK6vWx/JNTDpqRCbmjtEmJdFDK
n9Gz4f1svHkwLPt+RP9eFhL6qPrJxgUaqpx9RHliPFcmFDkb8SRE4BR6DFKDsxEP2Bio8176xO6S
GCMJDTyzhhdtKbTMv4lcqUCtAKGemJSc2W6Buy1QGz9ooTlWYqjJbGxvHnHycsIHkSyQltMULx1a
k9RFRg4jSXiz93l+BD9eDvkkznnF75xAPHWlM49CRhRvuTzKbj3kMIrKh1adk/tEE74J0k5uUGqd
3FufjzL0hH81gdYWuUV07Avsz2gQudq2VUC97m2zPH/znLpaKOG2iMQ5jBCd517U43Fv32dw5Or/
etgW+xi4no70zNmj4QOMgwpQ4KYWmv0Vj344nhIdZjubdRI+sfvhH6vNHmNXGG6YtmqR0x3nBvc0
dFNDdzgnDrdl8y/M5l/+Br5DSs2YgVpNjiDrUJmhjXcicIK6TnlLgWE8JNgVcuGL0CNezVfYSpQ6
Vi6j3KS14DS64R2cLRYn1LFZIBLp6FA4Iepgb3Fj9pXa6io7pyQtV/iHbcZN4Q+CI7UBU/PruzO1
y9tODr+noOpJR2mZJM03V50u6OAEE9qOt++qk16v/Na0NOD++hCw0ottJHIb/0f9kHhNZw4CeVFc
10DU4euyl+FIDQ1MlhNi8ChCK9cpYrkWDguvzkOCQjSg2nQY/7fVPwyJ1InXA0uF1y9aTjfWsUIq
kHy2c77LBxiUt243N2vIfJI8HzKdOfRvATy/toOwDpb1Al5eQKhuqeRdcH9uXe4qwB9c+6VLQJNH
2KkDVGBUXXQrEa0lvGCEQkzPoHzIHa1iwu9cXG9eWJ6d9ke23r/6wu5uLKSff/nJLY/5m8dgQGcX
Du67b/bNJRpIkCx6k47ukI8AOoEWDMY33M7hkCoBfV0ITJP8nucdtL7J4BnUpdfn8FFxZD9mpn9k
O/A004V6oC38pcBx10V/2foJzC+9euDXxotekbYUM9IV+tPXda4Zv67CJ13kIBzDkwSPQXPIPkcy
ODhPGeHbT0IyA7LyenQUsKk8ofgIHMsO26oR3ocZU2VSThmWGCL1vtmRRAXgcJfuXT+axPMarIap
vmx0HRmVyBSYDwC4Xcuo/J19xVZ+Oek+sEkHZKjfY7mPTrQ0B4RKqZT7Bk0AT6VCfUJRH/ALJBcU
9t6pjF4dcJjnMhozINK7dVTfpTQv5gaWyOhCMEj+CPLigKsOiEnpJpXWZlmd92zqFtFl9bnpMdH/
p1GBgqU5OVJ2PbmAGMuDf+bo+5E2w55VmznjgfEPxiWAeJlKyT2m9LY/BKWZrNArNcnd7im6ez4h
sQoIc8yDwnwFqc5Wu8WfAnzW5jiXUvgpVuT++4Q1h0mT+uvkd5PD+q/IyIteCL8QkTtED7LuuuRq
7Rc9S1+eqFcYIXL0L0WMV4EhzYeU5UvMaR6Q7vfpFEpSs1fndq7WuAhkZJj79Xww2OvLjzDopURs
P6q/4WZ0YsZyBFkdm2IiwWtSSVsYLdHwJqUR0nnqb2xe0Bbzzp9D1d0RYdXlkVR8T8CihvWXy04e
akwDGCkeB22z/Za/Y1SoIRLyT59fbl7TotVdvW4OPKbixvULIvWC2gi/0+mcuaF5wvH51Ti8eEeL
A6OCylcF/k9n2RQxr1/jwQ1dI0K8k1FNLQmeyWnjZ+rAq6jVXi1cNzfJpFEZ4U6T+1juy+PettNd
9dZpZmzrkEWrvw9l4OwAnkcimonkkZEw/ms+18tzGZ4qCKFYfKecaQ6rNpb3xJ1l1waESoIeMfzv
+hEIrQuAFbk039P1KecTIQJD3GGbNXDNz96LX+3O4Ruz+DLAKb15O9gELzeTBAkGWEOh4WHIH2UO
Q2nJk3Xnbj1t1UlM03QhgK/9OAmiCHo9mP2n1aS9/oYk+nSJvvRMHrq6OMJy7gSoo0TXgmM4pN5j
yGO/mza7RoQ9tVKduEGYLegCbaAkuxdx6+P4GQfQFeZOzFzCQAGQcOI3dtWNTua1OiPrAwOESjwf
a6z1W5x/TpfZPV0aoTcK7ifiWrkvryx82raITbZQoWgC1BYk+awrinHlzFTPAjBwjPiQxNQMNGl9
NM7JZQMDJgeUj7Dd8X7yv/pmnf9XihVtaZa8fH1ggahJx0VKxThUT/pdhTjYAg/n7L4upCK7VGMo
iXQ+oj8SPec706UB+W0zIWfQlqZ/oXqsfnDE9qylIX+/lO8Onu1NYv0kafkISP6FJb40RvOuTL4z
2DpNoXfvQGPOxwuhNYoWlZm5G+r+xz/TXnnjj1Hg7BNe9bPeT8W70fvLmfesP4lxtTaOf6ym1jEX
lpDepLmB+LwuiywYng8c779BcVJQBUwS0BljKhhvjceKJmt+uI7F1ItAGP+fXiZeKffcup+I7oop
Iuh+/28jWquqAundZb/ia4ZZYelG/gO11Qor1VDvb8UZqM6IeCmkxfyeY61i13esV4xpv8AeCEhJ
CP6GUf2NSuH6lKo3hgyrN/a0dt8GUfp7ClwVOXLGeVcpbMpP/vOPx84qcWnBg4EbPRmT+LJmlhTs
+BLNu8EiOkeBFpRmn8zwArjWCdsDE+HTG7tfndy68egYSp/2FsljLcmxzG5YKX1VhTaYiw3CqCSt
B7yUYGrjxvB8nUtrUgqK4/8A776+EFjz2Q6sLcq3jw64S+yulL6m+/IiRKlk+KMCs5mXTx6N7nUj
NE3fUm34AApmN9nAkPW6PdcFEM8RNsixgDIvASSe+uL2pB6z5mr3TuDjCNuubwcrr6uH3nWRUn/0
/ieRBTIKbiMeVhY50lkNfVjs2fTLoce9s1RoqWNNycnhvHKn4JO3dh2bQCCCJSE9weFmnZzYdTDI
JblyomY5kccyFne/CgSot+PdbmtVdgjZtb4ftcTHLJpv7zQmPGqBIp3fGMQv5f7rwbjCj/g4GHTd
4f0+oPqReW2MNFzTC9y1so7t0rD63g5SFFayIHJHHNXy3Un3P06wIkYrsFK4jh0V8lpo0HcOHvCR
iqYDXAuuIgIpCCUdZmJ1pDNNbVfECeYhhiiIYdz9uFNoo+JXmdCNH0kp1dQOIsbwS5XehFo2zvLm
q7gkak54SmTew27KvTz1OW2mGyIdfHMeKVy0O/rmVlrhHoYTBebVgvhgtOmszBspIvCzhMc6Nzt5
GZS+tV/YZQRBKaf+NspekJ2nyuCXVU1dUk6HY9/uGBrgs7Pa9OwUzUOtufQmffDM++bqObV9AIei
ZeTTjGNRr2RSUFPY+KTMaLj7Qc2oU/rlQgJItqIf0yt2WbVm10yF1QZLMO3rr+t1heMK8U7hs15B
kI5bwpyoMvm3tGKC3nTfo4OeBg0ZcY0D/4emU/xjNRieFHir1htp5lbugQWPlSf2DKD1WTrkNKQE
gbZZ4PbB3+smKhDcJCCVSSGCllpww7PoWmnqPHH+t4rbRjH6Sfccm2h7eTfxqcL3xKB0Uob3cj6J
HLwZhzlLqJoDhjaTd6K8xn/td5ECslGcs2sibKqs2DEtF3AzTMmUPKzB3yDMGFyPe9KFdrd37tWd
Vfgh19l1RpghkN9NwBrsKpKPin8a4vAy8vNe3NL8zDOVfXQj6xaUVjOpB/t5PM0ApIWYuNUtMvcB
xcCPEOVJf8J7Tz6klmv0gRUsSdTEOcnRwN6MKk/OEYGzjit6lO/9PZbCWScsNLqe+j8qTe6SmYv5
TgZBFUeBEN0j4ujVyXz9emQPPHmSNsYojG41l9UceNLezZG5Kwa3YR6c5z7mfyLGFN0PgVnQG4Yf
uVafGO9M+rSp+2PXNNpBIKX2WpH4yhKnP7r9U5CFBYBD3AqZwLG+2irPtkOtDzUAP3H3+hJhM3xF
gQwkxl9++iX5rUGWPoeC0HlWqaSJx8HSENIIWuc1/9UEc7FfPwFKIOKFQHmNYp7fAOM919/AMsc5
J6rOXBSKBJJYbpX3HmTNlQe71+xKrGrU18/kSMBdvuniwa/hHNkqfiRZY3AWGxQ/XUc1TW5myiE4
6TH+OWy/60fHiB/47aORVSozhFetyvj7h2ETeLMTUMDBPLCX2WZqoSseFwXRub/P6yRHbInqdxfE
rse6Ex3YaMNUOaVR7SUTC8RUOePdo3TcfAgYJQgZrCL9ipIHGvSqHPfKLyq1ZL56w1TjPxM74zr7
zFtNAvoMtiUv0B75y16Ib6W8EUNYMbFi44JW9/xKRGChc/zITv+BaeTHmGMvDYk6YoD9LjJRhBmv
535U0m1yYYk87i0rMFiNe+KsMOe6zLzFTct8pSe7xjVjY2DnvoCka2OIam04GmxlMe69I/oFLB2N
GFuOpb1FaG1dm65yWvldasPSJUj8xnacrfdDXHYp2WRXJD/jaXeyrt3YR1p/HCBJHWPziNwiyfVD
JFBRvV6hc/KNOttWbhz3Fj5lNvCYRKI3K9Iwh7KSKAYWHo8HJZMpasDgLV2ystXUaNIui15caocS
/nAPns7O1qkMQaqm+JtE2jOkYDirqI226pYbouhBKZHojoQqDTNutYWaNYcBmF0jC+7qbwtiS6ZO
n1z0EEA1lC42lO+5/13/A9gZAppT5AAzWUFkgxiZvyVgJLeCBjgovF+3+GEuKdFS47xDDyZehJKI
P6uyQ5SPtEo8XybSEd40oMR6nj6rNxdkqXMai+YcarYGfEUz5cz6IDoM/oUi7K0gDeWcA95oshsr
BofOprVFYFYkrcRbigdbCafXTcb3w9FuoWPuW0GA3Ee/702dMF96seNeTrS2FzsGq7YLlkKFQ9Ak
9Nxv/L5ufH/ZHSQm3bi6V7jdOSodCWz4AxiOs0rb8McJzI6Ut41/d9S6GS1s3p91c4bjoT/iq6af
8yX4Q9kttbivQBLWsPgNu+NwlWJ5Y6j7pieXOdQDDMUEpJq1Ca5VW2UFuYN5mWus0zJr4xJ3WR8G
ELNZslkxc2o/+bMRtuvd2XaF35HjwAX0upaP/MpcmlPA8LPuqjQwnGN6EyMX+IJ7EatoNrXX6g62
EmFRd8WHsWgbb4k4dLgYh21ysnJLF9xOdw8D1UO8eI3827vFmiBWua8FpIQqQ6lslSrgdr9sQvOm
6ShGA+BodMDNSE2cFueoHkE8+x0OnCJrnPKXoqhnHN0gxUL8K+RbIcoYg23dDfUoR+qNq/x4RjaT
87bnvkua+pNaiE914BdtLVxMoMPIvFsmIKbeN7O6DKPHWDd4jJywKNl1hMBwa+k+wwGKfXkS8v2M
cmrQf8bAwSPjwKSkU29WSxa5bn0Mu6jGrB2a46wxZE8ViYEzCTCFZ1bYPJIPQpmhTbwcIW033T6a
ZY6lNTeLa2r9mZMHzu8fqnM55Q2OLca/pJnuPVqGLTA9sIUo2tLLXi/tl98wavSZJHJwEyXPvPXY
HxSFClrVacvc++tGi+/CnAp6xabHpTJHtI+Wv5Y8RLbIc7e6PxCvHztEsGX3UwCf0GqOKT1qY9dJ
gY0KVkON7XCS3Oi9lve9h5nUmp3RboBxfBQMCdKeXoEBu4qBh9/3luTtvGhJB1gMX69/hQaduBej
23VzZT7rW+YwPASbYvxdYEN3H812hxMn6gnM9SVp6IwMHsFVZLPAlJy0+VwgEXI7sMHnL1t67gDA
zmjBCjTYDP6Xpw34xJ+jxvEm6IG2acnWlHEobwVicDYtCTlKbyHxFEeLMA5+aUq0mVP6f1w+uL29
JWg1UdnripQ0MNQFJv670AlBCDDDDpjzvKlNk3P8t+AabJunaoCa+nP7FmSxpz5zZmdhuZ50NjnU
0fKjwqUblcZjyFTOPPWPSvrZ8HDjBTNp1oho9NGOZJZfxr6ndKqyxMkwvCmTNYj9eDLHNG/ituDQ
re57kb7ibpwhs+ZtO3vbTEGnFTVw3QWt4xpRpqfyRbkuQd8OW9jBhELsSgegynex8Im2f2s/yeR+
6gy9MXTb8jcLFIkYeCxdKXcVQBLIPlaRt25U2VUZZ9Y/QKRPv2NB+PWdu3yLtsYG46MdVF3CkymS
c/4h551/zhKtZUMOFQAsQNw2q6LTEUTubHJOA0G7FDn86bwf9Ml+rL15FwTKHSRqbq0ybLjnpK28
9sgNAEoE5AHP4K75fJUG/N/xTAO6hW2rtIX/tz3/1NkMgDbRhJ74mLuGZPrMcTOueg8nZ4jSdGj0
CVTxBqVRwX4ab3eWpd0+sbsG2kFhc8mNuqdRgQ+yvVQasYw34CQG3z8+QNzy+FmDlZE+5iH2n95B
B044iJWQV7BPOJ0XzwJZcPxcuXeGXNDF0gUPKkTzgrUnZf9p9FHU8EySB2EeOMGUzZk4u5J9qn1+
r9xIy8h8Wv3nUtQq10LV485eng52uNHwRbzDTTuMBeVXCBLunZ8Brcq7ixkV/JhMNb4X+Xpgh5I1
gft/Xf7G4MCvjLe9T3LmwweJucS1aHskXsNRHYhf53FOdNG7+eIyDRiCBFk7Bj+fXtAmqgSQzoB0
rqmOSeKoh/mr1BjJ2CeBzwFXmalHSeaNqUYYWCR/wZTEbhXy3nLpodZXv2JQzV9YlKNFFDHOZe77
QqAjw9h4jqO1I+btLkUQ6jPeITdNgDKteA6YvqX+LBJ9a0B6q1T8taZLy+dMuLwz9b31sWMZhv2n
pDNVuVdRPlm9vbO9Cg2VvrsJkWmIB8nUeiTF5q1k93A1S0oWnrNWINUuZm2dz5sx6+ozTft5ZnoL
XNaW5xR9vZ0RHHZGtenHtTv9IU1zyX75FY4OFiIAulnIl069PTX4D+9KZOv/kyeE4tUg/7QuG3QO
goa755zNLOWd7qJlKl6s2y8mcRpbFQehgPQgsupBKdzGaHhrWOX7Q09ldpS3U8XsY0RTA0bxKhR+
htdSGjnzVwkQzQRxyQucsphS87kexe9X4K3gIQgh5fiekjh+8tG6+3erFsYsH44UGcPgQtYiS8N0
KEl6Wdmup1LRCiemRJxN7uc5YrP3SdlDjLpaRxxP/J72ZwJEmdGAGJ6yoeGggDXZjkeGbbExDisV
csiunLooGEQHHp3EVekS+3a/Wtzw+FSR8n5q8v/jal+/A2d82yXJftocnb2/HYCfHhK3ET9kds6N
xIWipbmRqwHCFfYXKlNL49wIqgQhtaCA0H4V7XpLxSOFPC5YgvCw0e7hTAL0jGJ6N2HwcSViaAd4
Py3rYUOiE3LGT3C0qrDqGddsRtiTvbT/s98IA2Jbv1kbj9B+H8vVjuD/ukT7nILCfiozIEdBPW+P
xCFXeMFJ7pIObl/nwfxNAjwGIQDi08JjnbPHDzQi22e+NhkmtIcXdSOaL6ycXBWpv1HnYjptEESH
c00g34eJRRZ9fngFqj5AgIzku1JD6a/jVziHojzSU1othr3buGjCXMEfarOGYyAr7LQD0J9+MZha
Rx7i6EG0eU2vYxBTQ++ROttzJfMVeZtjZyCytlcj/xATWgq1YTluNnN1+vgdZVGPRvUH3WHf+EC2
3ZW1qmsHEZOgI8Jln18iDTFnG4rq2hukgoQbeViKhKLIETSJZvuufbTOeR+ITmKlwoquy72m0LG9
DhIkMn8xGchkSomrJpQ+9+184ib6Z58fcuOtTLDl2qEoe1nD9d0fclWlSUWVmK/JU3zjMA2LXFke
hJw5ZcZvx0rrLcIl2RwqN5ZhOvm10zSqcX7K0o6gyOEo9VuMJ81QJdt/rrPZA8KbStI0DLPFF9Qy
1GGbDBT5QW8j2jf5Px0nssa3Qcoxe348wiZy5zQaUzYW13OW51LzA9SgDCF3yifizgYMwtOQCNvM
P1qWvtL0OfENuYRhyZO3PwCtB/WdZD52NoI5FYFD965/LZf2WOk57JcekvBL+IawMrJM+Vlr4RhD
DMhZV4DgbvngHSwc1i1fxbaR/CTjXcyBvsdaiZPdQr3KHn2QaeEKsHnlNZqHDuibkdcid6Dtkhgg
xq0YVtamjBDa1nxvuEKtGxcOX02KRDdLQ2TGU5mzdglXpPavsFjIxvSxlZYv4FvvD6cLKtid3Mfq
fKRjhFw9oPW1ji1oVpiiZO3h8MNEW5oGBfujLEi5YhgvDBkjC8t9yxzzonSnKsE+WwHKf2J+yDr9
ud06rXnspFciRj7L0WuZgDd/hqctbrKMaUa5zJemci57cewIrO/Xk67MXaz+aZIQOb9fT+4lVrHA
M0F5IK2PFmoHjwpzj0pSuq4YNWdJrR2tFLqVAbzJDV4+0DcUgXjcLOmp5kgCu5dZWPO3h6uwuTqA
hUuk7oh+cct5TDZbUSmxclTKJQ4dDnTnheq2nrE0fYD3hf0Oioy995Sb0a5HzMjbECSMKtlTQu5E
UBprB0845rTF4Jz0+AlC2TUjFq6l5WxrtXGvacGXtuK8vfUgrFimMSqljJ+7cEe4eDGb9/hPwu4b
TE0efEAyihUqRH7l8TZEaRCjQir98jPo/vfFMlMhd2cJgD8LQu+SmI+DjuWVVNWIT8W76U8pvdkU
YylwzWseI/1rP2plwpiwGq9oEHEZiDzcV0z/XrWRlXOOXQAyzKDgB6U0bJB9DGNuR/TAR/7t25JW
aMtn/xZcrDlkOEGqnZDkblUAeuNZJ1GDMRhEy3X5KFIy3UuKvw84YJx4tiKi4HSubzv9YSc7hs/8
7OlPSntyWzRSYm+kXU5H9H4B1JwZwm3gL/xwMxOscz6JSvynnMZufBiakA21dkcZ/OGBfomOYomu
l8WsL40Vu0Ed4aZkAydhIu2TI4Y9rxyOaZyJswA0Tcr8q/OieVxO9PM2bC33z3RSBTElKUxY/qYa
n07HBTN1dW+Y6oyJ4R3S4W4WyIsoKFcTKVwOF1TydUgeyR94QyTwXI3cGxDFeugCn4P7plzfBD4B
NyjSNy8OpdtrrQg025N63j5iXdmpP72uOUGS3O5W498eQC6CoHWYGvDst1SEaP4snwfVWI2W2pnT
EvreIir5C7T71vzQSPjIcdp4AcHUwaClczJ8KV7DgT4xFaJkZBrtp7NxdSRAlsPEQ473//VuBoAj
E0EPsopLZ+UFAJvxr3q5kRoBVG70GYVCGWxeK6UcLrkIXM0NQ+gg7aeJCL0caQd66LVehkjQr0zo
mOzCk7DNfC/kdsHvExL9qSBYrB3LL9sx1400YTjcf7pytj9o8yj/1sflXdQnn4zjmjFXat8U93On
RbJzYgv/1z/ZhgtQwaS/d6RQFTAK60S+uSA+8DQfMD9rKopZlRO2InLixsw0+vgP2x3a2lobVGoo
62yO9PB3oHl2vLgzBK2Mo/p3nd6NDgVjG1enqq41CvLWL8aKShFqt+SWlsZP/RN3VnXe80uvS1pz
sCm5ELCOJENeuSaNSGsvbsSgqLLDjOKok2vwL/w+3uHMD3Von2h/ElCZeJfDUeZurvP64g/I/c8d
WKu53m516tAiiBiQNDB0GeAijARhA14STfueig5e6xwqWhBHcMkxx2GN5ZaGM+UxJ/eUj+olzMTj
GydE6odEqF/aVsP33ZptQ4/gPWtJXom7XlMKZ9O8saPRWNam5xAILEnennGv2OpTIj7WVIwGC2fA
wfH5LZH40/vcfJ3LFyeMWxvbPcBvyDenC+SCDZyTWMfGH9pWeq99VNjHYkgqKhP5nNIhw2IPllU3
/t3SKP+y2dk8914HwF9CidKEM1+A/LIn3/t0V8zYVZo+eY7mJL+K+xvxG+vUYBzkfmneuLr5bACL
LGijmxWH/tiYFROHqwLpeMId5G8Ifl8SwaKYja3u7R+/qCHBiJePyDAQt7UoRgmRPpnexgLV9Mzy
7qmOU6DGf36B/hZPYJTxMT5Qu4ysLheFKz2fOx3EzAuQBSMydYMpyrqyn/+tG27XzgdwSnIEVx5o
40G97x8hBvhbP9ta8puH/rM5MNwfKksceJ9qaOfuqIa393e6fCieCc6ia4vNgvnxZxlSrB/4LTdw
5yxejLAop76zpUlj3URX/k7Hy2VIbiAA4lJPdOAa6ozowJzKSx2cvn2YHRDfpxhwjHkRk7QZqFrM
Z+Hdxybe6gV1sP7A8ReikNYb/YP45U7zsxsjablWc/ovnHHks3GZie2EazxxQGU/p8Wy5iKSRUcz
T6GloQNpz9vw3dPhSQ7Uz/msE+G2idIvvlsDnk9e5j15b1ECqF6vNtgUlaZFUI9T3X1yzPLcMmV+
akeaIlc1hyhRkxfIc9Ifu/hyLaMDybBOq/mOBi3cDISiogJRJglDQAjku7CNifZS7iMHQnh9kUkG
XMkVAgtQCEVgMtyEldccyIO22Rt+pmYXXaQWTulc8FWp1fCpTPS0cUFGSJtJRGGBLi6KBcKcQLW8
q4M+DqVKhwloi33uWGb+czrtl67k/4qHQsKMTLHIG8VkK2e9MQzbrUwGHRvcx6FugZIE5dHD/2aM
5BScb+mBY0clWkiWRWEolOPV3KBan4uBcSpZOdlahphHec8zsfki0fg/3nTQrCqB8LJjIiYOlstX
+47dn7SN0fzSoWpBBCxsvV4QzTGcBb9rAHBR6seRcwKRnrfw16gTOsLajWByA9AJcaNK+rJpAzGh
vP4XITYoi8bEid2MIG/R+X2L8u9vWpFT7+yCVzDsDb+XWjC8hYWEHPECP6pQot7V0Ge+kh6gRbjY
Qo9y9kC/RsHBl40Q/+ekVul7XMN0dmu8ZX/EvGsZt5GOIeTKr/pItcKBfl0eFmE0InS2kL4okchr
wxSmHzlRmEjOuvNDjr682eyIjBCESdr33fmqfWXQeh2vYt0UU6Oh1al1yyYQCJ7hNySgHRKDaXib
V4wzApcSsueFaX0PC+JOtRyT6jdRkqLGnCqosntXexXSIf+2SNVMScvA8528EYMwsFfz0C9yTart
xtCFsF462tGyZ1YRZMvEsI2DKvdj/RikCkRUzyAqM8wsBLExkfPfzfJ8L2L8aAsaMcX3CMauH/P8
TKrC8X+O7pe9GhdFwKPa5bvjVSOsOeQsOIACeoWFZkV5EZGv0Znj3Zjgx3qZf3aJmHqbNg+AApo/
K/X1zpxeasFeOZXpG2i5dnFrj/zzmn4YUMs3AB8IIiqoguGxp5PQy1DeDCJHGrl+rCrX7kgEkQSE
UKEDHZajkc6OL1GsA2ivGAS+1w22elfilITRTg1oUuTGE2ISg0mjrpdLgEQSqwoD1kEsupbnEDNw
RlLVfMYDpx/lu4Ked5FJrgZ8cO/WWE34SAEJAXqima2SsCd/cLqzac6SQykpj1GxahzvCjpvjfBM
Ctdml/1rXABIUGUGzI2FipYMxlFpD8lPZI2lMXZytU9y4VuozxdNwZ3u/z+SnbAsoWrfRkT+XWi6
MfGJeir2bGD3JoCvaa5cgQzR6kpy8eMfEt2Zx6yHeDGSCqG7tc1Kblgh8gb+VPIqZvuIWoj5IXLd
3Z6B3rPzwXHZGazlb7CRi4Txj7tOGVl3oEM1RnOYAAubzvojCWn6/P87t6NOpTMdcOE8mFrjREt6
+fHeRfOorzlFs3Vrc2eWcAqEXusxgWxwtGY8EMkAShVflpH5RoYW1aQZ5kgCwzyRfAiEVt0NTVS2
3LVl3Kk3iOcAJADpahtZ91CsC7octY+SRAO2xmsfwrBVAsL1NZNX0QikNFmfHhd7gXR31uF+xF4u
xZfpYHHg/q8+R84Zw6LUrSAP0LvSva2ft4h/WoRMEkELR4UYYG+qcApCfjc7zCWKS9yKViPTetiR
WIlIrpv0FiAKxwRt8lUp+tL6Il28yhS6p9FP/M2hDeYNolQR9y2nCe0lBzAKBaP5Ex0GCYGaIqyv
QsMDdje0Br0N8kZC2ioVbY94k9b6XltrwN3dc8YiWExgzAMHdJ8UCy+erSQahsqignKWeyRHfBGK
RIe8CgBq/2Sl9hPg+dVYj6k5MtNcNBbAZKKg/Z1VOoq8E3VjWu9nAWk5WGXn6v8elQLQbdL6sq4g
Lu90g2b8sDC8xgj9VyFjVirZLJWFozG9jI6f8BVh5YDM9bIJ83XahrAEH4HcfbGGmpO4nr6JY7fo
r+zfLTOCjWmPMTcQpp6Gbtb3IiMCumaFTmrGqElcj9au/dv4Slo9SeUPmOxIggvZmOt4BnGtIior
dJXhkjCnI/+AmmHkQRO3miKVKNI3u0tg2URw/ZtNYj0HbLD4dr6dpbbzSTCoeCYkhrpCo+cspQjl
Y0cpeqWvupva7nzgRgMStsZVUumuUfi94z70SdaBcOOOZSyDRs8NVx5OhaNe2K/fucWqVXkRgQ48
na0PTbTsRycLMz1ZkXUnJoIGqVJ2zqhu/Z0SfoKbzV0U/l+c9BYpoLtv47hfrHe5AZAK99EtjP3K
c9JFon5VnX5chR4Muocpclxq0lzIWDqOiKYad4v3FqzcnCYpy0EfX+WIVY4l8udIAliGgzq4IitN
WU6JsmRTnwyvRk6nR+cNzLh48hVxJiP2gngQXr8AjYNXrTCKr9wVqzhHxxLQbgshNT5TaOe7q2yj
PajFrcLUkG+mM4wNmeNUNBiisNlpolnOUr1DMVPnWS2ht2kIxzZmDKcc8bzr5fd/eFE2mkhWJlqt
GEt/38cm3OUD+FmjshNmNzDpoDyaGSb4DFuktyBp5qHxZ8I8yr2mWJGx4sruXkidf/adJl+VgyEU
qI7G9Kchtc0OgnhQzlpYCncpGksAWjsnL9XCMZmpMXUYtN0STo+TjwoeoJhVTuattuhaZ4bbXGfX
Fjm9PfySHNOFuf7WeMNVnf4hHl74qVeMOYHJACR5qHOzNqnhnihggSRjXONeoMKLFRULhi/c7CJo
StQs5qslKmpoJxDYsaiP+T4ZPDFJzH1NirkL+OQTjSgTx7EekUimzsLsdTsA1RhGWM5CK1P6VjH5
j9iCOg/kvK0YTVdZsf/ytwcR79RQByy+Xb45Ks2pKGFcDsVk5lbjCdYUbzARV2JOlnAUiQ321ckU
w6QR3uxE+T1kzhTOG2ABRtEJvQsQ68gmEvjK5E2v3etVTWkuRP9H4YeEQwll3bBLCsEOIWJ0Ye7n
3fzWfOuq50xGWGprcJ+TVucly+tbxgE4DgGrDMuqBN3kgkDxYhj71Ao1Cla3p8NrWC9fekGsnZbM
fE9JtHVP3aZndQ2qHPFgj0VDEND/aT1Ng2pumIqiirKnPkhtws5sh5SJIKul/FNlgSfC2/vRrJVX
z5OcMmQbpRZrNtGM9wSNikCQ2eZdyuhR/NTJY4M9OL/wWxsoiWd8RcCqtfUgC0/1Qstur0Fr+1DN
B693dN1ngunPwFrh2CD8zQUzHJAest4hNqtHBFkP1KmUQY5zk47VOoFDrSDrImDUsoc1vabmZjC8
xDqSJtz3LYCnQB0feCs+dxI7lOxW0+OXJrD0ysO0UKaRMc9CF2jDUTMxigxDkvm44Q55A7QG2b4q
DAxXRoM+flx0H7wCuqeBLG9YgFcMwA1/MBMMPBdh7S9MqMQyPsQIJe6+uj/nRL4l5BBzTEy6oHaG
nyzRAhhc39vVLBH6/fv14Zw26/1ysw+92S/8dOA8R9+e3NiZhKajf5itkoSpaNFVV+/Nz5mQvyHU
eExJz+FGl2KD19Z+sGK8/RR5BZNHAzK8YzOGO9YEzL+j4yJE0wwQMHFBa7+DQ1XRIClxkdlEJuB9
dnM7nFdkUYuFIpONn4biSzKL/65sTCcLhhDYrbzoF+n1SIkkBPRVy2MZ0ScTxS0SRKHOgGOaGNbf
Tvc/AfdVPkV1mqfaURpKJmoXKkV2srsreYreAOIW5YLo5CWk6c8nogmqtoRQGLaviQla+Z9hJm78
Xd+/rIwUwu+WjJLqrHILwhhX7VeNSszVuNqUK8rPp1TtAt7GQHV147tRubM2jIjlkeXrVgDLOGLz
Vzz5YLOFZ3/saxLWWyXaBZFQN1KdCI+GW4RIjcD6+Vt6+I2aQ3vxJNZVjpyG+q+Rz2PgtdP++HIh
nPZm5U4R0KvbVHOPqLElshhWtGXcbgJD7HXYFt03cY5o3j+sP+aRXD3gWxm3Y4klIjtRsUZzB4vZ
J9UEEu7kQwknUyO2vCq5CsVd+GfrckXqoFS1+2QBjnNEuZRVt0UvJR3Ltxoau+paSlvd6fTl6KDa
C4WIqZi60SVLmZAqHFpLzwNGM2acdnw6NPXbdATKRftnuo1g1T0nRT8sDHaguOHiMXaCVbUT9zJI
dBODh9FUUHiPXMdF1Bv+utK0Ko3XhKMxqaZv2+cUGGzhoPJ126TwRn7hHSMi6qRPNOgDj+ei3Fk0
qr4hi2ttkvEiJN18zot+hkyy/8TroKHwx3mnQYdQwOtbRapwE/3Pm4QH1DLfe+kQbzruv7kQjvpQ
dHnUhJldm+6mYeDaneKcyob6M4nTeDpUAsJQSd08JbZy+jBaKGDCjEL1GxBgbrCgWdjsxfjiIuDw
XoeXLCtDGo95q59S++p2dNsbZ6XHmUy//dwF//oYro6BTLVXiU9Lwzi8ZuK10P5Qw2uYOy8qyaeS
X+DfDQIDW4fER1qqcXUKikILu0m685/wKXxux0uuXTF48rMQHyuciy5cavMZqzntsk4nPlOuJWzK
ew6hKph9VIVaVjslE1+xnFJPTcNyjigIxRmpyugkbCttKj5qZ2Aoz31BYenSpHCg3dqTRR/rFOJn
wE8AlcRhnwc2CymQwXyNrhJZMMYElN8Ma73pMya1eZ1mE++MJQPTKlsop605uPz9jIGa2+yMnBsB
EZ1NtuhKmk2gYA4rNphwOaa+iAiO+T0KDTwT6B2GMO+iWDe4N9sNv0GqefQBOa9WhS44FO6+djht
jncZkl03EAD1wQcEhHpsPw+IHKUK4xJzc9DI6WiVfx0fwI4ZXCFC4ZGYMZHHjn+pLANwJ+LfAElH
Zt7Mt7iKdwVib6ZFFBsrs2Eq8+AJx81QA5CWZKLJcSiFBGfk2P4mYfgpFMlmCSQuYp1fZ+XQNlCT
aCSt3Ssb/N+Lv6KCIthe9c9GBXSMujW/i/EvToUk2CxpCeNwHSX0qcN7Dy4EheNioiX+IaX8q2zV
XeZFvoYVDadsVoaj8CHj5ULqzg7LFWXs+EZ00AJEc+1/Ew536fWFeqcktKadvLfTjV47adV3xjEn
7Qe1ajRwVwm9h0hNcnppEllBPj2foixPV0bYUww7qEQovQpr5SlN5ok8UhThCzQOiPZxIybY6lNj
L8Z0IYT80c94niWeUH/rQHD1azpwfbyOU8BC2ot6peC+UrLPPPKULTcZQx8v35lnRR469DNVYS76
YWVyB4w+xcevrreQeoABzuPzLKp/MsgxVVy1Pzg9igDbIwaMo85Xa0lkUYx60mQDGqZ16jYiU9h9
LWJXwZViSXMtMi3G7eqLCAU8ZRtUmV2ZS0Z6X3U0Lbe2fY9zwVKK7UTl0EFY46BCHE7u+bXNN+Oy
xG9nFhowHtgjiI8Jp2JTx8ToHGKbIsOrcXThEMaLHc4wfjiKEmuLRGqlo7/+H5xnHgSgVaztG7Bv
00PpTvvoYNbPJphKwuP15/ekB+ofUAZoGE3qIkiWAOF0C+zUbL6wdQiUn868itXFQGCK1PEksmz7
gVm6yCQp6Ptkjw6fzN2Zkb0PWxnG4Z1m76DTV36Moe9mNDHy6BFAwcDotWVFfFywfdGmtEZJ/Uhc
5OLRjRP5SSGsBtXA73t58LC35IJfp8ft3zkZmJPxp7sXT4oRyeSfYXCa/5K/O64wTF3y4LtCNLvI
nOW2rHHELMerV1ZZxbFJui0BLGMyfwcZlMtW1uT+aJk2RZDVfIIvmdu7b+zl95dmrEuDdlCt20+3
W9qfKc8eftzQqE0qT3IUEfBMqj4W5pJikeGBsJlGB7SuahIwfjjgkJ81GC//lcf7oWb4YXhTnX7V
r6x/+cYwjJdk41RIM8URXs5+Xy6P3jVeWv0weKWVwm6Zg7UEemXPj2xK2zwL2WBn3DRZUJ/id9cG
B7Xiz8uVlq8QbHWJdrRgkFlQWmwd3h+unS0/S/zS0Inq/cuOytVy3j1aV0w+BxHM3dlVghOh/DoE
C9EnvT8Iscfv2Xd6RjnzGzcd0X02cMbIThfmk/N49iMcoHD0PV+ko2wHEDnpZtX/WO6DzlvJzJcT
vQhpc6/GGxlMDQIt0xY72Emp+KMu5sbQOp9h7+KVrvx2i6MJQiC0T2P/GRnF+RqyKAiqRk0V4Wiw
isBG5LUDQ9uiQ3S688xQ4gyMuZhBG49DeP1/BHQ95nDNqJ38Gl0xyP2ZQlT+QMiC8ZL7eDf9qFq0
H8Tv/mVuwyAd6lsa+EvivRZPypVM2dugWxUjCbG8fIrS5G/dFBH4X/ZV15qzCPiAapjc75auBt7V
ojD3TQaNUop9IFG3DtvFN428oIC2AhjyWlCeN/qZY0DWzEbdqof5rUjdjHFFZufsDdbg8zxOkSfZ
vyrBbSu/JALaeZ34852flgofNuxz+f5TojKzHqJ+h9zGfchkk4vzCVeFNXfoPx+mQrZjQMJkrMYY
xEs5yi+RRPPJa1TUYwwuWeG4m7JDhYGlv5ttUvXecyc/7oNqBmFuiLiJlEAd3kGYeiOjsudPVOMF
XgMfSWNwA+YiBu9s6qF6e06Qq2HGVI/z/TFYPYUsn05cnXqRxJRIciSHdYGABLWkKKcnfX/5aW5B
DEYDEZldxRRUw+SwBmm3k/Bh+akKMFUpZhbbKXwqXqp/MdEbE7Uy6niOwUG0xUjhDWbYaq0fNsUv
HIsVEebl2MIIC6NUAtkUAlS+Rt0xbW+r5j48OJWev3gPHpxf0Rs+omhQXyUD4UyAIp5WNxcdUMcF
/EcmVWLNtSiIyNVcc57LhK7WawoPYAy94o9XkVi3SLA0jz+7mxraRRKkytLrjPvA313wY4lv107t
8owclKiVXHYMJ7daqW3rG9Or5lorqiox8Nt0YK+fpVR4ZGCwVgn/3UbmQvROk1RrYziclVmKqeg8
ZrsNAf9F6oJThVFLxOL5wHAGgAbk65Gy3SlwxnStNVkRx/sHKFjAviQIgnARbFkdKtyPpxI/mylq
83ndq01RTYWnlMLLQ20SFHRBuXqNpQR7GuMrtXe4K+MwwXFD1orRodzlQKoBcsxHX+ckhzFdsHka
gZFLNG1EJV5Ak+rnWc5z+m6IzU0SkoTVg5PTivA082L+WjW8GNMigWqDHD9sNEzsAelWinQSqS0X
Q8Gj4ocaOnr/E5qJe33bwH5Ve/NMFpyzHHOHz4qViqlBfNiR6fO5pUK1CeFXL+gEH8vAzfexOuV4
6L1LIBcwSjkyWbaP/udo/MV5M5bm9WWux+gNSr9dl4rQlLci3mNqv6mtHudpPTxisZraTtNNK60c
Z1vBTEWiKjE8D64wlo0kAaXYQsuYtE1NUtAN5vaDOPV4NmsFrzurSXkCZtYJfpejIteabUl0epjh
beOemq14xgvFtxTsHnh0zRNkiM5Sbb6lFGefou4e4yHRmxqvq4YAfic0XdMl3Oxx/Bf7pG7g0DSC
V4aEYJRAyXUZXFRdOq+Vl7JW73+lUWLZZeA1MdkYalDelLLXF21waEXI2nXsES6h+ALZ26+UZPEn
Jv5OnMxBKYHH25py4Xz2R3KUb+48huc0BEEwwM8/W76wKdws7t0q44QWPqBMc7KG6L2b2Q2UWNxW
iPuV1h6/ECLsILsIJkiBjClFo51ZeUZU5Uyb+C2+D130lg2pQ4yX+8IUgZQy/PjLd/sqIoGi6rTT
PRE7fZKhSPo6Kzw9fzolRGw4PxbzJdRmN8yjjJtJv5Q4mo0vXJSYn/ZBbuiJz2z+IdUUZmvguxe8
g8MU7eFgFTpEGu1olLKqcJey8zggYWc/cSswSZMAd37N5H//1DPv0GVnNR4Yw5M8J6AEk68/QwxA
tf0bcv24k7lkBU2YL6A8pms0HKQemTr32GJ6+jhWWX9WLbpynRf3F4WlsfCoBKpU1Pw93v2UxrIx
NSHhkxpL5QPe7tlW01h93Tu08nq5yp/q19CfPNKxcrB85Lr+KBseWW+O7xkebLL5Qop+8RNzmYsq
VDhRxfl8frxr74L3Vn50MK4tYFxJj/Q1HbjXL762ed8pAynPriZ1YlSg3VcwXoyjMJKXFlfAtx5N
6QThPqO0MWGF/KQwfVU8QTopxKfaYC/3c3J9r5W8k2bsapmdLBKRE/Wvh3pjMSLTuQjL4KpyMoYQ
GAyIO0kFLh1KOYVYYwTEuV3S+DxvgXI/QQvaRcuv0tpuVEUnpY4KLFPTfoaKuKd95/AR+vLUHPcD
Mt1ZhKiLt0REpTUskGpjjk6fUV1AxDWffQcMe5EyVoklafWd8P6kK00uaeBQxxvVj0sxzLXIJK0e
TnlrGkV6fkfefJLODa4ADBjAOHWpc39D4qn8SuJkJL12ycrFMEBTlMbZDdcOsj+A2R9EyIXzlBhJ
2e8BGPsxdSTg2OCQzgup0B0rn/I0jtxo8Z61otGtxRA41KwHLt3jmj2K9oC0DEJ71C4kQt3lGnX9
zphuq4xZMnQ8NBp2no4MDqA6++iAj8FiKN/qw5mUi0/cpWCtxPnnU3cjoSqe+HNq4ErGOkPlxgvu
KugisJX6TJZl9YQC1bQ9iKeX7dAbtNUyVwQ87Y1fd1I4JYNOjvR90w58bxVkS9EiULkDOQ/xmgEq
s9T1H4+vQ5B/oJHao6nd+lvGds3lZp6FXAxfZlXvHe/KiOTng7550Owge2MDOIuiydQYI7G+/nxL
ingVgrJudB6m1qyEiLV+IiMQvytSG6/dVmEPzALexnLEysqq9cC2Z428vqXPi+YAq3xg9tNiGJYo
FkuVS15+upVPH+Y3+SxcWmovj8YwWmndA22ppp+e3QEiO/YcsgDL+MNv/t3Qu2oxVfK0IKVpWbil
mi5ORZJMMj36rSU4Ptr7Pc/3CxEaDmgKesXiVNv8aaf4EUkSzZ/cLsq6E+f8CdOjlnmEAXqGKs34
xH6ska99oN9wU64iDXjZcL19QmwYZNSXLD8Ubg3dO3FAIjaA3VoypHMbHmzbdRDysI/eZpCrWQbA
sO3g9HCHlKMllAQERqIy+IjI+KBAGYqFNOuki1B2a1nixGKiYWr8PMspzl+lf+fAK8whvbXDEY1+
0PkNBSwNXga5HzW6y0f09qFCdV8A/BWSK4mSPWZxj6B/6MNg93qGBhzZGWz7oXNIkpaW1z3J9AF0
+1K4G4aJPiAVF887ViRNu1mA38GiQ+MTmG0QssV1uMind54HsZRHoXI3PxTZXagk9AKu+EqrceJ3
FyNdsX4o4+7GQNXSLfxkhhUzzfS6asp6Cv6S1c1H5vw2uILKeqf8ZM1wqkVTSa4+v/MqJYn1I+WF
ySRejEDlJvyCTVd27KbLO0PAWzjGfSKvZ2m71y9KntyYa95soBe9sic2CTK1ugLvP4xBVX82lQUO
5XVA5IeJEWkfk8ytZCVwPyuRKN7fK10TnzofeA6xnIzmUhcGK9s4FzZ7zvgVGnzfO1/WKoj5CKGI
iyaXvBs3CTlbT3vJqjgetAOgxl2mHkNQf1Zv5QYD3jkXcjcpLCcKczcDGZjgBzOHdyrnudPtaSDI
x6OAYxU5lkCooWuyE3rH5HXHBG9hdmOfPGklnpx1JLvcNoPVVo3XDbadfvgMoBu5E3K7651d2ukG
zuUyjvmEZheSdItI35mVpS/fDfJ5mPChJhm1HNtLrevUwv66j82bOatNtrn/OqAqk/YvX/ELs/yR
tva/SQRJY+0B8RBricaRMCYSBaEy6V6tFivsVsFEKEGR1AQFszGbP4iiLeFESJPf9ZXpsZwUQHS3
QQ76QbajQbX0phU+/dUf930c44iOlw2L1dZCJBeSq23EQb/5NPcClOvidNj3+sy/Cj3nQOIxDxq+
IdwJqZtJHLFhmz0oqJU2btcZmV/hCpmHLPhDk5kO5BH/v72A5NYy0kIhV25SKDuMSYgdacDWUWHO
x9inqLrkXVCMyWKMzSCy5MMVna59DpY79HLfNEddmZawOvGk0LyrOhUdlASGDhs4tGyzTlYtNvzB
BQTV1S8TO+zZijzj2FvdXCg3LIKct2yHRdGqKb9CWnqZADU9pF8DlH38RBSRq7Y8reRhQ92JJhKh
Xw6DhY34yUlXMRV/Q2UPt1ferui7ShkuEPiggRzSYFbe1OSc7erS6c9ZGvq2BPWV3tal7kWOA5S4
jVdYlK2xlythvP+jnGZxx3LTmwk9klGccFKdGHwIvXabmz3wbTyQoUiQGwY2IJytPZCvbaKDg2tb
xjC71JjhgH8jkBUzvePRJEdqSEVd5tpi9r1KeQz7tyn/MnAdv7WcxRWHrLJfVKxibOQtw8PUX/KQ
CF2GZ2JmANduWRSNoWO4wls58R5ARI9XYJTUO1AwFpnDGfKL+UDBL+s5VwRZ7wNxILjamlX2tc0b
j/uO2yxUVTfEZcdIG0ryBeBx4cqWhs5bjE43sRC8g49M5F+odkHJywJgpLkbD+zhdWb9yOj41ZA5
1fTwwcFYobxqMDJoqhmPxMM47M25cuJtxeDFnvRseNGPPSr6MHfAXdAcVPwE28KWaVsIlhXPvN2s
dXSyRTAt3L7DviSv4nqai9NCYGQ2mouGDZlhse4woSD0wMW03Gi2rc86C7nhut5oiHfa3dhy/6Xa
IPx4VIucph+/vpTrueGvher/8B+JqFV6vW0tgPMbSW08/ozs0pD5VT0BHTtHBiiOUP8qOZM1i60L
AC9j2PsujabxD57Udy4AhMHgCEOG945Jzg33ZuPBjwaoPVcTYGMQwGurXOqAaAqHEsrFQ2sZHGbi
blGMfWyx00Oe6obR/cAbsqhQjYniFb59cN6or9HaxwFN0FgvqkIlDLQRdSc+6M4i6d7KZfW8F7s5
REtU1vg6tKIeZzgo3MPtmFr+/tfayaM5o6lKkLPhyhYzU7B1SGl7Qrhc6qyerqPBIz7GACtDG9Zb
wRvLHl/zQc7PUES5w4KsGVfX7oEvLMEj2okdmWZHZLQBAvFWIVtF+PDYqX8+jB6APJwt721RAwfh
+E7uGItkh8ExBMfSydv42E98xqYoHzsbjMg91BHaJFFuyQE+5kQxgxQGls205SQPkFpwFI6+dDwh
Bfn18rDsldACYSEQK4eowUFEMZLmwGrWyMR7zWYJkjZoc2mRKlS+5BD+csc0gwQBzCniIuc3ho4t
Wb1a5aj7U389fIfByIDpAfWoP5BdESAuR8lE5dhuAZcgaNV+EtfbiPtNF5z+NuTjd1mqdIPPgssm
ja7kBPl81nsGcdDTHXMBGWNBXVVvPF39CliQhWnozY1vU92NsyJ2AsUvKCv1aH24xXAupOguFEkH
alPfmkQ03Cs8MP88gwcIYGcOgRKRGBCGe84m5mchHBAAjwRDvU4dEUIGNumxs62BZLuhSaqhfntS
KcVetGXhvztdvmDe/+j6v9k2z2bstCMelnAiGWB6ujLLGcQOveHvFg9ywSAv7+xETaVvGf4BQl8Y
kY4RnCL5hOi5uPnV9IGezkE9bc0Y8Bs8Pd8dWbvW3UXCP/aDp3PlnmqgBeazCgwx3YQYtuNMW6aQ
zh+STBsW2k6fsGkVg/z1TDgF0Xme/rrQa/qKe0PAevNQpirw296Cn0fOWgdu+k/BTm2O+HgXh2WA
qIRzDUag4yx3lMHPSEIlvghI8kepzQFGveXUG0Wy2EspIbUM2yyGz+jKwGbFzzhLlbXdOXJuVhb6
3/TzBobdb/qH9EArPMB/EUJknuFsqO581RCK30aRUOwl2jXsUXKKFyTjQjV5Kq4um+8eojYd4rhJ
/Ons3TneCG9/oMMvAjz87HlQDsczDW0G3ZhLIAUHTIkBRXEXr/2QkJz8bhtgA9N8TxQLpwzeY1bM
YUBaZmjiM4f52CEZ4MHAgyWDGuxwNMBpbrobmovQ9EiBKsBNPGCXpC2nuWVQIuOGTiVkIjXbd07/
OP0GS9/n2QddXxP/rFzIWVnhgHM/n933Lmkvb25m5JR/vaiGb+i/sfv7ZyLOGgagx5K53XFpwq6R
6MVldlesa2elid5yyOg+fKiwws3xblClU/X6sEozdUh/fjp/IVoO54tnihxg5bqSFc0fdlmiAjfy
bN0zoIH8OAGzO5lllnsrIYibqIkN7Kwsv4bdZGiobfsLHiH3pwVoDDycs5r/Afjlper751590eNV
l1o/U+lP75ofqmiT9FeQsp6t04UTDBVT5JJB/mWfjU0sw6Pw2xX2K0OQ21/6QWzR+bePUjs7xDRo
PHBL/GjL8VGDA/Sy9ce/zPb1KdCyNB1ZaoFNMt42araPF9CGliL50Qxqm4MafLEmWsUSmiaYnbsP
a/r/bR2qSR82eLe++n7JsM2lgwXweye+S2kRZBuHimdlZ+uhGwWebDvVGNuxhPEBYPteT1u2t7SD
gGp4p/KYWrUnptjBc+GiyUVmp57X0L3ZM/EUXe3Pwm7wYFpicL0DFhaYHdlqZu4X+BhSrBvC/gc6
9sCEr/vJMhNt06ismlPf8nGFe8nTwK2Z8hs/mvxZ59Bc63HwsoPscmhu7zPnjKHzSBByeVyqhTy1
GXTEOJo2V7CV6LzaoPF1sq7iyYBACrOsM+R+NoBhYfzkHUGv9mE+M44uuCOeqK/xyZHVqZcMCGqu
k2L55/rVuhuQ2Rwh/N8g1oRyoKxFViJk/zSnkOgtmyS6WSmqPPdP4QTsQI6K6kazJTtKcm1gpq+1
XsNY36sTDhKyGPRAc166yIROsx5c1ZXz3PRLVNNFE2pq3F+goxLTHwMj6MpfwazHvtQtcLow6XzT
hrcXO4IkfrQT4EyzYblMNI2pSg9URjkIEyNEwRff6hRfud0rtftmNGgRRmzGkYY+ibVy24pfXgqG
/qaRUoSFR0cev3OEZfaKxP247+svBYan3yFtYTe5KjZp6PECyxGNSYYiGCRr6MzblbyUXWuKnQzb
VeICQhGVlGZ53AXHlhgeuJDmNg0Zoyv1ZrkrP5860JNm2L6pQQ24tX7RSMXmqdEmBXan3Md2objU
tbpXJlNyZxGpImOFwaFeL/17rlx87MALOeL2Cguix1tgtldehXXM5zRGj/5pn+TzkgX9T9TM2hw0
xfOCG0i8VOMyjgjG9Ln7Ir0yQH1rQfOo396TAE8wVY5BMqCVOy4L/jQovBdCO9rp9+Fsu4V4397Z
e2xM1I4Dd3afAl9POyHFP6Bi1eaSFa7QdpipnRtV3Lio0OSCLJHu05qB3rXGr3RodgXehzcrqSeI
3vmCh0jhCW/re96lYQybiSfR2NqiOZ2TpYIrGG0Y1uOeCTAlLBzGNgJnr0FmW/BZ/5J/SwC7naKQ
3ue7wgjpDtAwMEf3gvdeY/FK83cwiNQeaWPUeXW59J2bayaMGpFPglL5JeXuxtE1H+TWQ/FRN8vS
Mvuy/gXrphZp21M/Gw5XiVrgolJZRNORom8y/VChuLqINIw6+Oz31EF6qKz8Uzhrr96SmzLAWpAg
N1VcKIW6BHwql8K+8VAPl/qEw3v6qYI101bm5R7smEeMlI3R0hGX1PLYalGXtR2mQN3tOxwdKesl
pxoBZB7YpI2xc7uMx4tqpWy+YStbdvLzVLEhNj4JRuQoyPKcmATYb571XXYFvQYd3UzbvhJjB+gc
5xCNBJGVwaNk3womjYlCH4luv7tEbhOaAFqNxi1fLjCoaFRt5f1JQhuX8gIuBk1Uu/QYeNYELQoW
rOcarv2vIDmjF+YCX9XOXRUj3N/GTl07P8lzv+BToGsjSlOiH12gf45V7NpscBsKKCKBBgeVN9YR
j9OFLZzJDWlEyqWi1IDQ7vWFouD4ta01kFtE8pmsRVQrjEuQKtsHn9iDfQDIUxuQrjTrTggLG/S0
gCrGldeb+Rvos5lPUM/weDbHTx6b0sOeWDwstOxlAz8z+kmG9RamAVxJL3NmzyKWte8ZUWwG84cu
3MZQO2JXQ0tHfXtY7PG+Vl1BErXUVEhMMgH9VM4wuap3qEGzpkU4km14LNG0SOgnH8fSRQjGlCjb
F5n1OC0Ni/zG/EMdqTTKH22RuOg64eV7BCGeEkqPUVDp8E7CV2xlQjd2qotq2pxQ6Y+Xjh746C/1
X+/YsF1cxPlR3WNG5aWY6cRp92mUlAScCfrARGC/++hyn42sioK4wiD22LYiF4Ki0jbxOZJplp/3
asuNIq1ykO6wsGikFCUbJsbqSmhv8OPmMWFnRpmv2L3i2CVY4ZihsUlEct0SUV38oOdS0fToP0KM
5DvbfsIirGvosVKlSTRNggH0fAm9wcfDdE/NIOZ8OnlrxopBhyKk+81/KB00/E5ptplwNfhWSNi/
6bI3Ox3/yF3qMzjV3FKn9ttefnPhuXhPR/l5q4uApzfpz6QT2EkhfdtZoKcx8KZsbcmGJ8qaJidV
tu6sVpfggdYkLvLDJyRQiSF7h9hqWoGjKFZmkpaT23/SOysxFbqbivskPKqh0+eY0jWoTjWx29jo
5jk9gAyEsOND1K5M2eEVWrh3sUA6Ky0H7aXyNQBoVOUfNAaMmDE9bJ2lr8oM/m3oLoVyVCGBpZop
rskAZpJmfuTrPTZIBFEGBqAh8DsbtfA/CqDDNGx9N8BNXyq1H23XWlkNMwEA7rNeVD2+4BspLPsb
62jr9WOIAyyP8JCZo0MzegWguc1UkN8wxMpN6CBCASxu3r/VAA2ySpKpBL8/yBCoXTBckMT89o8X
QBdKiDKcPx3k3zTS0vJ79iZ1jR+jLVffd5NhfzNp/pYBYA6sokCfRfx3DxxqN2TNZrpcA3H5yvGg
G9UnvSKD6O1auOCXtZ3rL0VRJQcp1JuALUzUaVUJr6xlqcvqjcjLT43UYx/44E9RwYnJNEeaIHNc
ompuVaARj4l24sJ48qwWcL3xsg3LZbWdDBBOBzOHKG8U2kjXdjjRKFg7FkTcmxyxmNeKcuhXwiZG
Y4WCQiBcGw+Fo5OB8TeoIn+ucABWxjlP6swzDk/iVCnLH17FpEjQ8JfaWrsvZQ0JK+MStJvmp+Yn
1u02bFe0Iuw5TY1Y/kdaUMpf52Qzm8Rpsm/csuKxQTX2M4MeUnwChjLr3XmRqwmpKMu0UztVcKdH
zJCYaXYiXhyGD18xMGA/qTV7yHsQ2ISM5sUIYcIw5caS/chXB1Auog2jMo5Fsu5GzuoTB7JeYNx7
WTGQRRsxsYVKpockirNMpGuPvZC/0Lz2bsGTGQZIPyPj09ew+um06tNmKOCKRVJM54X+302DvdxL
GmgVCIr9K6D3yLOuoTzh3guZjZ+5QkKR8Uo9DLAOTtbrNupZGV4y5K7Jt4j26wM3THabm1tvB0fS
tuct04S8NFbKVY4HgxjgprXvQo3fuhZSdwUzbRzjx9MXvda96KvBo+qUJ0gMu5DcC7gWPR9rGqOh
kHU76kakHvCQ3q+QEa3yeJBse/xc/KO1NR6yCQQYfboE8EmxE+9zMqOfggRI+x6S37F69EfItdIt
24ajPYXh6fMAFrPU5XvA1QRBCsgj6jHlox9HnCrOMq41wS3K9p9IaTmvrvwiq4c83uQjfhSjzBIt
cLZwHdgQqUXcft+lGwhv6dtlzZIK4snc9hR1BWl7jMuWNjzCiZLMUfGkOUdcGMZAszsqNpy59vJh
iJSZAMsnHnRte3+OepIE9uopnWJ7UPqyNRFIMV791mx8vuzEg7H+BpewuRQKunP9FnEZcjXjoJkp
clVrd0i9zj0KxqNyhp7rqHa1tbIRGluNXw1VkGbMwdZst02TVGK6gSGvfzEJaIjnUa67bUbwCIBV
GJzR5mUj4OK78TE0jLuaCEDcVeHfv++fSfaCUK/0ueBsBic1zcbELpcLfUarE3nkawu0/zljK3RT
5YI1a3n4eZe6Ma0B05oxWz4GaJ336a/PdfIO0yxZIiov7xInI1wWQ4HA59NeS1tse2J/QlmGUvFL
4PcxntBHcJuLA+KpGGraUJnvfoI3T9nP2Ev+19Sh4OUZdH0IjluZz5ZoRSW07KlxCu9bDE8TBuEU
s8joXBsO7V6siulF1Jlb2FTuI6V9Mkloj3QhHTRLgxlVFPT/tG7H6MCnfSx6StfwM/JAai+V82z4
KUmXNzx+KpwadbiCWSNVJSaRwK0AZzVg3mKjljlH1LAfcVOMELubbLr0SoOPxcoJj9nCRmQxgvsV
b/XsZr6PyUNC+hgNKsG9Fgjn5VfPLFoUYWxnanXHgYbaluU13IRuDLje2ix0yYjI05vh+B5HTATv
wN2wI6nFOhO9mDwuFGZwlWEoxrR5vRCn8lV//bq0jf3ES19NdAkykrEbwQaHJJFEzTB/AqIihFBD
lGYJpXdyGmUttGHprBejEGTyxHB62pZNrU+LjZOUEo1NPYt92c8VebnNgq7v04fsFGmjnRYkChkm
YxPbk2/Ml/j5BLxRL7cZfFb/hMWLwBLnK+ZIoliDg34qvdqszcOcx7FyPP1Op8saiNBHkW6I1Pem
n8CZwsXDVXNvJRYRwG1cjdX6rgT2XEJ/t192O4qu4PUGUfEK7oa2qIY5KOlGiKoirZlSqInBlB8f
oXbXaH1LanF5rsBySnlc+41flhhvjFaKF1qJ9CyJGzS+IBYiWA0oIo/hrWC7U20bD9wRg/mUGkin
BJhLQDfsgeGU29vWoNEv63zkcyHEAlWx/uQ+/4zrrfIDB6V1hq2o63uBH9p+wX66ZDaT9m+zmOVd
AlVvgCk1YWR9KdRsyMjgAvPk0a+dEKKA+3dDOi18h+085Bv4I4X45vDxIwoNPqh5Wn04ZCL7ZmxC
7kILQI9fDg4yorMJ590rU3tbnnxguK8YCFQmApFfTnFGEl1v0oB03b4omyM4jtctrqYE31p9Qb6p
uKCYWV9bsg7AGo76K4b2vRGuzBpFh+RNOfH1pq/HDKkkxGZvIAcdthFQ4liDpQxTnZFJj2Ibv/13
RDkA4MnEZ4+g6ur6NnrLfyZBVz3Wp2xoXYAjxdydwBP2VnjSM34aFiyp1nWTFZV4mowpyeAdXm6E
p5RIxTsICTna50+EX3boGtF6kMtjg/10tiAZdXOE4cteI4R1cZkZe78gH+r7IxyCv2K4A99Q9byZ
yQi8S1ekJpfeUg+JToGdIt0I/oSUWVOLe23L/S/5f6Sl44UB8NMFaTOLr8hkYziY6Rvp8CGgJmbA
xn8R9CuzsXF+7tg3+Zpjws7glbs/JqZiYAcJo3XnWC8AjzXErfriRxub2mtl8mU0KnfrfvecB5c2
Oj9AUdlo44wb3jpFh9kYkHw/2oqmbCbGuGtnGYY4mZcXn+wTZ7RWArAZNPVamIyUHKE6Bv8x5MO/
WzTiHlaTW9MhFmEciG8m6poOrsAZxHFjZPaudxFkeEDYrlj4muRAhF55P3W7i677hywWw+bU/+rd
f5QDFeO2E4S1XVCYBfetKwkh5x+BI46EonLDISkBfAUBDi0Ft72CjybqxsqyU6FjTbZRgbvYdVq3
PL94qy5q0/dpTs8colNreLeXIxoqtyLF/owKdtxd43tsUtDkkURrFWME8T0LwiwBMA53lhMoNZPX
wi0Iov6wGFVidicfG+uXNHhiMyXaDpB58Oq68c1wASLHUArsQMzvL5WKOnSlDe0F3kf3DVnzwYeg
m03vbCTSRwQetmrtdeBYKU4qKw98bmZ0qNT8qBlRGLryTvJWE4rXs5GzGGMDfJmYaWSZ8QqqqljY
ba2R3A6orBDfosdXJeb7WjYWoT7qDJC0z3AWEzf1k8kAEl2m0SiOJq2KVHf37E+yPXkxCfuzQXx/
uf5bA9ZlsVar2Fib3wy5kpoFS1aI7o1qtwik2kNZmILTpglDQqGVp5C7TqydjuAozKyK2c/Y5Bb4
wSzGFEFcKDGpQV6YI1SS/UvIM0UHms7ts7S4dXw0Nh+L3U5wpFAQT/Hz23ABMg3xFGZ9YK+KL2vs
f70Un+u1zZVJTHjrT/61Mdl+cO2IKStih3SoWy4ti//Zh5r1FUNrZkWBW84ShmSDb//FltPmsUsQ
OYxFaV6LFxomOnPkVyWSC1rY/Pr8zZumZUrUh7kGXGueGyrJK3Cy5p12GJZTEGgyiMm5uy1T22tK
1P09RahzRieFKyBpBdEJp3fms14Y4R/PeWFuIQDi8DuVD/jR9Iji0yo3fogbr6Wc0Vj6X5NuKYDQ
2H7GuDgd+wrGgJpiusNNsbGUfHpZpBQ/4opPxHnC1+hWXSTxUtPY3hys9hElOkwoFLi5gJdNis43
60h2zFuYZ/JXqrlNw91PS88otal2ExYdRT4WjXFqcKy2JQ2luGCCpGCOAJAjbBz4uwgMyXzwp5Rg
BUqdHCjKkQjIlmq5alvNfbFRAQmIDoDvrIHEMHtrCntVKQJoaxw8T0aW/Ti2qAst0Tdjxp9RJ4wh
ftBJvPo7hqlmJtNdXGhBQPvMGvBk5cORCBl9x5BDmWz4f7RZV+6whcwKV7qFRTfMRHnH0GTLqpgb
IPdvNW4xtzn//aUD2EaYrVV4fwSDrlp8AV/nQW4Ok/yH26LS2T6VHmAUdQl8jEM4w4JqTVAEcNpG
N2w5b4XXUSxuLYi36tNbATRQ3OHK0T0BRXs0ZnB73OcIFqYZ8RTGS/FNoNhZ4T2aTCgjWGejy8O8
+zFlCoNv6TGnGOGPMbNVuaUPyufdwW5PNfGhfDmZ5vgVnqK6fmAfvvaAcj5QLNusvI1DSnyyxvSG
zEkwGJX/IzoZo3qiCKAsWWZBVmEryJDupD4MsLZeWT3uCL/QK6Pz5IwXA52xnUicctSZuoj9way/
OOjxkpiRbWl45PTA9g4kprPsPM1h646VFEmdA64XMHgFbIdzmbTnTNTTCDvfy8DxeBv+30xcQv7A
RfmbVgKThXrcj3c8LgLwyA0wvX2+sYHcusLUzDg21ZpL3j3UH43qzNzefHLl3aQxBKZkNmI3sn0K
cW5kACmt5Qju6vV6hB39ZkgALf/L75qxn4AVjVbXNg17ech8FdSEmVVg/IDMzKD98SWzCuXPSkGt
miEsfQKD3qXxo6Sim5ObnrqefnVmPTdx3FcLK/dED7rdvH82tXxez6IAZl1DPaFljEhnG3bYsFmA
QeWQnEuXzKv0L0m/GskSgH+wvw6ZM28J9EBey9Eym6f/2ALiQLu3IxOU5XgUzlIVPP6DNOuHo68l
4ICvt4Q/zJa/EmKC0nASHNEWxw5UM72aN/tSWTa3lIaxmWtW63qpFj/Gb/TtLABDbBEtvvVQM66e
UbQ/k7qp0QvEE7oYt4xmL337x+z2XVYLdBmkY2isdNU7e0xiZAbLUg5ptzoZ00So5sOG7YBNe3Xh
Ogcc491S4RjEWquBCke+ov+7rrXV6iQPEiSwyHW5j7LKTsBHDBFWINws/5+aO696lfmYW51Bs2LZ
ISQaoDIpc3mf05XDljbbDMDw/rkKVA/9l1Z8uQjxnxgdlcTbrerpHWNSDgr35ggOdxLw3VY4zQfO
Ql/lcKSORmufNJ2fjxRHTCtPC5xJYIxQkJ7R5l+51aeeal0cX7/s9qfIIdi1RyPLU78ExofThk90
bMKKYDWxoOHcdRV3kUbU5kEfFUOHtH2uVdsvCET3w76yXL6zYvQynuksW+ZsDI+6pBE6d7Th9pT/
58slh6HqNgpB9yJ+yAYoLgoh4gYkhwinvBWjKy3qhWoErq4NHSnpz3opgmD7oc/PU3Y6ui7Qb070
GFdEoaZlGnLTLDpvebUWYdJaroS954CvOJ6+lAxq/9wMZP/NuGKxXOaDtvWSL1ZVM34einIWJ/bb
IYSxqur8lIluF+XrUZvMnbwQLs+fyk3XHYw4n/XswjssnRqdDEBb5pTahiS7jFVVOpbosB9q4eHN
MI6BZ0MRJXTCCatbKzO+6HGUBuPw3QuW4EMpaHNoFVwjBpi68Hgxt9a42puSngFKnQ/ENkcbloEl
/k0k3M1x1K4tcyXWUPnUhZeges4lM/kWTPUK1dAm2wWRwSNtlzcNiKWfAARIb4O5dRjMOARkKpPX
lcf+hCv79mPLF1S+qnGxGHsLIyq4pVvnDuiMP9XYENJAw+CKPRcW51HMmUbKJdd7tW9vCV3SYtGK
Y7h/KzHQxJchfeRnZRIfEh81C6gRLwDCguVLrAWafwPZcojQ3B2RavK2V4aIfJMlJ2Iv9ile9die
FOIOQdbxc6OX5qO/UuFOdZfDJvHS3zEKdIYAJH3eUGMFtM2EXGc4Qu2N0yH1s7buy43C1KuasLHE
NwfMQ3gBmzOIJG+1hVP0CdcvBulA3MqihWn6wiNsOJk4K5yLA6PGp7KIYFvNxfrkCJVw6WlykmuV
cl6s4znvDPqd7rGWw+fPXB0FoyGDFkZg7P67tZRXmyCxGAwyfl6e/S0Wkmzt3lT4aJqHv1bITZOu
8S1TqSsfws7tpfpO59Di5rVseiZ8e6xGuOTYk6W5/Ni49ugvgdFU9lWDcjgXHg7zUHfTfjw1Da1e
w1IWhbtg/7ZFr9BZPKMrDrwmMuo7Kgg1YP/j3wE2/LMBor5oZeDtrevgHFOwIW3gJ+FC0kuQY2Gu
2xSvNOE8Q3gUDS/rvAawXkreCqPMquIDBOOJPsxc9ukv2bXGnCAEuS4XTZ/Wp5JdRADL4K2XVndG
QWi2kIQProCgYP7acMlJZ3YHON2nArqUhFroZlTcvdQjNjYYKQUSLppnNfWiOtVIzd6LNyYqa8vK
SCHF1pR074GkjnGodd6pDcQ/na3Dw9VO+Xe+o8JzIoJK3+3JGMvU92ZW8Evnq+iHRc7oergqvwpa
y3X9vraKsmno9iPjkO53Qwbsi6KsI+Io2DWG7CYqlzk44q/BvSOOvXDLAfi50RApdux9Q8EospEE
nZW5LLFCnaRWBNNLKHYpiiU/+rgSLQRjoNxuPRxxXKqAoXNRz4yDlULktJNr7rLd5DDyhIOdWzDm
/p2Pa0/QPKyLDGUOZ+fOvLmMITh3kIrxKC1AOuwu8pBuSnzCA3BynfWfI4m+JuF0s9SgVG4gKuem
3qRm3a2X3TKPpfvBDpJrIlvwtiNEUGYARz+XhJaDWW7byUhuTkA7gQ8nOFNKph0sDll+OUIQcRVT
H7ytj5dvEuw4Vn/Htsg8F1js2GNxGmy+Kr0SujODjYE6sMpEqr7QYcTi2ldSrNf3vZphGqN8/DfW
b9SPYodnrw7I9KAy9JKk0Z4M76uKeHAF5sa4XWcWjslvh26UUIhTPODV67QLoRsZQoU2Jw2sc5tH
tb9cvWAwXnKOq5+rHzGxhMLB09+1uiwbvBCguyhLWwAo1A2432lwiGxcZZo3fGNr3hSGUk+5BpOU
heoWzrv4MyPNgGnLbXmd2FYAGBHytOeL/EFvG3CQRsCbjyenjd1l5+XmtTfYSgf5b7ju0GeHBAgG
dn+XjVGE8t5fOdX7SiZ+KcCw9yFiDYcPMys3MB82uJxdyeXSPdOtVJgwwoAftPc/bC6wZncBfLTv
+p3QiftGsqzCww9rdG3ykTdQ4jXRPSKd7nIvbEDUBA6p166r5SjL/szxabLBLLVJqAC4hTSzrwl2
6wGVePD325NNsEQbUATqiaiqnF/ytISAx0MOYVDkFHt2DdR9XLjGcD0wHJSh0HttKYYoYrnFaR3i
cl7sqBKZMBPcbIIP2BeI4/Kost7R3HGr5CRmDLi1buBKEjF9jQ//aSTHzdPKftyXnU+niakWSgnv
TFZjhj6R8gu8DMYyuoNNEdH+d+lqv6fp9DXnKPb4ZAtnQxpK9mnE3S1ivkStcRj7YeOHeYjQYXly
eazha4BqXbOtRAsuo7LZMGAs18WKWQOhWvxHZms5YG/JsoCMK4L0cUoBdp61TRkfSk9Na0Sga+6/
KCQMZqVeFOOAznk6OqtF8g6estWtLqHqLcCILF9oVVcs2ZsLwB9WpVrFJf6lzgL3f6U4sLOccnrz
K5PytM2FB4l9ELjYi6WqWq7j3zt9DWJv7qiBFJ5yg9Ux8n4rw7E/e298IFIZFOfTeEpeyh8mxqrR
Q7Kjk+70vQ8wRIChM/GqqKoa08uTtS8Ov0hNEBq9DazxY3S3u9Jo4JZxQKEpJMUwZ/VRUg3XcsmP
JNBkGsFoNYQ9tbcbjKwMKa6DeS11x0YjlcsDzfQXT+MxDe8OduYp7MJBO6Bq3WzbQCAf0q05Zs2g
xt9wO+40vzzFpTESsIO9Q2UkG1jaiLmbYjBvXNQ3cqmTNVvinoXHY6uMRgr0ybvG2jheOz+qWp7D
gBCJJDCZd7nkWSMfJDhGZzeEMt7LgLsQvga7Ym3Mc55moWo2Az2EOMVb8Rv+nzaYc7WsyCJaliRs
g3q+qZkP6sTFGcIZKEQsWIb67JIs8flHERsRhD4zsucC5tnUiyrROqsBoxt9e19Ekx5TFRQ8yasi
n1g9KunHo+Q+nvWrhsxlPeNpXw7kBNY90Tdz5PAjRcFcLEbdBp3Ev1beB+cjlkun/1IiE6ymi4N4
sq/a1DjEzws6E8Nj5Fqzp9Ofc8i9K+C0vANOBsrhg5hFHc+vSNAZdc5wDUAVgO3OVHQyYCE6GyCh
BCDb4iRb8aGA3G4CnX2A/kIAPXXLC/4B+7H0GNmKSX4T2eF1oZ/o0PFh23zMRK4OcukpwvRRKmbZ
2Fd4Jq6DpFamf5c/eED4C8seQKKAEcAEW8spoNh6RfvADom25gZP1u/moZ2fuWMVsopl9LcMBdBl
IkC6t+J5Mv74m9cM0A52Y5pLdBR8MBkLt8jyl5KFwzIFW0hPoE9+ho88ecU0DDfhEj1SV6YK6hul
PCTQGWkNTPEd6T0ORryi58npr8akbZc99Kwv9TV0Rs3GV3wNUyhBRwlIvhazPmJTCovoJtAB4UZt
ZMdmoXaJnit1SjKPIokH9KuZ9meUT3kDfzGkdf7DWfTNdAGAjPx3K4/klWL2RJhCa3dNxqiTdtcn
Yza4FfjRsqM6oX+A7p0xfeaV9tWkLQqx2dO/1Xft9lseWS7a2WSHXKjSbSiTv75N5lXvLQotqe53
iG8Nlr6V6DzAypFUIWoR2DXeD2WlNb+o1vuAVPfxZGqjRQqnEoa4wWGw022A+NbH4KIV2iU3JqKs
Hxo9Ma8xdvR/lnBvTE1nFoOp8IjFiUmJ8D9iWblWNeXpY0xzxAehHfQePnAvy5mvYYIqeKOphBhC
N4lRdInub7R/SLVyRpT1xfz0QCB9DByCYi2ZFIYP2GRuq8LN0ct8Qt+UFJP6mpvuahxfXRzuxGQa
zUqZ4NwmUafFvR2GpF5kPRzb3FmsJyIMKznJg60KKalLwU23qZOrkUQgkeOI5qpvTV3KP1fcCIle
S998CqSR43wpCCGVcVGQ+r+PfXPZ8gajgog8DhceaiL5+zuL3hc0NttHn0J7I3VaPlzO2BCV5n0f
PX3VhzSzWZ7iVtvB/38wH6AYlKsIaQY4ILssuL7YihzWML6TyWVvHxj4hW7gsBBWFYSBDf0WYdj7
81qCoj1ksNUQvLdSI48Xi9P3FmngSGwkVw3368SiP1Mb/kbzkzmsDhpwzsEesfaUNPgMexJqlyAU
6WcMyqtOvT0SVydXYTqh76TxJJOSIo9HKu9XOjx1Q0fGTOFT764UhaFteh2C5tNE3CUFZrRasYOg
Si6E/Lj+bzcxNdRLvBrCk2vAsAFAFn4ZmO8zkWAaD520GoiGmhUXXE4caN9AcAF6NOZ1XOgeqqGI
tT7O9DzLrVDyturQpUykje23FjnPrvoCTTKwW5X7If/KQ3EUiEEyVPbLZBUllqNPdvyM2bfMxoCS
wWN5sCVg3fzG9ZQk1hMwLr4rJWN1vXr0/ZZ2/gKzY8YQgayYyIvE6zuj6992QvfiFbCZEdq64Z4U
mjES1xENB1QtoU6gPI2ekrg3av9WtCLto/aa0paba9INuR37dIdPdbr9U6zWFaXrstPelh5jEQFz
5vFIU7lbdBxCdy8LJLexSpNx0YEva7EavsMDFMjCWDLiKQ2dmgIHAtkdley1VNhn2C3M3Mz5MtZt
yVJs8JIV67W2r4bJXdkXnx52lRYAF5arL/TzLPhhMIqmTJq1oglO8Ake3uA4S7hyBXTXGoCJ5SmJ
RgHnuOx3TE8TOB1Ca7L11dlYFFGHHp/VKz54tfDsmCfMWECRbpU5XHns6kbM1YRA6X9f/jLTT4Ua
r8KyfkZFOzX71n0gk8FiLtMuySTGSc9tm4bui5mADa/4yCvkXEnO4RWWqFz3Ym7vIdbz/ZBUX8ND
fQpOPd4K2VyiZ66YZHNxTwlyDK4ieBMn22U5yHQ1CM+T/tfIEC79QooRZza2IHojpWqEVGmRAG3P
RlZgx+SSFgDHg07baYoc3wOjhaiKa7u4JGGIChBbaBlWM0Pjrkf0vOcbhDdH3W+qa6Erj2H0CEN/
EJTcx3EEfpUnzAy/pMuzdkT42US3jKADxWWnJUPeCqBs31feD7rxClY2OA5tbNLgkvNyM7vXHxi1
d5YTUc3gGYu6sOTb90/82V+7u6gyJ3z/R8VaP1M/x+BbOQb6Lhw2DJVAjf2cXKqXVKmZGoVX457a
SEe8zqgtR1VqC58M3ek82TeFtx/O/OQtS7USQHeypM59A8Bs6I5UqxI3tFYjqYqFELLQvSr8ddhW
0VdittvCryKLzLunbHP/hg7AYzWCvwWj/JPJ76AZSSwvftEN++q1EjS29VPSKHawILgOYh22AsNl
lZa/QwkDIF2YaHZBR3Oq0WVSQEqfKh4nYPLtqdYdqPdo1p7DNOCfjWbP9QMCAQ7AmQFGVCSvzF7+
UawlGBqD7pJ6d4tDznyvzHqDnYkQdc/+M1bdT8F5j1gWX9C4d8Wwd6istpYUFOgkqZ3wrVSHFpDZ
UMBXAiyhVjVg7CJ9tj69aca46VBUWZOBF6+0gZwOfbK4/YJixvTNPjjBzb/GRWq9HLDOu4AnZ0cu
JTwA0WC8qxlYnfhoI6xYTsnGE16xecIIFIPxWf7PsXy//kTbPKNU8CE/F77/VZ0coX0sL/w61n/r
mpyJvU+pM+6gHM3NBDfMxjxwqMMweS7aFzbz2rHMLE6qBEomnbnTTuIe3BBQOyClIJcEe/SJxszs
FMSweIxPEmPNeCk8zNotjEaanP4Ikkk6/wXDkprJirD17aL1B/ZhoG6ZtmMsjzaiigA8LcEwwE0b
EkQNNqz613YcfgcI45l43hgq7m4qF6YMYUTZ153JxQKV+LRh5lAAGuvF3jtPbCgl3cYgJAsKxg6V
sUrCtOqjhmey9HxjMnCo8LpP8yOa0qhXMZ+qrLrLDvR0qBLRDIqno41Y8zhlDAYsY51vMh/NN+d0
r/AMUkvHnlVhfHoLBGBidsv7fnD/ubJMvWjJi8pINZhnzQqP89riJoadwWph4ZqfAx0wMqQNklOQ
pcQnOkJXWDSS+3lbaQYLFwqOgLI9lIm+cqYoWDYNqavzWNRisQzACF1YcAD+kXjQyXU8zelHrUq3
CcHW8vyvHuwg1Dv0RpRxhABGGNQ1kZgIxZ9e6Hy7tMfNhIB3j3ilX85PlrYDLmozQOH5Iu+G8Cnr
lytCyTnYrdLg4zwTt35G1ZRGPZjpgKX4q1a/HVRGjqWdTICH0/H6woe/99UoaNSr5adLiQGcT1Ch
dFFHfRs1mzzoru/I+PBICZ9LFWI15CFjp59tFglclvS1/9iiXZPvZHxuTpcnR2PsXzkhTrgxcbBp
u4yyh2Qh3LQjNijNv7/5k75Gy3UhgpizrBHz4wKqYe8oVNtWVhKdhUovSQDMut49kDgV8E6MrtHm
ndjNUl2Vi8Lb7d1gLBNV23YgpS6oSncUuMS6d1BrbgTiFbG4OTB1447W06mYU9t/saXjgAoPmL/M
VnfjgBAyHQhvJLaqhy3VsUesEKrkJCCTon5aQstUG8rMWI/UyskiB1ZFm4vvsPv9wYEoUdpbEvVK
Jknwhttc2rd3I+xkdi9pKiRe5SfFG3dxqxAfTyU17BAziRjgij8gp0OHSZa2xjLd7QAh+UX8a6Ac
hX/yfj0Q5GByfP+/y3lnmcpJ0TEDUPtt4RwB+/DxPICMu/2Kq4i+T5j2jN1mi+5izlFrGKOeWctL
mEmsSvLe34Kll3AgSBnEcUxsRG6eivvSzoWHRsnxEI/Hv606sJ3jmgfKFhW3ha/h5jlq18Z2aIK6
mmwzjo/ULdaXZ3DGL7PwYdwdc5zzbroTKWBX4xLatuH+Wa6/NAXWVo0R/nrX37Bz/tvyQ8lZhCmw
oUpa29sYPoygzrONP1pX1Z24LnmEtJdFbCeL8Rkzx42N8RbLtxSu72509lRwrgga7iZ34PD2IUnh
ejiyLT3FYaFNXAeDxpLlrv8AvBky0l/dDDP02JhlSKO48eoVM8ncjXinIWww0jYMGXFElkd8QCkq
sXlBEmKp2NDQvjdnUZB3m/VJS8AHIEiCbY6fjyHx/LIMlFBaA7SJvy4FPu/2mF0QR/Bk0E9kkDc9
SNf7K1+a1jbXe+ohtma5q1ZnYUr4ZmphaLNVTp31Akh87GAhMHnap7ZnPn3xO6Hv4ogi5Y7Ml4jN
bZHAA+1feFJxpHPpzPacuaTARlqq3GvGa2+GmmF6EcRvMm1jAFMG5rJv7mu300zmnVwpF+JNdzSt
j5TfgoGLHQiasobHVB3O81YjjqymsgHqESptvBRKxc9FHwhRxw0ezqnqGt18lCzuiF/qFJsm5z4J
DHiCR60uYDX1Lnp8nR2fU40tzZuvikTkyb3H7B4gM2hA/62tRVR91lOKitnvuoElWv5RGLrZ9hEj
yZVHy2Eegn2BGpOt2Pn7/GKpXmdooveCgEI93m6rVUwyn67vUHwLfZoZT71agUOr/Pl2kHSO4SIk
2S/Iwx8Ofvv8NF8jFduKdf6K92oDqDNpt8yoN8dsMALp2rVYUEVSJAWrqXTakV7l5JWfFJ9H8nk6
IqpuXp1+ZPuNy0LHiQhE5FOp5Y+CJAhHu1enNhynsqnrKhY/qiJiKA3yFG3rRPlJ78mtWwhv/E7T
8mZB1R2L3PxEz2zmIE32sxsOr6ZUzcD4eZgYqWTJjatxhYKaUJybqugyfuC+UdylxJOO/NqNwyH8
gmrvrVWyH5eJo242HwoJuL9PHnMn1EzgVndAVZC94/ODXqQL6Me031CXeltgyo/LAesVk2HY2viB
jpfify8gWVct7B1VhESgbhGGAJsMv3nvWMe9KfFvqfJ4KUetYcOzP2EmKj3NudnitoGQZFAVtiPQ
wVMVOIIEkBpkKWwr065qkjkqtk+6xPzw9b1rZ+83tpTMUEAzEI5UTss4geBYvKgnhkZT4oN5/saR
BFdzfwyyrK8du8AdBL6OedRbQixwchvF8AqHbQZChAoGVL5dvhU85/GavnN55IBdH9NunmE7sA/u
XV4WNQ1Wjl9/bcVVZ1ak2Zvyz/TF1OnprTmApXXjklDsnwCBqC/c6E7ikn+LspQ2IYKvTmH6W4fE
EiWtRZbr6kop4jEWfRZdQp29lQzilRMJQexinPuDhYp2u/TWqzUxOw80FGvMt+KRc98uvbx1qMqh
qalNjrf1D+Wyaxv/LxSqPHBMEAIhfF+DegqSAUQTcYBQYr+ZjzMyX8iXFDAHSOxutOfkSlf5aLxD
MvbEdtvdUJTDZIIco9Sj05R6qYn6XezCIGv/cgtrlsdz7uba232+tt8LPQGGE0vtLc2FNZjuldO1
eD5Jo88PGuerJBNGJTQnQCo9EwwB41P2uQX3I88pn8jmGgpiUnCdmHODlW4NUoLYq+eBj3Cr7U8J
yTDrH/zbUUGifhA6QOOLEAqzBWdF9Eq8nZQ64uF7XtIDTpEiS0BXZ/+Jq/mBb7T6cwNtql5tiDdT
be0vC/hOEyW61M0D6IHDXZYAk7hzMmLaHyp1QFdlc+Y0wKZZgMIgkJe3Y7RI+uFLdZf6Yyq89iy6
RcEdw02kEVkDzDJxd1DPlj4WrJP5WBPRJGJiB3eZtd9AioWol1wP8iXVk42gfitMkNou6WhEWRVw
OlKpGe5lea07teI8NOODtxIisApwz6uedeF2srNLCNiEPFKIvTrLxEjHVFxPp5jOds1jY8ywkomd
/0BskfQlDPcoMBixr4jVioFkEbxx48M2hAe1don2kmG6REfzsAyOYyIOiaDMEY1RY8ukMVu+1S4v
Te8K2MbiSOLtk6C4Ghm0gmgsBovJueTWl0SkRIxKzOsmrBr0hMYA0MAphIuoKw58u2wZ6mJvsCJP
aEVRYdHc+sHHWSB+6V11UuLr3pgUqfWV2dCO/IBoQEt5oURgRNs/N1nr0suVfMqN6Wd0niODoDQ7
mG/XAQ30Bi+9XVlM1oFsN8KTuVOXAirnJp6X5rLd0422dUesRtA+x51W4SQHf3vgPHp9GAL+HqJP
pp6jiINYg0/ky/uvKN3HLco8qONsDHmu0v6X1mv4Raof833ECK4/DeYkY3OtlEGQF68qJSHD8gyx
DM3ebKHcL6cSuF1WZtpb8GmqKZ1WAz015oGrXKhUhBltziW6wXX9BClCZciBnMdOrLJx6m9AiPhs
l7Pb+3lVh57JRizy8MHlcOQVOUS706IqjU8j6w2vU0Zp9UGGl/XdqYJIzMeCy6WEkOsWFLI+WA+u
GrGP+HA6pTgKmkAcu0dO5ii+24lu/KFk4YzcRa4BfjVEL8/usRwQBJGzNO3EVZdSN2LSk5hnYvWS
rUJ1M7f1g5p/RrTgnRyA4Es+2yvENUYVUvvLR5n50MPpHD/HI7InZ2krPDeVpYUynPZaVzzf0WOS
GiIeJIAuy2tzHoPM7OUiDqEUQwNmK0GrLuNTF3+AdsoHfyAVn4PXqj96/4D5zAyYqmGeCkBWW+B0
ISkV/AHcYDK3utdPPD2vCad9xv0HdPYZ35oTZGNxXVY4ybv8JsCGPDYwZEb5DlUIVIq0BtEUOwo8
AIsEvFqDsXfSYsWN6KrBE2ykdc41zb6pam/I5qUaekcuyTLVdYyo3eeIvva+BdVDQMQggU2qivvH
sV7Im7gmPWeBunkvYVA/xk2X7avNszj6m7tyqp3XVgnzagPORyTnziSNl1F8c77H+fhC6gH9lQ3G
RxRKttH9n2+8mgIIUJTm2Ztd2ySXeSuJ1HAZx+FENT1qe9zRn0grfsB6ngs3nop1no7/AI/9sqjV
DXmP/mQhQ9HL8mkWOGX3h2yoS1//LZzZp8gwiUm56woTEdSAH8gY3ljl1iS6rjI54oYaHq0zQmM/
LTK0uaR1CG9DNQ6Gkbin78m2ggN8OqQFN1TH1i/CfYN69uWIPJ73z/BfE2UF0VfZ1xAR4gdweFPm
KuMlkAFTM/+EELiwoAJyHOulrthNU0gaf3VveuwgURqRbAc8m/UmOgdxJ9iHBpX8XtvDjnMzVmv8
Tz29v9H5YUWwO6Qj7EdirRG6Z6sdYTC4C+/GlaCOU2q0NipRGtYM9cn0Gj4Fv810pM4f2OZFN1EI
t5BXEJS3Yj3Qraw830i2dYGMKNZOl/thNjYYqemHBwayajO0DApwxT2O1ceBQK4EHnQ0xZ6ub7Ef
N/eCgtjHwBUkKsPanqFFlaNK85rYkwHQmFQSqhoGumWyydOvNuvdrbNMggSIAAsOiol8L6bDEFGx
f1PR7sxDaJGZrTfTKEmva0XTdWcLrYNfWoKOpmzCpBLVl3yB1B42+bMO6TmvVbiPdKThleQH68bz
nPKsi/QWe3VTjVxAcGZXK28sSU0+NEc3J71ddB6EDuhIcyYbbdCd0g0zN4+8DpLnSGrR1vjRY842
Q+Ch2tvmWtldjUTUJh2Qbn+f+G9u62AshtMmtSki97d3G2RMutrTOA6Ggm8ar1CxBigoDZ6zRGK2
k5Lhr4FA1w35k/C7x/EC2ZJT6wPLaZss2OXHxFutGZtsfU3iSoGagfN/nOa3UX8l62yYXL5ISbia
s9llmrU8EvvWBaAZeBbJSvsdLPHYV20C0dw3CLO/RunSm//ZfTf/798gE8PmbLW1LPqa9TBvSaFa
0INmv4RD6c8eKTWPKRU7ixqFL0K//zzZmHXIMrMnF3JSKXZC7v/01syGAShlx/QrBNFv1g1vX8U4
4giWqVLiQnvhqSuhoQBJiif9BS0da2X7LcB6dzAeLs2yVSXQzrYrTKjRDHxHmof7vzg01ca/hafS
zcjMcQIL0WVm/XDuSj+a7XTZbn/PLTV4QXXxKsdXeg7JNPLrYdr7MOd3rTUZuD+kUoJFt/qTmSvj
aBxGo/a8hpPtO1D7zkrJMWbsbqnWEfCF8GdKU1PE2WgBF5HRP2ALK8uhm0vRCt/bHT15XqaCpvTv
6aa6CzbNr3j9vGH5Oqz8M07rYwHzPnpDKfrjn6uwgueUdnTG97dkBZJWKQ83Y1PHH/G3Ayn6kxIS
MfMR97T1o9aMG95bS/YZ2gaRrITQLlFraueG2TIg0Rga/X0seJpFxGMzZ60mzK79/uvJ8RvxoiEf
ZamQmk+OBecPYyfSnh8MDtjQneywWUafSx7njE1ykVGBkbp9mRGm92JSxzTzCcKRWaxDDv+9zL/J
hmKP2SYVfaPyxL7VtWf4hhIiLE4E6xVss2dSUK3k09loncZH8eISoDklMuV26TQIw9mU82yJNwfY
sr1H3hSIF0sVvMjCBUI0pnIGmXATXlxTBFV7tu21tOqEIK8YDMJ4yjxDlhK4/mgH7cmI+LFE3mR5
4hH4NGBZcqEoRbxGqKUya635HDGlRs5Uz+IQP/HycB/3X57858eiXVmNzdf1mHgeqa1WIaGlgRJL
P6MvC8m2YamXEXEe5Z7m8IFXlAGQrODXNBNPKl2KM0gRb1v4xBIBWQkcYfnS067oL8tnBXpZTNE9
i5c27jpJKqBvFBW8j4mqER/VXkKh39eTZuTODirq2fsIlPtZKG8ZswdG8pvlj9f2vM43ac0rOtGH
oh0LRWyh/rG/+pzM6pvbjT79ay0cnzkZcfR7zM0sulE4defUdznx0jBqub+/vNrEgUdV1fF50Cqi
gow6zJ/V623INVoM866mtDhXz0Q+kJwDwCzsBchf9IXPp2J9Dk86RLziM/t+vadlkb82EBmFbu16
k+xxxY2ixwePCMIadtWZERuztptopwljf6Sy46IBAz+abBU1aPpWCGHyH7W4Gr5GVU48srrxihzU
Obt1JIsawginaKWgLVCdB1roghL1DkIcv5X0LrJaMpGXb2I73Ehvgw6VqSjSM2/+Uuy6MXuuSETx
kOpEH1/8L5iyY1w/J37z8NN72GPAmDifX9/JJ3a7gylyqfJaDGHenVQ4t2eHe5su08pV/CunveOW
lkx+XOw2sB0B+WvNBbzFZrZgy1GjoP4VYAiRxvan1uEoMG6yy5HNrCp3EFGsMs4Yt5TqSwRSRpAP
8iSKEs2EeYX5mMHOQNXIbfJ0JrLD8KLkjyhrEnQF54hcCgLWPjm+jcM4lVyTQzjAmOTGt5AJF81S
4Qbv3HCK2iWWIJyjyNf+iut5cZ7yvO7FWfl+14B0KmEqhH637Nsmc8Y2I/MwhkTIAR0McAllsevA
26LkFw8eMZAnPWvYv8iZMOQ8lG/B0Lk0WbZCsVAJftAh8vyA5PJvOqNq3ZZE596St1kG6HP1XV9l
6FqAL4IrrXAZLTI4xT2sF9psTs2NtxTrYYAQ/oO6igXeSxIE2RFaDWgirL519oBndHrDHURlOeOV
mXsMkSnWgqXm2asBk8Of9yatj0/O4tomtiJgnSeyUOlvminK6FtZOcvOr34STYgriIKAyYP5ObVT
Qaa0Y6LxVDWKCUqRaDE2UAQdYRs8h70uiJH5CZdYPXsMpI4iK8+dXHbVu7Ih6gUn0DTmeVfk4V66
k7HLr5TLpVbZmx/03KglDb3BCQm3CsxLTAlgWSaMInWnx0DwHEPoDsnWbrDuJJ0h2Kc7YDNLMoz9
kt6/GhVVXlRSapwkw97R3HKXqwIuM9iCs3L1VUTkL0kidHbIt4IDRcBHUsCUPPKmLtwrYBYA5smp
DohPv2Bla7u8tdSv+aCOWxvEqwkdi7q17l01jVWcO8/3r2MORaTLqnFXVEO4V6x27pzoqF+8+jMU
7PASQJKOdC+0gRMw/GK57B73MmsNVGRAhHm8308qsrAkjFtMO0EjRmP1Gnrss+Rvc5cNseXdeKHS
1cPM3+sduQSz9IGS37Vrrfl2WduNyHaPbN6cVnFyE+SQOGnCuKhCtJgkfz01OpVPGZ7G3NvkAnhx
/z8BBoZqddx14e3HoJbpu2jdP2kVzr1UKBJeZxgaMH4SRqZxlqIkR3902XAV1LtHpTsuaW0UW0+7
xvCV4WckG7TLqrXDK7bW/WnEpYD3rzPPPzOdkUKVN4rTaLbVB9Om8DbgPjJDuoKp72SlXeDoQl/7
D7QY7IggMOnwciUW8hGZyk4HKGw5QDrFGsCDoxl7oKijPamkk1jmRlpdxoHpdHSKPgqM6DWCqOWb
wZwXxFNvveM1Qs4HpYZdjpGi3l+zf9LfhUIrixdKqb9IuBfR89s/Pfz5wjD3ZypCHkq3VzgRxzNa
MNPWYAAOtIxQadBU3Jr2O8W/8qRqcxpnuC3auwe6YAicJTHxfTEb+fEpm9GiKnM+RTPaUWvKHBH+
GlGc/xBsDUVdofEdosJ+yWKhc+PzGsFT8hx4Bbo1Iy6M4GjIqNSVOMe88fU75kUOjhG6J5PGNKIL
UDPJR7J6XPYPPjjtmXX5sOihUZsRcdge/+gB4R7mLh7YpEmsxX0BQReUO7ha0J2mH+bq+s7tdERk
GbMc7++NIaCXRF+fwVLWl8bjLF9T+S/PbgpG4/40QVgj1xIhNiO6N7JWvS4X5hbsQ1T34TOvUjok
Pf1/0bpJi6RR1WabdBANO17VXNU/CQKiFaDDAdeeudtSw9fCjBqkb0N1baPFMXXqZBTRBhStZ1Rj
ydFT4KboXAE/43JyLxeqQWzxo0fAIAJ1zLL7rPFs27EcpkNLKg5SksLbfrJBAGgpSAsisUiSd7AF
y7lBR46p2u5Ij3RpUSI9FEsBBbXnWWfPOqbnJxAicDvPTjolx98HwjzelIbd8rb9N0EdQkRWYJKJ
1J5GOhifpU/22hbCjYX4hrWExRGmqfjJ3SfUsLTYYjt045xGNSPrKua42BSVai4YdBqUXItVOelr
LpzQmuP7hCf4bqhqrgICCwEGCRX3fGYpecEb+lSQFzfPpF2DME7+kT+0syOV5LjQ0bv//Zfw4bFh
m4bLYihdiTRs8QnlIpfEatk6eYDj2S9XeB4WDqKCWG6UOzQkxiE1pMMayGE87XZDUAY4H+UnC+ov
LX15r+GRUWzRlOtEtyQJEi2vtsldkxjphMMGDQhgRSLbuTwhzXybtOo6geWHVfxCDUKiBeazoNGD
k1v9WAlIlogQrHssm+R5NtqJFSwHy8pxavnvIiTn7vglCmVwrA6MrrcqKf65ODwS6Psh2sUMnuti
vof2HmdcXhYdP6ahiMryZI+XumTsiEp1IhV1V2LSAueM9b0QdXr9QilHVRIRV1ppASgt+ZMiE3nS
Onh68/6QEgol11B8h0j7e18HpV40Zae8WID/EgntWQneYUYViHuE5W/92KdRKjuY1ef4Mjyp9KaZ
6CMja8hMJiojkwJOAaKXOy5PMaDoeik8XIGwT1+LzatFBO8uUG1bigWUmKxeqfdpzxzH9Wz8mRzc
lCmTcGk3tx6vbDlNduriU1UU5AoVLYLxYRn5+Bi42a62a5YXSUq1iNe34+2jHOYnOb4wq2zpVCt0
h0iew1IOIA4g8MyUXwlHmPtBDBPZ9LvXQa/GkmeaMvAaHJBMPwNT7+kKvyyot5tHtg4mZH4bAcw/
F6/T69tewMlc7CXgZGYSQJeKX/hP6sXXj+xpBJTW/UwJo3DSgwnuSc9Yo/nR3FXVIjK6smY+WPMr
Dnq7G0M1xsuTHLaWbxmXcOj3Zn+lUrXxRMb5fDhNFSvwTtqsF7CJrkyms3T0QoD1khZrpJ6MCAcF
clarYzStAKyEJUqyxryFnk4WhEuo/onEtJ2Z6qPVqi2tLC6/RZ1F67yF9isPVJWKlg+qck2WpFYQ
GEBLjVRJEHuV71emfhgJ+ZWJI9RWjhLsu+BmXsM4P9gZ2eH/gvN8n50F9+iW6ap8mptNGMEiMqf8
u8iCYLx7k9hcnUNO2FrNG1bMfvIFkVAtXAvWOL+k3GgX8iRgBoGcJ3zDKY1qufcl6gb7tp+Ni0yN
DPwrBCtKRFXnT0AaaRLR/z4grX0Z8vPb6YJJrzK9ku2kdTYLFzNqg3k3mAMSoGgDWPfUdUInZ7cE
3YK+nD6dQPBmqPEntoMfvP95AdR2zEqhhmLPJT2WtyO3gTHZc07Wci6Pww9UVm8xOUiCLc+2L4u+
ljIxgPlfOx1GzCB7jrEzBXG3hbX+Z4XAlAQnVphjVP3xxkEw0ctMPxus8iti85jP53QWjmEHWCvE
l6XtOt3T2TcsNfYw2vU62Y47kjUweHx67ARYBGNlU2Q4ZGe1DR4MvbF7pA9+C3dcN+L8kpyhz8HY
1OmSA3wdN5RHU6AF3j+kdlsog562MnvHj5PxtHZYXAYKCrdBAqdRn6NA53TBqdfi5kVqELBP6Fgn
F2HpeJIQttC0WiPT3vMB/4Az3yGB4OZ1vZm1fkA9lolNuCvLe6UU84Z73vOoYZNyVbLz6eH22zjj
x2XYHdf37S0RNQGtwQt2I9twTyKSjETD7Pe1GhgAoj6GVMbGIYJSc389pub7ha1Rq9gT1B2BplV5
fZGDz6/ZFUr0VVNBatdq7klHcxZ+3C+Y7IVW9/pYYt8QGJAdOLHGazMkRDcBLpDp5HmtOpMX0q4j
FEEJTFsHVHX1b/3klDVjUES6ZDdv0pN3qhnQW94GycfaY2imnhBhiWFzftbVnM8SWRg/+eHpHXtI
vU4p4SKU+13fBk9zhoQVuJTrmfn+m4hIXVsLtTe7yUYCKluSuCm0XskBBjcBD43/gbs5S1CtOue6
TMu4pgYgpjesrlPKeztuDf8QHODltVcE6/2S9PKXVGVyn/8/yZFnn2woZd9upN91KtY4UfFo2iC5
16RBukVa3KX7hsxG+WkXQQvonoLMnrhNtIMcGHJL63hsS3JCb8V16bDgh575ER0GrCU4qnH8uBdX
qSbcQ10b2+nyYQ3pvjSDM8C2eiqM3cRfOeIzNKEeC4sBjmN4nWE7NHjIfbmqUYYwa3BBw+e81Yfe
QeLS8LQMpi0EH61SzbPaHsZmqs54XvZrKGpEqZ6fkU4PVlY9VoubGBkVSt7wQnexsstD51l9nmjQ
HZJZXhPjW94nvFGkQzLCWm9H7vP+q04NX0/s71lV+Df295QBD4hL5dNlITyB0lpVz/NXMYHhLlex
ciziw2x0VYEgas1AyRkrPrMNcK3tCGDKCu6Hf+7hxOGttOIKRusu7kMYRde0ADGwG44j+1Shyyrb
1ouRWzc1h99y3KFeLPqX2n0uVA4L8x8pcvThiXkVBo8YM+INgPGS1bytAOISqnoyE5BdTIxVUT9H
9h+hppIKeLc96VcoO6H8YlnhfBNRhqPLBUhIkX5cFgcFnWM4NM0zzQYLpY8en4jfakhdwyG8I12l
kne7CJkOOSxdWmBbBssC8okiPQlnKo+/8Cq39BtWktzx6Anj8w/8TB0W+SbKMAU/Hy3v2N4kKvod
ql5k52MFx0WRTvqepJ4GFrA6+Zb8y/efr87U19KQeRmV+9lGU/+N4m3lX2rVW7n0Ixqar1RMXRu7
88RQrtzivv5Yay3VnRUUp2pupNhVRwEE/aCNGuaaRszYWow7WCCQvuETO+394NAWF+Fp22h+DcQE
FhwwCAIURzSvq7QUYZcSHQzYPC3Y6cny7Weti8K6Jck2iwTOgssg4dzyvcwbxKVDEmlmGnfL2Wtu
x+uSHXHs1SLZ/jl+VvSWR0Z4Txn3XoSv20Ed6RSTAFhxohmgKa6rH9yk32mBUDvvjFBjbuMzJnVP
RkpG74gvHHuC+xM6QTV4QWy1ErKDYrTJe8RrB1/MyeCVJNid/RGj3SP7uk3hIl5Yk/k5e8C/54dH
TpSjqdGWX13Qu0oG8c/4V6Ih42EdZ3n6MhhJ5e4H5G7HIPzBNjdBHbEipw9MgxwXT30nfYFKYD/O
JLozWt1O8fMIcttFv6aIMejbdWWyX+YQjZjv+WXF5qEGdvz3v1Jt0TbVCy1axFcviwzdtWV1+bK+
Uwy8yGhzW6AkyTbDehg51tV1f8xPL2eShJzGMAT+1HYLgrZyb+2LuD8X4Zs0YoJ3onbiJFz8NiCV
rkktnD/EDR4hlnxlwNlSJGGQAqhumL1oRdu/wIVate7s5MVYaOtvzR5Id2RZ4ew2OmEzTKnlshfO
GwZsDnEtUjorMxbY/0zg+0qt2mspHmAn183tzXJhsglmic4UE4y+3joar6Ug2IHCKbwYLM4pS/8W
vu7cwBkKJbCyzI98RZsCmU85FXfT7Tu7ROveqEbj4DT/mM29D7dPBBILmVfMfimatmIzIqXyrfsD
oSXUpb1AYG0Ng6VUk0OH8ilcp55awrnp/MroC+pAdGCd2pyY1GrvogJXOnvcfXnbhUfcPc/JrwDR
GzcO8xXOXJ3qMxSfehbzi4LZwKWGlfjiHYL1Qo+50LpWRosgLiEAlvohDQgiRQfVRopUOjQpJr4H
hqbE69rF1t7Nz1nEPc+1Hp+A1HyHObLG6az9d5ZlR8ZZUL457aorhS6YmdxrN+G8awXgv+oII2Vd
5rB8jUr24HOxug/hlmQwxn/KDB10pNDDccCIwLjP7K7Z7XbLoedTxaW8OwKUN9ZCG/ewTfji53cR
aKGvnmx/j+MVIp8+zSqjsI+znlNGWN3m/CsasAYdDBQjfwDPdGF38dWDb1A7tAmpCIx5IHrNLVM8
OSMcHV4LQqzeWkWJSb+shtDAtoKsC8HDAxD83avx58PhQ7eyCGH1jO2BwtLqwKH8LZvw2qDbcuGB
DgrZsX/L9bANj0vFQoDkrow40AMKdtf57dOKa6DRfGB+91DEbpQwn89FVE92qZAAdd5pFlYqilP2
LwVA65BeuxhU/UVNonMxfVcF8xE5rPrJNeV8oojZxsxkggxUOg3RIN/xfkxXFXbEkgTjZng32cAX
beugvSCo77tcaVUa6COkMCc4Vyw4YHG79DNmn97H8OU9zq0CdU6kOziGkemCNR3t5ivNieLzBUmB
b1p3dgReFpdSUycyekAJ5D/Lcp6NgKYV6XKD/PuOgMWBIZuSP+fnEC5xETvx35tL5ObK7C3rfNME
DOXA64lydRslHNHCfgkD770vjFZJeHEYblCwAA6VnfxMbOwEzZ4mhN/YFlkMvYMSa9q6dByiV949
ZGmVj08Pf8CYTsMwpNvIQzhHFPqUMNqN87bAOE5dUSJRZrrISkC9eB6/ZVao7DwldRvYDRVO1/hE
0hAEiGhtI3znnztbxgiDLrJmmT2k7LTkHXA1HSA0AczNaMItS3MTwMuYxZ3q1gJ2Hw6Vhgy1XESb
+GAO2BdTtlYYXXFMoziYJY24zIlMpIaC2fcO18wxsCpzh3MEVUeltj0YUs45jcagKmpbPZP2TkE/
UELU4w/QqeP/pu68ywzpvrvfM8voOOS0O7y0cJbUJOUYbUHDQAfA7jTQxylxkFcqgMjvjDJ7uOb8
E//m1FVDMisQvJFMnPzaSJAFmbc10jcf45xL4Hl1gRNyH2L4vgG74y2jE56AB+NMNVm7UE38IRhk
IuIto4x/aESrcfr30Chbnnkph0nh5w2fu8Se+pX74Z0o6Yejh7emHLUD7RnGkxf8aHEcbGKJl+jf
avJcitfqh3TJleEEXWLiMH/cOAyADr3h+kVKzJzHTBF8oJB9P3l7PBHfpTuo0dIu2Dxf3//m5IOe
3EVQZDodBxCihtdpvFu2xIHIFIizchC7pfPQZkCyFnAND0n8O2EJG+66VQ4H3jPTTPUYo82IEXvV
klaFNMmyXBoMmXM45xlV7e2QtM9EnjTaitoMmLPZO3eR03n5EoNgog+EOnT9J06AjtmFZ3FiDvIo
HfDnZdJ6Pub2Czd2Nn0FA9V1YpYVfzEGSQS/S7Ipzs4KIiC/2IaKCKEjdRoAS4IiEjH4wpYE3cDq
jNp1UUIzqHXBwb4Opb2TpGq/RjrI/eFSd2p3XtqWouHgTveb7g/kHepRusAhPu6sGLFmubEgGmq6
+i8zyjwok4T54fHE4rn1xVLoUo2FK4is5uxQK9szx33shRD+30ocFHoVHHb8A1LZLdN1yibyE2Io
/R038THXvDJdg8XQhoL4fbByRkQ5gZ0Vp+NPhHIlrNrtBAQqB6L0gCmWO8bHk1bnFCVXtYb2pyON
HdFbd8agnwiXLuZ1eAmeTLQZerZ0J+t/jyZcEPp3JhiaZpJjkQMH2R0B7F4GKA1Nf79gZ0B9bBAF
qVThFzcAMdBVZd3LoXDSY1J3pQg656r5mckuZLVDCOY2l9luFJMN4vHWwNiadC62IhUARaD61W0W
fneUR5ZlOZhY475zUKrGwfzfnh/p9r7BSjw4g/n/yTNhJDo63SYusDJtyQwlO3KsXIUmon242TGW
z0Edi+2G1pvWb2pdnxG0NRPvH+/xedhuQoNHsLFB5709f9T0uT/eKTJTE4BRj53rYQBauyOkHpN7
6pddmWb6nHkGMk6KCqepWPNyNQCHfJUOa3CevReQ+QgjOQYKLMTp+u86F+fWxJBAPVFcwZEGnR0A
wZCU8ETieSc4xD+uqYqJZopmjMg6hcOON1B2LJaOP9N0jwyYmfOXKTu24zyQlqJOIBwV8bCD0JfX
VnRfZ/3LimUzO8HSTgKAcsdTHxVo0w1aQqdCDDXm5axqrRVFNDQ4GbgaGMZjJ30EO0X/lqgDm2T2
yny4Bnz5DvBHlDeMFPLvNUZdNYLbOJNp6qEuI9rIi3+NU1Uo4BrWh4xCal4TZSG9dyMWo/J62dSb
PaDDeoIlAmftZBaIHv0kF1S/Mx55n0ksAPz1u0KdRg1FTbtjiUOGQFySgYi/2LvXO2DYYl4SVQxp
2/JXsjoYjBsVNHX0k3N9icl+oWCdefmxLmKtZkMQxSJ6PhohhDBCDxdWJrCdumxrT3TLm0z8R3pr
Q61D6OJFCm43dMUEwA+FqOfRMlZZCldAcNyZQ69fnqtS7vr3wnIe2GuJ1SdmPgSQdTbQ55r9oxol
RH1Mq7wVfpjKfSv4VuSVlXXyMwicgME1MqI1zl0yfURKSCl85CntAHcTqv+PFwbegTdrhmnmtyWo
IBhtdE3zr8dEbGIfSvf8Sb57gB4viZeJWmo2EgWzytw02b/pTnnOOLwUPxPJZRyNwEIIOFxYNWWH
qGrbAfWg74jL4CCEG73/CzJAEfGOLO5U6rmX0x2x3Hu6tn+6rg1HYgjSaJTN0ZOyAFXQd16bb1p3
bu9EpBeyGuclGHLylfOv7mfgAUcJv/8Xd7Y51z8uO7GOx0MxelbhRSpOAdPadHgZVBWpL8iD/9+P
OS0rLm1DMZWyV8s9JyRczs4iYtP+5yvE3azQa9bAtwGquxpqVgfAOpLULBv/FTlHxrxodmB1V3Fh
94o1pgvJYuQUJSE9Os8fOgtUF/EUFAwsx0fRlMXMjzhn9QVugTBmA434338kKYxjeLr9knV04NNH
7969sdDsco09OL7yyeN/bbQ5BO32Rd8INTbIUSyT4XNvSxU/lRRU3B/+u+gVxpXycNnK/eRux8yy
O0xGOL+ZvPWAwypFcM775UDOF3Gw9cYAT5iXzw8uP5WeCSsI7rtCX8McLl/7S2MkixqS8g7NrLmD
Oj9S+qeme0EEGqBe9EuQ1Yqx5u2Pi0YiihuRj1kRC2UL9Z0N8FFRyF38iNtlMjiM16BEb3SQbWgH
DyARdrp2u6ijIBRxNf1lObM9IKr7b2Zz9EuqKRuMvH79mytvnzQs/lnMpZ67s0hBFC/WUbSRqJ7o
SPBVakeRvRDA161JswWBXBT8KIquqjDHALwtnum8ii0UJNWXqi6J/1XETDRXZ5y3hpSMJpgLvH5H
MdbgQBWVtYEH+tx61dcUmZ9Xt26mzY7JJVRHr3WKyt6Nw1vSKtab3ktSihDKmzU8lQWQguKnGT3Q
FivTS5VYmhE8wpVrKk1OpOgum7aLjyt/HMd1dZ/s1+bc8dOxptuBkxooQq7vuf1sHqAWgube4tqr
w1ZMpbLQLXcFWlQDmaIUCvMrRlPa+btdHRFCHqK5EKTGGm0rZDHBKlTMaVq1QRTtadxdVYhZovwx
L1wzgVABiSlwS9XAvCxW7Yy/H3kFdPxmCTGICU9WVGUKJ5PmqxEmSIh4nokBCRtd94luOs0vfMmu
nko7pGJD0BLOD8B7a7rOYQdqqABC9zQ3jExV8IzYr5MVCaZuBLu37oVmZEJnUlUkm9Bg9hp1DW71
dTkTjKW7JssCIkYoRF0depTR9k+qfE+9F+Zde71j9m1N5ISjZXnCwUqEIDNJwpy8KN7mBMs/90Ik
tzdToaQ8BUYgi3w+oVLAinUh82nM6uYoyGmK5EnicUSrZFC/lPi92GNzyMkSHB6w5ZYnYdabsvT1
dlgN47xWEhDOWoa4sJdH+lSdDUCBp9aNH0KvLYZMX8kkBH8nE8ohYyI4D0fs1FviKAP0OseMS0Wl
3fJ3zQHoQo8cjry0/Rt90TWBxFlWEjZ8jyxk9QHkGMMcB6kkIEtnabkNGwu1T0pl8nLq4pPBAhvQ
8h86mLsO4wsVK/xQbuiJ46rz60G+LYiCZdBjy23BHbaXAErPZRyajAyHU7kR+ozJDXCCHp9226mN
mshRM3tOUu/pZToCQZdJuHgjNODnOrViBBPyf0AyV/y+mBskyZY/O1XwkDeWNmLshPD/B19QnYem
x3vTk/2Sm6DPFCaSQfT1Xq+7IJ4BoPjgh/lvOL/twZzTJXCMVEOAdJ6uhLSRsBRTVZeLTedMgUFO
256Z+rylMSNvCpQycmvL/qeXL/HWHbdiA9p11z5YMCAA2tHJMh1tZkK9K1NsxFDjKeG3PD0jvRiy
a3M9VYT6X9ROqYPbxsPR5CFlPI8vW/u2eLRoCMuvdv6ti8jEvmRUIhyTr03o2X03WU9RU68kKwTR
wC0UGkET7yT8hV7a6DtQqP2jN6cMnqteGI7vrdIstUBQYKAriTDgs4KGTtz9nLOdXuSNS2UEaGWS
yIOW5Q9oBzjd9xvruLs7mcofL6T8xkq2KnCMIV2wof0wx4NMrIM4CH3PxxL4sGn8XcXpWHIDkxv0
lNtRu07tr6PAKShXGiYnR0sVAPhK0UO/q9R8kheKs7VC9d5mqxCBDa8l5V/9dNjK4Iuqs9Ldnorc
c0zfQMB9S1HIAk1HWzj+gSFCObxHk64cIeDWD0c38KoSp6bXt1gqEs9lRecgfBXzoMh862GGH9Va
YSBHK7poyOe0rBmPTmwtngyj1mI7/qmY94kob/dmeSZYmLZaSQItIrHVTcXWIaGl2EQTpMycwkLS
TwLIGHEgblY/nC45iFmqtMIZ5/iRrnVf9ERgZtl/VcZ4v6ZT822S14o3gDMZj3LUO+mz0R6ZeqGn
1x+aEstct5rY4HzyYY6hH6EZhxh4G1F+uqEwQfF7cHm4BVQv+QXWV5Rt5vtLdZXlyyLcz++wdN6M
+//VEfGluzNF5PXwS4DZknDBi7XIbVhU4XSB3QHhT1Lp//ve+6rLZLxEDs2Vwc7582SD0mXe8dyK
XZjAk4wZ2n+Ht7VhvDHWtZ+wheW7QyjB0Lf3XRYAGzaJmnfUIKvn8h/V6BPLsStdDazyxdVlYxNr
KA1j4RPLqBplJrkfQ86WqOXtbFpNVtNr6Mo0DQUPMYX0nF+0fWa0Fu8CE8SIMFXNbcSzsRlm0z+9
QdG9p37nBbBK4dc02P2gFUiqh8iOAE+MtUHLVWpJncthOssoADnTm8IKzAutc8+J4Ont8jE6bb4v
U3AZvDojGehMQygqr9Ycy/NA74QXHdy5Ab/SOMlF9y/jwMhmnmmdZXZhwocp0SFOave5FJTedlet
6sw5/qPSc7l0PhZBz0v5fG56KFaeBAdJvJj/eNJW6HTwDwUegPf+cZrNrJHBVGLZGVhGmTxmL6wf
bxvBp12yZUwaVbdpdDImKYLtQnoP4NSbTD7qNQ6B9jk12TurAhnap+U0HjpUepPy/gFaR2FGMcpm
IvOYwXX11Hw3i4ucN5ozUmbymTJ1t7WW1jtCaUkbQVERr+PW2CuWwlM/+Y/BQYwAZBwlYTQCbWUy
M+bFBo7UxFkJDqKuP5uMKP3HcDqpk+aE3vPbnHA4PLy1Lnw6EBCvAy39UOyTigm9eud68sFbWhwK
lCPiguGs+OeAJmE6L7XidpASV1vKjmEk47w7x9oeXBLL0d2sMwVBH1MOLN76aW7Fj3xOaUt8XZwv
AgsfsQPsWG735Dpo6uHE//nmj4XxsiETyraThyOrruQBJoeoRBCEnCafeGw18VFiV/gIlOm1ZCx7
OLgCaFpd/aOTkmtgXjhY0PFFe2aea1krVgxdz6AsioMr4hBsHrp39wQ2QG9vxpOUxd2RoDpPcCer
/Lq6df7IqyCIXVveKtpjfGpnEbvhqapog70yeii4be6ME0sZ4YLY4SNY0RtLQwdPaJ5hRq8omPQM
S5QXbu1cKR6W3eu3lV7kVHKI3kI13s2xS1cFt7ZAUMH3PzSuctD+961pu0I9Vfr7i9Vd/xIBp25L
dHJyQUZ/zfmWJxKYaVfu6B3Uo0AMoTOT5iNZoFyIX6H673XAlUtRe9UwStlYYhdtaz709TXxFngT
4bnmSAYJN4eShUNnnsvKukjUHFRSFENu1pHgfi+nAPcOk1t6x/qnv5innCAlk2AEb9DCy/pG1kOP
YRPJ1VIkd9RUMjgirj+ru9LGmA6nsWU/0vMxnIzvzL5Qv2dJlqmcrbNQrk0qrOi4m1ZoAXEwnl4n
lF60fnwy7LhatVJSI/Q4FdJW2TdqTaslEaI4WF2ntpquKIhJrT+XcBWtze/KgjgMbCAkcihEQlM9
J4m7Dl5oUQcyDfqkIizkO0DNcS569YqRm5w5rJOmAvjiP8w9lMDDjLyo5FiHRsPZntZdJMAlbGo2
3rhxhh5BMMLzBOqjTiYL1wDVv5FhdDNZhZ0aPVsQn/Q9E4khCCN8l3ZjEnIASgcvdBFq35NgTZbn
viz3gAsEMd3Cs6QhkP8ClCWR2W/taBBmPKWNFfxWlaru5r54TWv5Cov/CSxLUgBekQ6abQErkNNC
xCkttsR+imI8DzvY2L8RLnvz6DT+dC+A2uLmkLJpzva5te2MKR+z8cXFbVMWemwITZL0KU13LLOX
jFSrpXQeMXOoH6CE2lnSYEYseqTjAuCA+ab8sI4OJcOKhtR8H3N4CO/msy/9qpciPlda9KyiKGPf
nGqvNXkZ7JXfFcmJBrgXPHKM1CASol/R1XM+srARzxwSaRJlzXdenl5FwG95IjzSu4vuW0k8VWqK
0SnZkJlcZWXN3Y8OLuX5AWBthlAPPiC/6PDSVpBg2q4DGKvk79TQ+4KANaYSraVPpp5tQlE7WtJj
1MWn7TyaEOEm7ewjRR+ywd08TmUYubJmwSJ+oc5TiOq8m8sqfcs3kmHlh0tese4/FcRa+QxRYCCB
2jZp5/CkZ8VqWzSVjTxiiocGVdvuY+19Bvx2r575i964rpcD6gGZEEOXWSbWIydQBfWn4xiGwkNo
6jlcvzySbg/NOfRkzv5ORBHzHe35CIWQCiRLJ5eb0hWJyVOzBHC0FoIoqtGHSnukREeQHoB61j0p
sRvtN6p+QXdW6uKHYFY+vpAAArGxddScVQNKkcoBwVfRXP48GeYhRH95p3ToIotyhlsOzxOjRv8J
z6FMDilFhTV4kX5QWsVkzfjiwBL2sDgjv059LNLwFrxPMBZRnpgGAGXTALcQZ/2XzXMlnON9vWmP
Pbj6cypNUhl80Dn/Cwb6S/YDFhkvPVuXcfHHcIMHNo21eenAl8h+jKEfK2QpF0kYqALZCHyxsKgW
16Ri7yexwJEJ4fMpL6DifxCv1ywMvRb/mbxaXKdgL5wbRi47tXnQIbM5SGdtqjYetqk66l4tBVYF
znbpzv1hr8i7/21sS4hcmqCGqlUi7BGxusMBmlIHPRSPtHBpDeEi2Btq4vdDve4OKEs5gH3EVBkg
wBNTLTooezxut4n7yu9QZ4Rs8WyrlxuGRdgEC3Z4PjpMp/NhZMESnBsynUjunYrkKL+zgIML4+V3
nXq52M0FohAL6tvKT3NL72C3PQPhYkHqL6K3xH8gw0gyGczn497rMbTcFF7VabBtLRiqEb0R26z9
kBwIlbhrVwTlF+Qe/hxrIfuoqryminkqR67orU9+vX4NrD1eZFJBCFcHX1MkbeHLgUDhCX/ML2Ex
sfQlf4STURnK61z/hdumkV8/1rT6H+gPKyCpxFO7CiZf20Z/e7Kga0foDtvDNXx9OX+01ysEO9Xc
rTrM3O7HkUxnRoTv4+LetQYbfUX2dlibqHsOXSi96SZrxr4HB0GKXXS9lawTXoHfnEsE+L7+PdaV
ua9STfwiTY/JgoW1/mreOIjhUxo5ISy6LY5NQqzuQp3n9+8VysN4u6VmclDVqk8Pqc0wn6G0rl9l
k6MWQPjLj5RgZJDkK2XiDQJdFq9X2edpdKbM1i4yq8JizhWcWJ4GS1PY7IhptFnWIT1jRST8/Azg
x410yQyl5wegepLaXdmZ4zm+akPzvI1BikTUhhDBONvsmI1iXRKVZ4Sfcvzdait5OOD/3tzp4Nu5
iU2kzTOTBHy+YCV3XWLAqyYPnzPmwAHQoQMMflAEWpLKddxNhMeqBThO1f50KrvVXvpWG9OMLg/o
QePRkoPkCo/XH9fBjB1tPy8l3TV8/7m58Ouql6UF7iNx1jZwljrkQ0HIj83LHaWiBtKKgAqC15zq
73sNugKbihIwwcHLc9TncutYKb7glj1/F07xJdDBRvy3mGGN07EsBX0Y2LMQJo/YOO9+ta/AwLcb
IIZWGM6C1YPXSK5oyOZ06UP//OuqqrddsZjRYcoF3oOWGoAHPSUkzhhYkXblPY2yQt2c58HzXE68
OyoThs8Go6C8EQI0uRRnxJXqnrmFwiu6WQAETg23Phz8urStrVcisLSpSz/fZpW4bAPuKJ5X4xEr
hFWeTkmFMKZLrHJcxKR6qvdp9ekFgVrCGwBF/2A5st9uodKTsr80pltiEL5U1II1f+CjyJXmkOm9
b0MgmnYsiVXKtJ6v3LB4LfJQdFEu3bBNO/9Xgwon5CjWUk+YQXEWQN4Vt4tU+IsgTqJwvIMHLm8V
OmlcS2qFvKEeklhbpUN4T1FPAI0k+LOsrZejM5LPJgJFYM+gr53y1OUBBWmjeAFeynbBBqLbchZq
lJSuRxCE2QQ6qoC7G1dKz+1ljXFTu/yq7h+5XSp5GY0wmpvq923ivtrNrlMR90CexBGIedKec4dC
xfyxSaWQhABuGPr/7Mjz6O4oTIOZifZb/fIdwMqX/rxcVeFmG7w94o/ej2dTpKjXmXOcEOk7x5gu
xd98uTJQG+7Kef13j+zZtnQ5EevL4O1Ptktl42uRC2T7NmyNmUP+GtkhZLeBenfm9NpE47yZTYwn
Xv3V/Zzr2t++rj5mmjYwh8UO/3Em9tpBph6RnPTWW9tLML4aZdoBcVJXhi/fmmw4g6G+IWDD+Di9
8BoAMmhn940Cu6NIdD8oQ1bEjISZc4xRCzyToA4I4Pi0hzPvKaHikAcX0RCCXR7cq42FOath4S+2
k1ocq85Ok8lQBtnDqBCE0NVnd7lDAp8sDd2fzrqSSReQgvwYgShWN4wz4cscxUdC7xpl0vS8PFIL
Q2Q6t+2r0C2uBEwh1WKjWbedT7ok2S/YlkyMzBFBgMkXrMliqZJ/CptNQzmvilmIfLCFQ9R9hCpk
OMCvMmHDp/KOcevJjcMGi4u4BMzXILIhS01MGf62WAXbrPMuy79IJOMaX+VIxjkzbnOb9JJpLqrw
8fneKjY8lWCQiFsfLkbqiMJ6XdbcfXhrta/dUNyjSNgPbVfrqUEAZvru1dPq2utfs3NY1N3/y+74
oEzkcCcqSIwwL69QHxOZlaUOljToVXnEty3qPaJdHpDimCN0K7GE0Z+PSYCBUhuASXwjkKvqUfM3
2VWPgDzLH5HHhKkAGlmpm5uy4tKIJIahmmezIKIp+39m0P9Yjw3EFKbqmmeQWFHoYpJ54JW0thJs
dJ2NiJJFayezSZUVjWGR0GK/ZQn/X1yd4k5mkA/jw2QSWnZP1GBHSiVvme7qq+SUI0/DC0in+nIp
xEvxQevdUEMmbkMd5GBJufnA0VAO284BdAOUPiPXOqx8/lLWzUXQOhSFwkrZeF29t/vI2WA+y7Tm
Vp8C8QnnzApDB+S6NkyIvethm3e3VzxawGXJflGtNq+sS+wuonNf5S9qfMQP+2bB5hkfL0k+ktb+
UyW5MOSetRG19x25HIu6axuYWF8FbzP2EW68Nzp2KcPVwS7ewHGMw29J8eTyBMtBxuFAPLJinuVx
I81pm0YG7nmCRBRPObsAUm6+r3Nr56+FEypAl/HMxkQtFHwi9W0dAcU8pLvi4FtZVeg1YysWqxg9
VzylnRjJAMlnp0vG6YBPHIJH1iIGR11eulXRN2cR/OSVFIlVBOvMYZXdr2QzW+fh5L5hFlthvXxW
NK7LFWQ3xeH95FjjzeLyz1P2NUSIrVnFovw7w5UsAgjJz02xd11CNUGbwCi2faOoOaOi/s6U2Uod
g/4NFRcEx3xbD1jxn7T07xEEe7eUiISEs5/B0rTTo8JySm3SBxW2wanCER+7/c/b2pZbNzTI4V7O
ix1fDjkuf2/4VjMp3yFCaefsAv1GbmITAeUDKz14r1+DVgTmXwkroez2PhOcQCyK91psTJIN1Iw7
LpXwCSRHWH0cD6ONQG44Wh5lBBbawu7jYHP6YJSk4qkOGIubigDi6KdmRUpWG8zQXSFYso+MNxMf
W6+APfaoYPhxrK5r2Edx5wu/Iwpfh2Z3seHrak8TcpDNJ0k3mPyuculMzau7uSflsAoOpxBRiOpi
3Upt/tebxoeWzupEkaI9FWh5qD9NXWY6fuS5oeZMwdAZf1uXdm9q2E7LIqAJWS0B2pmHMxl6nywC
1xlQ6IQcn/QIKfokSFaWlX4YNeabH4uuB1yKgO6X88US8YxFMUkIHjx1mjHfJfiZXvkzAqvhiEtv
A8hqqPiqi/Vy+xx1iAXPH3AttoVMTM/+W3JWqEbcsucmB78VM5oMS1DILj7VGW407uR4FzfBn9M3
Ykw8J/cFPIgoVW+XEZ3Hdy3hniBwMojrI6CamfdrdQ8g6/ao04zUTN0ZroW2cpoDtzsD+kA5RQ4X
9nHW1ePNnrbmtq/P4RZD7Xq1vOSP+taz0raFnK3QCNykw6chubA/LfnLO06AmC4bk2XWjgu2u9r0
BGgpuGB7yuk1Hlgnkd25aCQUtah1ZKmOyhqCZmWE7vXOJjyJu132Cjukxey8gqWa/uEJr4hs5dZa
pjhkybPKnYWTqOPtSbHMihMW28wovisZlNJ8TyvH9oJIVPy1be4ZCgfl2v6XCYEZCJxkfnOQNeYw
vtbxRgpxNpu/ghC/5GI1oeziUmO5EDAdPV9Tgx22+th+QHWLdkIoHFoICytztQGv37QnCfjOUHr7
mqRnRFFLnpDeUUoPeJMsZStLO5GP/HJzgkPcdHc39wd6ijS+60atMl0lUjuhniFB8xzinHDlwQ8t
jE7o0697UE6VUF/MHMce8M5oDcfI315tlFkcgG7yee640Cds9AD8BA/Yfp3j6m0Q3hFiDGNctg+7
i+yAwoHkAkBd+bvu7sruNk6UwMhe6NVvXpKFzY5CaThwDoMgHDYVPamwGQtMbNURNwUzTblKK0VT
KneWH7O2gT9sCq34LjlIN8lRTxTl+ncxF/VY2Hbyh9fLSPNUQ2mUelBxDW1Jj4zgDjVRsTOuoXQ9
y9en/3CGGDK16jAZXErBv2Ruv3Ui1l/dBVSUrq2oAZClnA65D3RlAtLXepCjrlqgdL4goYOIoV3W
KYpOrwaXH2FSsI07+zmssH1FY/AaiH39Rxd2bt+FgWr+nFqbl4tPIB3wyoQAICAZfNV3dOjzjYyb
rfHvw4S+JmrLlXB74O/289/tN2g3BXLxUmTxl7vZ4KOSsAhjGAcfo8L7148ya2Uz8jaGsEIleKJv
9Fgg+765RPkwU7/ink7J/aMzqy9jLMYu9gwJ3RUh3n/EYOb0HHOZqqxUjZiJJpv9juUiHvGWBRG2
3PMpKqGw1lTbnC2sRPTBAqqG0eEy3N7ofAYmlFRRor2XYOZLXdZxo0ldemhXx20s6QhZCdH4Dybx
tCDvPVmjdstUySTODrA/fGG0L0q1zg41Te+XCAJ+VAHpiNbsLpawd7lqjPgj8P9iMUWvEZSYoThu
c8ln6dMYbSkt6eMuQRWNs2U+g8BjDGbM0eYR+YdI6OrxSYFzLrDAmvqdAIiC6rwboAtNY21RDEGq
BXMTiTsssLX0H/0b1HGWNS/9q1k8K0k7zDmbYVBA+eIe5RNXPFAzUtr9oSv1if11F2lOio+idgM1
x0vTSToKq6PHHAtPMRxx2otgby/1/faQ9ND+r29CLbdnOqvx/lqGYweoImPSqZvtmmeu+f+G5lzr
PGf6eZgD3GuAe3V0fXWltUoG1wooexOk2wAmuXgZk4jSF92x9n5KL1gJXAn18Ijc+CAxBuI6WqdS
j8uDMiOnjYQuPhncInOWt4u0+TFoWwzf7pWcdam9HuYq3qf4I8sH+Clu+WlHKQUJZCKVHQGNx4RB
SP5swVqsk1QhtBXfP04n5slmdK5xCFVDtDra448JZQSmYbrWm9ygtp4h72odVLXM4BfUdg4dNvIK
HnO5ROL7odB6sibzRsXwXR3x1oQWsrMe3PQfYXsvaXanrFaoEJFvl/zhhwKO3oZgp6Tt036xUY7h
RAalCEI5nQjpdyzgMf1mlaqmiLpmWaD3SJxmPdghjM51v7KVnRAMJRUQM3mQJnB3a9FhT6xVcJyy
p1rq4wfIk60XumvZYYr/3q+IMIfwgaSEaQ4G3fV0XAAaiBfX8m2nr4WTw8T2ObCzsq2iMisjxBrx
qvvaOgkbAJSbEk371E6UoRwUqwKAagqy2hSzXEXpM7EvS1qD1te4sSfXbSufWSfXUtHuztQaSexQ
jcww9dT0a37oQY9FrLGzqFimi6/SocBEulhPO7wvITY1140sXsaREba+7ZbJFvOLBz7xi71OrKE7
X0wKp0duj2ytgwzoKjSOt3JWGu87QYrLLYDEJ1/eT1M1O0VjJ3xskWRgE3oNE3LoH+8doMfdjEie
P8k1ZI+e9n3Zcyzlo/1gxJLTVj3vNbp6ZLTFCFIXdpYQB1DabNjRLuFMHbcXTUmcdMjwqBV/Uw3K
x+SJlsAYYr0I9ymXWINMf63u7Q6gH15itV/khWeAWDBxH91OZQmBjZSatfQD+rGo2VLB64BLE7kk
4NizBa3OQUt+TCd770TVU4X/JQSJU7xGUb5ioS6cwI+PsU5TZCxrGeI0iC1RzjkNPhjDD5kLHn8w
sn45yTFskHhR3qgTgmgNXGS0czO1Zqp9Ukeh5dmMJq9WEFof3soEtkORy38ARvnyxqQIkohbRrpm
HsGQN76JonoyluB5OOWfJgvr+YShzKD1w5XWtmaD9hNPJJukI+DzAR36V0N3TG+PsnkIwqCmdTHi
Q6Z0va5O2AZnQGo8vzGdKArV+LF4lptrsopkDxOuX+30kVXA0IBazmNIATkk4vvNA2JF0mNu2Uh4
9eiN/BnXSnWbjq7rMSXuKjm7wFYBkayvgLLkX/6pl0IPZYoSY9QYZdUqWO5b+v3ZtOW1YDh+nVk/
yl5HbfYoS9GDW9H1FEmZ9y0AbLmpwimaAiD/JazzvBsJi5Ln9QLyiv3ATZU52wkxFruCDhGrl0op
YEkA3rV8t4aZrY+I38MpOo7prES8HeVpLc+f+bGxeafr+tXSqJ0HoGAN0J2hywtR+FnA5Y5ysaAn
zyUZ+AC9YZQutMUGO9cRafJkCkBbIh72coAc4qXp5oLA6kJWieoKwYdHrVwCp+oTKjB7ZnAQUbHB
7qCj+d05O4s+IJB1A6lGeDIoX9KzR1qjhxUSmY4NhR4rJNE5iZcXGqGsGD8IQqzCtDqxT8/weNLu
x/coch2xgxtTjcoZN7slp+ELX6hIeKh8blvASRMxv5fgff2KeCmMG6zm3V55JZ/3t4KJmBf+5Y3k
I57rBIGU2TvrQMRJsr1IQowe2A3r5P3Lu6GXEOMwo+li2vU3+hQfo2h4eD277rNfYmQNPZ4Xuhq0
qCya4X7MCLmPmqVQMQ0suBCE7LHmPyyc1t1Cxnqt9Rwur6z+dMybNnyGB9UO2XlZClrq+XHGpH7j
LY4rwmEFnEoez0lnOJyR/TL30kMto4YcFK/xfL3PrthgH9tVkbX5MuwOvSitkwnEUsDDhdeyth63
7gFRQIkbH3OmfRF5hSspQ/yLkMavqBxdoomIL8TbWU8gKlPkbansi4ugA+Je7TrCi+077PaMqx6B
5t4ggPKdyrf/93iT+BaVAb8xWsNFGdTQ+/aIhZEj5YShNasHuA7O4FwUnsTYgxZq4kQJ1gR2utsa
A3U+T/mycho8itvSWBZB+S4VxyaDqDQXzY6qWAZlOiij1jhyILnEaq/Io3/FxAGONimix39zPzJj
1BG9+Oms3pLuM6ePoxZ+ZvrbBmrsm9xt2slyB8GC3vRjqeyTp7c9eNOirnFwlugnU9qOiZDyQOwA
QIdoNS+5E4BxCapOroQM9AHQztXj3vJv2M2Y4O8Oh771IzJBnm2VeCeqygUKYRJNR5wL/06P//Ui
/xA2T7eI5LaFiG3pQTP9QiQCguAvj8UnSAT0iyVxBlNgp87uPKFkZ92+aYhTJ7Av/E9ZLXCM6ePZ
/aITtavhM+ArcOfcoqPNpobQ+yPw18WjE/D+jlShEtxbYnYNqn2Js+Zlrvq3GFJsqvb/hsNdFbxT
aKHc5xbJfx4frTXN/36ZrGS20dGuXE+p5HGzjHiT9HuiTXdyA+Ulyt1I3mdAYwmIIp3Vcv3vE6TA
Lb7xMZUwsKr4XUf34jN7hxXL5je8IJxZ+7f2Kw01bQD8anFtCbazQhc5z+PIG3E+h7e9fwcs2oKW
KEFMFM0+uD9xT7mx/rdWIJ20pR9METQpBfRQl59sxSWPw7zJ0Tku1mb1r4UZ+GQzJqbTKaas1QGE
qKBUHAenCdZ4OpS8tz0pfHR4YK/QU1YJoUMcXeGnhzb6bp1DtrCLAldjFDjQMiZbjW/u3gnaO07B
ZKutEYrVnlrf5xeUiSXlGgClYWPIy6vvYQamKcdAniuboJZ+SIDRZch8CfArhtxN3uN9zUK83wOB
dOpNK4UDpH6BoM228TzkCWffHV4EzSTJXDjUXWCBwztBLDhtuLFMIi56m0g5zjsz81E7jqVlfvjm
p81q+jeeO3CPVhLKEQ80gbbdvkAEO17vZBcOMgJ54wCsZMZAmXDlsrUXqdNtPJSXUTk4AI/+8Qsq
vCjAaEbedmR7Ol/oZhZUH6dCtn+/HK3FMN54hW47MR60PgSXFBdoPTdAjoPpk5aE5KSybZTlZuxM
KPuQ7owzh6CQaKzUckqEM31AA4Fm7IUl9ieOvStHVjwni+b2e+EHAt0OKjqFqeogmEcxnzISfE6f
1+kjxjAyEwwry9yhWIKIHeO9BSFMr9KbPfHSr7Yh48iJ4Mm4lGsFkZeZzmnkC9P+tVZVsy+1pQT8
sYIyP5qRe7pr92oPmfrb39FnMO3sm8dGBEyjZGS7/p54Yn6cspxwAWNFYUlQL2IOXqGTaWUdZ/aD
XjwAVHpTsfvtvAKZ025fI52eLamz0jCRjIkdVGpMPtah84lPCMwy2Ds89RcEnUBk2jQvrZ5ZQehg
2wg5mo5MBsd0ZBcNhi7fQ29ID/OgtCtJJUcSFJ511Q3iw04h2nB6xq5V9fVYA1hBJoVSLcn7f0ky
f/6UGSYj/8I5fGimp6hzz0YJGCbAI2Cf0kTQUwgn68FBOEFIV78BHwdSf5Ut9/s1T49n7KvSOlxN
XqDC3jO5uJ2nRQyrzOf/ln2BqFuitVXCb6kbMPaG9WtCVwcZao4D/RGxMS34TvmNbnDOn61vTiC3
EfcutWtzo1ne4XGVaGGkvh0M1xvKDElnzpz9yMKlYMEO0U1x+Xdj1LQUcLB3d5Uqpd872oCNr49Y
swNqjLd2CqGdC4OVg26vn5dK0sxqPoFR5AC7eDoucNPUWWD6iX2kz+6PB4OJboko3O0yykiQDZTB
9jzEgTVzT4tzcKDCAric8bUp7TMwZqkmBdHRfXDTEGlfsHu0NOC2S+1osPSOpxQqJFCoPQbfEofD
oUe9SF727082E/sPU201UZAN21+vRZPlhrzfuxBaXafktDrSYobwwblCnL7gmXXaIxWwtLnI0xUB
2ZS8dqKkuj6fkQX2hT2f0gm4625luaRhrSWIJ+XQHQOeatN5T2LEfdG4vGQ9hy+R5CZG95asNaxQ
u1JXs+HNWkisgNqoq2MLLHUOGDmT//thGGPY0083v5FrdvQkevR9XUyiB8DQv3USZB+dQ2mq73WJ
ivWhfyq0gTZJQCT1RAQN15rMhHzAEzQNfl7CCkiv6l0Fufywfx3XIthlcBPwMHMVcpUicjGXjZIa
9J/53W8b4xVak2GHFmSOdVfaNk3JCh+4rBgbQ1nnBAA49i9qM4u/rRadW8vBDf41deQSOwGEIMP3
Bxi1PRHK8bF39Qt/ijmBQVU3QQvfm6IqfjuEolDFBMEquFH+H43KhGyppi155fweGitcjducqzkf
Cno6vPnKgxAn8j0xZlIuFutIMNsFLs8Lolesv/2e6zY5wqFLi7a2LT6ypa57D15somANAOT5krwN
bE3bhw36R94eY+832Blq8YnSYdBh83LABkTg8cCSuLKtcRlXFpZKHX7A/mJ0vPaAEzGEl9PBUI8H
EY5311fJJyfp/IwviOy4OM/dTjLIbQ9u1a3Ga8GlmYgQ2xhbZTMgoUTLVduMaUUFbG250zaIrSeq
FfFotik9jqfa5xrA7ROQIMsjjhuvf7+j+0s1Quyn1dFlq9A9tb9FJhban9O2kt0ZuZRBSj4LQXTx
S2mIa1PCkO0Dq3TW9qPmUicC40HvuZg/zjBDop2dy4ZNW9PPjFxFZuOHp0q5eZfuiAH/yNFM5BbO
qPUDPkL3y2rbKHBIc7sZI3z6Z4I9Y20dh0wZWx+B0aGNDRcafHxgRJtLZ5WXwmwkJxpuz9fdlB7r
I1Lw9PHh4gzFVzewZgBC9UBbjowa0s8mGr4p4W/CmFggdicxlG/Spwwnoc3GfA6e3Tlcp7M9O2Ix
uNqOg0h0oieV8HILwZhgIO4eR+1kqW6dmdWyWZpgJaujepKXv/i3UkLxLXkGQd/t1Q7C5thyX+Ed
LdGMKoYMSLzjudIDfaQEDoGcMyXOQW/9eKeGA+RhSd6agEjFLqwx37aaEtYipVj9A72rF1LQGa/L
rhPNZyaG+NRbH+fKs7odXi1APDfQgHKJA0N1CmddejAYWXpgew5cP7P3Qly/jq2aDxcdWepy/g7h
ZEmAN8Bbb0U8MAO1Krq58RWqY/5XKw5/Wb0CLFV8MRF1DJ/GQfioiYCdLCOLKj6UIBhukZAx0bTu
cB0qWUfSRchlj3mkQc0EmQGlHqYHG0Q/EHvqKXw5fsAXg1v9fzpNsPDKzoFjCmjBJ8gs3esveMOt
CTPJQkzIv32iYPGXj6iCvqntaQXsVzrBnYif6BFYgQJ6eOm5zZSFv2dW5O8xW28P9mdl3B32ksLk
AGAs/goWW61FedpLjlEMkAxtvGnXkAiVBkR1/8HUBSxXAaB1YH2S0va/T26oG4wk4SnfcFWS+vhe
MuEaqMB5252xATkB02/DAe612ViKtLnyWWpFof10ddqSfByOnaQK4jbrrgQuyg+15H9WnVxhL+9H
bHpRcXWXgEZ7jGkzdUPOFB4BZXAj5pxb1vy9qCKEhkrhUV1o+i+tjRmkevHnPj283GvZPN6ed4Lc
k2Aqldb+gzEnBLSynABsQruDfdyzYUbdSREHhMb7KWaqm7/vo7ojmGVc/MwRWpbrnPv6q2RAO8CO
v8jx0lnn3MvHtF7+0d0uLPP1FiE+pefxDCfXyUFRom9kpUdzv+1Owk3WPk485OLrUY4Yk0onfThI
qPOcGdPRTjGr84CW4eEj5yYKNJqAiFeW20hOAgedNcqphyxkSvG+tRaetMNzWSxKK5UNSTWtOPam
qy8NU4CFbs++uYrN9WQrvwf/BKxhiEaBsM9qZrf6vUa5ooT+cSSq9/6FMyd32tHggn1qxXNsiugH
zSGP6ScvV9+CzfSLCV6ExKSCPm3ZUSdmOEAkkzKcAaWWsJstLxoqfcWbtgkocbOcoC7RhI3e4yRw
9uTY4KnbTcMwlZSt1qJtYbJKs33xWzcZY0HRgTmPEf/qKsiJW8IepFcoBeUepMVgJe74jCwf0flt
/PzHOWMi+hcgW8ibnyq7xWxvEd87E3jxxpiigN3f8kGf6zOHbwlKRPaQArSiY2FPR5wPkgGpbZe4
lY2qeIvGtBe20ALuAZDmb8j3SokXEY1GbTya5RxZjkuaAV12FQKtpMjHWUwWv/S8A/0NJ20MRgE0
JgD0SiNTGavdNa8CVceiGIPzbI1t/N15fmpdyrapSJuZkA80EIo/a9YQjiMjaZnbRMsO0jw1c0jx
Rh+7akihqlf2X0oXt78LAu4iWlD45pSw5M+idq2KlAF6vHL++Q8/KXQ4W4NGBzi1AkH2tUz+IKjT
9tFEmLUztBh47ocnP6VJzIKmnf7USQR7BX+wyjVx4HUerxr4/PLVMbGxfHiKMkz8C53CwFCIKhTK
/e7i8S++leSbsL3bsRFazyACrIOdpxEuqeAxG7dtJuugjg/wcylQYYZJqsOlP/0A/yuNNYjPWxsM
O+AOm/k81eVgSIl9B4HxlUdTSd/Pxkd0x8oiLBbacNAr6ZQDZhU+jeDQv2bWT/djiPLZSKVGONjC
23jUZeUKTtyLIdFydpdgEI+4WavhyIOtJFxsrlykq6iOLinlKV6AXvPM7tDEF/20PDB41x/i7CRv
fyNiCQ182zu7xKLL3v+2HogqBTh6hI92Yzfxehy8IUx1AA8JA0Fz6n7Ob5suYtpceWg+wfkR+2Zs
q8u5Lsag4vBoTlVdPioREYrhfm+F72yUMdqZkYcFOaK/ZyNSUUZRJvSyXO/rVuy9fvcbGagn5HPf
849e8BxAfHugdwZ12nmr5wNAP4+MLqF/FotD6MW1NMA2wH8jlAth+2EbrLrPgJe+hrD+IoFCtucX
LpROVpzFXLTYGCVLuarvzFljic8iNhNFIQAXA7tdTlJeYidMWnpAyR3IDGUjuxVp6NsYqMD8htoY
JCzZ2oxYYehHIYT3hk7x+PzvcflGiIUnRA2IQ1gj0VC9hdSxTyaF88mUX30J8BaTk7dnALnD3lI1
uwlC6f2fWiqr+eeeLg9M/Ivg878Jm/4YrR6tFoda6yTvR58rbvdmPSogwOeo04d4nfTvvfKp5C14
iHcvQyR7vE4O7fcEzi0vCJs6HgHtUvh3e7brn9rPpNnVkI9Ko5+EZf9bNSUW4EQ4pjg40PqSrjI1
/x9RVIsIpHpYDcC29gvcxfbwiXKiuXWuc2Dk8ThyHriVOVA9/rnpT+f8bFPvtUsUNJZ+bfBvxQ55
FxsZIcMjJpIoQmIrPjrXSen9h2hTQArq+D3sI1y2znq3mkuJqedOykqMxxQcajS2YQNXGmAyeWwQ
OznKBO9xKEbfvvcW+axOD57Ve7emk4CdMd2YAv3/DZD0YwC683Kkg1NQ14nLFzFwXic1Y9KibuMx
ac7e0Ql1q/DV6R2Th+jRYQIF175acDXLfLsWzYh7kqFKLvBoi8aY5KDM8xmCp28wyujkQWXXtV4O
4OeYR76ETSLssF4N59K6vCAfVSleU4GuoqDQIOLdbL7upNPVOmxG7RLDi8Km/UOAlbh0wP8h+iRI
wNkZfaGVipOd36iYGQFLRoWPv5zuq71gPT3TdJhNduyLn8EtlZmkvD4+mFVjABmpd56iJbm+McNB
DSrlpgBjrI+lF+1LnHKr6R7terxIZJWoEVEco9S9h72X20/zgKPHpab46bj9fSEKWZBB4EUHal9m
vmZJ1xNsgiL9R/65zeUKbzT4nXV7kTbHbfhIkxBENpDgI9pmcOpeDJGjN3Sr9F/UDIrqU1HSlDWq
x15NX0D9H19umR6EZ+FWlZ+8cN0UtfPSKOzegAVSrW72aXbBhaqlDn3rjOZEDQlFfCZXiNB3QX2n
GAvAPh5poeF6n/Mfkq3g5Wv56aHr5oGanRXgBuqktetzmRJLeX6Wt4x2uAYzK3aSE52L1N6HKrc0
TdYDb6HdMucUBPc0BdhO9OpeCFHoo02HxVetyt/x6vFeokc+TpeoOpRQn630kn8UowZ3yuiGIl8Q
rGD2JZV7+UoauoapivSmPGR+fNFhnkWXI22yVLN4nNargp54UGI3z0Uu05xcfUjy16M88B+3neZ3
QbSSVPWvulK3wRkEwpNIUH4Js6KTOGVVb44ygGCVk9iXMzK+Xqi1BU600Hwmkxwt8l0pJ7atyQFf
GWdB7GuvTmw26/aAPENjvJZZzkxVpnOMopAkF52TF8TBh/BPL5FzVc18R2R1oYSK1FxeDU8NHKTk
Dyf1G0GLdlOR6zjEuAGkQsgyXiBd965LUfgyY/cp9Z9ikvbCNMVwM8U6efjTURCSMjrfOP1ULIm9
peS4rSF360eyXBxyn0v7KUkv6MkR5StfI5uUd+B9oUbCcPqASiEKUYzy+8C/p00YCa1mbHMQzhtM
2BpfmEETdi9hhNnWcjMXVXKV+Qkl53BT+MTbdZOcnHMyx/78FEW5dJOmGg6rQ/kGMoXocA/TplJ3
E54GqfxEO1Fxwjtrm2wp8hkyXl+/gTEe9deDNUM6v0hlnbnUBzruzwuHLnEnmd2pR2DkubXqUvO8
+SmFnn2GvKCGw4jDhYlR8bLuYXs7YQcE5LdFv8Esd85WjNkegKGv3HPAgdELvfAHbzxsNVJFOPFf
lPED8RraopIsZ4MHMR7YDMWL0P5zD0WJx6heTMG4bdoVatQntlxTb2iXb1MtSYCTXof1OMVO8Imn
QkHlaEPaYuRTemtN9gjfkT5tcnL0aKh3TVJGjmhY2vzereGECaCTZxmZNpSOubsKdhozOdxe/nJ6
Dh0fUtZfS9pT5BbXbpGgf8Sqbvok1jvqGi/TtfosboQCpko1N/mCQoOvGvKaNNmM4DlyZ1EUY87m
ErHMI4lxoSTL27u0loqxR7MJJG/hdr+VoAFjpFGtB0Iv1UrFXOS0qTs4gTfjbe6rdLAYSJDjVGT/
D9DT5RNiDcd0BZOZABYRZCcc5hEZ7+GKCP2JVZwxhMC9y7OYgi1u7Cgbd2GrjoEHKIXx4eCiU4DQ
/Z8FzyiY0WCRIz/wm2nvgd7O217mfQgnuJCiSOW5tJyfrx2/vAHFCslgNjYiiIwHTkFYlKyh8aDY
tffTrWUmRRH4J1gjRuXOoN5glvtw6tflMwqWyQ4Nqtr/jphspLhLHvD8jCpAjmApt1l+9NJaQDRt
UR9utFIdGfyCYDCWSjKi6hhUvFIn+J7pcasXEU7g3/qUnxwrtX71AnddXQ+ez0oIs6m1sSHRi8rl
nrNm+VZjcPyjbjJxILGsKTvxhmbBODB1Epq3y5pplBGi2Emjdh6812U0hYyVVq+/OIbj95+SKXGZ
fC7fcBkDPSJEWNNaCDe8TNbaO535+Z+/L++7GG0ey56Pp4zcihsOJHXpqxK0XoV0V2z095cm09sc
oSJmk4EsQZRGZPjy6GyVOd5dwH3CdHqEVRemWCCWZIPOfurrWqcyyluvI+xTray0xtpMkA+xY9bT
biqLlRXwmIU0dEPpISFDixuO61p/QJQfFXPxNZz8tpaK6/PXPrCtH5sPiV5ODG4q5nknmGppagMr
2d94Pb8OSCdjSTu5qqTf4AZ7IEx3ithAgyO5IWBo48B1T6s89XPtT+X8oM7mvyv99NGcK37ygV/W
jxyssKtPn0qyIB1w4Fh+W3aT5HEd00cIJhY5mdlKaLAj7VU0mUoODTKH4stWZs1EAnUgwuPqHUOY
QeGYGANcSNZ0UUL9Kj0vHsWrp0CMmnLNeB65X1JHk9+5oWNvgB7rrt615ZX/i5G64jFfWLlz2F3x
jYlmSCNTy/qXNPv7vqiaWN1R6SqP5uz36PZY9C5hVg2CDSgRYXGxwJr57AOEmGtrQS3S+JrmhUTs
O7tJWujpMkq5T9UCkHn02mh54ZV7fwpVgmmFv5jJw4jWSVrrFQPmmLZw08vuYvDiWKmSYD6oJAqU
7a6Ep1gmNRqr7R1l2TvQdSYU1cOystpQLs2Krkc/rB+NfZghGsat0ppZTeXdDquv4lv4HQWBbWMX
7biq586nEubehNRNkC5RHymCReO0baZOfRqknmy4D+nQR9zbEoRqdLunSvXtQKDdLLmoM/Jcp/TL
7LYTF0drh+HEGlXd1NYGpXn/bJt9FpkwQ4hH8E+OTnrR3iMV8gDMlvaaJqvCJhC9j9hLLmvIu08T
PSw3HOl7H25kyrPDiQb2r3PwArY1EMt3RsGVCRE+xx0nSGdCLpnL5vmSioDYljQNcmMWsmBjfKSq
nTcKZrZjpgdtTYtegoe9wJFqCzptEPjPb0z1fAfb+wp/gMGhLRuAMVXacbQl3qasRgP/6R5gcDby
2TFgJhZnR+q3ZVtUzqM5rSumFTZpf978vfYJsyhcI+vhLzPib4yI7orCCme/effH3sVlLWbk40zh
gcgCAkbRjqrmqTFNUFCORPKMsJPDFoguB9qSoE03VeDaL7d3/XEhgUlVo790jPyTENClcLRdevzd
IINdVTSsILElx/CFFpRW26JWBiNhwkwlEhTYe15IVSHUJFxQljHJpweiAoW2WtQ05KUnqobGDFxE
mkrquPz6q1/BiLX7IaCbVi9iPFDo1M6u6urlQZ+jNpsxiXBpQ2esuBHr6xLgai6Is9Ln6XEf9VUM
6yd46yGnJcvyhIJK0ZQFu0OStJvdY1tGVEU2pkcJO5g5Z6IGWly0Qx3jV/G8SNwdU1WE/5L/AXKP
RzDksZzkLqS9ailFRLjAVos+StEwAVCzOTE0blVpbWj6nZP1WAM7bVpFQfAxcIvmZhXxoDUEsABk
w9iel0u8aEfYQc/IKlFjKRkkbL8kQTorCiN38CBJCIA91eT2LG5/paK5E1KSTbnG9CUUDrnKziob
eH9C2maOp0GgJEpDNPYHYHErZd7Euq0i3JwhA21nqz2Y4cXhEg+1eow9xquIJ0E30FR7CvuG9/ee
WrxL3wMTllzmF3AXJM6QQk8beEuRXSBe7G7x0OPFStvXX5HOY3Z7HzYV4sVeRcvNRHMZBMI+PYgi
fPNHZ1y5P1nn1Kkq3b0e1oFA2fNWKeh9bJP+2i8E0Gwklohur0wlmhcQld1jG2qtyMuthZAUcC/S
3N8IPeR+cTFjWlHVTH3VtNALvphvU2uhcr0p+OWAx9Y3G0ExUY6kgRc/l2mopiZteghJwpFycHbM
5OU0vnQxF9m+IAVGHpt1jHHIHlLKPMChZJc5e0wkPezb7oTvoPa+s/g1z3TEwZUn3oNcgKFjR4jY
A9SJtlzcuPmYHJHRT8htbdBVQhMiYxYI81lCaFU7BI4SNE79j4OxrH3Ksdr3R20H6/GV5TjfNNjR
Q6nqVSz8/tyBkI11Hm5X0uvDKCEHhYZu+uWGlFcdqdC1rprWOk/mgvK9I/4YlENYBerE8Gm8sUbS
6da6lvbA1Yl0dwWMVdtpGDAvnjVPd1GJ3Vy7R9H0DxmTWwxgZCu1D22rWs3HvweFV2y8OBYo70hh
qjGmthk/UJdbAmX5qD3xunFlqOdi4X9U5RBC3aEsv02uz5zspdAUpgl09HxPNEkBK1YlmoEzucaW
2gSd7IBYDwJBhuvl9KXCz/HE3E/KwKcRoNRFchM+4UFQPeAeGZljW2/hkAEbcYoXwwSw0y/1wrsV
Efx7U+c+5azJIi64qcH+55eUCHbZnC+KJTVLolo4L5KAk0KYqNVdCf0fiDzha54waci/gy1grfqn
nITf5ccKR3YLt8T6eO2gX4V7Is/QOezz6aN6r1M4e5XXjNA44P6YDJRn4tqdR5V9BlXFqSulrkZb
LQJL3ZScDqMnTdwIjj8cEo81i8gW5OljNDhqjmsnyZ0FRxLsTAOfqiWWC+Gvo3T6s+7L5zFYR/Ir
C6EY5DwvT8OIrgaOQSgYD2u+BAIMI7b0/8V7H7vH0E14Z5W5Iibdf/3ARoasYER85rsB1z+44cli
uYPSAeYPcOt54ZKhEGpFCHrLiJ2ycPeQ8lO/FM0vzYbkY4Fcjqs87MztQCMAsT/0U8MoJFs7lLJI
4y0GvtyG8/ChMGBgOazmQstxhpRNnYeP4t2gvWbUJuR1JaZDnsUYA0OiQbZRD/AEKXH88MuaqMwZ
IN1ELY+agScAtP9Vbcf8TEanXR4oHa/HH3oNbZfTmL35W4Nmk6Qodg16yHRaAc+qiAwKTUbV1zr0
N/SA877eKi5NQ4uaQyd0zdXltVMg1mJrUrgP4V+PIQ1+mNcevJQpiHlF2fMZ2jqaJz22lZybJFtR
tN/LxW5r+COIrxueVp097IaL+F0+3jIcAO0p0eS7LTn4m5v9+N8CLLdaTtNmG95tzhdhsPxeyNxi
SQxPs9h9/BcbkBTQxJACCEYEgkABFAZdsZreBnuiigywjd0BRSEzXxv6jp+F+W4Gog/7kps28dLt
k/CNJ9njZp5PZNpOhIWiO9ArqQ3tjSW/2G/DzDCnGWo/OvQYI0rGYxaVNgfGWzK8Qk7TMr4/UV9b
ZdfeoXIqzeab5Y1odjuEx3d9BFZAkOgnh6GQC2Xzgm1OTyKdFrbCAlcQRy5VG0E9+o4zgnIHiMIQ
NGqoxJp5zajsCndzW1Xo49aOuSarYhgxLcvuzBjYr7/gC83kxo9+yzF8EWoHkdU9ZMIIX15SWRLS
nHLt/nCfXGkZDnhWl9w+AArVrUkaIlJ3zr0D/ba8/Q0WeD83kQPrpf4dff946KxaDC2vpE2wVFk6
incMWl9zCBE5uQsooIkPJQ8O/1GfZQxtpPhfTDirMYYzS/6e6FG0gUyVqkUpeDKgNZg/dHthowKv
N/Do1b7QI9UHq7FMMuUztjVB/6hRa5XqINIawoujfiPOZfLgvA9wdgSg5CoZvEywr08LT5jYWhYj
oilZEsf0APP5kKWpjBfXDho/mNIufnq/mKlHJve0mslEBlnBPKD81/JmBNZ8dguyDO0rKWrY3Cqb
s7M88+ze9fc3YhgpeeI2BSAvaAxKM4iFIkMI3RxA7BhfZbbXjcLiRme09vLTft8330f4xVIDnyca
HUbuySQtss9fQgbt2yMEHgUvDpDdmhncLjiYNc4VD+ygiK0LiKrKthMq3enM5mVG1Q8oBqjPT3/0
FGyf6gsEW11R/2j2/1jm68abpQtozs8k4u9QXVRC3OhR1zsg8ynfZAN9nvDDCLTHVA1DowmGHf5N
wi04zn3tR+OihlmT7IEOE2MHlYK0On8fzfb3UEBMqD+F93zohJCd4SUiiDXgzaSURDV/D31GMMpM
gYIR7Cc3qLN+ic2OAvZxBg9AQpyEELnsuD1hIpzsjoGqOlwASmS5XiwvUlX2x3Nv3q42Mi3n1O/Q
s+K2N/817R4VfaoH14Ef16FP19krbNLgrBvswbaWDLwLNtfmOFr8q5GjPJdzGHB8wssEP9PWJKU1
sIKVL01uj9jfXUYP6kMNVSbcA9aBO8OzZHtms7Z4dpJ6BG+00cLfQcJCMWUlPcII3XNOCU6ialii
D7zo72NCpSOW5XZDjhLsls1PQD5kaLomno/5Mhe9z46itPUH4fYJs+unD8xAK6hjsJASPqroGOJG
M6M9cvuuGhfUBBZ5F0Kka4fmvWGKEFqzOwuF1uuAHICu//UeqXYbY6oRlDKPlsLANQ7pBuKwbGsw
DIBJOJmSgp7GfJ1NxVjfPv93jTb12BFXlhu1QtSOsB5rfHjBBbL8BrTcq2um5/WacsRx8o8l7fnh
CmiT51RvjGDPXCXHLc+YG39xmpXHXUt3D6bcBuJjh8rQgHJfZ1YNUw4jWwErFoe5ioM5IIIoegz6
Z5QwY0UU+oD1cYzogdxgXytxqukGcCWmNYuq6z749kbdYTmLaoJ39YFKPDCMQ1B/c8TOXxwaJs/F
tVd4of7kB4X4DWiC9+h60BXgxVUDPbnF0jOaOG7srWk9holtb4GLoy3zRaQRCvjDhmVylD/BLmxv
0O6vm945794pn7gNjaSQH1kOBtmYlKSga+Dj3R7/ctJMo4Wij81zvnQitdu/6sAK2Vn/SWGpdM6Q
3172kKHDWLdYC9tD9FMCd/IBd48m8ViaXoWtMJUrssB/9kujvEe4sPbVQhFVPeUQy/QtwjqOFK/P
SgFAdr9vvUgtrP9wIacLVUkdlhAVP+OyC0TlfnqhVTo6qbCaIl6P/CiAUMtzjMhNEZpW7MO6976B
FHWbj3c9DYerbcjU2HF9F+eBh0JjRna+oSRtcd3t9uCWdzXVskPZZO354ALQPXxto28fdmvvAfK+
aawOvvyGTFICwXYx9SI4+ymFOxGMRUPqW0LJaKuUM+a8kVadlO34xKp33ZjRpljbNhf/1dAj1oMJ
ncYNXJxukXeplF8Ih7y/9zBB/6gfaP6POEFt/mDqZDORrxjQWeiZmrKP6+79v0nSWPvPv/89Ejc/
YArpwmVH2eEUSPsIKKiSQMHC+vcrhcRQCu21h+jP42ZJm4ExxvKZaqvM1I22F6v9TxvvQgY7CM/f
+vF6YIaUAfWyjPSigvR5R+DKUHlakNf0yDVfgfIr76DOtlKtIvoUFKhuGEb3p1HXrGpnMHRQ0AU0
gALhVLDFZI52s2W/sw7n+HdNr3sHvBuwvT959M4aW+V5TZLpLC5w34urjWdllq3emZLX8wOtDWY4
4VgotwB4SFal5iB86iwW5ezYfzb6iGRtfxcx2d9ixJx7gV7LbOgr6UmLWJAQbw4p+Z5KNv7eAzsP
rWHjuDYHHR94Mzdc5RyEJEEv2WpPgzn3JW/oYUTJZxGAyE8KVslYnoKj15ZHB5C2hvneXLcggJ5w
sjIzRx00yKJak3Tvh3ExTzxm8RbA49aXWtXNFo/9oXr3XBryh4BjeKjwTSgqb3uiwe+j3HQACUhy
P0YadJJREZtA6vURMpW6V89zR/iLiqQlDYIbMvzKs/ciPu3HUsXXKLr61HeqeWqX5+tqZEgAZLFY
eFV+pH3XYprdzjYmpL8peErwkFfI0LZBKAKmcCpqwVJ266G/B/ZvLrV+yYCKA6wHxDOvu8TXe4m9
pmoDambOf3WexgCeRh10N+S1Gm9gqbNDOiFHTJyKX7xYxT8F8vxeQW8n0Zs7jThF/YLBzkM2Khgf
ozqj2ng/z6oYs7aCu30d510njdHH8s/Rp8eOa1Kn73sE6dVuzLBvOJEoiVckQja2QY90F4m7LkeU
BWawLkL5Y/jtnq4Emj6WCRhFGwEk24L+qi02Eg25KZvNJbeQFqXjkLHlRtTxHUeqQdCKT6ZukzKZ
tFOKzSBBDXthVpVL9LxDJlwT4GqXQ+k6rdV+xq92XTyzFc8agLrEbmGzkD9R4LF94fhlzZ4OYfWg
GVBlBLnPWNa7lFIvcU9CT9gl/68cxaX+sbL40abrk/TeadShbLv1DK7e/300F+ZvLMKRhqalo+g6
HlfjUAvMQZJJ3wiXMAF14Ba1QaKMhweVVvKw7SeWa6qdE6AMUkAju1BSlPy5ZV57bhCfeGx3LTPQ
Bpn81dLLNhlSGrVuxP176KcbX/0LwoclCmqm0sRjtui594RvLOKE1Xbg66MfevxdsgF3vRIQRCc+
Ywy9Yw70UkPVbIIL4JkSgR/cDW3ssN3qTcxvpVppu0qybCjF71/GwHqoRe4BKPB741f4Yz56WW76
MhLGFxvOxOzEeIvPscqWyUYoFB89PL6c4PIC1j5gyhBWj8x3IrzK/oOMDseKjK6EXYqFFUZ1Qrdi
ziggiYLn88WTORKfgVTnD1P+qhhiciwdF0KyEHOeZry5EAvWobb1j8RPiP5LvWSL/nmDjsFv/Ccs
CaxI+7/utbcG7jUvM+gs9onsqM68960yukXDvp9hXfrrGxF8TSgor2qUGhXBxSNCxeNYfOrQcwzG
Qz8zNBX2YgIjyZm9JzXL6Gq9n1hBKl+xCiMcBki74GfchEHMNs3qfGNEgmGn+MHJnObQSSCtZR3n
Zi2AFiJM8Yz2P1bs7YG9d/A9BRTNfvxsYWGGWo1l9/c1fHQ1XdIXdz0Uh73mJbiYLX15IUEK2GDt
pBOUzy7CaVbEqQESXr7CSqwon4MjberKXMoX8O01Mk/SRx6AY4K1R0pbOkKseoShrbh863vME3fP
ASmZdhMFY+erjSzDlL42GpLpaqWJrstRN2GQrR+bXzF6y+Uv4harb4vHRAt0JPexHfLkTZUrPt16
eQktQIQh98GP+zHa/zcdfeOsQOnz5EEcW6rHXLBQs/JuC6llrPFbJN/yaoYtoKLuiMrdd1YExpds
xh9FBVYiMgQxy2BYZBZUB2ElUUlA6LTe7lsPuks+TVw8QMCpu8Mp63LZ7/ptSEPdFh0WBXeB0+xQ
CVHvq8pqIdSdLj5HskPw699sKnYw4aM6zlve5fvYtJEWXGwQBYzbuh7tBwY5nOLf3AEU3AyEifS1
rChRNJ2NV4+7jAMNb7n+3Tib56msnw5/o/FtkjbPqvCnH/bV4ZAHRqVrTluEJnUC+iKMyccOpe1V
kb2Aa1nMK/pkCWmhTknXvg+gxMJRgUPF9QjGL/OVTvSGKfAMjdgTwlU1DVJkkIZvGx6vIJrcwVxj
y30WkpnF1z1sffnCpoRA1uTSnIgW0aekvrnqLWgLGckTLAfv18VxgwtWdXhjV14yqhScg9kTX4tF
YTQ9BJ56GtWXYGj0Hk8C+TprTUV/IWuRjR97ld3XlmV9YE4rZKftZsc+j6C6JLxMaaoO1fNAmEmK
OtZ8w4kf9YHQh7KQclLyBEdKADVDeC8e6o0RLJ3Ac8/QX4SnRHZWZpHP9DEY1xbWCLjdjdrr+XKr
51AKbHW7O3nPDLLzmL7imwXIApo8KWREQtj0lhsf/BQCRgc9qjhcFDOWowi2YcqWj/VfvK8DNZWm
RZ1pjN7g/A6jd+8YF5QXBUHapMnqprughvue/ZkMTytfoXo+HQ3hdKE599mYIUzNQFmzVoVzl4Tz
CmDNvL1XdkGc5s8OEUAdxbZlixx5AYNM1pcBwVvzs14cwzz0F/zr2KUoXDreNRenBlztZQGDpIkF
CY7heaehy0jgH9O/sMApXlIxfj0pXdQf79fpz/upkyzAN3I4BOBCQn7mhm/mruuAxzBKMVUw7iMx
Kzp8/cosPYYXDkPMDMXzNEDPkJcV1j3NFZTdQYWPcvbSEdAiazWNxWCewhQGpZ2AiUT6Cm4iFTZd
XamIIz8tVU3OF9gEm/L559c3IGEbIKwVGItiW8rs4sjBoJBepT4LLPb/B78vzx2iYJdnti+d3lRN
aAT5hVZfQTp8LEUqTzdU+hEkLc5K7L/0FFGahu9CldrNKaCSxq4BkVK3tBtrtbvyxaHV68hR26iL
N1EI+ThQPjH8qUqraEiR2Q5FheAuptX/RA0w2tMOQHJW+dttLGrQmfhaFOrtlMvkSfIJoRTQZBJE
/o0SBFd/xwQSSCK/FklR0f5viF7mr3Nex7TSZMHp3JGLWXt2YMp9r1QNM2EaAFdCWHeTukz7StT6
1i29TOFIwitGm4q4GLMVo0ru4G0qfj9X0JVZVwndo8zxnueUh1J3s7Vf01IwkeZYK6diSJvlY5i1
VWRZ1Q5oqIOMwlRHoEGYvjwvITBpxVHWghnP8jQHzXbO2oFM7iueqwQNpvHLA+SjMnlVkGl7y/EP
W4znyCp3IhFXa/PhOjwxkiWwn3o7oUKFExH4OE6I/hItd6tGlGZK1luLZXXWLoa1kb16/n6Qmzno
uraQ/zW9vRcamVzwZ/Z/X3Tra65LdAOef/+y8w4HJbD5sxc1vbHYHP9v97A87qdRsdnRwLliEBfd
N2g1SMLZjiNBF0ZSoEequAu9tTlztdD6V1feg3nJwnaylCzObK3WuRiEATi9s6W+KXxSTWjJlHRi
imS6YYhjBd96cyfr6DocdkxKwe4qQXYKJsqBBrjSq5IgybUGNf3/Mb+TnNJ2/VcOoL/RYG0pac3P
Xn8w/SmSrTBLtC7iuKcZvhbSacs7elsFrtcJgOEn896gwUVcqj77M4Ajj8GBckONSUcR4ZDF6rs7
1pDTxJUVhpAAfvBI4/l3eufG2C7vU8DhH6kIOixORT2Q8kBjGqb1y9c9Nw6NzRHOZ7Z9rsL6iQFf
PtRDKVEvV1UUqef8smmR58lWWVAyo0oWciKb0mCWhQhodik6qN7CO40wSr0r+hBivweC2DF34sb3
CJxT6wxkNqznwGAbdGAMfGxq/Q/GE/nCSkch9z/Js18QGWWAxPBAsZ510z6WRGzLi9cunlJd9uDg
eU0K5CgANsvxuiOf84yFn4TWA2mgwh6kjo4s7m6QYss/wdiI03GPCdhUhja4a5ItZyLIdR3k1OX6
ANy+Vnj7NVHBN+PrHmf9aLouosAsPW/5gjuERDzZtKF4xlwNZTmorNAhA6KhMaX770Prj5ceDYDA
9EksxLhAckovRtX3UDrDCWa+eYSIjroBpkTTPdIUO1wmlfMOScuOy8kpGzEmjO7ZlBBUvR6hDF4t
i47QA5HvdL4FZr48XuPk3vqr1ccdDgINP2Pv5RyJzsRSpLPvXut37fXcwlK9iLEVFaeAGENPBn/e
dmoLRIAbKtnNXyMqvO1QyD1ahRs94QXSM8NibHsUPuIxOn3nTKa6w1MXR+bMpZLCivhsEqrZlqhb
8a//i7Zx8j+eiHkki/6atEfVXB59Eqo9jLchvZitanbfLDjpKoHv99s9S2xCrD37Wgu8JZqGncA8
8i5PKpLN+zN+j0BKeNCQu1iFaMj7CNv6be9/Ai6WoQ2v7mQ2CnWK9hlYnDzqOIrkW9MUyMYf3yE1
6R+FGmWNc69xENO1WQgg1nCZlshkD0vhbIaN+YYcjqWKEvrKnxX/9uTSwNj2+W9lPEfi5So0tmSb
UQjXDCTxUQPkSnRI8UDD5qANLHUV73+SQvfPfVV2bIpcVNjUYTjuEF0IUt01PMktuhsuWC7oOurT
gVEGOQO/36oEZ0Q683CVGVGD/55Zyz0hGWbUdZYxNk+MlQ2T2xzIJNukgzvIg6iwW6/POin+CTnT
YK21w/1wIe2iqqu+/sCYUiqjaD62XrzZxqGZ9Wi1zzMmXWOMabeF+4ZR2Pn5zftdINHI8V4YClO0
UjgZa8ME1uwhdbbsp3nh7XPJMMkRjoG9Yv5GnhWs0SurRp1Wd5vOPNZ6HAnn8lO7mquScC6jaT1i
EjYbSBNCVgqoB0uQzVxz9NKJAhaO/9+ipnhIAdYfhpQDig8ik4wUK4zyyRPUtS1Le2NQF+FPxY6/
IKaj6e/TxEpFsiGc1xxk7BofExX5AV+1LjORNh+rdXHaETbpaci8gKo/Bb2IxdgGWaBFlHhjnudc
pyyLr8dsGo8ERdksHRc23vMRcKBg02uF4x5fHG2s5CUnlXk94lSPxfoDOMKoE7tBQPv6/GCqRkTK
BHcqhV2ghyYzbW8y0LEBRCZoksRgK6lv8rq3b3u8pTl5QzUtRuolTcxRvDsqTbpLxO3W8b4/AXqK
bGFkFjrVW8LFDsjn1U5vj3vbx7XiQ7ZbACxoSjIUfKJ6PNY27i3Z282jKz1E51iHKuCXYwzvuuzC
/ya65xtq+aa2JkclYzlIFZfafpiKGs3tyRQc0KMvINXpwYLdG5hC/ifOS7hm0EZyFMqrVBmaQP7/
C4/BQioJBFH+3zFQOQJjRB4zzTdN8XgtmXCKVCTQqpx+5RN23+zppGIzr5U+7TKVroxY/bpPMb3o
vOXOu4p6DPlJQAPS+687UI0ERNnQZmMqjqHy7boWcuNJghxHJRoABS9q5LW1ZRqkU1n0gKa+SF9l
HKARf4EioKF1sikAlqusDbKDc/VphZvN2R+yk1L5/fL1/2wWytXFBKG3GUpCYdZ6eZE1Hyg5tv98
WCj8uim/g1MGErC7P6jLQNtXvWvZMio4cDOPP38aHk1pmJKtd+CSvgt+LJc2i42/6IEgzcuI/yb8
B4sy/Do2ABfRANgu7xjlkUNxnkL/B8eg5LDbBJpCGKGNbUcQkfuSG7TzXwqNOIAEVLsCbIboVfC4
5TJpajZQFOHZakT11JKgdA0Eqo65Xq+jBHG1zSbwetTSL0xrCSyDU1PtN7+jZkAmH5Sj5r9tRlXN
JyZpBVKraAmleaxN2geR+bRHXAN8+4po3/ihnnNVPHLbsBjGkc/RYMnae3mUlXGtP4GBhGKW4a7b
Pa/7/lkdmN70cBAlupu1FiVU692FvWnyuexgT4DXrNL3BgBY+t+IpKi1zLBTXdaQNVz+qJhEaRtv
/+XmBxVU4pbWa150EwMAloArB96JnpRT97hUt0f3mcbCJZ4SoUfWRC52F1nKsXdFmd5XD8aQXIc9
bFHvneWeOFqHFCUdgodHJ2jdPEfKNxCy/9EluknpeUK88Cv1cEmFohX3WaeL65DVWTXHNiSiRV+B
auA/yKCe85xzZ6YQ8SL7vGvHWDb8f4Y6wod79LqyP+UnyvVwX1oI4HY8OsyR7uM1gHezCiNOD8Ho
/YSyGpCda8MJ97/U0Ct1yEoylYdZJyXAuHzwpXve7qmAjcAy1BjrP05GNOKoM5hCPa/3AEkRvQ6Q
nPW4UCspasYcJhyBbM6uTgtvF3GBxZ8izc33Sd0mGLUk6+AezqkgR6bf8ndHX+b5EsbJtLuWCqqc
57MVaYAKERR7ujmtIhNlHqBwQ4xw9OZLPhB5EiwNpc65j3eTv/9wznVb7ZLyB3nbUkdE/jeJY4mL
YPd45BHyD6WtUNKd6+4DdoYRHcDFzqlzKO63vbfbqF9Rh6lbtmUCX9IlcP/UxFbteFzX5VQUjfHX
GRpv1xNzASd2BH3JgvVEiU265ZGko5aHstQ1qnKsCj5tqFg3Wd7l1y+bKCOcuH4ye73wiF/Q1P6s
joagAeQjqCYbA45j7TQqvqvv26dLOHMQ/7d3atmR3lyiRVQdkntmcTZhafSZUnfD2JvkicmYDttS
yetEsq14QzsLhkNW/5x8Pruj2ZFAZeb5sV9UH+cJbmOqYry1Grgz6trYYHo555fd00zs6zDtLKom
IuMXG9fZF2dFowvz53B3tuy74YKIVTnHO0ojQ2KmdwwWNFQqTCTasSesLQE+kq+lGZ9yoEYGpMYe
tS6qOtKcO2YayxM21wAzQu6FVkaPQwEKwJUOcgF5HZz+CRNsUkkspPfxS3Ipti61CIu1A4yiijDV
kTAuwxbMC8wL/E3OwZQOurYWbIBffFc+LI/1IQNhoIdMn4/o26Az7Mk0rHCMQOsTdHmbEBuyzKzK
OiqXy0CzVDr8Gb8dGJrd7OEQj1EOml5Kkxo1eZnvgmOhexxhUDxjGOCwSX3OwUcfKV7LvYndV+pP
ygC+PtLKM2l2X8oiy92jQMWu4r5mrZ8PhoPGQwPuwEFaMSgCRKwvupwA6ojk838/k88oeix5Br/W
T5GCnfuKMh3v18Rtz1ypwZCRzIkeen/rLNSmXZ1zaEj1M/iMCW8hQg56Rd1L56OxjzbYK+QwOU0+
VthfQqR4OKjQuz6KGnVGmyc3HkmeYszzb0SXeYmfQbUF2vP2M3+Xm/eGPcCk1bcewXy9aaOcROo1
Gv6v5x0wjpZ1R6EOhnjzCSs5At6/mT6N1fFUHWv1XwTsrx6BjeYRwedtABG/wa4dEwgeCcu9atVF
HNeNbBQNJhOQ1pljvbR0fIGl7XUvCDv6b/8eq06Fd9R5/uD7EJODTDYSrRUG8++bKRWrL9HTl4H6
IoxiKgc5ubwLGovNfW8RU+N1afVnUaGwisI8TqS8HWJHGWT5+I3WAC5qeqLdeMxaI/HQsyZFtf5O
NeWeThPhQAAb/wL3QYlA0kgExq3XT5DF1zY7Dafm1TcsnuS3l3LFnZPa+OL0ypLsjKvbXQXg11gW
E2XKm8rdb6jikbdXTYc7YHp8CviidX89vnE7YY7JrN/qJxRCPi67C1W1d5GgPr6epEwb+46Idl7I
R8Z8OunKh/EWO2zfnikKIJZ/8MayiuAC133oXX8bawf+hCpPovOImEOSnU9hdp6CtRdFTHCSpQpk
WShElsO7XlNTN4lnRLmUVLtm7nZiJzC8WRzkjm2L2S3t1CQJFzySaAQWC9Am2lCJlvhP31shvjHC
F3Idmi/1EzH5naZn6+RsEKCpYiK0xPH3uCKyIOWU1FzWjSF6y3kKy1vnBLwGbtW4nO9PqGrIgEl8
hs9St1zTEcIBm17fTOEWerWWhfi7JMDkVeA6XO7rEoGQNy5rF8pp89t8HGOBMD6Q30hd1jxdiRoQ
52anYG80Ez8Efmvz+ckaAZnOlqim00M25DogOrzD4cGFsDX7GyJs6R8q6t03lcQhXX+nCfv72k3D
8z17moSAEaZNhMlN70IgZZH+90QJ4/GLbYr9aPKJ9j0eFEIsTvVCxxidgWGicNf2lu+4aFy1Py+s
4AGszFQiz7HK07O2DtOMMcO/K+qIj2LSuOUM74cIL/HOKvyXPfQKSlZfxacLL8ZxsrzQdSXI71Nj
ZERciiKUQ0VLts2pFnYSm6kSw6PB8dKKnubwupgzjYhOcOAV3tHewxk1KYAP/i9GKVpklb/ib0bY
KxWYDFJ/HILPIXE3LhYJBMYPXh1lAnc8UwFbwTYQN8AdAvBz3ddaU7ELe/TD6YwyTIrVMOyWr5Ya
eonfCXjbhRpqGm7gmtH6WHoeja/kMj2xT/fJoaUFOGastJxbrhvtrf7ewYiYQXzUDOe6mGO5nlDF
o4hbv+s++ec1lvTogDqQ6l9JM+wGE5+rpMbxoLJV3YQNNEU3JzPx9X0hONW04hKQsLTwOucDHZWB
T5HsDh6R3/uPEfDRp1EiaP5pmaISoKu1T6otoAnx/V20isdhpTxTbmnYHDovm7na3SONp02zgfjm
e7IV9InrVcNjWEZzo5K5cvLMJ3sjrLyzqB5bOCtD+QzslX7MXZuklmDMQ0M2qZ755Y8O0FBhw0wB
h14DzOdwZ2hvaQ0TKEwtgnFAJWXOoVQduK+InecCYwmWf8XN413mOMdEo7cyT5Zg8Ekllk9QZHYM
p+MqqMpjfKrVNt/OR25lNj8rt/r7qs18RPlI2O4CZQh+9LeHM/vGLwgEaLZWY05XKjnZgOanqymo
Uhu7Ly7PUPqNoi+cYAxSiTuh6tIVTCjBP5ecsVIquyeMnBA/tD33VaRkijviTmOI+kLi3d5o/i6f
mEHkkHc8Tds59OeyG/QPSe6n0ydjVgE/F1sJZWyMnLr/X1+DSg7pjoBHogcSDw8mZPxaVkjwkYRS
vfuKlf4hXCDR3pHTw1k1rTvWJzPl5ko++WSkqtkOjk9Tjc1oCuaL9+lJ2xFAg2F8tu6JoqQv7RzH
x8yJ3J9wEPiuKQ9lMaTxPsqrTv+fCPMIZS6Y4UlUbOcTKMCNhT6uM/eEMEtFtBrI9Q4Yom8LKnDM
shKHheWysWXuhII0j2Cuo5wq0Oub0y0dK/PTdAkyyFwCVYkoCPkBPZe2p1cyOC7js5JiVWCaoK/f
azSw+xvKOECqNe8tSbDPzXyiJtA9st6TiQknW20ZQ7TJIVHnsUnhvLmNBryRLMIzGIBvGPyj55ZN
msghzRInD6x0NPbBRxqzSyfZyUXHiebNvtyuzt9umR6YKMWCb05AffU+6HxzBcT/MChiDen6O0r0
Y8Hy/9C2dcFipCNFdh0SHKF1xDel6zx9G6IwoJx0dZ4WM0w7fkfEuadYn05MzkCHXqceNkNCgtAq
WzAVHC0paYFdcyIiL5baN9rLxK/pujlPboSyNq7leK98yx+18V/EHEXVahqPqMFQV/rMDm6K5kEL
sZ8GqXupWebf1TiE0O4EngxDfGp9BMV8gBuCGgIxeajFs3HVuuo5ARnXQHowZ9Yc+Z0cjzkp5Hfw
nvulusMeyEWj6NkKhneyGQ7I1br60FR2UqoW7UE9s+aeVgEfdPirzzpxfQWxqJuWhuZl27xRg52P
93jNLcvtejoxeUNsaTpBy51I15E7+gbiP5IEeoRPVc5PkTXCO4igdDTFEHsAG+t3AF1KLi1AUYe1
wuXll0DYNNRiQo9SNStu7EFHfK0t3sHETDZYsS5toxQ5pcR168L6q2OpX+saW/u9UcpN9emIvkfz
d2K/wexO9HHgbQMRQ9Wy6h8510H/eDQb5WdyWf7Hm+ijJDWVS3KBEaIJphKptuRpKTxSLUo21n6R
2uzqLA09ireI+FvAHOJhHBN2fsFIvKqX2wA3rg3k++hfldlBGz65xtbN1WuKFe7PcF8u2Xkahqc5
JzS3hrmvQ105WyS4V1s0oIUk+P3NN/J4S6HlpemYr+c1G6KHKwicUKztCwgM4x4uJ/mLvBkpTU7+
60sq3NQaToK1yj+e3jf4Qq+fm5TZBKFWp6lau0XoKoFhhTwmN/+fgYKoUoRsO5H9/uosze4cQqup
/hl0C0io3crYxUPSPJwNk9V+W0KhvfgrvrykafpTszIGKAx+5bIG1NeYZdyrZ7JnEfO89/oYYP7V
9K49TCJYCnEZPMA4n3D4Qdx7+iRwdCrQ7XfpNFM3z3epNzxUHOmqiiRHVOBztcTr8ZEaAn7XUaMV
FLbCDgM6SzvxukOJx42RJcndJDBkuJ/TKQ1vsBK7rvF9Rzel6Y9jM5nfPpfTHSkfvSA/njt8fsDh
JUaIzi50jltlcR1PRx4M6L4ZJpwxDr7iJ67aK3sm0iEPMmTNGslrS2fWYnj3gcGpubZGSGdA+cqr
BhZzqW9qSwrvFItcBzq8IE0F1zwSXOaZislkZ/1TTBUMYl3oWFOiHbG2PEPtbR5aawVUnzhYo5IU
b6TU1hYKQD5RYStrimphGbtCbbxQRkslfPk0qr4gsIYfCseW5Yi99K11vHOLI2+zN1LVJHBO3gqf
OZFwDsAhCZ0aXSezz0R3T+o1ZKBxlTXHSvUAd7B+n1NQVj5JuZanepi0QCFQJfAh6sUIYsVR64wD
Z+xfgczsXscNEYTC3UHDdKt75qPwVo4XAeaRUYhPyYmEyoiUbHusuDQmevReR6MsAH8Z1SC1U3zB
iPhtIB4QGiT3H5YFW/OhoWuu9IqzFnUAZZV0ejLeKnuH/vS92Ooj4nYfl+Bi/8vw3yzV5/bvo0oP
RDynMSFQUbFE2lecZUgZ+vrnzJRXWksD6BV8eRdOMppiSfRQpop7daqyZn1ZwkMw4MFBYVL/Mf/J
L6nr70FnZQGZFNsHn8CKFz1lQa/xuZjZ/1XrOON7txRKAb9yV8fzVdyubPPvREaNbswvLp149VMN
9Li19sYZDi84N22gy7dHyjIPTuP7oNFLr5NTtvvqs8S1EyObj6HUeK+UwQKmtVpIizn6ZwR8kfSq
fTsjq0XKF8X3iX3CpFBsDPq6BInah0XwNUHEo+BqMnpMvUFTphydX8TzFJu9L//i5DU74UD97Xou
1k4AXlJ2iZusKyCjpb2dC6dyE6NE/rjVvVg8WGh+Q35cPKn9rkjbJiumPHsZcn6UcVaHWFc7c/Ra
UAYReDhnWMMdlow4KnoixtQCaWvUbpDGt+I598CgaIDZhD2BDTAFGWTzF97nXP+gmAv8xT+RBeeO
8iN+wfM+OtTN8t+cYsFXLVkwaNEtRse8rbX7ugX5hR6Y7eGRdZkjIdTZMZDGWEVU31Ua881orfuy
24X/YaRbbEzl67sD69cJ9Rbp1Emmf0PIXSbODBT6k4SnEid1eUFkPSHdmhx5cbqa/n7XmqSyxMci
aVzZfhjH8XZn+pC6DC2vLBamr93HjcsDxk8BZjBKvvLxAwDqUmxYYJ8vP31RW1H0qTEUzrwmOwer
cwilMxaqoXRUdlRZemibZ6KFOIHCjA3ltRJ1mT6/bdFw1L2ZlkubYKM9BK5gjxtug1DmH9AIOJnT
ImEr99FaAhONHprCokZIYMPH+j1kNPPavIfHhniGrt9IAOWt4NeHAZuTLvDiIc9BreJVAKuE1xDw
ZJirS1Yb/asnastyNPcfJDL+KSh8SOR0KZ6oVdzfuWFmZDCdit9A4OERAP8DSG8Se8f5ZY0sMJq3
ZP9mLe3UI/ZyewIzaisppqIAGmMt0EU5xlBkCgGreQYFGnptd9Rm3d39SV3hdID4j5Z7gvI+JrHB
64+rP6nydVaqd/6a3TLy6+YOjcXkEiTqiU/bzp4mDmiGdQR9ULvCY1GzF4ycGGbBcBdl1ILGE/xX
VuxtEliaVVvWlC17ZF1O7bpmf/ceDEjRkDn0uiPvKeK9wO86aw7/yu7F0pWlGem3qAPDtwP8Lbqh
Owz25MrGK19u4JzwCBLU4y4tgO3A7lIVWr2Q498KPqs6ih1nRZseaXyaN9zWRUXaJbsjEhwlCQw2
oSMIeU45ceaATcGMSUhx8NIVtVouX/JuERyIcl7Etkfoj7i/+Oi/EOSc9OVbLXCXM4c/qgzyf3tZ
ngsTMBlQCEMIa+QPX8q5MNh0qClUGfdKQuIzkeooRjFYylbcaPac2LU13OPPxsEt2f8omsYJKQ19
c2rFJ5jfe1leSX1jwd9zHzBNIvxoLE8XEZkgglkqTvZTM0ztFDEXrwo6Dp6aFoowQOGFyciy23HM
oRu0a5i09QdueDmKfYMg8l6RKb3x1Gg8HpJUSOqorVtQ20dNrbIl2l13zPn0ETrN5gB+JCT/viIP
6t7kgT/3fTPee6utAwa0H077vRvXVVmTHqMKEzrhVDDF1r3r0QhvVfG6vIyDG/IXrUPmS2GRP6o0
5QHnZm5XKoMHC8kaxCBwm87W78IA4nFUu4ygKrW7R1AexSS6SwbosJtBfoFhTpHnjt6/u42uNRwh
xdrw+pI/IjVWqzlNXtAv8U1aBoYx6F20/jDkhP67fbSDdnMsfrWQiHm3eA5SHBEO0BVrhh4N9fv1
n+/c4m1mxM8Xl3cIaqNF7gD7PCVADSK+ChO/3GbQAXYOvIskD8IJqeywjX4XLv87y1SXUqo3hbaJ
wyVTUhDW5E0CbAypzUqlM2FYYWjIn8/Lm+JHbZ8XPw0T1BPmR/Mknqm8ac9XIOSK46bbmXorqzao
ZnEyCZwfvmMigJSazZkrRsaO7InQNJaZq1xu5NIvw4IE7YyDZv9SB3NEEAE4wOOUB8rqH1To6ftr
OPeCNEIJGIN5In5zXG8PXKHT6GqmFLsPXXsUpAMoG5w9dJzCZRXhPUXexh8HtSrHZ8LT71hVeox8
gQGFraoRQTKAY4RprQsxPq8o+0B+lhayi71BSs8olQn7U2OCgvmp5OJOB59mbEndFZF4rr/Y1JDs
B2EUoppVJECpzxNcPmTvO3oCOqui2YqBvTl9odb3bxFvVs4KMbaLYqXfx0lsEsl+UvU+8IGleBrb
Ixkqld7fDBa+FqLHCUEWHb5Lv3/p+94yH9dixOQecVO4p8lHsh9jBg4/+SmhjvH6fSY0KsKJgFpT
Ca4ru2K89jWJ263/zgpVylpQOKJYLRcHewVjfx21U9vhO16oxfijpnFJHFojoP1DAsH7CW3+S62C
uQnH9s/KLeuUsmXFywxrtSX823segjdkSK2j4HFzehWsFWyV3XkP3ChR1jUiH5wKJxTVEakcu6dL
oklhDQXETGyTiM84zFdiEfCTahkNLTixC+ugVHxcLTGNlnEGSrbJhVSr8K5XV18LE7+f9d72DezU
W8bNRN82EnJfxNh/WU+crXnic6mZTvM0fsm6VjtYj6m/JlFZdTRFShoVUWy53jErXieMNFnYDw9F
aTGmkka5ZkyvaLHvHLUxJJcHqg8Loton+13vS+lDTr94614UfmQpDjARds5TUrOn1S4wvIF0bYsi
eLVPcWc0FGWYqUmQFMJYMCD6Rss5+VIchPOKE5nd3MWLUqrMSTy1OwwOAyRnJYRTAr1biL4a1VX8
yw0xWgesAMaM4Vg5UK4YTcQeOCQ5AaIMIcOdePl9ygER71Npvs8OOzijA1Dw3nlFjaXFE36aOgV+
2p4zRmMCLnEgtXGRcscSXu4tANBi0kawcNeykvspi66sqqUSnYojvyODD+sESYdY95AcKSUQOT9F
6U7Aw0aPvQ/Gk/RwVCaspE9e6RYKpUD+gSTilZMAzvPX4BMJmeLgQ/SOJuPgg7D8OZYswoqPnmz3
TgxnV7VjfkSvkMV8r/8dA5eSQkQDbREVYiMXU79IhObO1D165GPkgTHVLdisYHtcJcv0GmS6PVYX
MSvrcwmzp6cyVMSn1hbxrHy71pTBHZcI7xM5ALVl9eUd/MuphhPrS2mMHKD9vwhVKvhMc7MThlbL
Ayjs+0di2fF3bqOFxSN9bXgR/jvG6NJsBcF+YaC++ULnfL3dMfw9ge9hZ+vgeGsmdv/u1qEvV5k8
dBU8RmaquSk8AFWTucLdc4U4tKKhfj0tDO2bV492TaEmrg8LleTtuAGHr5M3q1OUW6FJNV6TW9eG
FWuyFhukqt7P7Bmn/o+lLeCqPQwn/PBYj+VUAIez8LmRZljCvMd2ydBOkpQQH93lS0bqZidkKCtT
W7n3bAkaR1frCqcn8iM3E+3UMy+N2IFHv7JLC6HUY4kAvc3BTktMmZ8Exz4eykczKaNIeRaNrkgm
FvJ64ZPyEkdc6AngDND4ZLfDu0viKoEwCTIr+ilo8kB2uJUS5t7PLjJVvOeUuO5DvdK/34W/q5j4
lbqtTl/T0Pbm3+4MgSOvwpqrvM22s84cwiBnUirzUZCiGXLnH+ejNqdCNLAFCb8ZzhNNrYr0eWhl
vdZMVLYdtiNOmj7gvsD4Bv0bE4uQx8Zqi6mbyb4jepK6VJFbJWZSDrKEYNF7ZtduykhA2n8bf9LY
XA+1hpjAcM6VQKI35N7KZaq+UoDmHscuBFCT0Oad8GIqD7/NE856bVV5kKWikWMP5VjGm4VZjSr8
Z8jh+5fWdSq+C+4I60GsmHTlt+9a1UdMhiw6gKDm/FHx3e0ULfdqTvG6VNzxzQb2u665qanfcf85
bhb/8ENoBwXsThIcdZAqXRb/0Cmje7zqKUs2dXBy08nIfNuC5NLEqycP9PjrNb8TxKw3Dick85Mh
FRIs/bljDGC6jaBNqw8caov7A/viap/SWzsUPdggnHzAwiDbGEfLv3VrRSQRPCWuc81wAxxIyTKg
yDLd5Me5juI3qsVkr/5cOl9fc18nXRO43+kDk3m5Db/MMp/ytw3S7nNHiZ8naFQKMn7FeosCU9Wf
U++xWNIfGEJFpP3AtfXVttvnrJWSVyt2trWUbGt4vHj4moMkXxRDbbjVraNsex656uh9+M/mOEV6
sTwjuNJDdqYQTW1XjoYBtjKS3ygl3JyHUkrqcePJS7o0yT9G1KAHR5e3rtXCDho2ye8AbtDopcYU
CVH+h31o5xheMbXViNMyluAs1mqJWgSUn373pvMHlZkv/CSB7IfvjEnBnHs6+D5F3TteBQPeSPdu
MkZVfq6ZKcMC/G0FVCmIk3HApV3wtUsBEXSYv2/jBSWv3KOX+uq934G5FVt6ZrY1Du0cPtyR85PT
gWY48rTOZii5ruA/VOCYG2fjCCTZv/6dtl0IwqsLNRkXAp7cSJeV2QcEvWXw8q3gjnVAjcKnsoOF
EONY0lxHAQTTO13CzL2svEnkqMOgfa9njVfoh4F8SSXnrST6BuG/jm6nukIviN2Vgcm6KkYLPEVd
x13Jb0HWsxSvuuLUgjwOE7+eLELHBIez+j5wgLmvEGIiyHyHJGQ5jxP8+TSDK51+ybmFd1sCFu8+
qSoq81w4WB/GKLYAp8vTO+Mv8CgMVk6kOxSg8teyxxmX+d1r8iKzUrekJBUr04HPJkoF0WCWZ5IQ
D66XuffYsnsFUCG49jI0Kv12bEvadOkV9KTVOSXYiN22B7pL01wJHHOV2J09iZBSsW29uiQ7uOIG
LaO8VHzloYfgDDnk5b493D/WrkH6gV2tbuMLuDTKgnyK+tNJPkYYTssmbXUlRAaex2/4JdNLLBmE
9JTIy5AQTiP1USmi1FVJH2SPxluhXGBDKcKomobjxrTYBOxc4jhHVmqnobOR85LFw0v0dffvLsHn
F3lzTymaa9UA59i3WBBi0SaI4lUm2LK4xmUfp+fg2Ofh4jnX0iKLp6ub3JZyihRnyI5fPVk2waih
Z5tTWRmU8YYN7aSE9V71dynaprxeoYBXcktATk0+4APxckfKZ/YC+ttlYu48i9CWdeUGytGl4RnE
Y/Ae5kxgv/LysnZy4cTfXfAU+Zdv1ETMG7G7KODfRW4wSeTCnzRy+JaQwnpJmDV8ShmKGvqBIJPF
lkypKUvkV9/f9LhuiYG4EE9BLEjSq3Bg6mJx4VSf2IOiPK255lERM3YAjRrxPR2Sjntu5u7lZV3M
0ge4nzpm6hVDM61GK0Z2O1Mzx+S3S868hRTrhyOzrpgBQAkz6lkupZTg4ng+uNFXvJxQDCc13Xly
jTmGvb2UcwZ/MvpIroxkuR4No4+esyypXCAMPRWlQIbZNw7zuiBe9JjsjcIKY7dEJw8ocdJnGwcf
pUZG9Tj7VVJ4/fqyghbFQzQZaSNRFw8DvMxIlfr1rIRRhRkrWmJWJ7asbbd7YQy12DZFBxEfOftM
r2qJDAulO/4RRDCBLgrHKLgbkkE0isPml0Y8AdpEg5nJ53OmGDaf+xcZSli+WZrTGzjWk4+qro00
WZ76eRgmoczBSMiLrNsTMCKh2fu5P9y2EnIW6v+dNFA9zptyAG0TFSx/ON5HyopLF1WZzdDzK30P
QSwmU2uWc5/ryUxsnKzkvU1bplQj8LbpjY5SUK0r1KQ4r1cgcjhJOsN76uDRoFyX7Wu5VmOjOzm9
lTcMxurqy0k7pNxAyr3P2kotqf+WEGxQF19e9iDPWuF5kkop+PkL+2owvp+88ZPSqmewzSwJr3Wd
izyp6u0eLiKKFaqqxAYr76qnshZ1r2vCVzQSkV5f6GIgmXM0M3x75anOzpPtD5DgPQOyqp1OkGZI
ybRc6FIvcLXJphq3n3jdBvLIz//iQA5/Vg+orCwqZYeRlYdvGiE1dvr8tRBo7bEqYiQwFkdaViWr
bogJ/cN81By7RdrlnFPQ1xErDINXT1qSXqnmm3LNZwpeQl3/6Xd8gX2MsshfCtcNP5YZ+IKDKWHb
u8k262Y49RNk479jaKrsZGs2d3+IC8Xr2wgxM5VV/m2p5FsyJHZ8FHzZIeLIvaHI818Sj8T/P0jy
I607hyHcu79EmNzm0ALf77ZsPD9Isu0qiaDh3XMG97EZYGDZ2cBkC+oo8UnCoOVBdzOCjHDgaE1h
mGnbX36N30LbSpBmio+J7vblLgPO6zAGD6Mp23xmVnnkGh/o2Q8jcBOZy6QnT39lhCKNBSU99GUy
d5RlgkgxsrGy6cvR2DFJFOn0P3hopVzomZRORAaZzAAquh6anZIbqVvw5z488pcO/FjpuZBnPN+x
HxZ9qyiSAsCovm3mnSWXLqj0NEoYSv0sP77G5x6miZTJnAKw4eAIanlnXh2mwuvetXgvES0yxBXr
F0qp3CP9GgCIzoWNiBzhL8rTIV4bG30FEKKPvpZuLNnfS+bD5hJZpAwmMY6wDAAk2rXh5FsbThoJ
FyO+BH7OssVG57psPtf/ulHPNHNimQAVRWDeN0OTKTVRVT3j8rrr5b+vJUgbl1MTCb+hMFQFrktX
HhHQioanit4X9RVPlD8IqbCWURys6zdUPkgU7X9HYqS9UAfGmI8tozv2fn6XpfrMCx8J1SK0jdNF
/wrmfQ9FOHV795tq4iIPHxbXf6TODQ+DB5V/4jmsIVjY+Bh2MzESc067CMBX5gANRr5b+1rZAYE2
7RhqorJ9eTr7LsUnxTZ6/xwYrIZwYZ6PiO6fAarSTDVffwhunQsRwrRykpiunS4Py5BuAmxKlHtp
mdaOD1NHg32t6s5PP5Z/B6wpTWN2vjAV9oFu+OkP6ETH+7l94D0pfsRNYb8VseG21DvESsxAudxj
fxsimMBK6R7S5bfc7IbbBMwgwziWnoyKQgyFrRjg1cGjAhjlRUM0zyRbSJy/t0dABpFY9YiGMKzm
f6MNmtxrdKXqeomsg7W2jearX1iOKNnibLadW/nvm7rrOeGVV1jaY+DfLwcuHn5IK2B0X2inyqF1
umZ7PjwKzmtYM9Y7vsOSq+bkWYJ/R3SoL2EhH+ofdMERW0nK8aOEn6c2FWi71KXRPnh8SE33S9tT
GmOanqBIfXpnWlNaAVTVzxOYMLiFuFwuVoSB2gj2OvWVgJuLO4WYc8uu4IWkOwTx4gMQZiPkR6vY
o8jLfhpezfsRVpSsVlWUTSe0AYeq594CR3a5ULyNxgxM1chXbInuVvVqjfQIIxqaQd+zUArsx0Xd
pge73vZScaopNFxAA5sfykDrSDl0tw6j/Qzfyr6LT5Zz95XRqj8Emrp7i+LyoAGFm49Dv+48EpKf
xkQ9nLwEwR97KrTJp/bC9nCDvWEkc9yDs2d3KDrMK6wa0icP7JZw3oTjLeMewCaimXJ0HHbtJBxs
H1/dWFKpBpGi339s92uPulp3W+s2l8qwoIW8n0/zu0AKd6VDiPE6LdN6fgQscybckIYr6ljdQGDf
HHnvnX3NYR9GWYp443dDOspqC970h3rb5R397psx7l+K1isgmhHFdWbLPojlwa3WRLmccKNmbKD9
jmaTv7jVOOxsWurjwMzClmxS0aihwGO4pPzJpxYVfe1a7zwbFx4F9fs2xDqQvAELMaW90XcK4ifC
PcviA+Hp6KSqS60Y+VfFJte6lb/97tYd4/8qAL0yZV3gcjBEyXaBdoo6JqMpmaAY0BefAG7SP8Iq
4hDNdxVnqFoLDFrclL4zxCYvZPz1jfzjUzC/Klb7K91TWuFh1jUjuU/6vFuK4mah18gGAw6wexky
wgwhF2wuwfnjsPMXPRBD3awFb8kj2qy7G96eVlYXMifVN1uAbTlBF/RzpK81AQqamAAuYgdnMr21
fFxL/o1H+okeQN3rPWZ8cR5ymcxBMu5369rqXdTtd4CUkjaQj3n8sUjGLx86Nj+lpDlEqo6oshjp
kujM3tZ1CW0g68hjzggyl/nvLF6HhjSpdaAd7lBFYNwDXSep5JSvqnW3tJ9pQ0zuQAwSmJOjx83Y
18+b6R9IxekAHh5mp9dyrEX6T0rworCk2MQE4QAqrO5J1aiSGdDgcd4eirUbs2OHtCV0FpruDgxR
2i85kpv9Q0ILm1TNpGplln0kMC9nP84dMCPQJc4BOBKNkrk+qWgAH4+2x2zDA0Ltjm1vkeJehyBU
VTbWrtU/eHt+m42VR2LqYqWkQPxrBgMXAogcEk3eD0GN5SmDG8Hqo43LKnqTIqLIbEbpuQPAshkw
SXnOyF+wDFEUtzRQsvicWcvrgXwDmnuAYPb5c1p8zuEFRbUQKb5WYA+PCg1Gpz3ewlXD+bYSPlvM
TTaswCXXbIO8LZXmAxjuQCkm1BIcs5YIAMK3NxjaNFyUjBL93sDZvpaCDcfITCApq+iILFDuH4qe
ZsCfB3zid1uujXYI/TFIzVlpBPKAiC0OawW+vEucHRtNfAEEr9MRIhimanRAw/Dw+liHprmkEMOA
mvJbZAEyH+zb4A1JDGVEKm6v2gzSpdz0Asn/OEMp7B4TDFiePPbYLJJ+nzQKM2MDido43sUKoa5h
j+MiXmUJVNyBtSs+0hG6kbdIDSpKJTbDPmVwShGBmvf+FMuSqe4RH2YqnAacMpyIACwphtX1AaDy
oHq3ebS1S52weCg8bMmwal13jeXkAFE65xsJgGnD+SI6A0MUZJ6afF9aDtHssn8oDaNs/U7VXUAh
UKG4v/NiUQcsGXosgTVtqOpQUlhWhFbKm5DtBy102SWc1PImX5gVjEw4QWajSCXmD9A2fJnNFEL2
3eZ4W4JSL7AFovhCHCrKN/lly+DJWbC5yuWQ17n8woNTVbR9DcSLpDEz/RTIxvkS+Q9dkRhR2BNQ
LVWCWJOnqzaBmN/VPrGK/JT45fLRfQ5DlZ81XklK9t+LHx7kcgEBB/3AlpWVNy/CSE3TYGg/yg7l
MmX2BKW2NYvr1hb07W/8URnplUgJDor7K684lKlytViaxn1UITlBG1qQFqanTepMqUsHZWzjFzms
01vDZLssF2CEPakUMkG5dknZKuE+amOwbmOnnmYEab6ZJjIdZyNCbtMQUeK2FnnR5NqsGvJNjLG8
5ocW+hdhUB/OZ5t8lReKFOQuC8v5tAlNczsGuO2eyyrW8rDkKAlk1ZJN9rJVzgkbkFw8PPWJuf0I
xMUMn76v4VCDiTBdnEo8mEP5DHC8R3Id3k4eKsrK1E26S+u4CFh+no4lczAbVt9nmhuJ1ZPqqziF
A8DXDBi8HR1CPKDxrYTK5LPJ8pu3aseYs9EMJZti357O36KCJk1PbXROmpeQrKzHG1Qktv+wciWD
Kz2XewVy7K0f1rBxcel0WPkwIV1Y4Qw96WfnjPQDc3474ewbEzoyBMWw8sTciGX+ppCyxo1nCseC
ukCBlgWCuUKOJXIQF8Mp0y2523KDe9hXGVzQ/ZCsxHP391dmG5FFrOtlk439UUl7wWa1Gyq4hguY
ZF6qwFfzwCiiRTAYMQLrtcmjgxKbk17888iBPM8Or6aRe/hhvpSuD8LAQ6tkwL9yqIQO/emtbPqd
T3ze6vhI0HLKXjcHhSfIuwhRXP2iWAXaRWPlwATmALesQAhdIjsbSPsOdY9cJT7U1hKA4j2Ly/HM
amQb/qRAYvZIc+XAb+yPAzCmFwzYZnsMXx2FEgLKv0UI53Y/TPVo570TjiLr32mraYmvrVGOFdSl
C7Lm7/KeghkArMqtd/pSjVp0PquIREUUkaSLua2lBSg2e5VwALP+Xg5tlLtsTYFEQkkDv6mgJ1FO
zM4zT347UBp0W4H+3LSlIGJqp4ia+hQyGUvV+zzJ3LqZ6lPHtYF4mWgIbr7O/dihXArL12Wm3JUa
QOG7DCKGvZuKIVLJaZisO+mWLw3IJRGkfvXrbX5RkeIMNlHiQZjbA3o3o4rwzWGWd5gZSwXkjtgM
MnwlPoaFTPEyIkf08WaziDUWMvuInnDzCwMeMwFjCqLg1dFW3mpIbkgAShiRdmcgWNwR+LUwjcNX
VVdaFDAOar6yWdYSCfCBc9xxjLNuz+7XBTT+rfq4cxDa0UnlmWC8Dy+d60zPI5CGGod/w7MVdCCr
CUiIxAPpiyfQY14dAIUKUfheAc0qJbHvJuVp4oZvd/vEaNwblYp5GKNr558V6aGWjQu/bpxiXL9P
dog8i6NCzWcIfUEIQhiwRunWZRgd92qBcNwkpOx1sWkWLKAAeZu5k6VU6A/CmcE7x5uN6/ei2S/Y
cJ9qv7oq2SXuSsBay0uy/Q3KbiH684EaXNi4mouZA9Sn8Pj46sYmrxJRgFAMCpmsPi/b9m9adct6
KOohe+6nV5EI/Av3PHqaYNsTSVhgHSAx/lsA/4ssTHyDjaVO4e8KaNU/QMnWqlQYFX65YGvXN0Mx
WOKhVURSAmwuGbkQ/mJPP3BCIj906ZMSVdVbglidXTCJMEGkzxUFF570p26/JspgDB5fUhSZm27Z
hC/eGFXeoojUrEu2Dhq1xZx6S5ztCoMLJHDarhZ+nSYqML6tzjXciGKv02RoUGdAT833PG/HfhQ2
5c+3rtL32z3o7vwG/UbrMFvBW3OMk0MAmeWynuJksSnhRzZaUkK/N0sj9xOZFIKLfY4PHsMeaqLI
vUENYPjVZ4LwG6L5k2aPexMugrtVvltvB9xYB432VpB/MeqUxKOqRq3sOTUEfrX34dg4h/4YPvSh
1uxrVohar9ouoc0mq9roYegA2s5EdwK5LB0x0z0H5GYh2Q9tPaD3LWMpDmGdm76sTeMfRnD/DMpV
mkTAZavLSPRrX/tg/OWCDDXfhldSFOyqsep/zq7WshOyHMzIPhGXhM1Nz1oj1WzhAImrxgoy1cD7
QzzBKd6vJ6n+hOjk4adui92SE0fIjyR7D0EoQFprNSlaProeh3TMMMKqkoeOgpklz97v1pfH8kMS
0dDQpvX1biUTBn+Q5xAnP+0cItmYpICBUNxVBgYNgl6HoI/5wVdRFgsuYwukY2cp+AIDRZWIZWS2
dGdO960+2xMe2+TprZGUStDqU/dwchXV9snnM1f5ytTBWs5JVRQM+MkD2WOONRhv/jBg5zdPv3by
1BAFixYf+hvXtaMn7NFBR58DPLKCVMPjRNuQ39uuinaNssrKatro1TRfBNARqdLxcry3/jZ574vC
LWLSTvXJV4oRs+fQtoZOhHyq96YmG3OE4ZgpkH8d9/wDrLbWBBX1AXerqFmWlAVsEgeezz3ZOr6d
wF7Ucj7t8eWXUEm44Ah675y6BKIUiwEmAZiFru54PVtqsT6r/Y2UHF31Id49ql5UjCpXCjOLwPKc
pBExsjs4Bibziv6nNr+WLPB+DukcYsYPWc7sb53ftTjXVhFdOgYJB0j55Z7s1OgSXBxcc6Zbvzx0
AjzInWfJEztmaBIz5o4ZiRet7lRKjnrAfGXcVGTUjxJoDx7ep1NAwJQeBczqsh74RC+NU0ZT6LZl
HlGEpP6M0KG3g8RNWK7rxXpCC48Rdi4lqbXDWF5/y5uoSNbMrj82bxPL8S7XBxy+21JOCUwKZtwK
IFrF68MRmAILRFW/vLEDNJmxVbFqXv1GFNhEAiCdGYL3iTMWkP3y3Ccin4WoT+qe+EEnHDWcWA0U
ndnkih0cm6FWUBzJS6QehzUq1//uQ0V1ALVSjNv2ttsl5m1VhW8+MLJ/A9fFR5ZPHblMeee1zU7N
4dWr9wIP7TOKc+VPLIPXGpNTdjSg8fHj8GjN29nl73SHkPzdIFfMu88N5uXDMPCA4nMoaQM1xHd0
MAZw2GmhsZd5MEbFXmQENWSXN2Q38rk+zXKEolXAM0anXj+UeWttr8KOO3ABbXpZx/R/ofyfqRku
mcricn/cqEnYVT32DgqjUUXfUXxtija1oRoKfRyihEQGOdYIxZYW159RkddIvY+2Ub2Yv5buKJmk
YGOYkq5cUHGBLOeN1Jn8DIvj4p6CIuXjy/EW9V5Ni120YLXalsb1SsOP+c93aJ5uDEiSKUMfdEZ8
GArs+ES1f8bT5vKUi64AoUPlJzGa4uBn8qpuBO6GzpCbemkMNn/7Ufqkl90lIWIU0Uvx2fJTuNDh
RXZlJ1k7APePZLdXZU6+seRBgsBdZBhzfngicGA1KFI3hvwvBV5qmByUD9md4pOeSckbqhO4/reN
Z2Woi90sbynSWTp4Kqch5XA0xfA6vAM2wi8U8dt3OYyUUwazT8Yp7/FYYQWN0bg+1vi2lJxlaln7
hzd/gGq2GTN0sH7JXSgsHfXojysa959kB5CL7wpQzWrjAVmiy2NkEbbDqbmceZV4WvN07eTTzB2u
dwptnrP+nsvS00uKHLH7o5hKt8mEJz/zImHFo6jRVAfIO2vYAAeBDwQAxlcKBgBGj4idACUJFBzX
ZHIyyjvgVTDi6x3RcheVSSeOlp9B+TOHbSawRefHycAPA+vly7Dbqg7aF6ljltqRUT8HsBVHjzoi
UOb90+ihYwoKY91wyEoKZXfgS4DxjNSFJAD0nAaqjUJewVgS0ltKiIDxoRio5tg45biOyQUWLGZD
BcNEYx8EeBMrUPaF+fbrIQqOxRUPwGkB8ng9y7tLpRyE/myXULfUpFbFfAgHFDgQ0dr5T7U37TRf
GF6vqDJt3oy4QXVI5bmP0ms5dVsZ4SoPqmGvLv5gryluxEvYd1dmha5ZakFQtIh9F28E+3Bb0Zwl
wRN6agWIR6vC9xqWB+sI6PFQnPsu64Yr99O09D8WO1959oDN/f/vQ6OIxmD0EF10vUR0740NnzDe
kzwtL0/lWu4FQqePF/+no3Q+4p/JdP1AkS7HJUGbh7S47IxAvz6IVzcEnXsQgIC7jZvAPrb4QPuj
6qb3EOMtpy9oOR63RoYMWR+hXJU503rpP/xkolTFxm4+4hvY+aO+6KGtAuS1cOlbI0nPjrgLxbZC
MPZ2FMgvs/euFelhTNGgb+1o4oOacR5Wt3Lz6htelZsPYE9CjcDvjEuhEzyQE0eIXzibwqpRc+uM
DpIO+sQ49KkdJwsdnNZbGXroqgD4sGmjay+1JxIvciPBnC5YbjX38O5HMt0evv5/yH1fPuwxAS3q
K9mNAuaRDbIiAYcJMISKfH2Gt0eX66fF7rMvzQXcfM1a7SGMJ5zh+VfyWsx718c2AXIXIcN+BQ+F
7uzXKO9/VGUtkcEp+SJCnjJ0EWb16/wqD+nQFKxwhkc5gJyCQ7fmhuAboU0USoTwKnoc/Puu2oYK
rQ87FsfUV/QPpHQ7jOMvjBPJOB12WXAaiUDqI64judfMesHPMKi9Jz+Hvfw0HD+wbXD02PqBewMj
MUvkaxdTUEADrMY+gduyPCK7Ng0M4J+C+xo/Ogtrxart+jtROyE5oOBB+SqtnT3QWqOm5D3ulvM3
3r5xob6pHtR9jqy2nusbXkPqmtKHEUz5A1coIr6Tnx+8Z+Xla5Tp+O64oUysea+mS2QY++Ob/9ro
vsb2v8FPLOykwUhNTsAwln2w0gMNNM0CxJHQj5kTHfhMVMipW7C3mVzLfTB7pLzUp1SxqTYZRZLw
jcF/etM7BDIvAG1Dx229gCOXypC/XlOlSUGjNPXhCv/QIZkddUTLBzgkd1fEjjJDOAQHY7dpLnjb
5Ra0pKpu7i66iDGbRZlq0xIAiUbWH8kHlzFsfpSz8w+DFM5VRg7b3157MhpxxS8XDxEvAnXeo89u
PIBBGeBK7aIbWRC53N/bcjacF3XU7AZM2HzXI169wk+idYhUbpJBrDkg84C+yLLZH7CYRDpI1h/K
M1jcI/5soSDsyTCqrZ5lxRSJh9XHsidFwRNA84PtRXtjhZZYzPeD2VAZlO6H5eB1Q2KGeOOxxLlH
DJf5pWP49OMYRYVQTPzGk28WWfPMWnsbpJ8qFYxeSahOAoV0BbkCIWwHdw0oXo58KNqFL3s5Hl7J
Ll8wHj0JjM/JFWc2PHueXkPKdfBM1dnkPAizL0kyYjLFhjUD4jd/cnpllTb4bcxAlYnoFP6iSL7V
bchyTnyGNu1GeNuXqtKIsnFzocP7q3WoSOX/oURY8kWtKEE3avhcBJE/cshpbfM5/ZncXh5L0d9n
zv5yuYuSau17FdAjgaf5ZbmyvHE3UAEHS5b/SSgFTacSBWzI5FqNDSYzB0RSKGIia32kaiWUwxbX
xcHoZ7PaHgip+8GhN3XARImH+RQ6g4t7R1Vyk49KKvPJAiz4rxGOsfvM5RvDcehpLyT9snc4+/qU
t1nr8aJtEllKPmJOcvbUWSqpKNqQBGSirW1e5hP3EaqCzoesS50uL/ay2hA2UDcG3EVoxdQNybx8
VIr9bAv5HDnrJaVFMT5uD7bJDR+OaTlv82ijao47pipviDmpLATmkpZs8Ojme+ruLUdPkdOFhf5Z
UmvZPgYoJ2dflnzshFdJtgTHNAcmOq3cpB4U4VoaNBGCZDZFFbhfs60TeaSF5Asw525HH1FRUxdb
oaBLK/POoDxsIwECbw2i8WdNtAhDyBimpnCQ/MVavp5gHGYg+boBZYVzYpZ5sKxcKdycD1xd2DMS
DEyyFjxBq+FNPFYiA2oKwA2awLwtbo0Xi8p7pzjX5ek75ZAZdjtUyEkKtMF7+Egh/8b3tO87FIHc
IP7tFmNtv4CqcpLdTNVSauJttzduGelobkDSQaeP7VdqJiJU0vW+2czLYqNmEXEPuQAQzbUh8NRi
rmQHYQkt5yJ3dt9ELFurl54ISfX0S8HVasz0dX+UHeNwY+fjg42a7e6V5tIkyk9wCXwuYvg+pyPE
/E3pBRQpHMquCE4sfvohd2a2dqg1a7udeuthwsHstKdM2ABgi5oGG9ryHR90DataeOOZ3IrQlreJ
64Wz6A+2yn3Onm2x8+/DdS0dn8nqskLMoTFylueMUAPF9DXSB8lGlqaAYxpWr45e6Sk2T1Hckn4W
oXuH29voEFiJLGLOqVqkizTKP48XMjCLOw0waFVo75474YiQcHzFO8CZLUGyvGp2c0TZfVYjAHYF
Sf2cv5SE+YPO3W2vjs1NKbb9WKeai9AMlrXotACgfqyxFUkdpUyjhkXFpw3e6Fk9HuPuXa5tGBy7
vehb4hJRDwMdBDiXfVHi9eHAxL2xX+Wd5oEMmdtHTktviz4y9RgI1dhFyEDrx+bOM+5oYNzzeex4
IS48MCqMUkMVxvVTtLOJkadgRlCuRkl7L5E81hKBiFjq0NeAuyqVuk64nPAhiFMcmgsbmM6BA0tJ
ti5NA0xU+5k+fTb8yATXYjopwTSCjoiOFTOGL9QsYalk81q5wt7MtqrrLjZrV8tHV7Ha6aVk3oq4
yqReEgVI44jE2WuJ2Bs5CgkXOws1TWOSUPilcb4CfPp+5ZihII2HHaPiq/5rLgbtJgNGsNTo6GUZ
QLZ/ffyM65nFKW8gFO1FMcHh93kwzMIEn8aA+A0GSTyiLrShfCKlgwIDzAJTQoM+udZXtjm2VExW
XTY2nH2JBwOn//qwJxQN0KFNwOmcPbG63dIj2Bglt6NhI1OsJVRH/N6GLHdN44pPk3+WyNGS5xQ2
33FWi71JUkMjHtWP1x2t9ATYK1C03nOdILKCy5l7pJw9GC2saCAs/RRrt/9HaWGoDlGDAJ8G5e3m
ajQl7LDaywAqDT4nt/FxgHm8sDIQBWlyjyRi1Mgx2B7pAFy6wA1XnmRbZc64Nxjrslpf88roTg6Z
avpDUZvadmQ4NoJ4B4FFyjR6Ego8gyMCmzLg64cxR1HDvaTJfunfKHGScU5VYT0vRTw8yOHFVKYy
x87mrHq7wDv15A6lsm6i3Yl4IY2yDD0XJUFmcSjDgr8Y8c7mr9A/pUweA1EPIjaxeG5tZ3KtTC7Q
U0m6Yqq7r/W+BIaxPryBksiuualveTZthqmBFF4N5DDOsT8a26sbvkrkE1JX4wU9hLzZSIB8E3Z7
5gSe+TE0pt2f1iaf9w4RvhegdfVygD/7LuDY8colvO5SgIDUNAQNrbp4zUyip0bR/50yAKcHpiNU
hKpmZBlNInXM5/KU0GtigtR1PHB/dw33eooa2a+Kfz6wkf5OI53r3o77N1AAKqwdnqD7Uf57Y+xk
46SmakpXPDmmkpBW4RdTrg1WQ3DRsKodft6PufqS9zgSCOShik01U+0CDgY1G73IsfDOb+aTxFHd
2jT2fSqCGJR7xEtFKiBPiMbpEOgg4KuA/jf2XghH4hSqC2fsCNGogV0SJT1MInJ5E6joHb4knnIh
Bo8xcap8+1rer8SRltPnTa26tyUrXIhUAgF6bSPXO7Qwwpvx4UAIapc+UgZPD03RbC1e0MKEt35k
ZAhG0GXwo6VDNtZzqp4/6aqen/tp3KTnnMqXG7QmHANphFswJn0xIxkLAudeKveV79exyRg9HD1S
uESQ5aYVjZozC4k7PmJuU5zj/ypHvHozxyUx0t8GxpkHVFPjkEwShObh9/Sy6f+AnmF4MZfITH5r
PZyxxKFU1nBG+NQ0aW6p2SJwxuw3leRroV6La8yFTmKcXZnZSXy8eXvFV77Xsikde0pDHGlLWyZZ
J1t1NmSfGJuOP7QhVaWXKuIu7CmHEjH++gymwZ8ttwdG/FUnpms50AR2HxwJgUk2cavYj1QrkZX6
ObdyGEld782OxvcIsISGimiJ4HZ6wpA2iBoiutP+Sve+nDeEFvdlxRcPz57BmTdTg7R9QNif/sv9
WqhnDQklZdwnl3XswgjSoSZBQ340Uk/1SH0VFSgyNh94cxVT6skIN0Mlo+zuN0wX/K9zT0/KHMHA
VthV+JNW09H6SD088+gdufTYvNEtj4FV4N00dLxpb9ZcS5M0yXIsLEeCMlaqEC8x1OtHWwSPUAc7
FDpGtaimIRfpvAua9v/X43OnvmOqH7ied3cVLKU/zRut28al6j2SDjkNEm0pLHN5aiHKP+PbS7gn
scNlZXZl7J20W8Q8Kc+C0kYWOyOQc8zyaQkNqlYTRp7GPOzK2xRrIlskkYjxkeErs6qWEIJpNMqe
cZRORNFDTO/MTwwrjQdsHBLJe/9avr1UaWS+xOkKVu3nzqWp4jIeyZRZx8A6sSErok+vkhh+FCsd
sRkHTrdQY9j2LMm5/6oXfncpsceM3fhWQz5x+rSLY3b74fSXgpPYHuH1hYxJZYZydBhPSWKE0ELb
XMn766u1Cnxmo3Hob3dZsFVD71XtyoBcIkDGPZp8Qch5HecL0YNAkDCLhAsDBabOHOg747KoZv86
y2unypKTCbxrIs6YEJzC4M21Ott9NtSwYDTo6RU1XGdHdkou7yJij53/t3e6HygrTuIzlQZHKi2I
GEgYpETu4hrKXZXN4HBASEt/Iq8kM9aJm/ezZbCvLI+i+EZ4iXBTX6+ifylEjTrKKMLKh85iOGr6
vTA7KV2owkTnz1ek/wt4IjQMbE6JUPaQ0tU67qb27EuZ0/zsdZyAsgTyZa3Dp8f4wsjdMFmVdUYd
K27bhdbcnnLGoTPvAb9/0TaKf5CruahKu/g8D8HETNc4+pwYB8SBCFOH+6uFVGKmKFk61uAikkME
6rRVtVzDF/aKTffRR8olB10Vla18hhg/3IeMEhfgBZppj0fSBUog2WH94PCRQ8umnISsVXA554ZI
cXo/UiWyTxTp37nKyupBMcZcPZFfXbyvGdG2bN4GxlnaAEBN9HXbHhrts7kMln7EaEpN8bEOMmg6
ILdRL19VFVnyMVjMQkfXzPHBjSCh7b3Sb/v6ZnyWny+bctwbuCWcNPgUmLUKUvfguccVYNsjZqcC
yOmFRZDuOzsP1zxgMQbDo37RTRWdJM1fiEMSTsNKrE3Ru2TSmYzrEGH8a+QeTXHMe5hL2LmmNKJz
XllaEGKnN/8+70w26hvXQLXBXjRXoyopVWYWRJHlf6dmRW5CywmnyYDHP747CmFRuQ44dqHEK8Oz
Ij1Lqm+XMr9rPZUZ4pl40bzIQwxU30Jnn/8xgZ4lXSDPPI7GOpd4PrT4F/Nla1GrnrwLddwc1bqr
Dufk0CV686lUwf4/tCK0Ls7vf+wTA2zU7/UHfS1vPTpXprIspCa0PfTLRnvSF285eNhmm+yp1oam
bW1weUy5Y7DsI0L3k1OquXnfU94ev+Fa+a55zid4JjoXsiz9qm25Rb0rzphr8g4KfVyYw6g9Ez7g
sbi4l6pqbesmFvtjnFUA5AW6ULPysa2R5RVnkYzJeheNOOsxRR26mnHlhcFAbIqUSJZDluwbLPX0
6oNVJgVBKM1GsmaDa/2Z8D+8j4fldpxcMezFqeljmfcc3VFr51iluy6iGn7hqGGmo08Ieq68UXIV
JyRpY5ZUHyqv4FYIH47bMroszgQ5bSqNzZwZyj2Rk8Wa0+1Z85NYk2DGS6p4JgqmQ3z4ck0Yi6La
Zl+IOCI1vvh+LOuxR0WeLgmzoWta+g4vpdyMww1qTiQYQi3STo38SuOZws5h9qx4nLWtpi2BdPEY
jAW3xUsPCIt1h+e52Zry7uccewoYT5cpNxi3+dmqhELMbsj+1WoRnElt7vQ/fe/w7tz2UVETT3WJ
81HeomgXu1y9rnOcXrq80Fu+zkphjGR+CcSJ6yGkI2M6Uhz5z5ORYDoB9T7R4aKdbMt1xDVMwO7J
IKYXa8PZsbUc30n6dtXz1RiinsFe/YL+FN5TPW5EzrLO6XF6FgW7lETOqOTzVQkmUYQ0EBJ5wAbt
yax65U5N2g2Mzg/KDMGN4BSSTsF6PTciF0qV/w17eWWyVAZdkOlxbkKFKGq/Zguo5JLaQUlhEzfe
jokT+QKRsh3qe/4juSJ82Eh7DJz6w9iqOFX/ci6X1sUHUD4wQ3icwd3ylL21mQGRey4nBT58RzPB
u49eEzF3JU4WlwJmfBdmgXscswnm35SSmHbanr2t3ISXmv9Ujpu1wyiUspgrK0YdNKiBAQ7RPoav
wHleJnypjwDpgNJ4G8Vbl6cY2/KsHBRTEDyh9XdnMhAOjXyw2hEFGgxqUZZvHNZwm9sF4HOmgAOE
EAYRMNnhgiT1/WWkJ7xOdwDjK7gJNiNcDZMDVi082L/g1WjKVeyo7WuJiE9/Vv0cWSOHNj6wDEX/
gLiO6ObQWDiv6ot1rBqn8MTDo8rQjI5LrRItJG6evFYkuY4O7Kp58dEGLS6Emay70x75kmGMEwTr
+VAkMEf48TS7V3zdUq7HbxJw9qHvM/Groz/eXMqMAx9am/eKNvnma5bAUhGzWSOr20TUyOp/fvHC
uyXJVQ7igRXYgL+LTNRlWuebMdeCOn1gNyzQVmNP4NGzlRS6KlM3t7tF54FDRZq6tqLEeAyo1mZJ
kafxLdD36jhb8a3t8vd+fmhT9qMtomXbtOMrI5eWRxMXZqAHpUmaqGzaoOfSUbKrxXU76fcxYkVd
ANrZFlQXYmRN0lZROIR9dbNKlfEBXk2Ym+GelLuEyCfw+b3JV+C3uS6ih+HPyg6Z88qKpSqmX0L+
yu+aV7GZrC4pWnBN+mCMRRh2OrTS2ZdQulcD7SPXs4K+mbEfSJd+fwLvZLGRxkcGpBt0VhFoISBg
p6tZLpNkiQRRMqrEcCqIPeeUDxIXI8T53w1dgiRBqFOeN9qYr3wIGtzleyUCm+Mxb802CldxVcPl
z5CVxfyZ68OTaksGbDNSFBMYBgjQL7J5JipKqMu5KrnjEA/dc72UjTbZW2AqvhRYiyhiHo2LoSP6
qVzKRzJvgPkbSu9umhG8oZcl+Z+DcDws0aHhLmsq28j+z+H//3wj9QvRYVUdtakjg2eWoFNMLA+A
P7YUSFV63YfSC9nzU/p7Dxxir7dvbxKjY51SjsSs2ffO+ihS/xYhVzqlzu68Qmf3FFSGDpsr+eqZ
40LWk5/zaylRFc0Bxk19bBTMN83/YiTmJoeSz1UIXu/iUUY7bRFf42p1zwahcX5cu0vFlZqgC/82
VoOdv9mUPjDwsXTeB9YTEg9BPm3y+Dtbpb2pk4DDi6oH9uekpyp0LMEyuwFUWJhbXEXYtYwnu3x1
+J722NsHU01x27E82EJuH3ISpCuYl1/9bh1VcBYp0Ym+LKMa05gdDEnipFzDeZN6bk+VwMuKOYD9
TUCbjyCupT7c1dViCcUXfe/ZZwTgvuvlXh0WvFqIecLnXlHhFYUXjIA2+Z3UgsAMTJ7h/kgL6bRC
lLQui9iOB+3XoNjb+q+AKUxFDpAOio5qzDGFSWrFrjTqfFWIWBjKm6BHwGgx1TkR8xi7ou8eQy53
RvRDAGXRy5wlPauN6KchppZyPue0qYNkoaHy2Vhy7aMM1CuT2nQDay0ryeW6O1u5M+zzuc3WFwde
JWhjsHEq+ESXhRYbsqBf4hM4Kz3B1CKWl2TteLVSkTzviw9eBOpG+NhCPOSuWiAKkNIJlbUlqV/g
aM28W+LX5kyt4+DNS425DRwtdhPUcrA31ASjdBp0AppSEPcRax2lcFjVRZGuzOt84m+VVGzQV/d7
yPveCKBkU9Y6TVuW4DIixoAb6ouzGigBXtnMhsdPXgj5jRehmLRHqXVQu7lepFLF2lYRrz/IvFmP
khhCSwCMRGojQi6ix1XgJujwq4DUawXhhio1tWnJ7ZsZREK/w5Ldn30vXxGree8GSN/Z33V47Iuh
WkFCt4XYzp5Oob6f2Hlr1vcIhHtC+58BDsiU4ylavapd1sQlferAAN3gAYZSibIkdc1P0Ry2/k/X
3Pjhz+o5/fvlByKkkDqcebf/YSes8ybmmSv+IIgqgWW13kv1YAQB+tvRWrtg+cRNQtvPj5+qUqpP
92yUWODUwKLMd64xd6/hboFSo2Ch+UtY3vAGnE3YN2otEGRc3NY2PenzcUfjeumSLcGQURlcIylA
eZx8N1SIzjnTM/d0RF7rYazjaSkz34DeKvQZT7iOqwu25KzHmi6rrhNDVq6MV8GIUWIcadLeX9De
UQffHhhjcnjYNLY2DwGRX9VxJ3fSv9o8b8R1zAPVi1ylSBIErTNjZO2hX924t6ghpV2PMrA7wcZG
Z/SB/SHRV5yR130aqS3gvms9ACQwI5+teesDmzioocpVsEO1Hcw5uqXXFFzXcceSqXcQQ5aDte0P
IBhurTuFQb5BfPatiVAZU+G5/bR8NFKd2BPv9fgcCx17FziAb1bJWUYXHSHDzB5Q22vA6AsUahbE
We6YkLQknWDUwBPWLjzvlgIsS0XK2c/60NJmgzbdH+4NX/SqyKQ1xi3sc6VjcQJMbNmZopV3+lEu
Llphsyk9Onk6laNvHgCoVNlopVRJCMAclI1H6eWTZaNGPJQsglnseObz90AAQx2+WNVvYPfQn/1M
3F2cRPuPdJgY3uqt7VaI9BJBA0DeHpnk1nb6A07AaTDqepPym1KaOZsHyvqMlWdoQ08wtqje63Z8
wjBYUzKlo2ozjoZMYxzCL4eYpBxY0fUiVge5oyPweds7dMhqKjdYCi98N9FjE7UIvG3JqM1so4iG
W/K7c+HVaaezUmSzcU4tuOOQvp+HQqECYQXpigakf4BZps5B+xD6l+1d7oiCZxlejONPPEIJk+Tn
KkGOXJJ8v8mS510SMrjBPV1PEFtSvWKkl0rG7DS9sqEZNrs+fRIXbNb3ovayGuSK+tAd13bdAAed
iX9QdnYQwrGCVUZ6XJksKEa35w56QA9hq+RwrvIY654UdMBxvoyfmwnWWW5tYqb4I9Jp1StODxVK
6pwxJenBdAi4+Y5y5MhDVXZEa4XBOtso2GcSIMTvDlZ0xaI64Ua7j5vusfPqIP2YY8LkQxAoL/I0
lFk0W1B62MeI3FfZOomCKRV3d38dM/ENVGs9Fhl5qr1tZEHaG/yFpWPUmltsWacfxq8pvrWeLQ2g
OIb8zM06PGOWMofB33KRqSeP2Ipx8rmHUAleGTY4wVdSClflM2jVNIn2DWeUXB7+Z2VIUkwqFo7f
Ie8fl3h1vb8DGNf01XtAwlHSCvbyVJ7uXv/jji1uAN6K74J4oN7sddUsU4EIueVwOf/rBGU5sn/b
9qEn3BYxCVfaoOZZOA86WqzuNtm6LSUIrVE6Sqk9SoohLegy8tg+4+zXGQn0f2DzpUE5K/WWQR5F
UYm2HjcdP9CMdNpaknY4sGfKWBRy4Auf2yJoXgT8D3wiXimV1pu2Aj/0E+pYJ9o0ZIrgQzT1CCFb
o07Nc7/gZHpv4KD10zOHlsdKjrhMPW7apiG/KXiwU2NTkt4zvkYrq/sZiM0+z9bM2xHIQuNvCVzT
G4fFi2Hstllj2ng8xye/+WgomnFPFu/N5dBuadiYlmNJvDhZEUTCiNvwKzaAgdRANKTXxeLbWJS4
xAzC4EYM/iVVToxx9+Fg0ECKZQeWJFiT8dCI3QknDmrxbKRuSCHfhOpMBV78zolAD6bfbTKrkC7d
Lr3/nT6pm6hHEYYpt54HltvyaY2aZvdb4O+3kMWhMcDchDyIDFMCOUChlQxZ888wMf+ggDsC0YyW
86s9phhpALSu+64GmmWET1QPyM08sJYKWsdCpGtKn1ItKgUCx0Vm+HB68kWyCoSrzb2c5qvSPDtk
PLxA1pqmX+TOWO5hEq8be0PQRnZP5G/osxCALAi6uuIKtu7nWpS4KUbCv1RjEYkCbhm2yL7zSP1e
/SyXXsefdxXfqPZA/AZVebba1qnV5Bq+Jic3niD9tzjt5JIAM/aiufoW2ytqyQVIG0ryZ6BunyTl
uZ4UQnHkbaZKCqqWqn6F3+GRN2hCL9N6CW0iwhmEb7DI+rGEFauBC6nMOrhfbt6CPC820bHwwBIU
J6I9LQGdLqQxRVqxOl+HfH20mCK25I9TX7IxtqSMjYMMzBGaOjsCKP1rxEPh22uvGceOMVIDqT0J
edcsasITltyO+22WRrtiVMvCfEo1i7vQ/qGY818yu9q2FmaQoL713Zyz/pY7aXJtq7MR8fdxbpxL
kJUHQUiAyEv2vqdyeCiYbQ1d+SkPx6CyZDGH9v/AdLFCX4CA2tYZgLA03tDQ/h9bAf9IBcTcY9zx
oT9EFrhiUQsLrvWftfIgfV/oVDB/6LsK19WmFJJdm+W3wmFScrKl9mODJ7vzv7WiJx27bn1tZkc1
zJY2Up+uGZvcvuP7EEk21E8bFJkUbRkM0xAy1idZj5XwuosD3pYAiQ9YtNVy4q9mgpUm7zhNcI+o
Pqlyb9wZ4wDGPb+LOSH1a1st7pDrDU+anGiCNwpoT0EdnyHMbx1tpny0d30YggvbLu+VcdgrsgJI
quwH0Pa1gtUCD2hMkK2cSWvsNeDuT/beNrpEPObz5Q3s7UJ15zks36x99xJISjqFyuZQq83e7D/Y
/aU/FdKuwYzfOyZ+8RERJZQ4gYKvLE4tORkokCUktZFHw3TQmA7ujiOmhKUuEPB76G1AUyAXH1Ly
VoWuA0/zBuO5dgmfkuaKxVEFzfSzecGkWtAQ/j0gXqD4qD079PcBhmxOvJwpdpgesfeeMd1lfaU9
mVrm0IdNFi4VlYLBJO2Eh5YPolVyqZkdeRs7DqkUj9AnesKnKH2bOO3poXi6OHT7644BW0uZftTZ
0QwXG6/XaIFG0lz1N3oQX6hQUifVsP0SE5U+o8+sUURqlEejEGJsqn1RubXJ90onnM9IEtJ/CeJV
osnbor1Hxb8fHaZ+bfrPyUUgcEoqVT8Zbyza7pjonbxerNrW/VSNMU9ZtSHjh5h0wkAQ+xdhxOxZ
eUu4igjOsL9uQyKWKABUxmHGFJqe8B9hzUnJv6yn+gZUGKvVMJoTa0D7VSdo0lEOzwlcifSmMzVG
GVXDOFic064X8HSlgGZsDLSpRxweIlAAtJboBgkMsESTzyxpBkbCEcsD+01EZVmQOPQqmWyff332
TJrvRkEOw4H+0EW2LB9EYsenPTzrcAv80Os8H1qp7CABiI2gRwOLfzs9O5aPxhHi+UUD4awJx7Xg
HsuSFInJiVuYxJ9RYpO9U0HbDFbxJ3GxSdnhG6Pfd/2ORfpOAAp15zDNC2WJMbEHO9Zdh4EmEcTs
LM/Hqtau1MsqNXroLACosPyvdGEonGU0VXAtm6PlvyTCs2kF+bWnIoJD9Ln9BHlSiEWGemlAvd1D
kFW5xnZoyvZdF9vQ5eYnnJGjolDzPwdFy6qjlZQgu+UhM10ZwYcv7YfmeKRfLlBfh48kDHrXSVAu
J4x+CguAuYjTWyx/zPl5s9MVO1FzhuSdmjFBWg0rQtWl4TEF+/TAf+3cNAnE01yGpND5sxLeeVev
bIMEjfcHzuaBD9i74B3PTleqhJ2UBaFV650mFBhg+pDas6qgEpBPSoJr75O9k5TDkPK+/BjJhkdo
2nRu8Hxcwzw2ocqfGpwmJO7xs53tRyAxcVvaaDDh+6exAHdM42Jdk9wjUOon01BktmjJQ2ipWe/A
Nd3HAD/CAZlEnO9UDQOIquYJOrnrWhTu0Uuzkic+0kHHTZL0LHuJnORSTUtVdkNbFGAlPI5bED5S
jUTW28vw4mf3e4DdLh1AKzZAXFxKuyb/N/aJxaDn/n1Q2hz2G3+6RCs9xjmjuShpRMWWK50ISc8T
r/9dChOkzLDDJlDkCfXM94qhJ564tmeBz4wqiYu7GPHXNPWGwX65pXkEjL9DDlsgNekuDUTOubP9
YRcfQuCkXPUK5RXdKDi72OnYBYoEzXcxWkjuKc/PvvnBZOGalHsDVb0haqw2wvFBk6bhubZmqzcv
pEP2FP4eG/af1+WRpV9GE4i67JBCxoZG2vVBh8ZXMS0PHKhgCGEdSnSusXSfogKgc7urc2hOTr9W
cppmgjR1VXESnEHhP/cmF7w4I4dMJ7gycpFMIzdZrUXhCJ8Kqe3+W2DlqnJiN9C/1djix0xM9Df8
ZFIjWt1hgZ7EEhpGNxUEwUB8jXOicEHd5MJApq34k1j5pOuvtJSb+fzob6VmeJaWUptIt5cqua0h
rnTmVsrvNhRCDIdWCp0C/HOXw77P4cUdzvKjjVS+fNdttBUmuBzfYgus0rNoswpKmgvOOLk4TRtE
GfrxPXx+UgRXFotALqsqJCI/nvhZ/c9TvaHG9JLgJFV4okjOCQtrvfiJmqkqqYO/Pf4E3fWBTM3M
tu0I1LKcYQYOiLaQ45seQXvfOqtt3e6tXZWy3oB6v1vY+UtlXwmwQpP91o5J+K2ZIhiFk0/fnuCz
3GGIoewWlNzKXppvKmhxi7hdjzD3L+zR8g/dgIC2dcjIULxGMkar1mMVMs8FkYqoH/YpaWkNGxRV
0gwy3gucL78FVAB67lsCh1Yr486R4PuPgxFJKoBOp+P++rJLM4gpeH6J62A5QuVCun7k10q9kpm/
hKIoP0zi1PoNhoWzN2ZCYYGB6/VQNBgiWzFf6YBpwokshzb+kDAEm0R2pQyeWTnhSWJ1nGjkE4eT
HudP3JiQjADJCLFy4r40Bnn+RRNIBRgBWBUgY1eWcn0PllHrDKyYPgBdAJyifaIgvsnhlNe+1+uG
+aXJzbhmrjkOQ4sHbEXbDS8Vxt6TR7vqsx/XwJZ0ilvjcP+bC4wKG0yw+76bt8jloVUaWCjJryOH
yzQkn94s9FxCpixAC2uFbshlmeMt/GnpyomGkHSu8HmOgLk2tGtYKcM6nWoMdWzPfY4niCgq3p1A
25lZOeRZF1FZTuBuRRNqIsZvCFqWbfm0mAgGIyBPnNnGsj986TNQlnt/CR+jndTirPntR8tcBEs0
Scjrx9FbeyYoIvLnFOh+hkAp6V4zUtpX9/PfD+je+e7CTDHG44u+ux+qrS4mAespAwOYytgrQnBW
+onIQvoADaMYq0cKx021JILpPQQ0l4rK3ok+woajWC9QpZznvzagXAiTWsAT7jl6LbMM9LOgyIZ0
AYnl8zlzJunIAqXHst868hKfKPhJXC33JOgNd9i1RFqIXxH6qh8AWziXhggeQAQRIk/zzjvYDs2A
xoMhW0f/dkNR/arZwDBsAAwRLNoENX6ueHtU2CoFR/4Z/ptohY0s8XCV+HOqVEiNA0JO8R68RjOp
2HH98w68Ntb7BGeY57ia+ZhUVMlOVVgyuBT6eB8y24reeu60LVZazd8UwPSrTzRyTpenITtMMl5P
mBKFuyQsMINN+vI69t1SF11N5JJGVRT8ncgMoWg/ORXPhdLj5ZpUIL1XD4YU+rikceb5s/9wpeDX
5kNQEoFOx8bz+cg5S5NuOQGIccvw0/ur3hr/pFwGVUV7twrX9nsJbqYuAqSA9Ir9ciHPmlnrTRfj
E6dS4fuDcHoH4WV9Q0GITUsX8ksm53AJvazIIqJ3/k+WomLIjxDW3Lmbl/ksOi83HC5I+1N4ZFXV
8/I+cvDvbfALlTIwHySiAKWRiKPbHfo49EphFMJBvbT8A9qS339fPipnoEGo93FQoTtJABoVpiz1
RUXW7pqdSUvVl5lBFOWqAAC2MS1TWdkE94nn1oQSt/k14pRZlNf0RVDcJuuWh8DYo1j1yjeASccs
pQO/Cc011UeszcDVF5yRz5UOB1QApmWbGcaUZy1G6AG/gS4DwavSo/Dd11PhzB1RMwFPb3NKp7Cb
Vy0309/0mz106BrwaUoGzcZiQkUzflYnNrVvpUu1SmJeSMC1wnNqO3K7jHEMRZUibibgAgh63oiB
h1rcLczOzFZbseJ+VQn44z4i73MRyK7KNaKlbDA8XZvcl+c1Azl4526bx4jr5KR9k7w+5m8tSuxi
KeB35OoFzjrp4EWtP1JmKZlIrNRKZQFtZLq5bjSyssuL4UtQeUXEOz7wa2a1DWlov9KrfupmT6Lw
DtywpBLQ4tu6dWRCWz5fyVJ3r/FVBYdT5ASr20g6tNXmEStR0noQ4j5r+KCm96nm5+0m8r4W/ztg
7MU0kTeMnfZ9U/70aJRJ4YatqzkflIgxP1Q3Q7o0wCMm8ZySeeQ3/IBOBzT/CgpOEyEotIOcLww1
Ab1UnLUAX/7iRzSyLhAWXpFajGC+mvy+2MTIBlgSIYwB4iiYbLA4SzDSFnIqu/Ya+yfOncpBCLUD
lh/o0zokQA8w7pdZU+eUNr+kNcTP61s8PUF2W1Sd1qtUzZhXiPIqxehrdesTQcZxUWvN8AfwOX8e
17bIrVuWSi2lLZfAMY4mYhoP59Gy/IkpLFEeo2MEkqr/Gaofh1WXTGmN6NNsw8mKetGkYFOuOOTH
oTIsQMJ3j076LdqKb6r4qmJEv/ekvsgRe+eV4hiQ68kumyCPy7d7T31h+dKt+W2tA2leD3twa3sL
3+eQAFp9dOPcijkJkZu8rpcS7SeHLRoFqksECHzohRW696+Uf95fcCQTg9YqGhx5tCjUTKPLdTS9
eHXFiyB4y/7PoNCdwTv6WQqDnMmwLZhrIE6e7gZWzFK9BDtYkHyUzwD9X+De3nMLqLAux6vZFkbe
sXf55FMVWGu6TxU3W5n7T4JIF8TX1Nu1MEK5aktmvlbxmTWGmrEh+V9Ib32zNQWqksyUcqvZsU6/
Qj+d2t3CX3Vl3TuTi5X/aiENAUqKEF7ofGiEvy/1cH7okLM+eAZtE8zsA/+Kf5s9jlZNCsV+3nzf
gahbRV6bKxgfPQNlOng42ifedd4Vu6kOsq0L9bAvPdvQmNQ57+aHipGuUZFooZx1KGyhqFiWXU1u
Iwpwn3PIqHtxRBkIj4ONM4iFORranHh8gx8sgLjhzpJ5X1FDuuO6Fy1BFwrowYOCWy3pjFIjE89t
oKU53IdYveI2eU0Cm95x2qMhGiQ4ojLj4VHd45uurWqEqFWvF9xFnFoqERp0Wha87iUZR6ifv6TO
qYl9S+a8c0tXA/aaVzih1tgABcQD7/5i6V2kry54jLG6t77S+pBNEBhqnLBbkvUjeyLX+32nuF9G
Lp8zv9S4kquM2pNd5qaytqBf2tXK2xVseVOzHlqbL37xLC4fcXfDt4Lk/HChmSRo0D6iq1uzi+aL
baa551B7OGOT3JpMxsVl3Dhdckh8mv7VxxZtssd7Xr9EYMLk+KwoGpSpjp2UvmtWPLeoqiZtci98
nB/9zb7eKXSOX79c1Ea/qsCL/gflUVNn8xHbuwMAMcxKJBCtESSivervFij0bun6F6RcbH24YA7T
afWcQf/WoVnnMD16MmvVLhxielUQjTqt8ef30HduKAKrvREhAWvbVxKoOPwIHfKNXTEIoDN9X8Ap
Se4J3uBSTMgPpNoe/d1mlnlDIBrNpeEcJTIJw2iPMbEjPMgVqPuLT8q1ekvjopjwVfpNZhirChnj
zcPGIHZCYV6DmH5EzpdK/VrzJlHJQaapXFYZCHfLHvLq0reA3EklWkJTeTifDQRCFTfaHsylCzra
eDLu+sITtPNMNY2Y3zhOGZAUrkMYAIOvv6xWdcKWt3pyWTiSMNgzl0Cg3d/Nw3S40lAW//jxPrZT
SsMa3IaJFvk7PDyNx8C7YCcrgLrVZXkrA9jqZxkkd0nvjYDdoykeshJA0046/xfAc3nf1o1r0d6X
eBKxFyf88MjakcDbwauH5/wFSK0x0ibA5+IAk/3vLMCW7+aUXuLMzsPd37/qyju3ltPvt6KEIkpS
/I0FVHt7JpEnv/pke88aPViqfPmlw3LHUpMcBXglYHZTo6ao3H50w5KIJYBZB2toWvgRnhwVxAs/
Im843c4bpOKM5FimNotrB9teYGQnCzjO2XUOrsqdU7FdJ9fNpAL5vpz+F/98r+r0yATZYhcEp07R
bp5+ljELR0muKqFMzVaCBU4lRqdbQTzMqu/8DIfREiLdSGmIWX8vus1TIrzO1TIu6g1qEjeiZeHS
grCnAkw+sp2QnqyhU3a/zfwqO2MnRn6jmgJuJ6nB/csuzaPcPsKE00JI6/JCHdmmQRJ3T8ZkYIp2
RokTWqsRytgq8KVTm8Vqg2tL5pbodEoOwnWjYXY6mF5Pm5UtIqCRtZlG10dB1eymkT9USVunkqs9
OdGhUw/TLG6eHN9DmywRsW9cHlyhIW7zoNi832zyiUvyo+U0KCDGKR1ltwMVZahir0Pc6ENE6ruD
6apzqYHXk88n6istxoedsdQfRaz/hj7SPe2NPUvF7smyYMN/FWqvaOKCPu0aKbYLozU7N/663f38
MVg1eFOa4lk32X6e7D3wbX5DxURKibf7NDkmYxiPIVIbb/2jQ6W2CvQ5kxZ32CxYK0+oLKELNF01
aS7/uV9JZd7cuBgJlYus1e6H+9rWXKOEV/I/PVbtm+3P1p5cRUraey03r2r8uRuyL7h3HwuXJZQ/
qgCzThvghUnwYL9X7s9jGt2UX4rskXE6B1HccSNSKZwtAmRfBPtSloQwMCmos7MpkqXhkPcjSpWK
yhoYxvi+bGm16qJrKfxMcrPTPIRLfX4/PDnSxpQc/qakDd6rAZuooJBRn/k3WLfId4CobM8tcqDq
6sbfC96rAEyLyRk3HH7WhDvF+CSQMBSDbEvNYC0h/mO77F8rv0Ot2U+nm9e49GaeXKz9GNYrp44X
MgxqyAN096p8PvckahRs4p+3/waHeQHHt+VRcOdIcWorsN29ZvOf1mlq3bd+NILVCEo0eVb/qZkO
59CchnPFw+1OXi4+CaC7B5hwSHpiE5RN5KXvcFl0EeKQZoLan1h8YC8JAQ5p0gHMjSE7nJuPahLe
1jwOSwMe+F5ptBIddsOZHPSJAfD/UIpI3f0uINtRCjiR3DkRoMdBpKsAAPJ9y2PV1bDLCkHvVEPN
NY9cH1V6C7w0TNxExMDoMuOIhV0cjRuUP2xNJyJsDGc0NQLhO/JbgTBcDTk2bCLrSI5mt74/FJH4
GMHgY9C6IPPLvvDYszdTv0q6h3GuoPMF2imsDzkX80Mm3pG3N4ys2NcL6MTW6kd0618fUyqDUR62
F4QoqnfFuLF02WbFg0noLFS+gvHDD7E46KIKkRp+obuSbOx96Mw+SIxNmOE0XD8XuzKhZ1zLa/WA
0EFLmZ0GJquoREOVblIMi8IU2bF7crR/Lkp/TXak6FlmyDMiC3ccHIQwhig2Qy6Xh9Y2bcgJzNBK
b12HIbNIuKLpAI6AeJ45j5CHwjme/3bbo99pkcWAuBWHbwU+WCGq6fWUJVi7vZ3FBsbrM8xc5Obq
gf0UDiL3lPo6qx8afWMWd+ka0SqaGcK/yEdJigRNihxeeOw3EvHNkjVjFYs0EiscDE7gide4bNNt
CR5yEXpUKLrh+qhynpmoxcIAYnhk/82wOPB0bTe+kY5KDcmtCfdFehIYhK4WCBBbxhSzzC/fjnuc
X5xucIU2ZSlfERXQqs4QIrjnjHqF+8Q/gAd+A5vpDSJ3Vd/hYpyA3oe8O7vu5TEof5m3bW9sqPK/
PGzUNCutZFcdzKN2lCEt5a3sobKT284VBfictukXZb4F2Us+HHkWQutzeqxEvMhkXumswIL9YCB4
723ZWnFx4r6otAfZTo9w7PJ4emk4S7Vsbxv5Hird2iTv+1aW1ITS6QeM2cnH1EkzybHtAWisZfuh
oZykkm0zYdWkRI6k4XFsS37jrgiRT01uzitKq3TDhqocP0Ex0MUnQ9NRLknTYymcDNLMoR/xBlzF
FQPG+rYqYCYvegrU10QQ1I9+CkIa1lAi0Bx37DpFNhI9Cuh+4l89etJjEk7aFGY7FF04kb7ZI7Tt
9lQNUvbVOOVb2BJc+gGnzcZsVxUgQUut8XaFDIKz3LYNDgNsz9fILq8QJ3GmNjDPXjTLTyuVGTZ8
i/yrPZ6W5+MpEIg0nsg3nXOD42TUfOn4JaDnycVWyNCt5zatJ/GLfqSDbdZ/UrsVtX0Se9ChCWZ/
JeXSt2QwOBNVKx96vQ435kVUi6UGcEmtv1wkDwD7SxVN1FfUGmTqIJNq+ufxFwl5JqSD/UTghHv2
EJ9Y2eDl0GyIBzeP6j81o5SxjS+lLLhW9Lgu+kfSILcLp1hlyWuQSv484cjUOvcYvjA6PTMKf7JM
jahm5H0/Hy+b8z98HhPCGDnhCrls9E6XbBdS7GD89ZGQA5/zvZ4qOdvqiyXFJKizEHb8oDxa8IVL
v1H0Z8AIsUKFElGei4tytp3yqpdYTySTDwoLCoXJJyjQ3JQAFchHCD5QvFfxGd0k/CVBwZ37a2ZP
v+a1MQPTU9N4PbyuN1oubZX2SYfHRv5mO6tNOYGSGCwfnCfSlpFc/aUbb4hcBatH0E+OAZyQmENn
yZYmn++sEkneREy5vWf6CMV+H41fCJCogSdX1J56otRfEgj1BMyvYrd1B0F8ecdMcP9cRWlcrSt5
inBw+JBVru3GipAgARUtIv1VYtrXy9UIIbWLTdJHUgF8ZMJFDmXFyw2yKUDITYdZcgkz4YZpSjvQ
EGRMrupPKSoTgfagC59gaNlUUuLNbGk9ZxhzIrDZPIq5HZGDE1mfsVLVpp95xwFuOiVOF9S7+/Yc
rzTKP0KeXiXbK7l8tHIfMicSyeACwv0jDxPjeEE2fAJZVsDdbogwTgiadxVW1WB7ol0YnbzPHAcq
A3ygtiMwFRSKrb0/g5F4LzravLym9LayB+GXvfkP7EjWINybyu+6xPuKTizDEsQ7k9QjLEJihn5E
Sll+5lL1r0cFA7BLIeBTtE7o8PgmHgR4I+yME/5WxINhb0PmD2+wyCD1EV5LIfrrs94zIH9fs+g7
3WXEUECNmD2f+ne3LEa/DUjE3GK2o7S6KItnQMPRa5tSPe3J2guv730vLRYqx1k1fqb9WhXloOo9
1B/ahs30nl7PSQ99EMivSdUTItdErp7n+jM+5kecKHchHOl7fuly7eibdRjb73gxTNhofCW+aVFG
QuL5H25LkKP7j/I3XfHUbnPLsm5I0tOYIhS+g0i7bJ0CZPKsqHLk86OKniZ5oyjNVuv0iwJiFnWp
DoOwi3lUJoI4Q+6FAGI3XE0Vp74lfhFMSwGjTk1r/O7wPoO+e2mexi3Dyg4WOjMCUB9d/VZPQEnl
X4LMA/4pjg1VVCnK9OTHqJMVwHc+93DvgQ3ERiV4ytCOMkWSxAuKqdpV3m+XOgnUw7E6jt8Mhp4d
axM/468idvNtsQugqix/87x1I4Ru84cceOHf7YnhHJNAeasl62KdPoxdbl/MQKKuZsEkozCSvmCF
Osg/POa6TqCuqoqSvwnL+Ym5gEBLFMfWtTWdWyXfNTm7f0TS2b7VHZmU4kpnvhfHwSawRR/TRCAT
sULCit7BVd65ubkBkThE9YQuzhcaxvxdPjruMez3PijzbRPoHLNvvRr4neTCs2EdemM+gBXIuxNB
8IwGYjIafpnLJjAPTeykqZiCPcOGXTxW6gyAb0cYkyGxjfSGcjA4LDkTe0h7qj7FmWhCbiPAIq6w
zOg5kG15uBeHXGWjxFCmBFeR55teEe9RdJEFGEbEUjBcek2Wk+/fPIAA0dI+2jPSVibFRjGdFd6o
gOcv3mByIp8hwXg/nJ5M+mwdhZF48q621y1bM/JnOUnBVibOTdrtXMSQ/fEnqx/9fYgMXUK69Lv8
4hejyltif92d7aGIlw0J/zdPSnxQqkO9Lmxn51wrwpMh0wwDf0OHLVisTofHIQIzA7535R81Vxxa
kQqtEPljkdxaRrVktTnoDB/RrIB1FHVMYms9qEFY9MVzPUJCd3ZCGKap3FpTXRPfSIEuduRdrY1h
6O2GLHUE/OuULK/Q8jtA0yfNUBCYGaRSe0f2T7S7mKWP8QJnk8pDIeOHYmsLAv5IzxE5nsKv34x3
lP7MxKlW22ExmcO4LGUQt/MhPXdVBIwXmMS9H/1MN2ApSfTtvUrP/sAeLWPlqaBcskfWEkzSvY9W
Xf6B9hWD9yuaAXbqlO4t4uoA5mm1hl6sXh1m0CjC866KNc/ua+DfhZ23k3M/SLNqu6F3fcmGbbsq
nuv/DN3yNAcQ8pacvqCBw/X1AkbBbn1+FPkiHnO0/POGMQ3PJeloGLRoE0ri/5I5Sspho+qRUMGe
EYXUJ8v3ftT2H+PEtTL8oIrA50KBQeZ2jZDNxR1RdWMJbVfrXI9uU7r+zy7mQCdmDQg0GZBvbiXq
Y4AGt/8E6Vt53/QD4w+NON5yqcMRCD1ZukXKBQJ4FTNt2NFOuWmdmXcyeCukh6lpu7kNhqCxF9WL
G6HeGwtuqUXmb3zT2UW13j3gLxyw1VFZXtvUH8IxxABoLvKYRavzONbC0g7pVb39afoJ67hGf1EV
I5CtwKQGksY348fMdyjWfDsA0u2rvm+jWJMzFXEUroalq74VrOv0TwQAm/PTUvct8LfSYe7L4XY4
jv6jttPB07pHgGj1svPNk1fzj67xPA2S+3R2Tt8tLlZ+m5AbRjmV7JZAx5rS/hXTHCVsWeS7jJoX
X8IMkazMnSaUvhZW6yior5y2da2huCw1k7S1b0GHXOKPFBaAfiS6VStsFCLTCVd3MYpD0OqlG3Uz
9d84r0yeX97QzuIxVuoAc+ayzn450Y/gRMikFWBlFQDGP5FYRFKafDLZD7UYRNf+mF5OKI4rIFPR
I8U499LKQV82noJsWS42wHt2A4CTRobxpDuK1FI0R2PHipz139uX6ZCoG7XWcuQcNFpswNseQrsa
Kk51qdqwKeQ8gH+cjb+PYlLfuactar7T4mJx+9DiFoAD3MZyh0yX8c8YfmPMx4kIxrzGJfUdX11j
Fq/k9lZ6dW+QQ6hBVgfaZkAfnX3C71qrHzj+P1e9HN7yEQCLdO4isWLZo9KTEr35WsE/6T0tRLLa
oec5NsKj4734pEqFWpPp8kC1LhNwHtDjw+dwBaI3HxGMbNk5X4YcFV7JKcwrs3+HG84yNg+ymaLe
othkPMbT9ItBVyXnbypWq9OFUx6iKaHWG2y8XR7xGT/nA/7rOJDfk1tFMXpCE3Up+ovInWWYJQtp
6J+OV8IxFgN0rQpxujyJf0CH4Z4VfoEfkCt+bC/D9k0kzhYV3MJ/3mWBOfls+34qNbCQPV4oYsUV
M8sSGtrYVKzpGGrQLqZLFlIVV8PTb1CNIwe+/Zsrustre7l26hEX78gfTn3Wfnmd/n2naau11Esm
oR6pTwlB/SDcARpQEY4MfNApeJHZUQVGAaYi+E9FXzxIcwBmnuny7Cc/m1C4gvSZ7oxE76l2ja31
fuoYvbiFjumNv1VZSE3R3ubsC4cjE80Gogu+QrOmIBK+tk5niSPbsOxaOQ+fBR5qme8y78lRN7gL
SFXHM0jxtXNTSFY4IolIvdVeVU/0p39LhjuZb3jcXgReofa/YCgcAVXgBcI3QiZkoyN9vyTB62XF
9H2oCSuoXswrlHeHMf4AInkkKhqEivO/UfTF4A2lXBMezgzHslBN0HnEWwFJxFszIdcbN3bUjM01
1QBXPihpZAmQ20tF80z0Hh7Llx6eo1J25ir77I6sIIjXvTPnzKDPegTnMk+jVT7bX8+kWiOAV4nV
N/8IkkNrDSdragMXPERR53gxRu3ib31NRhpwDwBE6lzKQLeiGsJ7t11VZlAAAOuvFqdkVp5pO7+u
8Lq//kAMk4gdESiZ+eVb8LwVm8gH+4iGbAveOhOcRKWMO/g44MyI0X3gOnAYNf2vocj8UJ6jYuH/
dxLCxxtX6TVR/ayImm0QfmD/xL8/uJLpLJ6aF/RH02SiJtMm3yE4dYDVUzV7qo2z3nUwb3erZoXZ
axbsTAp75JGlvvKnvCB0onQHgMcIFknl3yeoh83mOppAHoEXfpuc4mGF3NQxn1MakbOWP/w7rqLf
vm3LBaXsd4RqMhKkP3SwKX8hxuhfO1z10LMEu9p655D0XYG9iOZvAENcRRhtFLuTgrAFc0HBA4Ui
WYp1m/WlfHGW35qypPuIhRTPS+1gNr14peeUTZkjhhkF5qaZwpHyX8rGVYMPao2/9DQ9lwXGqYkV
YLuR2CnIRsyrqwSws0YbXEZJXNN3Z8vwRifrduNQgLeRTFwxWbHZcWb864nFMQWb/pwQUzVg7JwA
3ByfmGpC1XWr4vgRdFRUcXZo9ojNH8Nvv680CKPY9T24vFwgVVLheViMkfwc97+EDf4jdnareZPU
Van8Xk6hm92Xtvg2bcyrlyUgWZiga2LRwoUfFrdfQo33qkEOQjdfZQhD4D6VWiPoosbWSX/YDbIg
EFPp3picKvyM94fYABaJMszDv8Fyhbj7vsAav8KkcJTldfdnLYONBbKGnTRKyucC9fYaPbvxxjHh
ua7Mgx4/isljI8a+SHOaXPNLrTwczDjFmtRkcCmfh/l1Cg1wzGQNRcLPvAlw21RttZeN2gartICY
VUsJiE+ea2DqrKFe/HKAO2rcz8jlJU9eICNn8jT/qpbkrzS9Nk98VzZY8HoeTBUU9vIhpNDaU1Vc
2YUPjWzRhkqAnG6TtAWiwEnWKSowrT9PhObBzqBsbJcjO7FSd5G/Jbz3HdtraWMckG2ZkMBdJySF
h8PQDwSD5vZS55w+8Gt3pp/1XbpVDTdPa925hsQpChLIkW3IzBHueOwY8uZwAiN/M5CnKeipYfml
7lHW1EZbn9LjMjVawatQysclbDnlCsxTzF7I60mYXLQKjICLpk8LhS6nweFFVAKSNw6SnkxU+lwc
QXiaWAk360KphpaRR64NBYXtR23LjT2bwgnWMf0oUCxrgxELwzrXQfCRgj8d8KjBL2coo17nZv5R
/K+YNs1Qh3/dTlJnoRgJuuCe2644wIRPYwsl/DC8GFFNHy2CYxiuFv+znw7ZRpIPWoE0SO4aQZlu
6JZUZlYwGYzdBQomkSRpNvnH0k2fQsthQcVQh1kwrnNwFtg8uAUoEw9xWNNikhfBTDbfAmRFtd7R
cA+qn4SmFvMrHlKLaUVcu++A5CvrFkGLVar3mGj0jjNZJ/iSCK9mPogr6s28blPcAGBvNmDaA643
sEGEQt9e6l/TyQPBWdMiTN63zuBerm1yk8bvQR7g9jfbQKOT/i3utEJv3EbVSNJVdCNtkNr+GN2T
XX7PAbTRdS+/+S2ZYXeFQP61FpyQY+MQwvbxbWY26SmKiffpeO0LF1PnDlPYuEMTUR0wLhs6QHdG
mIGqgkOAUr0lfjj/laG2vYBM1QpoPXc71fmmtAcLP6OpQzsLL2LNvthBQyZkX7vPgYFvyqFNqZ6a
va5UaPjIAANlTlvlvUeoR10Gant+rH3+JOd+/8B6qd3H8L7EjXecK9QKRK3TtdXaPo6h62gDgnqH
UfWP6OL0/a4U3nSixBmwd14lwRcSoxbj5ssNsdmiL3hVde+JXhgkrgLyN5edD9oa+oo3rf03ZQiF
uCuquh2myhHel8S5heM16b3uUG7heTOWIP9GymGgcXvFUGa7+7vzGijBn+kYDq6mPOW1tQcqXzHR
X7rILqMyU7tqQZ/9s8bM1ByTFoMIwpzS3LxeNQChHH0GOK5s/yvmL1dw/omhqu6Mg4/cRAuU1Hc+
a++6aSLTi6WHNf+vNLpOOHPuVQVO+u9Ix8dUT40yGToMy8CoO+diUk4g1hnuzRkS4jUyp+FeWO8C
GO5mk/Vv2GMwmFYE51m8DUFw8naDYY0XSYTzqHdl8/z+7PLcGkItSo1iBq/TbzHerqHXI5V409LY
6VS8rI7ZVITmv59gQmgzy/zYfd4gubWEvyeRuviAruO/S4bT9NPUyX3Z/vAlJA4RCoGhNKCW1ZcB
kj6m7up53UvsmLyUKx4pgnzagpg793hxaNyMJk6OzZ1bBXhWMZkV6W+HRMNpuVPSpDm63mLi0y4P
yDJHyhcKPLtoyZFD7qZE5lO5Fz9GOTY7Dfl4kJi8J/WG2AGoF2WDuvNI+Dr4l5vE+75gI1XUD0MK
YJmcFBDNsjQ5q0AU62gOiZYSDPgrmGsQyFqrzgrc2+Z2AvhZaDkAJpctuOwXsHWVt6ySVPnL/Qrw
KYEzBhW3ERaQ1xNdwIp5fesOlaKjs/OFg36fRdt5I9fOAsY7UdBQsxaVHO6bWMV2nX8k5JaeBbSc
KETAXd5JUKbHgPL6BaPvt6kXA8z0qd8lt8soYr55+SdjQdSATS8VcKMjLtvjOfLSVqXHYJog/a+p
luaRqP0Wio+x1j2iNEcWizSa08xorv/sk1j+byZNkr0u0zvSfh95g5PrpyhM03EXjKs3c/N/OC7T
OIlRPbfAMAWrmo+DfTiwVomn5Uzuq2H26G3jSsd/blI9QXVFT4HDN7nzzukyZBQr5kbC+BiwHg47
i1g8qpixr/5FipFzhh5yZ9+KFJJlAI3zNaBYXmPJ6CBw++l9S9zkuoCwozzdygCcrqxhVYHBS6fr
YMphtkylQ39iMLOpgc8Mgotna/w4juBljUvTGfRuV6cUK8RdlMx0Rj/bd3eMe6k2dxyP3b+Mn4CF
7xyy/aQsrrx20fgYbVabsGKQ5WcIiNDWB3L1tBoT/4Xh/t+I64V/tRbwE7paNit1FXbyv/UuyO1r
UF/4Bx0Kp8OY3jVwVCND94vghmHI1zGsWlPlqGsuhtV2r80gh+VMXLcmmWWPtFWCXYwjr1WcJEut
LHzCnrJ1LDU//P2ScQGzuQtmX9QdhcDrBRefX4yO6KbT7d/OcGc9FiPlrfpE7Kr3G9iZkEA7vr3y
TtTx9VucfMp7PXOWyf5XMFzOJ0J71DC2dhn/5CwVGnqFceYK70HZ4kf29abrPc+zysZC5kTXGOLK
9MoQY74fmPAX5UGviqFxyxOkQgiViJPe87d5Qe4msbQNm88lpSAcCeveP3ENgc4ZnyfTyph9TFDK
OTLZOR8fosq/7XSqKybG/u/3gFFGwJcXkIxtgTIDPh9zUVqR/dy2s9G93WNEzciPOnDE/PpjT5gZ
w6gn+Bz4dNjiHqTt3jF6SW+vSSEVYAu8hK2P6rvUlPLcOegbf0WMlIbLKhFatJ3yULztwlTun33O
KIPrGkSOWbeupwtCSGPly/Tnfem/gddFafinNJKl0Sq4o3H4N3/0hgYKXo9q24rCfyZZXUzqXEEr
qBgFN7xUB8MiXx4V8vVE66f2sGG4gWOQrHu3mlb7s4uPvymTmZxqFwkC/vA6yowV1SndBrXv1p6V
1T6NgYIFPzpKLlwhJ942WiUqYYWxNzGsCt47Gn65gA69TS27kr99bH/oimAKbs6sMMM0NjhT3p3L
T5ogBVcjuclcQGeoX/oOg1Vmd3VqhSAQXU05PMlsONv3JIhj7lc/kiQwRkNPjh2fV3Y+QbNYrPZy
BO+6XXvfkRI2LFGfm0YxZZb+/Rhb1b8LqKfge2Xvrov8bvqSfxmIRksv81Em6FSKsih6OGTr6Frd
rV38RmQbWNeWteQ3+Uk9n3psQO6EDJu89MHMeAJothXUrUHhtwfH7snOGfAxQsiIeRkNlTmQHCyX
7LMploJjxXaXJs3DECCfyxBUep8N8EscEOfNFqInfuK8bm895maGqNlvnZ2Lr7UyupM1bnQ/stet
isYLxX07vcWZO8clMQPZFzMHODiUxxGSjMt/kCGrDkZSLRJjT/5yth7YHM7Xgpm2ZOwd/9YjGxuU
Wa/bSuwy7Frd0UE3xcKU+jEEWlaT8cHJb1xI9YsobOBMDI9XwFVWUkxxlEUyoksHaVcokrP21SCY
zJLsgYpXi5bNchYaygKp8mFeMiMjwSqCOj2PcVVa5JpJnlNCOl5hpQlmHcdUe8f3dyTNQgBwnmaf
z5GZdj0DpTZJp2p6YFqiu/OAwu9gqXzM1eKpxgx2HqfyByap6B+PUiDrwB7LSboLT3FGHQcklw+K
NgM6J+ZVe+ogpitaF0f7f5Md1IWhot3JgeEQDFfgNuPXJcvYcMN9ywqb99DtZi22bzrhDxwxCjlL
oFGW6nygsV9/lshdjZ3Rgqi7empXZ3sxUYp3J6u/w+/2WFPx7mZivA7RgJQaxjnIawuq8qbYDOtw
ak8igW0hGefwRnXUOufCRQSinXBlZF/foZoJwUzM+EZws4gJWcVaekC9gG+P0Yu03c4whmSxh0Bl
E109LorriC1UieGA6IQW6yZ2SfadDcYX+GYLvSHwTUh8kDShebYAQyS1IVYGiTSOiDTNiGBEZHgi
Pz4WH2hSeo6baZj9rI0jch/khHN1DRdNo9N9ZT9Y0PIZdo7K34hjKTlFDZgF8UNeENv7cKIF4pNm
uEXCyCwNJI/Owui22KvSf8xNLvSadguZE8vG6I7ilflkLkxijzDgLYmw9g+a1B2aewaWplfkZKh1
sJn4teQjw6j9j7jMLds5quyGMBVH29Jt92Vl5SBsTPW33gGLbnaMcfkqWv+tWtIm5xUDOhOhofpw
AqwinUxOysYqob7bXHJ3YU6bt3b5fpNAD63yxIFjJECqy4eXXzSu1Ptvnk1ExmiIeSt37XIhHrYZ
Si0bAXdMuof43nDKCO2vMwdbeP3/p0TDyXAPlvAImceAi/SAniddJ8rhJqjc9dF+NQzbagDhzHfJ
Kxuw10XXFaQxkIDImL07o90spUIvKquPKG06B0rUM50YkBQchXsiCjOJTBoXfGYw3CXORZ+FWig2
sK05veC71/Xfh5IZoCFc6t+xMRtfUQ3gumWZjy0QCRR0xAFMe18v4UjqLf6ZeTvRNd6lWQsyF6t+
3UCr1LDnH9Rh9ITAP8HALd05gMzyLfAuoYWFJmHoXx4bcKU8k3XZBc4XtsE6R1x1WnlR1eJVL3z0
w3FWPIDTghYHTEaQegvG13gam/C2J4SbmJXsdTW9v0IRrD2r0Ru/PR7cqscTqg/WBYPwN8tDJrVO
ENqh7u1YpMriZd8/2Ra3dIoLXdwjBQkaO1QiycpSPtwXEyuBUDdJCw8YhPDb9Bfq4g6iA+V+awr3
1CvxGh/mQlAIg1pOxGVhSBN02bbmESY1rMiLMiMSfyqkzk7n/wXlBzpvUO9+vMWbWFk1+NU21XbU
B0hbyqJ52/EZE+Ra9B9aX+yM+JtvcXf521xHLgKO10EOdYo9+Y5Y+Gt8D5LOksDqREluCi0h8Dpg
N6XNrqqquR8B47S54B46IoqE2gTu2seHY55NmcYd3yQJTabchrP9csY5AwNkAmJd30SXzoy37bkb
Jo4N0ERIJRgUp8clNLH1hJUEGv9jchZT/PPTUmJ/+XXgvmRwoORMYE3rsbWkO1ki540vIx9IenRO
YqFWiQDB/Yr4796UwVR3BrY1/AUey+LhYlzX5lTc24OYFq8/HqS/mPV3vvwnK0WNy+BueXw/C9VQ
zY0s7xlY1j1YmdzVAFZTRUwEq+jT27LJ6hwRg/W/J+wd/8cCnXakk2Wmv1mvDgCa2KTv2WH7JbWx
NUljrUoK5H8rI8rPi7hiXJxZTQ3xwrmLiNs+JRUsSEx/u8Yvic1CEAV5P0hLCV78hU9nBDJW7qA0
mUbVmJhsV5GqlYHmIjHxQy9nqL+iX24UiiFxjkKgXoR/T2FKf/SLWGvh+4MatbPZOpkqurUIAFNd
ZLVIQ3j4slL8Fx48ojeBe5+XYd+VvlRcybN3byRXVjPLfiqD7H+Qs4KZylNpc6lHJ9UwP+w/RkDw
nsSSj0578ihTbUFB9vJAsT/X56/AFYE3TSGSn292uDzk8boipGCbRWfZ9pv69zqwhynV6TtfKERp
J2J2o5LnAb2nJqJjoeZrBDL4BFKG2wMqwZoKaJGz8efOBjXdRZCF1WNfcKJPKngIEKpUGk+vUZth
wQt1GEqV6/vIAPCfV12PQDpVjI4gFX/p/AveirSfZQn6MXyetwPriZSRaOCCFw3lIOiTVdGPJAFo
raZYnHlYeVAW0meWa1tB/M/c5ompq9863fGjEqqjLBtjFbX5HNrxjtE2sOv7thFrM+tlPbIZOL+J
37x/QGxOGn/lnGVWvudFPhC4nV0IfB6sgiiSFAQESKxmIupMtdninS8k7goLCWzZdIuAfwtAF71W
nDbS+PVvmXy2pZm3DvyU8YVOjVff/zpYAZwqqiqPjFwiFBn6VmbDHTFNWsPvoOJFxsm5Tn0WyKA3
9DSWQjPxCJlrz4y1d/4ebNuCJwjefD86gSi20gnQFqYos1yegFEpn6g2r92ESug+Yrj9odrKbt7Y
yVptg0GNBYsgoQ+MnBClwcQPUp/WvwW5LZWQosSscHdMNBvruNTNI32xoQJVSd6r4wuSyl8/dbae
zswX4ziFtvorXgOZTG4QCVfpX+INoYbUbO2y4FwZS1hCwfnZlrUkAh5GTV4XrkN2Nm2AYnVJrN+i
glmhL2j/6JOHg59QNWahVE+FQI68HmxOAI96t80CowAUoOU98NaGh58cX68YW6z5pg2G1amWkbRa
0SB13IY4TbCs1PW/Km/SiApcB+g1mQq9ToQ8W0wxVxdzvp+g2gl3yE15tUQdVuUabOJmgIdBVE97
VQ8CI8ypv4JCwtsbflNac8eBh4HFsDN3aGwyu6lqKOiApCIOcFJRcmvEQiyJ8ZW84X3Jsr8vX3R7
acjTovHZ4MhwO9dv7ghfwgoor1K/zCwZ6HqzZWywyohV+2tN9gVYIT1ffnQDvIpWH00aLsyqOs5H
ZiTK7WyNX8uD30eGvJ5HykfmH3BShq45C9exYNwpu+xy48eagvjPgrXw9/W5tEbdD59K8XMBLWS5
a5xyuFUnc2SWfFpK5ZeQAcelPAorwQuIeRZ0DFSB/6JptdVwDJFbE4vdt81Ei5+TQbjVXalswMF5
KTX495JJLbDQACj99TpMRJEa4tJnAai825sORGLHigpgP7X7s815GMg5zE8ubFOsn1WokfpAPpbk
UUmhmRau+ekdpJb7pP3OmORsozHModVnrqKHu4HS4b+cpjbUBtS07e5EZ0W2rE/lcdHQe+vlhZRr
N5vXcjPo5bWmnrSPlcdJ7g5hAHJ0LyecDGPerU+QFQPrEJMctq0fe6jxh9H0IlC5aB1gqPGkYaNN
01ujM8x8SaKirdMFnemQXFeH1a3KwE1dnP5e3XN9EgXChwXuJPv2kzq0sVQuCDqno71PgEvynOY7
ED1nRitCqy902ngvwCpJX37frRT+SwtCLDblHSlKPfu7gEldwc53Bb2ZIOxCuWMsyXaqC0e9eFVy
s5/bilprdR+2T835eLzJMiDkEAYj1FI3uiBYL+34XiLlpmgPQ6Qmz0qms4uqYGLoUSHn+q3Qa0Ph
bxiS1Wxk8LoZ8yFvWPZuLdzl9O3PiYq4XJsz6Xw4+75IQNHI+rygk6kmZQLkXvqHR/TAPlUyZgry
Cbo5ZWUo1VKePmgqIy/lOSViBWrkm7eAQUKomhLOVECNIpS5ufV9F6SsZunmqgDhQK1acMmQYN8x
KSWUwt3GZ7TIdOgzDtQ3kvwvtPlFTOMO+Zo9QSI+Zsr8aiu5YXkDRTF46tGzvZh2/GY5l/FlIxPz
bN0ZDDQQdYRkhDLukp5TocxThkGZuQll8AAScgvkPolx45hvOCCW1NXbo45JSQhl+Uj0ohXmBsRZ
7yut/eVg68tqNm/xdjNHK1iCoxecc/fa5sreAUlrCsy77PDQ1lYE8EFHU1yDKxyhnYE2+fNFOKvs
SOsH6sr2oJpG6agpqZeW4ZhynrMIjDnyeJxRsGfsDma2/WPzqJi4jOg6FPnC6CKkgdodSOQj6HN0
VbUsef3f0el+e0kQ/1HSk3YNYGLZz2LBlibkocLIYFPeWdBpHluz/7MjIlCJcVuvsfS05uz3YZ4J
9z1PtpVQBGmts6XSabSLS2QMHpAzO6ZItskNSzQQbm+qdPSZ305BjYI+IRfQXKGXlOj1ksZoL2us
uOvQaNVziYko0igr1neL6Mj3LiXBD0IXJY5Gdet56zgzMdRhDAVEPwiCSfPNkeAzDH+75dRM1jap
nFOIenzdR9vSzkn9nJY35tWPGrrkLTJhXJAHFsGJkITDoASMkFoQKCJB+L1ifzjwwjXbUCIpHNzt
i8Bkz+J784J/OgyxxYJ9DiwlkO7ULAuvgehGpBhHUZSpLbMXmCbS5T77O6tgbJ+EuaVouoYFnDlH
R39GZIsfKdaMnvB3l0fn4hc7LDT2XihB12MlxRslIywlys5/Je99L95df6sDgSCq79bwwL7vlbF4
UTjnFbrsE8ZDMpig6oMxRp3p3qiB4SPOuBnjpe3tp6ynMAN9LvZxfI8VXRHhKnqdCFEGo+LDtM6M
Qlapjwz4/18WFjm9Qm0QrSf1hEEQaPcHaDkqFlHmOzeNa1unnZSxXgJk89TgFc4KBMOzCWVWK6RY
USKFBb4AKVq4PclE6i3uItf+L7B2Oef0Jz6ip8iTXnxyETJ1rVObOPcH2+pYUKLIY5UF1+fpbl55
ipGYBantwSzhJ797R+7s3FAV3ah1S/V+6J42JGo9W+QY7ZNIXoj3XZyiBwdGMHtVqMB+TMEdZOlh
eTR4k9GoaBh6fW3v6D3+Fzuzky8QwNb3TmG4BYns7ug+ICuPCarHdOBhwZu6wKORLK0G7i9J0BvI
bECq0aYJlc4efKVDiZbTFm4rSl40PcI3TZI3nSNA8uyuI5uPJkm6huPY1q8cBQNI9yrdqdOZBkAf
l44B/k3Nm/ALDrpvtgxGS4Pgt2t3FTHfe3mdePJYeLJOovewljDtwFvPPGlLResE5UhOPr9UKafC
5f9v7MJm0tOMTETwllvfZR3Exic2BHI5aHeNlnIRd2sDlYHuXRkhdaaSHje72/LxKMXB5tBK3zLy
XF9JiKKhvcj9l7mo3Kk6lYwqKZo3flRSLjozu58bJ1tAuJxa7696Qpke4f48IDTfll0YdBjTYZPk
HBZiOBpD8V6IjvI18vA5mVdhC+I2Fqnw2NL1TJFoAYkDUjZJhYeYQvp3by5PhNJkim+JdvOvjH9k
XaH1pzJrDApvieRcFSjBFQpE/mk2TdVI69CNKQAfn28cn/8WzEBXkH8dAtXYzpGDDXrRxM+j6wAs
Y7HCD4UV19Q950D2lzhULeqP4NH4hbW7xU0mePexa4dp6MjeG7JXLt9u9cElLEpaCZkDLKno45lF
PiI89yyHQaR2D3oVhky48frnd92bhMYDyz3pSYIILHbIoBWnrEtIXKUWkGo0UEaLpl2aaIn3/oOO
WOrE4nNxBwVJYmjlK3T3FTq08xNtdpEruLIpurfLGDJxHNSe7tZNuO6/5yNZSjREfwlM8xCyZH9/
8a5A4rfFc3vhoNAT/HZQBvJi2FF9/5WHkeWwiaZH8l7gnngzl/EuT/VD88ujb6SrvjoggaWxm5to
2CsAibwyyy4fymFgT2nPhdbA7M1PcFcdklUQ41JodqXCBERVGrYy3pszWNOhNwFMbXE8jRQWPL/n
XO4FWmdBfAR0zA225aBBIA/tjdGWLWSQZmZFOaov2mnbvZKSWKX8QxPFGgrKhw/C1BTE56P/nd7o
5g1ug+6bdQm736R3bZcyQRv+/VB7s/WC9frmE5xVGEepMq9W3WDWeVZn1Ezd2D16hamAePLdlskt
DZdasV8uFpDGg/Rnr1wqSbVXLXmtUWcSNzFGxQTcNlq5ZAfERvuncwu62E4s+Nq3z/9Vs12PZBLW
K2KpXvxDRvP4maLi+zlzxImb2DdEEzIQEgSAkzmBwm5XnRFmWQHVGN2pshYiOIsNCgFQWDRRIOxG
UtWqfL2yaKKCopo9maXmXsxCn7MsmzmPicqpDTLIOLluSe7tCuJTjIMGSOaTvvu38kf9za+7w6BN
4E7HN0SKC4hKoy6+MkcYVQUbKcE+UDC1Sv+XaSpkZKBcIqrvXYaUknYBqf1SF+pf+zdMs7OfEQIu
J2XLuAGV7dNTXBd6WPPSDZQhpUS00Y2b1oErqylRZ7cVZA1LARBlk7EqGWKJI41MnU09QtxqkamI
lO0XgBvtrAIJuYz6dzluHjLnyBDnxhWdffQPHbioFHEbhe5bkiX1q2DFWaOAd0Db0Ot2BAR7/pNf
Ebhfu4ftgH5IE0OcwN7/Lt74M8r0KxTryHSRjWEpErpJ3XoypvteHNBPXR5dRdB/B5zeGOCxXBj8
7j4oMGP8JrChTXMh57EtzSdHx4kr3wA8VaFqkUFcyXiXHhkRhG0iqdAWxCxpfaYk6mwQnqzP54+6
6CHLXOj6bbCnBbgaEmRqusqcAgfSpinsFPXEsZgrsF0aRD2HziePJqGoUh5K9EtrxNQfNyQGHoG0
Pd9qoSiY1KAvpjafvjBO1zga/Cxc1qZE9uOVZIdCslK4jmBBA7S47YrEPWFSCyTDhZRBrcpfKs0v
y4zGGel5qM28sMGTSfM3k0Da1+sWtrNEEaHOXEJLzcK9yTyTN6eVggU1pQd9BFeqnxyXqB4/9nnS
XFSMKUlCmFpJCS0zgm5NeD4DqmuJFD26RSPIGDzK/KcDAQK6/Bb9ZcClGqG3NvFkE3dxwdcWTEL/
z1wfYqwbFVFO1veTdMslWGLCpRbPLWwCL1dv1H4zNV639iOxa86FzQt6bdxhy5GaXuFvV4UbVIM6
8ze2gpJjRwyQjLSZufWV2IdLzAwEIDbv18A6xSH0OnS9Wh3h8f2G2vHq8fS56TmJlIYY/e90szY5
p2kVV3kugPGqE3jBUBDXXEJ8eH4mPaKA+k1tfBkCS/tg6c/iSE0+MNReJzc5RFTs0IqzL1yakKoM
EljBs5aD6leIn4pm2yjVE+4kx5eA4/0d/1EhdNI9a9yxQhP+TAtLi17XJZtQmB4gtaov9GnUxo8c
mdewLri4ZW6jhdi5f0RxWST+TMbZnzsVvwdlz4Cj2sk7mlbPGpap8otk9iqCDIGyUqrya7Fp6Om2
OSIuVcD6lE0HihIyill3FuPUV6I8wSklyDxP7rPcaEgfFiaj1qD3TqLBL1gSxVyATPKj+C+t8R0J
7UCTJFe8B1zQpYRszuoz2wq5VduGNsPFDN7GEviVKRHadh7N6lF0VO7MWeerYH62P5hLqZll9j64
f5oDO/HMvRQuv8sevTADBkgDHybMb/Qk7lwDqVffjDGbgs8HOzE3lAi2yNgID4igPQfS+utM9jIF
u/6cX4dNx5uTZ9dZf7L+FFlwvcxPZgEdUf310s8/yelf17prtbs5kSw+gFdUYJtlD0pApdqGUXO/
+ihhUqrDQJO5upJMxrjofhRcNkqYR0cFCZd5BmssLSwnCCu2Y6xCbMzuU8mF77ecZeVFsSIJ7hcr
uVFiUhaHqJOuLftN/I97iOe6Z3NbXwUfkULFJs9f5o7FvwxNjyiHVpNH2HKLJ183wJ0613U0McOI
BigMJ5qROJwWkFSB0L2DENoR0f/h8+QtJYKpK0DqQrIIAa3VDX9uq3JPiv8/UpcwvVumICfAbR38
7QWFpypQKG1AdBC7EFvo7hV0B+1cXl0lvqCVylXjoW1lauYpAeLY7v6MWU4Y566iA/SVwBVYBjE2
/r1r/ONOWc91ORf0Rs22vA8LqtTMz1x3a2T47gS4HA40PXTWIEnk/kauzMpnAGVnoG8fEHIxejSo
uVCg7nfwjBRwIakr5FF+1GluIyAw7JHfJMZ2lyn6lJLGpG2lpOneBl0dzPcFN4lUm9YN/c3sfmuk
NTsC8RrISRln4XHQkzDoa7id62jIOvcMXk42ORuyJ7jVGRB6bCVbWhD+tPHubjqywOJFHKIBR5W3
GqKN0ugCoK6BZvVl2Jd+50L0B8dXLBIMkzDbxBktWnpj1C+AktfeAiS9iNUw324PqpAFIvZhhBI5
98DGrYP287/7rDDyRIT6W3ciiEhyCtkCW9AvaFcP8Y0bW+HkFB3reVNLgD+ix0XrC6SWdk61HY/I
z5oSQ+VADTH6eRFc+FIkSaSChQiMMLAfd80vai5lqr1JFMSFe2DBoOLTIuGs8stDqR8SH9sl/veY
iOjvYCWz+JY+MAXTSdn3kNZPm1Fl76vHRsjq9gD2cgQuuasjVqp9Yi/23VqpJqe0YtIG2vkUjtJb
aRkEM8tTG1s3xOUDOt7Zq27iDuxxRwomqo91s3Dis+gniAIvufXcNiDcEVMzCWOl+NMLOw/6V8/o
j8QKf+EGEqPE0NUontBvgrA2sDJPcjOQIYvZcHdsVOJFWNJukIfX1/8D98iv6gxNOvYNwXeh5+vk
pCqdHJaLcoQMlfmA5EsQVZkSN1MAt0XkTrmW/XVpE+dsdS0S4ty+Q/OYTC36VMNdkraHHoLr8Ep5
/lDKYE7aWdxe56zyUhdgNLFWBap6VwaJ46Pwu2TDvDxJxT2TcwY2zVW89v1qifKA7SJz2WmcR9eg
B1fcqiqL58POFWnZiI6GiFhGEKjLEvK2KDSyBYh9t/rxxmGaBBII3Qc8uaeXdNz1tbai0AHBNxr7
iHxMgj15Ok8eoykQWc/ZCHwPwxeAo76ZrhYlx+MUKlRuJILewMsb/9xmGBm/ixm8fzTRzVKwqem1
a4cyH7XLmXD8P7GTJYbXjfpCZQl/kgGJfkXYwS5OuGnygi0NfqICZvQDs0h17bvH7RpFiA6Xg0E8
NxD3PPf3PVRaBolmEqhMsuH8AHy2pRWIe68MvYUSsARUvVzCGqoKUtGlZojI6yeegJpvpu1iTa48
RSvBYd99ltz2rrkrv+qtrI/MBvpYpHLCV8B63zSw9CJDqDDaAM2Vifjp/MBOtYYpvUEqyrzT8/dU
WMBFXUZBE8WC2/LwSf4W2Z1DWnyHjYeJKln4ZZ+fISICwDkZNvU+iqW/t/OlnJt5dwUfUeY6Yyre
9l6oEPfI9tiD3dP+vm5eEz2eMZdyJXoC4iv2Hnm27J4KttGhoQm+awQ8ZzSFcgqwHjQU2VSp/JW/
FBAebKfk3XoLw1YHEQ6XQpSSrhO5a7TMNdKHXBhb5sq53MkF2m79EYAs3D/kxNV1K39YMlnUkRzK
WKqewdtUS0DSzMM6JDBseyQMEIDBVA2ihQL+gDpECu3kx6H7ldMTXTQAF6aJA2QbZfpC7B9qDyRL
f5frvxW/QvHbrxd+qCZFRitgIGO5/fD5KBsyCNoZz3HqGrJodD5X8efAc4JdtozVaM4jaANA9dwK
lMLYSgMnWkzy5biApHm4sYpYzIjmgesbgZ5H7wdExMLxnGYXGh2irUaZ91EUj+le0AaUjhSqmr9X
jOqAe/dCELiLq6eFHry0dK6weYkk5kt0LZsdbC3tBdUj8xONo0FKFFJTZCcEY5hiDL5VgvF1h8V7
XB1YAGshwivP3cCC4jONLou8g9y74m9jYm4VCEwYeBZlOYiAufoQdVjpXguXI5S+gu1vViRCWkww
YVLZo/8iVU9RStwW6IVt8sZ0JpJUfQwPLqpPL1CH7FKUL2F5BVB6IcwXHeMlisFKKKLlSYHLNRl/
Vh4q3fBJ4k5jT7hwYpOmS3ZJE36tTIomDg05wbkDWrZYMB2LxAQbjIiY9QJ2LIf0py9vlzPLTLz8
S7Mnvo8u2T6j+1zicfXfdXrjLECKH4rRJ1K0IAUGuEYRWl8852pjs84kLKg88s5CreuOysD4S8Cp
XfgyGTOD7d6SOhxZ7eBK+w6VxvGgrKFs1SlLLha+T0AIfqAkomf3NJCLU9hFvwykzCto7gZi71KI
uhF93KV+BWyJGjB9jeCu5XU+hKtc2J90KFPvufx9uwjfPnZqBt7PZP6ZBFFr9co8SIqqeSnZO9Md
SiiI+Leu+aYQvRAldG2z6KFuIQMPf4D+9T082bc7jA1iZDG87nz++MyocbRvFgicJyC99fIHZxad
9jxzFFRHwhtPsJQgeXYKFsLl5tyMpHn4tharnW6fYj6kyFGkr8andhedgzGibRn3acQvTdM/PuwM
F8DmXIOtx9dO+Fs6UMN3VXoBc/jANYF6rFDoyz6hsP86ZioLt0QE/wAFMdiBEZUXu+PVJI0Jkg4q
vMKYX3ynAi4+FVxD1b9VuzG14zNCMMhIktxtWB/djbTJILj61/WEjdpeftIU8XYyzOqORUvRvQRL
8jylt2im1x35fCVls+SmyWvnJK7QMjKrE4ZakcpipfVYpJ1uuvfSc45n6iYyv6aqhICnGqnzTRS3
1F4xArFiLaizUDwIIVJgCDwdB4yyk6pxO1Phi+BzkG9hMUCRf1HtCZ391nw5JtI4DgIMRAONjkHL
LOku2MPLEuxMOB9kW0wDq+r/krx19RfYyGu4Fza4T3PYHkvltgfvuFzQG/hhXoqaQEWkTP9Oh3CV
F0O05riBUzkFJ47N91IG48vT7aRlHSj/QCO4//7NvXl7Re8gkGyZRbcNkFEaiiIIbVP5wbbxJq9f
aqNpef/T6c+UAusjpURJCdpxqDPWbM/JjSaI0TCtktMhynDta86L1lS+4/VWQA/OUl0vS04MzLbq
XSul5/6sa2o/qn1WoKacNoDb0UhyOOlkAAZuqJUznZnBiMYsnp/kkkREIbkbuFJxMEfh4/khyo8T
JAfLCGdxFe3HJ4Glu7HAfqND1CduRbpV/CTzAIb3vmLGox8KFBypIbPF5VOfZmXd6PvFHL9UH9sP
N4l5qBxgY9Mt7I2NqXZICPKgk9LXZbqAZ9plbiK3LtMIxxYcT3zqeUD+U46wLuKUsYle5JDq4dkH
wBSZA7qm/sp4UeBJCQ6eMc13VdhIcwx+cZ2DihjVes12hB2gRSp5hHAzktpaU5n3zSmuCMoIGtmU
IYKbAVKk0Qs0uD3pLzC6btHwRkrRDk2Bl/nkpOzSD4Qo//kTAWEEIqJBJNzZ5E+nqEKXwvqDU11T
bUwaZWpgyLlQB5NewnhKbpbH/Y08QSMr3BIIVhzs7uWXtyVR9done0fg6XVojQ8c49l3zqFb4v1m
qDMJrzbizHSP2cNzCrkZUeJsLTp9w+l0RiIIlwxq+l+S0AqPVe//aFbu8df5Zt2QvKuoyYAE64Vm
x0jAw2L/7qbwCf4cMN2CWPy02atNZ0huE8sQ7lLb0sKEOSu6qwxUZ/TS+s5tuPs18E+IocU8ROeV
8nxefZUOYM+ZPioCaWL3fZk63MOi/3LGMRlwAfjq2xoq27pgXWIA5ewrIzeYTNW/fLN/Qk7YFj9k
Ua9RUtkzX4evYVCIgzagOfczEZZZn/TCei7SA+Q64mUgoTdPISfeRoFV2PkU9P9Mv+PYStDDa/9M
aj5XTHic8PzdwE8Mh/z8sf0N0jnbJm4e6WmcP1AuV3KPXuvgh/vTIcv0OmJe8fj+rZ4ADgp51/Nf
q5DX3d9U0T2EpedR5JWSDifTaSTaBW0jBM3GwGH4MMg6IOnoZDIt64CmJqPzBQH0w++Kk5D1AmVG
S4D5qmzlx1w/z8mSrXv8RFtiRX0NPv4EYer1KmdvLRRbcNip5AkzDAShjJPy4J5GAyXBqz6YRFJe
A+dBg3CnPad0sShAkszjTWpK3pC5Omw8l+DGJ4C9eCIC01yvUbHz8wJHB3lYIK1WrqOz9ZPjPWOV
xouPOIQ+oCpZFDTSbRBBwQMHOqhng5+yQvTaTij7dwXNNAe2DEwChn1p8aAcpRdi+m9amnsPgGUy
ApV4M2kC65WOWAkTPwBVnkuCPhJQgpVR1AZ9/38FT0K/1m72Bn+hNjg0G3rzgEmtQAo5hDU29/k/
CSd1IAOXaNP/pbR2W066cUklKMOjKJFVbJUtXdxj3vT9k4D48avpP7NLlPOlX7ABnR3LSnxLZm55
KjCJkvNq6KeCQj+J0pCrX85VyxjKSQMLby49LxWRQpTwMv/v2vgIcGq9ZV9/Z6yvsIiIk8LCNktq
+KlJ2sJm5MDdSX+uEDNJjazVAeV0As9qK2uBVCeezHIkojE2UOhC0BNvo6mtDQbUAXU3ftulCRyf
PXamfjPcDuXPQl97FiqQ0w8tDbE3AntVZigYXIfw1fiVXlGDhZSB6ETgQXNN6dglUwwgdqxP6bC2
lwarNXNPceUj4AVbXfnIYrsKb0Ox38R6xv318YZW0wqDvG+pwzVXFZltiNtYrVJgoAywDthR1CoK
+O4/1D0pPzIlMU8arZg7giL2fpnyoc/dEFRVqlVvFph9GgCttxpdgtMWtgRecRNvtgrjMC42FXgC
58QTJ6XWw7Gr8Gy5KBce08gPQbFCloFcls3OITbwasZmwve2h+7p6Ij5UnF+BpkbTk1uIbfTmjQp
4+azbxwxTn4vlf5aMQSxcyvmTWiYCHd/fbCV6S+cBwBGhve3JSleUSjjKgu74D27YvMStkdZ5JLO
S1X3dRYUqD+FGtDT/r5iKtWxt44MmnmjeAhSeMgfxRIyaKhwZp1NvG34UTA3VLxOseP4WGbOvOaz
81cP9s7Kw0NRK9kvziMuOCPxXs7R3M/4l/RM/+eK5AjsJa81Y7Lh8uryX/oPzf0ol7VJKE2prlkL
wN+3SvCIYjyJ1pRPEP3681nSiQ/+9nY7zFOUdBtw+U7I8T8IjJcQgLiGGnAtH/MphyWY88+IPW2s
uX2b5Wwi/ZGOKy3Fj5pOgeMHX+A87ibSlxvMTf3BxGi1Sx4CeczxcmF0JQAfvbUNks52fqIfCuHI
lrROuRqgui4zP9fqKSxJ5KcDrtHGPPawFbT8BU7yhpIzHyLgobb/DDLNTNhvs1c0HNyjf6kAPpAL
/f/pprBsdjtq8nfnA0OGEY5wTG812YFk+Z7lnk5BzgE6B4Cde6xw/XzBIx7RZ8scYPMBg3zYWql8
LN4z5pYRKKBcOJyerD16VQ4lg9cVMuGqYbnFGpAyxwyeKOw/JuyJuq+BvD6a0xYqTCq+2r7JQ0Pw
7UTgSFngKhM3JjcAX98yJ/ebRyuVeNZtFc2Kno2pptYOcDL6/Y+3K3BtGzZC3QM+TAYU0QGKjpNu
WAl9qNE1S0z4dyooPTovCduj4dFQnchmZZmLomNmZt9ac9/XTIga4JHqOfbUVv+1kBTtQV2J3qZ4
pT+WuN5+sisuENHzwxraa6VxjVHa8+CdONZImyS1NM4G7roemmzffZ6wPdYPgl5oaGWjYbGpaGuO
6UqklPGczzCOxz9lpLM7HL5+2sfmps54Z4cOAQlelsLxeOs10ayeLVMIj5SwkzcmX/8t7Eh3+J85
8hYH3JDR7P4GEAoqL89oSx6NN+DfpF0zhwQVmWfhIb+3SVP98uquT6qGhsgXdM3idujT5GWjmxUa
rN4QELv3V9EK0N/EV4gJKbLNjx0TwtEVzecaOkUzxYFDasyuRkMPsyloo6/HNDm2LyiZK0Sdd35J
b8876EeIbgtr/xy+UpOekirp7WmnVzf3RgfxuBCrSOKB0RI2dQ9gtBfoxFj/bifPubK6rUyzyNWI
fDO2nc3vEwXGzJcmzN+oKVm8TZttOCXWp33D1HFyMSnzwtVoQunbVTG/uUpjUgflG/ellvnnfOMR
kIPN1kvtuuOrzsasaXMfM7x3A/ZIJjBAB1gRX/GpmY952wpDc3SuefblF57zm7YCSgOz7eVVZ8+M
vLQUR+rLcGKEVBmorI3yPhu7aw+WmmYYE22mWIXmIQs41Nz+aSzlChikNesPXurJnkVtbCWwyTif
OARrei5goLzs5BZhEUzEEqOiOAN8R1jrSCqU3Tym0wqdeI12lW9gk8Psf8/CaSKEbh9hhO5xAk5z
qlaqZUfrSmT2gqpyFFWDcm/q5Dnkz7UajITW2qnPrR+WtFSICw31DinyzO9MT3Mhg8GSbbufZ0lm
1AlbZUzOyEEJcZrrABeWnD7OE8apn4BYFkYcGcYb+RdXC+c/diSI0qM60c/Yz4vkL5Fv1QPiWwYz
i8tof33grIT48kBpCM6zN/wFibyGx1dzbEm4s7FPMAXUWkuhG5bBf28VqJOQtaXt31Y5pozBhkuy
rdm/+DOFl+TAPRoqzSIIGXjhHAT4GpqZyfxcNoIGTI62/nCEsjhrhTUjJqg6s5LBcSmAJ1Ds7fnC
SwGC04VZZwqOUb0rU95znSIL4/Uf/cTKEOtOwBULhLkWzyP41pkPUP4z+V0WuYc+J6nbBd4jF3Wd
nIaICLcfJtkHWwVKb3zJKgoZgLWA9l7L2jLdDmec6xloFog4NMcolTrW42l5N3CIxBZGMWz2TlkC
7x5wz/4+p8ld9lrxDD4RL2FFEBlumHpnXUH5bYJ225+mFsno57gS44D1N5Uyy/0N/HJ0fU9LRe3t
gbqP2YMpG2LrDaF9v+X3eQD9nem9LaXNENWBM+i2jMkm4qlSpp/IyokR6Wm3rQ3W08OyxoFB0W5n
LJGTef6kPvFXMrB75fRwocExU6uGDZPysqXpU5hmi73E2/7zUjfJatqpqUK8oR8sWaIFlJx2iY+b
Pa7L7oL9nIQsFQmOewEDmyL5O/7+OC7L4nA+5OZngAgFzLrnTQk/ozsa1hf4jEG4AO7CqkHccin5
QG9ze986OfobVqv1bT/YfyYoI5Ob4pHX04KNBDknbt1gxn1JYDT1cwH8CMzVka68/ChWureavEmg
aGBH1yyEcq2MCcawpwhra8kF1Xn6Olxl36QTE5jek7MW5QVM5DQoRlm88v85owz6ATcspjFcb5rw
xA3/GE/9tiXqgFak0DId3BlZywAc3ih29bk05M8BvGatfOfvSACK33OoaCm8z+8WjCOBqJYuXiZT
LHh7Z54NguVXCfYwciE7r/hNGybnXhrTOGY2aSGLTsRzuE8+dGQZf8ogpveaU++7lgHzRdegQflb
7GyIZt3PxWLDrXYi31iw/Tf/sj06LgKxaLmrxZpX4wMSrMPdu2jVU47L+DDysVL6c5p54DbZCQj2
UuIPQ6cZFmdYkK6NRyvr6zEyWe0az49/oWF9Wme1mBsCKafEXYCNUhZEUwnU2h2C0gkVZQrMDAFE
NOYQvtN+weLhP/967Fa21EySOfnKuH00phuEo+OW/x+pNSG7CHMClc+wUJ3FkmTDcjRTYVOnhYzB
OMGzjl+022ayg6Qv1HooFLtLX1XobSip/JgvwRLuNGfNO4PwYcsaTseOgJ//t+/YHp2+bCYofyEy
4ZRZiDz/cktKRRzjSrVl1Hb6g+3gmyfd6tT8ltMT+PrJYGJbkF8BETaOnATLdNH4Rn9LEqXnECrC
gUHC59NoqgGx7ggaoR93N4CySCnxK3oZ6mdlEEXJHqyDKmEG/JG2t2j//VcAUez0mwbptnEXpyjP
ZAgBT/yQ28VlPxuwtqIPNBIkMp6NIR1MXIBHZQr3kjs089H0uTVT8yrwHq7bd0K1rrtywB6y05dt
Yhc0f/ou2BRP86VSDis5ukJj0HmIPMeanhM33CKujnbcxij/UWpazO38/Zv4Z8X9sr+szph31X6f
gGaYljnnDoiOSNOAFSX1BqxbBpHWuDkHa3hMglQLNnlvukJ2xVyxkOKXbWkRFf2Gis9MWg0AXPsE
SgQrGvqg3uEnZ7kTgWdZ+7lK3p6Bp22VnjEHPoQQQQgIeND8yXkaIMN7NF65hHmOzyq7JPsNVYFF
nCY+hKxvTxIlMCMA36Mz6VClJgNVszQg0y3egdLGn9Ihj08K5vKgALZwxNwCEWn22tkADsBls7iw
DgxNvb+uc3OEVsKyBLbwn45WwCG42pY2fetpSwTbxjM9ZJk6Lj+y0tRGFy9dO4RTCBYrxpDAQY8w
2RXgd4hZY268d8QfBXx0HnxlFDrBq1OIN1nLIrmSJtMt9T3SsyBo7McsgntYEgNfDANblnKY3Tdm
X9uZsuH1fRiEAEVzU58DmexJhcTvwRFurqVXnpNJ7jWB8a0h4hyfEdql3/g0794y8JuYpUzpZXTQ
oJ6U69EEQr8ZCQlQkoJ9pYdvd1LcUenvNFeL9nvXvUsqokVUuhkTwarFteMyNb3fyKlSJC4RCsf4
ZzRQQVQYZCKOQMeaVpWQNyQCLxDC102ZCt/t80ChpgLOeF4un1mHU+FTp+gaRBtM6tpNoCw00Mjr
vPofzzAiXJOnmb0FjNAU2Gwe9ehEKGkjU5l4faIMNhJ+azgO2t96+lBwZjfERmdfOwK9Uu9CfOgu
35+pNWFA3fjwEyYiIUG/7VoLYj5/mj3wLL2GHJVTmFzZ2PmCt6jLaq91sobKaELAM+SQ6SbTkoW4
/LUlCsUsEZvd72mbiwtc78jkNPy1JMTHxODU2DtACkZIueAjoKK67RlT9DhORF+yxZSmP48SNAvc
0niwKCzLkWlv0mj9/gWNQb5qG7Tpux9vMizN4UI96mQiFEG4H4ey6aZiHuFSFLWJRA5RCSBl5eh8
JAxgIpzu+2k+zRBR+7p6jkE+SXAbR3ETAEU0mVpj04IS+iQiCYpW6D0nY0CBTSMkxuUiP/s8O5Bg
fC0MMVlKpFZQ0OHDdFFSeuv4BAktLxkfDAloSA45SRof81H4QwfvAMUHNCOsMIt/E0Kjitx1Fy+u
1191Je+0wi+VzBv81653E0Hty3eyLJNlBzpCcyDsZX1gahs2pq4o1jXPG7lpgJaTA+6OiuquWnjJ
QDeJZY1ewOrl0FN1MVY68IakQHFOgVisjQQdCSQJ5m3PxwLmYW1hDzRmWXEdzD2tUQpFTkaBs9xU
/A6u2wfMXLbWBu2hi1L1RmLTQqUvynQi3nsIi0VvpJeiUsuXNHR2XgZT+srLPWhumi2cONbbQ08W
/0e1qama6v3ow9HIwuK72PpclRBRWD6j0Ycsr2M6t7JA3TH62E5rmKLFb0F5FrzpA+abMquM6QkC
RFnBiTFB95ZhI1Mnd8UGY9u1n+HpGaejy6+spP9R9j8hLXVmf7Mo5rjaeyIjBtkKhC0cEdPEHDl9
k4wRFxRpA+MjBYTKfO6Ew5k6J6o6LaufMxtEdL71Qr/+EeGYNcQam8xihRyBD0QaeegQr+1tFEvr
hvcDnsTTQjzTyUXQQ2UmU+lHuS9J4LCJcWf4LBBuzmgmcBm1kXu55LkQSFM6H+ucbC7JXMlt5dcA
TDvYc8ErTqSys/+x5kxMTANSK6DB/Nz7Fk+beQsJvSHQAsU3YDn8yitQY2ifnuUt++GmatnFpxs5
MNB/50FbZiWqKhQlgHSmk92uW/lkWfLceaQY/+yf98+BP990Eo1QXXrsbGO9kiSxVH57R19UV/lR
8jrhDmZJPbefHHSD7X0iDnnbdxJbWxPt1HN4CxTjq2jOwL81IZNN7JisWcFxnMTVCzQdVlTzhsOI
1oaQC58xgUuFWFfvSn1MBZoxSf5lLxeh4es3Y5Dnkx67y9hMq+5ecz/+IUMKSKgi44Mka5DG9+n6
vRH+v6scmLedrV1g7ksaoPYOJswawv0a0CBshIGIr3qF2CusTIK8xcb+0CPiaDTqyddl9GR6auFA
JZqmlpoKn3tmmXCmM6RWmakSstuHLtNa341P5Q1GnECy9k1jzZrQwtzQ7KdRUO8tr1KQ2JvdqkQ3
TMUZiia7qy3mwlNOySQx8MdTwjI6rZPM//OhLyLRJJHgAMkv+9moB12gM6J0Ms3ey+hMitMV4l29
Oyhy78k7hz0uBtRCVpLoy3MotVwph49qK1VEnk+mtSp5daT22uU4ieiyW+B8M42mPaNUNvB9vfKa
WYZubGNqpzxwDy90GYG484qjMqfYIymYQFA01tuTEK/8kHa+FyLQf62o/tih38mRPahxUJWHemgX
oB3kQyvGrvwIJkfFVfr/UH0PYatWmFfUxPYgmzrdZ8U0uCBtheZ/hjknVOqo9PTXz0ggcc6dDRtp
4TQjysZdesJAoCda3jgYEjXSrklksBgiQN4PtTqv4wp1lqIATNPskibHDHsF+XBrxMLqXfBsJk0m
wQBbU2hhx4yFAI2iFgGTyCIpwoVSDlLMM5S+jc4r2NL1NHSe083z95Ud/zJUm7EqUkuLn2aBv8YM
Ozok26i++z4PuMKpVUuZQSCPjvtyCw62Sxcq+UzAQ6N2W1yHa3mBSToFVRk6KwgA9lhKzpHZm7UC
m2DzYarunoJpKw7vDjrJ5KlV0fnYLbJ/8XgTskJKggzEYykzSTsGBQsaHXTZ0I6usDOow4tNFE8R
WkfNeD2xVvCF141cueJJsAIjBi8lVqi47wq8LZe3M80cn4wblQF+JTFrbHHEy8n+Vsmi7aTmRYB3
nwfjAihIQ+x7HdmJeCeqBEYdsKQWGaP1ek4RfwmH1tSlzu+AGR/jM7SqK9Z+oGu086q6HiFEjmJC
lUYcNBJjf57h+21Gd/LIp/zl4eh+5NeWLbaDTzuElpRlC2K2X7AuIyKq2pJwgboEP6jM0gYRM3J0
E3zeYd0WPuqy+o1UghoxRALEbji9CBBdJBpzWIII4dRjremcEJbji8tFGyGv6FSsZ04/nsMNlIl+
kKzW3VAGmAH75bpNrBNszQYUY8nn9xnM5w9mQFkWi8Qo+TCDFbUW5EQZoLLL+sNIPvDJTr5CGkVr
x32o+wxJNuykNhs5cKB6PaMqvbVCNGGhhfEWLTSFW9u5oAUEmTNfVs56nqHXhxtLY/YopoLqhftD
PWWaQPLtWuFXn6fnThNaP7HqcwB5TTeunYGH/pFgzE1sQJS5/Cj4ML8woSgNaTFUi/XF87HYCux8
zooVudrlCGssrKM2tuMaQTjeigFqAGdb8cmPQxbjotTxHZtWuiD0LlkgtjPRRKOkoFIcVkFuz0BN
Rv3va/ZDm1nMwr2pF2cSnk3iThvTpRlvpeFYESKFDwUYmLlCutYajqtBClMJfA73cuMx1EPeKtuQ
8VbeQA1PxXBXqyP+GLUemaZLFyTUoYKMrfMfEWHtqDIZMyWINqWJp4oEw74W5S3ieCsvbLCIPOC+
4uLYE6MO2ohrvJtg8sugQVi6JwYHpZ8URKWTwdkvmVXfjthLiuRadS4+g2F76n3Ixu1SXQMGflTD
fBCIT/C2hirgcNSup1KBV5WWLcdBWw/yvXFt9TTg1YFnfiUR6xaIAjYE7t1HuMBNIZu4xUP9+clx
Qs7vKPIy2dXttAFAY+w59YHV4Qn755i18WetZLj1imDl4PnUyGwD22n5gZ9Uh68JSxFk0caglL52
/xAuVTNIRkbHDfl66iqUxV+i04V9DgSnxlnAMKmdB4PPGV5e4UNmvGjzYSUBM/s//nvVfFVUuxJ7
P05eaXipL5d9QnZdmVUhrG9kaHmerK+ZZxWZbHS8Hff/kgRgny0ZFFovS1U0rOmjHrKjaSpPT+Tb
0zdix7s3/Lixuqk7x66RQ8ebzDFg2R15hHNo4QTcV3+wj628Ceoqc+lL4cWSzMfjjAey2w9yDi1R
EOqI6MIbLcJ/AqcTzwGaNmopChYTqzM8Jx/gkj7qEzHgOSaobQGmcoNiGaDOoZ45+me7zciwS909
BbXMvTeMsCmC2KlGysSFBxn1D4CVO90P85swxWbGsCyl3ghG4CibfoAzRp7AmT5NScGUupyDbLQy
iYVA1hOy6/XUvfRH6s259MF8I2aUXwsV4UDN4aulcJLk8CC0ed1Cii9R3zknh4sTZHZ0sjlHlEXn
f1raJS8A3LAjA2wnzikT2w6Gt2/xN5kJfnGa5h3fmnfpW7ysDBUD7lyu363c16CbPSWsgEyPMzTu
iEiaxAyZHsGws5RvBpr0NaFrQxU5CBhOKtv4Moro1lycCczt8+sZxIZkZ81avVpd7v8+d90KI71B
6fmPZnmezQ/ZtPTYNPggKhE6PHi4aFRu6Zh4YA5b3IMKg1mK0aq4nulHkM6SXpdLFAiK+sREpNQ3
xy/LrNckxE1UXpo1B/8j9+M3r2z0B/RNUJZdgly2S2bzvBZ7OhK4kxDKCGFzlcNQN5qcscH1lDVG
fOuR3YG0CLhA7tKSn2pfSyaDMCpGfgCOdx7aRG2EOJmZM/EuoVfrFmtQH573E3vZtf1T8eibvN51
Zne72HSUq9fmVBgGmfr5iAuqwhAmDMAwtrmlovvUN8JVs9G1+g2GlT6ikJoDUw0Vevk2hXmnivXf
Iv2UJAjGQG606tMbpkQq120EEeQNoWOom3s0cNrpGXIWiN+H7Z63be9EzqWSukDSpIyAAbddaMBh
hFzoNm8mLILRRI2ENUYrMEPwrBd8Nv8wq5bZGqw4F2P/aUqeDtGCtnGj1FrgYVqTUaePe6Mdms1O
yrCSNGnmb8S5499IKG6je5QDNIAwcTj3YH2gs7ifcSVId8ceFsICu0MjbHnuV2T8qY24Qnumi4Vi
xvNy1BY+TozrFPSJogEhg8CQwXkbGPWjZQV/jKnBtAzYN6HlkWkrOctvVDGvYABdDliq/mPKfyzo
rvd3irqTt52ID2fHN1DvsZtCJZCrXf8enUt12Mto5U3FkMeqBQ/Wbgbhm4G6Z0RzceEVCtCBv4R/
rnhrSRWJzNBpT3sEVj5xsZCOiIWdl80/8G1I5Mbf7u4J6KdX670D0EmEOYfVlKENnsXC2twGRBRn
qNSIJhhiQwRr0c11mXM8DaN4a6kPOFUzqesjrecZfpw1/EEL0bFvcMghMSChOgzcLGSWwzqMI20i
DSgEEXuEK3KM5es09Ybl1N8YJ/ugEsS88hNhPzYU6jk3Rx3bm1pEIrXU6jBPUx9OWXUrmzQtBBaz
YBGFT4HlSohlO0lvee6u5mXsF3bzrVePAx5ttkwBy6bTrEdRRVdnGZOco3+FojMoK4dU/L3/QXdu
K6LqRSBcMyyRefJlb6c2rptHM/f1VERdkpNP0R/mEbd5LEJkv58PXJe3HPIjn5GyckdIhzkocz+m
Ti6JRAzTz3RTZUPDLyTix7PeYOBmhbHnOfAkHYAYdn0bFeV8dwj+zXxujRTQZ2UEOyol4XsQzUJo
Me+C97ukmEZDZ56/hdoH+kv8Jn658e8B6t7bV8J+qtCP+gHhBJDVrREWjX1uKdqwwUq/W77RO78N
ofL5SGUHZb3XsyLox4HAYtEP24vPT88rL0gpwuIwnOxd3sSIGyOiJnMxoGYNOci37j7SiOmISi9Q
+kLn0GNlmm9w5t/gcLeHTWZnjQI70dnxhJpE7jktw9V8gdvPf36t+KHwnZv45q2STeRMffeYd8HA
mih7Ijwc+qrZSFjn9NCTIQzE+dbXMY5vVwyOxoNlnyIyMEprQOQ9Z3FFhL8UXg6B48XYQORGXaT2
8B0lm+zlp8Iq+HkIP/9ej/ojNlWAcN+OBdw37eD8o3b1u1eHPii1lxwqp7RNKVg+Xg/2CiP9XzH2
K6R6nbcHsx8Fkzs5fv426tntt9GSA7GvVmvJI37JqJNXL18rjw/HpfMAg4M8aVHe6TWQ2BXp61H6
51GY1ZjYgUAs9RlUZl+b31+njwfTwoOQoj375sFd/20SGz5VenZtriwUMZkJYjulRRtUrOQ7IdcQ
xS5uwsxRDNE6guzqr5c+Y8j7ced4Zr0MSMaf8KSOPkrHimiSpo9ldSrdrwDyzip6/aoGZ9UUHpRr
Ql/kaIXPliBJNj03e9R5i5PC3rqWpT0mgarrhSiZ7fWemCaPoCFK2e7pnFGO7KDe8AAyud9Qwflh
tZyl6rUpkZpFbzlo+cOUm61iQwoinsw3ztBjLik3LlVYbWF67iledatYE+fzplEPdbErYklRX9rB
x16ABPG+lO8GU1nEWJt32r54kYBGeM/HnIiCHMWIjXRkO+Qf/keHUzAgouySV6RTS8GSV5/gnzUw
AVgOJ+JbeEosbPoXuA+ePEinqgXpOGf2ZtwKWP+zgFgCJko4DLV+H9axwQdlxicCJDlCnjhT/isf
tjqr1yXRVC5zQ8/Vsa3uEGSIOYDJFsd9eyUU7NDS7avcbAP/mY4Z3cxKUh0u/7iEzxtPV5YXClFH
jEnv3WkO3XwFhEAxpKojOYqhsBazpBt+if6a3goXdFN+qCZRP57BcpZ9kaazNOzopO3R04qTSiqx
Udwq4gXli8+nOxGg75AMx/6GHc3BNmGnY1An09VFTMPpsLoMOKVbKGm4+0ZZCp14utHHz1/GtSRK
fAo+hovNR+/E2R/AV5HrDngSJDuDK3KyB08AWG4VOrSZA37igLCV1/Z8/tCVhHCIGxVkO1dLn2t8
tze2zLzOomhBkyTRo5cPKJ8ieWls8hk6tbdd3EmMWmZ6bl8z0xpYbXif3P1ebvncbxtvbuSA06iC
yrXHU309zlbaCesz5CxhHCfuxiMObMUGiXfXPeI8besyG6P4yfmA/jth0f71dqsjh/kHIuWvpJ2b
hlT6JpbRn1KqE6s3HbHZBYd1qYEhoYwTWFIQIyX9c9/IoMwHjVhZOy7U9Rq6Cu8HHt7NjzMN9xvT
veOuuv+3yP8ds9zEFtjDa3FeJ6RzNHnvPYWywUGIuR7iexdbE+73IYFL7hkJdiyjBIufGjv282Nc
N87WlWIch98jlTEDUfiIEn2djrGaeW3fV8yeLGr0WHYhfKPLHA/anlYB5svenN+bsPfwOmQlNux6
1g5bgIHZtJXj+L4SQ82TytBRlGU1+BmCRFS7rk2CYpyDtnLyN2harB4AEpVhZRj8yXKc2B7Vecw0
MBpg/sUWxt88F9s04fUr8ix1Qj3+klXT8mbB02Z/tssqTOC3XKSWBAqMWp4pJ3DSLNJd3SMoKCzS
CbAmyy1tu/2uId/IJhj8HlYInMBmbe2txlptaOyR/fFyrwr9NrpBfsoaODZAowneMDyGUR41RdpK
ibtHaALMJu5uGKFcaL/+eUwMHJbMy4+00apgM3hvb9wpcZFavCnMgoz9pbbxdJUcbuMJ2ryNe3WX
VFB7ooXJm9fCZmbWjIb+li5VZ1K0Yk7fHaCIgg8x2K0fi8i7rVc373NkzK/jZ/RQGlHfQq4aHiJg
K7crMZRQD49PXGc43gP/O0LHdnxYXUfYcSxJWh/3VOyBXpxzMVl424ZeDsbc0F8Unkdljg/TfAsj
iDbixvqUxtPTFbF7HL877EMWWyLsQdzOzf+u2pbpoBVRGyoyLJ4T3Jos9+d56O6iOgXnVgEgOryQ
bognifL8tiLab9B5XnOR8nidxQIyzVt6tqmxZapaNjZTm/tMcNg3nOwVtsSxm3XTMI0/n7tBa8ng
atiXQahd+GOSGrCToFoFHYOtt3UubbUJi66Mdb7jKygZrnDT6EIRXHbBonxdaE92OIR1NljFqejm
wfDShANMoF3QgIbW59uRaPImgsqSFtQLBNKW1XoaGN6rosmsacpyJOUsmzp10CkSyYKDZujpW29y
6yaU6Xv63a7BhbJE8ecWAh9yVZfcL03mR10u0yuoNgA1+Y2FNQRTeLcjV7V3pt17mn1VUWsllNiN
pBK91wW4TQtdG3M+YFi0Z5JEUDq9MDbuNpyFI0Xx7677gGQDiSmsHjZlQP16B80cEkVGlG1i2vvo
wt6GtM1b0jBGkGTeJkSif3fWQtqFQUi+Sm5LG02nom4M1dQ1dSqL2var8r2HZutL9reA0sch8EgJ
oekYoqrFZQnsP2FKdIuu93vDvpkoj81EeA12M6eIU7VXLfMEzfULiJtclKGKg3gq2hKqz0sQDGiZ
rjerBto2U+aG0Bp3VY8hD9HFOPyvgt4Tqhq7He8hpGf7s2Ei5NSYxWFO8LADDc0POTRzYQS0A3uz
zr9guTHkIDwi5gj7Eet6klWFHALDuQEj1fo4IxoyXvBoLvlprHCB+6jUdG2GdjKmaa/DqugChjU4
Ow2Ot95+wXt5nWemSij4TvwiJY2tJCWPkzHICZnUa4q+9GI+Mb0mXLoXF+WpVbm/GWFSawr2T3Gc
P7jgxT8kLqMHUIxd6Y/sR+o+vui/i/BmDSPLOXY5WhRhC4epErLIcgeIvdNeqGwJqtlpIL98vowo
8wiQI5lk2pKhf2BAg1Q7vv3RdLe8dqDWRCjTwkBj6AfzH+XJ243/b2D43iaRoLYkSHFfLag5gf4j
PWM24fwAp2Ije/sIFDRa4LlKOC2X0yS/CUbiPyYyFEGYJ1pT4dnijRLZQBFmPX+qXcY2ztgzMeNX
PTLoxdXC//06AV1bmUT2pz/S7yyF+HuI001DtmXtSuii3QAA9Zp7wvif5zh+EXNlWGlFrPhzoldF
ddOSRUhF7ZBkfav3Ls7wUp9v8KueqcWUbNhdEz4bO0z1yCT0fn9Eb/BvxfCPkMcVx6gv0Avx9hd7
ufR8bkIgOFVm/IuFy2c07ml8lVRnzFf3q4YCwTzVcRcN8bh6i7jjyf1V+4LiaO+qcIoCig0AseP6
fEguJnzf/9a7wNCX9gXOop1iBAtYFPBHS2nduSahFxQZmDLtJSD7OcCtzrqTX95HjE7Nzm8VImL+
ovCqrmfxgUkWHq3rWSUGz0f/XwrSI6O6e3nZcLMWeho3WdxPDf0aSGA6XlP0EoOk4djVBbTTwLIH
/DLW7Ykz0Lfyq7wkB+M6HSOQOb66OTQHLiMtrJIgmbZsViOYX1R7ens/5eImoKoI9gsAAWPuKoQi
4emQPgEQWCmk83OsBwhkcaG1G5DXNKESdtmifpLNle3RoL8v5N+wZXtwqlVezMRPRIR5J3eTQX69
H7qsZ67a+8UhgIlJaw5g6XuN9uwyLFbJfZaO1BthwOE/+y5TGyNJXcq83ohmhDZnaCVqo4Au/Piw
MFUU7Kk+lWZ9yAXRuiYXmHveMRGfMSVWN0B50bl+Jyoi+9BCdJs1neFBvdTCOJ3xpvzYLGeS57VI
0YliMV98uAKh4lR3kO2sZX2qQ8tjLOrl+RDPe0k9zrugkZLtGWBSzTUKDamMJGzMFt8RFJjejG3B
BHMYmf8phbvtGwSkRDiBSTSZ6TRQbVZEi3cQDjBZCVcLkcMkBBztGr6nFUwUaTka39TIbMmzbIO3
QZeqY3Oi6s2CSL4nnjxzRJZoeZt1wXvwv6Bd+6nYa16HJsXQUW//FVl6f7tQKTNLllelMH81THLO
KVwFeZBqXyuUiJSaLsAV7z1I//faBOCzCq4qroga1OzAws8zD6o7dFMZQzJldxJSwogsmTnr9lNp
uQo3B2aHylhg5XJ/ynd8L7tI/CkuDjS3VSQEVzTXYuz5UBNzwBZPVuz+A4vpKBp4GJMnXPxxjHSz
mDegXzyXMCgwmmAGpD4HTog4GjiZHD/CxDyT5UY4kpX/AMOgnlcv8Xxaht0nQykkt8JCnbZyT59K
5/Au0DvAxfPKJzUdA+sR8ZKvY6yTYQwu2nIeIlbvUUZHB4ZFJBNCGBM8FgdSra10drhRaGhqaAKa
h8ZcvpyDkv4in0KZGBqlXeTSFDjw6nVPWmlx2dkkuIvyo42JJCRuALd8GyFfj9c6QkXgs+g9Y5fu
TCXbtY4dqx3D0UDwG8ym+4tuztaauRC8Ih0VCdRtPefZO4uu2uOh+/kassFfeDwxQyCHqxV27r1C
HSJxGcP1kREudkaCyISeIrAUmRFtBjvYRdJ4Vm/BY0C5NNGgK1EDjo46jI8rUdDPfZ8hHyy/EhvK
h48YI/UJ/VJRgQNFuALcqX3e2tqqDKyzjfn3pYjh9R0C7Oq6Wjz6Vo8tTBBfMLIRgvsP1vhU0bjj
hYtZbnqkn68kevEow2yjPTvFykT9wf7/29XcN85FIJD+yP6RLe2c4T/SD3OQIzX4rvD/9ZyN9hBw
8RoDAmjwGw5M1B40ymsgh4bsq/6XYkMwPTHAQNkcuH2SFsYvUENZ8TiGdIE6oYWD6NU43V1TtVsi
/4Cla8ao3dvBdrAvjwLJ6fAuBTR2DFL3U2Gna35p3zHeCWtcikA02mnX7/oPwJDxg5c3rQwkbntq
jh3NRImaBlhOFHTJEBVgT3yjaKSgila2DQvcvkn8EDYot5QSTq7Z5oBTr+0yt6Zky+4YjrO08uh2
7y4BwCkTDgUCm/juxSZyezVcbeYME/uCwdgxwfQ0LjI/UXtTBffeH+mf2AiFM/b4fcKoteTIlt5B
CI6rqcPkL+wG+UhjfFxe0Q6eETY1JPPpSVjHYyTM6F+4ws2Pnoq/JtDFh/5LnXzEf4V1tX6WYm5m
cZDamSOqvjlq8nye5fLD96t2nR6pXLZpBF0LUuSkVZCkC5/q0WEKxg6FDLCI2cnpMQSJ/Y+LbAN6
hlQ4gHx95Y979K7W5VDScaGQQou7MmCZMfZk41i74jAKnH2OxnLkmAj2RiRcSVWLBqllT8UrLk6/
P95ZRSQZA9O95g2JmdRWc5ibA1mHk3xsk6dDPVTFxtiTeeNJwNE/vlt/0EKBE2wpfRGENCKicjs4
I1PGaBIEDNUlUylP9aelcpIRtFvLjvN2M/sdSgixhu62sHXHWbUaD1Vs/waX+w7z/7zeyYVugK7N
k9Yccvn3H1RjjBrJ8YIDJhrsijO5AS4glivfIGeg8oMXgckmnEYz966aXA1kXDHADgaQWkHNoroi
ZN6FyMjumhD1+PdGCJ0oUVt5xwN0WoSBD6rFUFvyRxuxv4uK6NKxnbAKt7ozqJy4eJrXf5EvxTJs
Cs5+Vh+VbtP98LHcRifCxoM5jN8bwsp+H3O3WX8qo8Gao3pNJsAplOYpSTeNRjEi71MJ4W5x5Us/
J7u1IqwCcFHuBLL+SgokqJxd9qm4QEGa0L3drSh1RVCOT0pMyubTDT8BhsBQFSS8vaFHPzTADgtb
aovMxUjLwgScLXTY2NIV1TM942h7t71JFw7c5q1MXL4CPIsbFW+8BlRHSy6J6OXfaOgR8We4H1io
LKlk/KWneIsckseIEFhEkOXg2wFMNOfdKa9AyIHC+dQC5BncrnMu55k2SAVN14192nS7Kg0GkSWL
nA2ISqRGSYfuatJumWEB83WO1OhGu8YtQ/L/fA6vYerZnq3JjAt9xo5z1Z4n5tEkDGCWPIFCjA2B
F8oV+k7DPEK+lsqxvASfKed8SKDZ4fU54nCkEX6eftiGOchpz9ek6Hln99NGUhFqj2pXV7QFzdYI
5oqxe/bKD7w6vD1Pe2s3eMka9gf2U3DueIDwW5XNQKXfJFXRtjTDZqcNzJpfr5qTZwXX0d73W8yB
IpjAZpZRPXavEbL6HMF4VXR6pfYbyCLksOdssPeqTiAOaYK+m9iP5YPEFuCw0n8g903GfHUxjBbl
MXhJ+LvQ8CI+UxkaZGZQiIvdnAEjUv7khJemAhWGQ0AnOAUYX9CbX6dsG6QDC8tAXvlkwG8huaOK
78gLFti29puppSJNObipWIKkSFycccbqAIB3KIOk76H5ucoqBfNe4TZwQ2GZD32rXufV+8mf0d59
C94wFvXeT6JdzQNByLVqaTGBTDVw6oRoidzcYx/YLFQL5qq6svmgySO2Ys0/KPp1moc6k87uxMPX
g27iwb/CPVyrFuz9LRaK8lRE4IODXbMoeZUgJ4kUcsj0ErZOnHPEE32p8JFEEaHzsp9CJGFlIgjs
mPgl14it3pXC0dwTJVxRd/zMsG6JPbkamWtgCIFtD3po+fIzu57VSEN9WjLJ9X7a1i4+0R1duwqC
khd50JmYS+FMPm66Q3cmYDSvCVUxMryrN0nHyZQJEqGdC5yVefw9l4qpphbSYjEchX504wTJaE92
06fp2jV7JiX3H7iVIez8Cd1SR9oWfGzP051IKHjAJTmmxlpXu3Zx1FcHDJ5xXD9eBiOqchaL/d1C
xTmm7dXa302RZwgCIt8OsUztBGRHng5LYC0OBdjYLoK06XqKo8GyAMlb+T/WxYsmfAkWTnGC/Y8L
/d+3w6wShoFynYdF4W64WhnVM0+PiKEoRk801+D1wDz7yq4+L+2j+lp8EjJXXxFbk9NyAH0UVVCV
gc4E1KQ4iCHKQUF8aQIV5B3ZqWzFlEfmuHEJYDxyUnmXMWVB7o/2qt551PFehGKQa7oPnd2fmIqN
Ius6bES+m491ikt6C5D6S2PFwhnsBvLJbalH5cMrfkbn9pEOH1t9NHwwaO8jrLfki2xKok9D7l80
LlyKAhDa/2kjc53tEduz+LVSbjfqHYYtR430K/K6LX2uCiI6f1CBxfMORhJO+dHRErwFaab8r0yT
6Q8Ha2pbHlphD5haBqvJtEfEY4or6bIFSxdfrMmJ1vFxlTOT1S8z+jHM9noc0drjLOlk6/BkGIo5
Idz1HE6Ur3/OFZ3VpWVZ8dW0th4hTWLM0Eh7wHxFVgTAcIpq4Ie7ShGWoWw9Vz8eBYpyAr2IxJr4
yGGtaHphgsBRiiWyERCzMNUmj/a1YxyE+kL50loNssOSHpDHPw6gk4S4cLWgvHsFshGboZogHhom
boobQT1sz7fYSbNMn526rGkgWIIG9fF6JBe7q+uxZ7pG6Q80pm1BEhtbUCL3chH7ACs/rWaIxUMq
W4Mc7q2RE+1giUhZy7BEjtzaUIM9dQR5R3p2eTmXj/TGL/94YC+NifWkA0wA1oiWwr3tmlJdjVQw
TrNMOvEEHV3DsJOXPsJDYIh2Xo59lNcq36AOxrUqQg7Ex5D9cofORN6tmITSvzkl3e/2Jvw3/wpm
8BZDKJL8EAW2dOfdPaAILv2zx5dMZsEtBFJ512uQa5cSGKqWSYk15b3W3O17hoGDtyF4Jqo6nokB
yhdmVk3eLN9w8xsW1RSe3db30CHBxjXBuqsyo9SA9gvB3gujkW84BTvfAFeE4SjH+hbTF2S/x/nT
ee31lIoNXGpkjRV/7VeVAGiqBn75SWbzpqFH5G7YQZLUiHmPq4zGW5wVdq7p+61WI9PTLJ9iTG47
OIeYkaZgJeiIDPgD48P2pQHtIfq8LW99msnuDO7Ge04qP0jQT2h5ATDb13pYDFFeiMOgvYyxP2B5
9WokKvx2J9PJa9xRSZ07lK51M2U5gLo/6HV9DtoUEGjijWv0dcskm9KmozHM6+kwOGnQGDA2ySDy
OmQEgR8iQjekMLfw7Gv8wvXSi5e4uFdk1WurcB3VuuH4k6sNHj921neTcA/YfYyVVUa03NQlL08P
3O2Cg05Ij7r0YeZmZtIkxM9emD+z9iFL8z6WHkgtFqYkki3VCYr/9AegJDOEAsmW919Q5xO9/c0D
hq34TDdYzc8iTC5pQ8BBFK216Db+6d57VQMXz5//+RF6uXlMuG3qM5Ng59EBxz69cC1h9xmN2lJ1
1gnnW2kCiURxKX6N9fYmcM8stWMLRsfhgsdWRi04mvSdC8DQNkgCXq5wNzxjQfPzjjf91aqRw7YP
ih/wFX72hlbw46nLCBi0B7dkvbmsZteQ05U7st5fu28TDE+uB4ZwjtLu7baW4MWPZPwRlLP6wasd
9Z3mu603Dpn1a08fYK4xhuVtz82G604phng2CGw5af+93RITmyQSusQgYLKCNmhINcfTtXnGvwba
aHAQ0tLk4Zw+J+GXUe/yoiGF8ZfFqPd8f7tgmxBFj46Ird3GAAcM7xIUH7kKDAg5CvrIi4EdO49V
UHfLB4H5irdPppQuXi4gUVQf7HTo6LufOgmYNZiZjadpCC7bPHH4HPsQ//Abt7NEzykMB2iIto2e
lZXt8B+3lMfSYG4R26X0kPT3aYtlaqtoOymyF7t7+Jt4dsQMHaptLZ2KFusTqZ9k3dvVhBO6F/mL
Yz8bN5WGas21FFyY2Yy49z3IBcU2PJFNEmT/zQEad4Vtoly63euzDI7YqPsMpVDuXfYSlbbqtyJ5
S4haPtT/VwOskDUkeVyikB3gPb/yksuD7t38C2cAiIP9EZSByOC6PLqfXu8HsrBaQYp8LSwvKhJJ
o5XcRY8IZkeMC494cSikxrRwO5iydqKoT6O079s/Y6w1hbwMI0+ft9L3C/t0EYvQ9bhRaA58dwgn
4tHhTPnDnx2DrE6Ew3XLT5V5Q6IIOS2fDXCelKz9DxBadaH2sHX6aEK6EvgPRp3Wh8TSwPUFSh2P
763V67yT6YvCfoTwuy0VsNZ9jo+spEAKrU5khc3cjHfeMm2Gn7QA0aoGSrfyVtiQitFEG8f/rEo9
XwhIyYimvrvMHuMvImAcVS3zRJlbAiIgSBSRrWjz10gYJFOPnC2hEE+ALpL3f0ScO6dIVW8K/xFQ
CB7+wB/bYAvgp3eK7b8QPnqcLuH8h9dl6bGsYe5h+cRZ3ofUqtQVPDjVKNtKvwmZl5hldRaD6GpE
S7wyVYwiP/NpWt0255i0En98tCftLkglAGYD1rMSzh3ZkB6ncSJiLkM0ZZnvyzHeWC9n2n50coSC
LzBK+40QgOEfgE4AG86fGnTvB9PKRi1Vif4hyh8oj5kP6BEa1Snnzvuor3DFWhGShVvkN1xLzzyq
zeNnWXrB6mVHXXUjVm1nD+ytkXGz5DXTPwz+MgTKzgKTmNPlIRbN1FaSTHQy8kIEOOL5R0mm93g7
Nb6kVFp90iNFNdkYHd2S44jQfDTmDPnodqj124S/SJB47CZWtGlm78qBvxwV+eFsoZSwf9bY/GLC
UDSpMKzw1wk2MajLYggccLclVXBvKiDVTNblweW5rxt++m9MHhy55DTGe8a0oc41kYuwc4Z1cKXR
Sj7WnWbfEOEWC5ol83qv1caOYkeUjjTwNmQSF4Vs1CCn2mK65K0FY33bJ/BbqZJRec1ELujEQqBn
4Ti3DZofx/PckiuryQzKzEN5WuCPFUbLi8rrNEVWtb3dbm5wy9Yjupa7FF2unDwwhRKmN9aaRtVX
FtTzpq+YdW2UERPomqhoRCoXrxJ42n3yLwMk1TGufxzEQsH/+o7oIRn+hkTsck0zF5vt7XFcJlP0
wq/z1IjV5h3xyXiI79P2LeH58RR+jCuBWeB9tWB3sfug5NUE8FkqdIrwbNkFW1ZhvQLW2sqwm+pY
UsZBonZsE+LN6Qp+ciHMo9UCEDWFM66n2U0GR4fZbHhXzRpM98qoiinPaModmBHgcy0YUEzpJpJb
YrTuCKusve1lQr9O5RfSITBg3bT0SVQwiLp/BI7zyDtQ8E5fEyLrtcYOfUeYusqmq93LsHGiq5pv
BiZUtmTYgJL9t0dPJ4ffj6DJ+8scjXoos63x0sXWON/f5gBMwpvsK5KW+VXd6lMTw/Np5itH8bke
rfBntdkay7TYbBRBJ7+6q1YO1OtEI0yBt9Wj8z8bbdiNOGee3uJmqzOhtsxO82w3L3Y21kean/+J
ASdiNsg+6BmXGpalvwXazmPmeqSL9iIeLwTJyNOJe0GaJku4yWO3a/uAdrrY9eHUr6phoHplDYPV
2g5xzPUZkDwLifz4j6nlTTOmM9OxIYyxEuaqN5VcYspqOXFY/a8K8tZZP7LsxVADKDY3ioHJUK1g
IO3igWbBahGz0ei+tNl9e9Hv4tfXbHUy4JZ31RZq7+Uwog4Zl5U+xdXv0FF+gJd3aQeFvydDnE1p
sUULlbfxH1EMb60xspNqpzCp9d8Aj7zhQwaNwSux0/wl5d6mnjU5uX66WJJT8Zzeo+mK0uHOUx8i
DmT6Jzs/DXdn2alrXZlD1WiyeUN+t62Hqzn2/nB6cVt62bwoAWaJ7dScxq3eNrUJTYf/RQFngqMD
RTwLjTihEkQTMor2VbGLHcFeuaizr9YoCs2dh/SK0D9WLjuGTZcwjzRqgRxHcVBC3v/CMVMKtPMD
l3SIQ9JtLz0XXmrjCHFj94s2NkBtsyw30J3HVTwYrCij48zd3lYhqGfe44r/zCKPHd/5x17uSrxs
zhmUaBEchM4zedEEDpS0Neati9m0bOjeqp8hTmmXohDGDjFbT8JWoqle8qXo8e0ZGOu7ajdLEXaj
b+AvNjUEVl8qc9VgYB4EKDD4u/u0SJcsmcnVdaBglYEQdxYWHOqrnQ3gwmkxg+vIVP/jzA/f85df
BsNPxNvEQmeS3HYYEVKYLEO8stw3eZD5wi7tD8kq4sNHS76RMniIs4y73t0YG78vecDFFABYa9Xb
zJkAMMi5E1iwxp6OEktXrQl9VoqjOuQov3wKGMwi17ElFrI+jBr6+YuW6X24W/B5gS2JNeIWuWLC
RhR1CF9JFlmzYLSGAJLwT3U3ywjHt6+5vtNbiuDwqbf2yvaeaWmXLnv4Jiuu1W/jzVsitIegLFGG
twvWuWCmb+kkXe4PbsX9cjzf722+zbtvpBRGBjf0O3sMyNdhw+HLNgSB8ZzJqHZIbk6u54G6K6mr
MfstzBTc07f9R7SWhr1JDhDJAkwCOxJs3L/b1c2/ICG2y3janQWXZzvGKxwPNNgk6PmzwgjFXWtB
Oqbk9Fs8GFmbx8lWExy3GOvsiMJ4NWXhki72McHL7YgkYu4pqWYiB+RPXdEnYR01CE94IXiX6UGn
JVXT4Df630dw6243jbW15NVReOeKz9H9iHRYWB1/SlyvL2ipkEPKVHYNKtLRY557X3GefZjkgCch
6Lj7vsYX//binhYiGPZ9T0Yzz5RBbaXvfU05wYEhTsWLL4soXFklzWGYAlvG4DGazXqMCsoQX8mZ
6obIGo4Qz+aOj350MgjWh9RLh77zvTUA827JsLCfPm8Et8BrZbgjAe4LA8SM5JqBYAlnAR5b7E5W
W+YAdlAG5NriUFdWru3gzIazHH36Bmhpreoeiv1nEtMIEM+f9Sh7SBSh0qukfc7N0t8eK3oVeiAG
L0ggkMQeDkWAEY0P3wMClOF1KaHGxRiw8H6x02q1HJBaA3G8e5/lUnM+WBzdgouKqKPA6XJTd1o8
2K1/3X9JYX86LvcOaLil+4c/T1MBD9XnLKwNQmEszI0WXjdCmCgpPC7xxcJfv0/Pi8GBtm/kb9bU
zoCnG/rdLsxJp99wvNyxLUxV5w3BxX2o/RGGRTMYdSBXZvDwv9u0CTX1M4euVj8zrtKkdVwEEovq
7+f/izJuIGf3N8sLFY8487UrfaCoDYntE4y7nM3dM6R1xIk3FruO91zJeywdjzxBPfCnBw1h9Za6
vm5NZplbqqmUwRn7VHzdXCPh2fdwfpnYuoZVkdtfqWjgKD0nt+99IHyMZJ4ocBVA54oXcJ+husTZ
X+7YPZKoSQdhhwEW0VkkbyRSNUn4k1Vtfe6R25BrYbo7PNTFsjK1fa8YmT1YkrlHZWbBZuMNmIgq
mhzZPYgYmPT1TOEDuiS/8GEiano0cV8thJWjOsgBgJJqf5q5gG0ocNJbsqJgNlZrexEb+wb3Z1T6
KV6Rd8dgU1Lrm1EsoryIp2tu5B9vzjfiH53AqkVdKiYcoB6uLTOHWfXGoCR/mlkffT5Wxt5m0fs6
CPzOU3Lb+KaHuXHWdQBE/FeIQsRMaK6eV6YuD0ikHvy3+sHPlcAFiVsiK/Y2Q9Q2QzgDHyq/S/tq
9qACN45iKR5WIptV2ot162gN/9GoYhmRg4ZRxl2+P6tb+hC6SwXZln/nT8IGPPZhh/aibTu31RzQ
ZhWlHKsG9DY6qONkNaQcjIbX8K9RP+/uMHOnRPj8fqeTMmnaNnUzJuu5GCKzltVGp4JLlN1oT7aw
X47boX5LhAkvY2uhpLW76kyuihvjmcHa3roAXiizmXg7PA6Dj6wmrCpdXPk3ikqcfjkl8a2GjDtD
FfIWNHrRgGbcb9OUtRVQ54dZO6flVExvUMwWrW3KL8izzeMDy1lN7Y4Hq3/+VxM8SczNB7XfclKT
V13IJ0FVN4lz1QtCzQKMhk5Sb5b06k2A55trcyVHfwA7n7q8iaNZ2uRNv1OHyjr1ohydD6Bq+5y9
iwS1YwCFzB5RP7d1vsBYctRLnEun/V6q1GQPEBkuKsLWZYTEqxZV1vQFpkKHhinYsA54roTXquWG
3Wq/XIeNLdIhi75H1xWrwg8PyCFt6hr1MGK/NjAKWHD7X/ineRRCfuxxgyuSj9Xv3aY6sSD+4gWG
+tGmsbbtXRxnk2hkWQYp9sTrezGyV42K4qk+5+U+4iIykCGl9xsoQkQUKnNP16YlFFXqFBmlZ+qL
sOV5ZD6wwMSxTINfLdW6NnyhdoaUkcoKZgM2PY7P4oL3ztyo2Nyjh21uks4lu8/bX0voI+5g6ilB
GcSrXoCmu0zSc/sqF9hmMP4UixOQzmSai3rtqokXKDmUvzcRwsHoaEtOObuZwvJ6dQnyDw7EhoJb
nK6SolVip2DbocxULtxAEBtyKYefWzsdLY1irum4JyBw8rTreYA57DTaG9kVYKtfNoixwCT9W8Re
+J64ixRuMc3vE3KU+0JRYnxbkFO2w2xK7gZBLWiganMPmvnAq3fK1ZLsuD0z2DEbcffHi0ndfsiF
3Ujl7vMvGd+jg0eKrBGI3wRZ3/T5A1byJJCKn26odIKkzWjtjlduI8yxyDmPFUFmx8y1TPztNdsb
eA8a/R1VwkcyhLRTn1Old9wqEEvqES2Wyw3a6gaPafaoQNKEMOw0MpGOJFWzdPJFXVAn0CnJ8oOI
hhmJTDgsprhaV6mi+5+GhD6SrP8z/KCHJ6Ct4vIheMeVk0r5fWcZO0u0xDKG3CvuphW2BJ4yM3k2
S+YZYs3gTjc15S1yZmJoUETyeBW9zGHrAd+G4cac8ukekxF8q3OOkyY2r0hM8Zt64mixDzA4k4up
qrFEgKkyV3j8OOxIQruOSF8ZqQRlQmzG+kvQYME1ZILbDWKI2yXAsXvTP7pE9Ukjf6EDVC9c142H
mjXmQrE4ixcl5MxntrZdpuTymMh3tuHsUr+aDKOteSPsoKfSjZfe+7t0g3sgF24Uan1zm9snIYoI
ks/4pKbWZrNp3LUe8S+wQynw6NVv6oi+ZPNDqSYNMvKknJxyrPqi4l6UE80TS+i3WUgvVJ8KOeHQ
2lGPxRUD+K/FjIlE9mJHVbSg6NT1u15cgunlRcpHWtlYENX1aGCMrJxkfZy0guUaIJuytFCUcDNP
wYUfjfsCYaKGx3/oGysfZjPUqU6Tidv0Kq568oUGdDnVtDm29lTnNmGCXF9VUbSFC8f+JMxqpNAx
wlEmmgPNPzBMZdI33v0lRHx6cEHlTgj8ymHuXneo/2eeUpzAPJfRZT76KS4IUkhkw88aFHP1H8+K
8MQcxGPfjqOXczSyfLBm957FLs0AeuJV2pKiClA0AlhZSQbNE9LTHF+WJjNiOpNu9U0p5WPku9qk
Muxtz1tzK76bSFrTv2M6x2245co5Dr/9iZDrM67Ytl5LLyzMN4Rw6fttctSxqK4yQqhxUY8U6uO+
zlc8CTJCu60FNmlGAenPSzFKfbIw4ncxFKxMJkGYupGalT8Bl8sH+xba8zI/sNTlpL8yjmmU7p2v
Usc7cvr/p1mbqEracUSwY9fitDkwG3avB7JuPX/91B2N2aG+qiKdtIQoPm8Xq5WqzttOW6yG2irg
zy5GbJvx0E+a08sBDiGF4P0iACEsq4LAOfsvI238CzOcY9RtzX9O9bdaX4uLHAGSyUAZZkWgCOlD
hk3ZQDOqZ0QBDRprx9gxBnlndlCOiyfidOgu7r9kFpPFZ/00gXqartNeI5qtXxRiD0rNOsZBgOXH
xzR0+ipUaIUQ+AS5PvJYNtxY6PINM0c23ckmLAz6cloSf+jD9kp2JpBFKrAViFgDnMCl7KIa65E4
7rMYArEiU64RDMsdJgkDCNpDAactKjKqYjdUq3c8+CtWknos8+cCuCOuJBO/nOPdvdRkGj5aLFq6
iBQi6g0M7hBnsFTN9tAkPXBpQbfivACPJhQlV+fNdMHdkfhdkjZHe4Wv41bKlN6cvgpHxbYq1JQH
Lipo4JPnXLyxQtgOGrUGiT5VfLZbJIec4i/sz83G1mGB+YwbiyBew55hNKKoZloXWj/+WHi0AWnL
mEPmmTiwCqisfhRe7eHOfFWkwsHplIHsNJhiFj4byKEWOXlCdiXClt+Nx7gOFgRQpUwkVwvFNxhB
pk535Kzv1Z18Vroci3beuNx950cyDlID4+1h1ftEyzSqhTX3rhHtUr+whY3ujP9gDckvW8fA68iU
0FI9Yr7RxM3HS7fx4cHPSpy0rz3ppHveTwFIr+ObYfo+EfWInh/knK7pRqX9eEG0cKkgqwql8YBF
QbiAf9dI5emA7zsADOGSteoMMrMHG4BmVfQcwmowyavlFm+mGtNEXn+H0/8kbCcSluMoZNsOhjpU
QAPRRCmepr7wCTqh+tv5vLHV7nocHPGUY6ounIfu+9Ok+jjYO/VQRYt5Hyx1N1BNRl2sxk5AOinl
NJGBbbwPzx71o17OFgWL4FHYDaU4tI0YXTF4UuvC8a5r/HqeCmQzcFESE1kQZY8LonBi1wWpOURQ
a9zQSdC/qS0OAiF6LlYChx/eVlWmmEs/mfSx77J2NmqoJ9MMbZ3uVW+4XEIKW5ui/A+AuVxJfbiw
z+req4H5Xpi0HRSzcWU9n7OT+qE87mU2qvGCVO62E7yeoszXPae77TbHPEFaYAym7f+Y1PhcC+ea
A//ORx3ab9yD6kiJ4TpkwBZ/AGbT7SymnaEeBysPYHrG8NKOT27UujUBfRKVPc5x2EjESF3aIzgn
iomxPEQszlc9YFG3m/Tyeu+A/a6xTv6QnTdbTbNflk9ilXVnrQS7Su/JkL7iX6Usw7E6//QgMP02
0glbBchGkPEJ/GcYNUN/mer16fzWp781W9oMvBAQQuu4R0Vipie1Ov5d4nHy2Xa5msCDAvM74C3M
004pzLEsdXzYMQ2jTOHycWuffDo/wXHjrygAeAbmxmTwY0HolOPsdpYfIk1H9fVe2yd3Haj+mZqI
nIEXmnatd7RByX6KJCGi9CM3A4KSdFidjVyVAJJjqzX2VQEZbu/PkBpKa2dqeOna5ZJ42cHdNjWY
DbFeEKdqC0RKOCfZC2e5WEV23FC1QLoq3LX26hUfCGHo2uK8jrt6bNUqiYqJtIe38g2aUW5hUTkq
FsRXaX29D84xWCAeRYBhPeDwCHprgN0RXBymGg5Pudfyzo3yMYxGTkD/qOc1jNuvn5SAl51kdF5O
EBQY43MG0BtUgU7a8wGeIoG/FOEDQiDSaZ15xUgCFYX8ubp1tfoPRZHqLuawppeOvRdBr8bkUMmA
oeMS6qUizncc38nGviPwX9076hm3Ju1RdQ7UrNlbF6JH9hh3iJw9REdlBMF78/Hk9qXK/cdYQ3UY
dXubNDSR2TCjeNMMwOGxQ8sNKZ247Gt0jquWoqRvWIWYQORGG3yi4NmBALFNmKWFAhMZJxUB99Wf
cQaFD7WTGJKG8Jer187Cxc5I7o4nKCXAKRcpuIAbVL5MIywX+E05dAoAsZWO0i9YDTaD3PtKzUzu
PMZmaGbFyKp3oq3pomWc+Kvhbs7+eq706YcDyp5GHq6jBVmO0DSwAPMAq+HLc/gqbKWBazRe6tiP
aWJW5PhXWHj1AhEXeoIGDhAs/LkFObeS1T0k+eaSVLTDS+v3ak7TGLnLX8Tgk+j9wImtxmH4rOEQ
5LiARHcbZZaDofCg2LCDpRhRVUQ4sD4j5Fb0Zrq3conrfEkhRLrDR+ymmOIYvM5wmo/XcwWz06wG
TnYNl80iKNguefBwdpjKJ8YuvBFVWOOap1+WTrGXOP22FvoFktf7xKlRGpHPpZ7LfNRjAQCOwdgZ
xM0w7ykeP5g3Zltln/qY2d7IKjHsP9INNDy79t0P/iD2V0GiY/q/UPVcp7u+cC9akUKCcYlHGROX
W7COQSr5bYgRYfVAX/wv/YX8NOYSaLwJnVE0KErZEuF1XLcOKKnHH0k/lKCO1m7KmdUEDkErGXyF
8l2TF7fhSaYu7z+Qcx92s/CiVLTW9Ik8N2dUr0ImoJ7yjebhOkiouPoyf7GWmWy/iaXnMx9b3/wp
p9/t1RQGMJ8L5Dhd5PhkB7RBKp5bHNdshcpmEdE1LWPUpjyrtufs2DrIgkhXKjjGDzR9UDpVIkvX
lfUBvIcw62cMzD9sL0jvyakSG4wyA92qWyuUm1PnfxNQxkD+5TzQsCrMHw9X8GsZKfnIZyiMLxOE
H6969X3eW004Rw3Dc85QAXHUdsoEQQLXincQ/jPigC0x17L7e2gUOV0clNkdbcteExDNHgv0UIfE
k3ds8SshtiShRBB0oUTb/i7sQ7UFuZZSKwyTC0rV14+fvNHEP+fgBqr4VBS4gkGrBv/YvLtazN97
o3gdr8F9E7p4s+veAexwEZlhizgAJp+KURBily9gAe2E1D+ddNh3voqRaeWiynRIbMU2ussEJLV+
/pthK/H2mO33jD81AiPzKlJeiYzdpc9AsXTT97gJRATi3545RWN6B5xiiPAmae8IVBJHrm3QdIKf
MT6/Xf2ZAJVKPsXzwMCynIpTFomtQpIFXAqxhWbDbYim8iBhF7zMTbdPG7pZ7tG861+W0vm1G/SC
JOgAkiRzB7Oe39yNhQ3w2YmQ4kuLsOZckawwlGBkAketilUM9AT+q8eND7DTO7vvQYZ0F31o70AV
0hkkBmShPlpDAjzhGNZtgF7xqXC7NlrFGA3dAqXNLnqr5cFXHSqbQmZrzJ7CFgGT/QZsmmIQjU4Y
dFxhP0/vahowaEzNv4eg7wF4qkcWCgV44KrQjJyfHnD3TiFUUJqZsCMVFVAcanK3rOOjW8VrYPya
zTsD1qa8n9Bd0AQy5XPaOxWf0ec88QFFPw/8mI/oD8Fm1wzknGTEpUd6pU6PgHmo5fYS4h8X81qe
zj26QmD1fZC0fgC/PVF5t/6HAvaahA9fdD3HFZGQUB/1XECzWPn2RocRpHPU0ildoMNv/+nNZo9b
9uNCExHVBFrMbhppwnFNsnAXMf/F2JVIsqQgHGrAnkyptCiVtaiU8O4VMZ1cMCNNAmdIrr7Yd05D
k6Z88nTRmXkvCvB5FTYG9EijM8ghqzJ/pnsStE+rd3tbyxQYrw00ZeUdz7HxBl8Kp/pBrzYw2y3a
hwnoP8Aj3FEciK5F2l1mfpaGcsgormS/TMukHH7W6IcAgZ4X5uRhBIIlIWKft7FXmzvTvKC1LS4j
LvArnRBddz4atxaQgK6HE/L39ctUgwtbymZK7OfZzanWIvfJjCUSrCvYPRZ7dryPnEE+yhlOOk8x
aGOidr25gdNsEC/dCk8taC+Fm9TK1GRi1HuVRVG7BhSIMTjvIDXZcac+yOpjS59wmwmPfZhFECiA
+kU4/X9Bu2DavoAk8Pr9bi5/QFm01qluXBRYPZBLWacTaXKwRFtQ6TIZ0jZYwDKQjlQy7Piz2hid
i772RycQntTRkyZugSsOx3Fc9QsxLWyuuQxXAOs83NSE13aKHuiBMwfls13PrCHmtWMjCvD9kstM
Z5lyjQKv4FfUuPXVsxY4Bi+ai7dM2z19jTvAyBIqY1MziLCE/Tg3HLmaQ51/Gy2w7MWIg2lND9+2
yMRrGZoQ62OJT03zDYzizpbpzC+5g8ci42PFHFZy3uo6EjcGbToDRmLklP1yeBtg0Nz7vLRnl+LQ
3bnYbCF07NBrqxEh022jfwPSzaDVIqzflAOAFMr1xbUMzN2uIt7H1te0Ng6GI6SkdYxrOuwmmA7L
5yUjC7TxXzCp2QP+Gm/45HQkA8yrfxhLIYiB3Yp7bZBLbLglT7cbrgpFk9ZnWGTtUUL8fiOuoCJD
MZwnIb1OTLGwFRFTYeRL4r9LgEdhDH2EKtiP6rJwpTiDKWIBliZkjKzFwk1zQkxmWMdcI9NBot1r
CAIhbYC/owM1nwK9IPhMYPpqg8REhIFoqgd3FCm8XAKL3XHHV4LOWBwU6xkeQa45qJcLniAdfFqs
DY+WLr0IrRY5+EdPyH6vV59vVTRizTBBnYdgk4f6I0IDTMr5m0tlnEzDtUtg80wq2scyKxUu84Lv
K/f0Vp9dgCOgmKv49nEqoXyvJTKFRKHc1slp8fpjmPo17qiVtEQr2XbWf4xNLqogUN7/ceJURC9G
5+eXQEsP8twvAB0yJtlgthjoi0ph1WFKyLpH5O4Zs50X9q1Rh2BFAaN0w2p1lTB6pnG4G1YZPR07
SeB4j/dVG9cy0dp/rYEysrKesqqd4jZxDsQHSDFOdK8imqSSvgAo2GveUIlyvHwKLhhIjDHb4LI1
yeJPHs8PjIb6lAWogM7PRgQEHTdRg1Yhe0pnNtdLRw0KgxPLguVpba3SWkCVdsew2qCBpfeEpjFa
lY3KSCdDLXWRmmrQNN3yU0HB8qOrqu9YUzV5cj88HFl++yJVhXoQ6Bb064HBtO6wI5W/EEV+zMcz
Hqgaf5kl7tpb6S21vyirIJtnt5FBnNO+gfCmJyKUxh/KB0cXOHGAameEMWRMSXbpxy85ZAncc6HO
O2cTSssFR4PdBzO/9lrd+NRko7mnMHclXBR3Sl6yGGDqzk7657+GLRcaPV3T5HesjHw/agUyjBvc
+Hh+vv7isOHchJdEvPypK6P0wC2D+EsoY2RPONrupE0OX/VW+FGTLb22xSAGayhdPphBoMZoI6Bg
0RU6sDQs4/E3U8dOjDiAnl11HlGirJ3NivH9LP38lCmpy9BaiZ9EVkdQHmJ7ElVNkv2MwJg4j3R6
8575MRRWHDb66aejgb9TiRUNqrz8aBAaoU9Fl+CACHqXPet1SZsUkaablelEaQPJfsJTCY1MsP5h
swZOdZs93ZAYeleEmuGbRU43k0yApyGN2dtFoKIYpwB9MBgBf506JkSIv0MX9g+1TBMos7qX3xl/
8rYgr2FG18hGQBj4cU0Q3wwJagIFXy0NomGM1n6RZEKsIfSwHJoo1fzu6r4dAM/3E+s838iUrEEe
48SsSoL6W6moBUVgcdof9U+4jI+swUexfBf3TyOZiCmik7E7jiH7rqJNmXGMgQpw9hM7EhmU2pgZ
FgN4Ubxls1fKJqA6PjyT05E/Ztd2llVFdGgLtHJgQSyglzIcM1mauaBIvxbYH6qJgQRERrrPH/B4
oRhfyq8ELfSPXadkY5D2Fa6MObW2zTltavzmmdSTHj6bAQKd1a3Szc7uRsWaGlBSqhfC6E5Nee9i
IMjQywEbfyqLTCVIeYWPDB7KhyeTsyoEU3iBz1Ev1gDc9wGJiHlEWOfRpx+X0LuSIjFrTfVYsBkR
erp7ZEhV2C0QML91bbARbYVLH36J+gaJWxJ6q+8vH/XuABU2iPjA5zRTEAkqKeBQPZ/iT/tea/B1
po7fWCVN5iKYeuQH7d/bV87vjhQ/w7wuNod1SB3SKbLTEP9JOW5GosLD60wtkUjBoV53mHSLEGsF
2OZWSEIYPj34lQncuB88gcWQCmTscgkYqXqNfUUoN+T/Lce4imOOuoKrWUbqvEc/b6JAjz/siwtY
FlqJtnduZXhU8zhqbsfaXFCp0jE3NAmEw2swAZ6o6quVdQgIo1U6vqbHzDKgLR+yjQ8cb/YIo30u
3UbH6Snc50R39+icCC4tRphT6FEFvDxoSRSCnAx9ZhDZNry5Sv+v+50xswbS5TtmJi5fhLSW87Ag
LwiuFnLE3Je5icSWioRBV8yw0j/NHN0g9zQ9Y7FK/Vjr2KAza1cd8lkeuCEwYaCRh+ANCwKSH+4w
MK0It6Pgl2nHXabJnrFCYf9XXzLh8RrUK4D7PnmcQEd0+Ysate3d3cl3ZdObHW1YPdAY243sDm24
S/ZHkhy8TMxwBZsYrCj2QRpJmxu+jZcI99aKGh7rmcbJxcgaX4DO+CcIH7rhRsUhMPQiutiP0vFH
0aZ18HfojZUd0L2yc5XMeewt1hr/wfwG68n2GwWC9PKY/Fho7e5jvZUl/+Hb5VPM1961fyjbjZqY
8CT6uuHSaThsmL0soKiDklEUbR8VxG+Wis9OSB4g2lRXCjhd24GwfP4ASv5bwwZGdUki+uxKineg
kY2T0W4VnMyxUrV2x+lS/zczSmT5jK+wabLXXoyUspyxgzPYANOvyecINhKWhcELUuzH8I7+bnOn
FrB9GNVJA36I8wW7xXLEKcx8m4EQcNfewy34n7JFVPqxIleZqh5P/1zlQ8LY7AdQUj9X1S2c8Tj3
zycieVTi1uy013IIbsHaXbGrM1FNyzADopF/LMquLvLeriV5CUKTDqx3V8jD83of2z6HApa8KJsx
AQsxz9wfA81ttRqJcd+2aIcvmlsW5nVXUCTgQfeTgFa3t+Q3h05JN1xTD/6kxT9buIlht1M181v0
MD2MDEWh1HKxN5T7Qws1gaFvksyxfg9iLXJbS1I2LJEEGto7W346hKfhx3CjrxMfDcn6P2H3/3a2
y9r+i8ibEqkJb3qPO73ru+gl6s3YGzln5/Cb9mRtp/xDylq10AND32psDc2gEKWLSwtlsnzu9AFO
is0okGlaAnyNwGDACEtHHrXpCMJElGvTXj040JeiLkIwKUT+/jIJUIln4jAiacXFdPZUo3mzmIc5
q0rGyD/L/Rix359kwoLWMUI9m3t3sGPDGqvT3jCmNT4MdDj70iApMMLtmk1lGSuXEQMFtnYX/13A
MxidepdXD3jPPNRhgIdMyLjAPWXJpjzgcAHVroMf3uVCwv0dOpWLaLD14l28iGCleWQlawe7ORRO
S2VL5G3+tWAY2prH/oVEkLSITbFGbsIvI2wvCVzTEJQ65SNU9l5bjwmA/aps5mSbQMpISb17rKNc
hmpn3vLlN/TTp4iL0iQtFc5Zo81okzHg+AVhEaDapwl2/AhZpG5Wc+u7vgkd/GL3mkPio/cTzTXj
kEdpJrjET6ckc3nLQiff05wYaqaIVgB7iJSCldM6m5bwDhIFRMjZ1Hbud4rPmWyoSdhzKGNZNgYV
tNLPHVZkLfrs5n+A15ZNDmpS5vcg4uFajhbUFfd+90+9qGP6uLo5V7KQXadcloL26dERZokCVlmg
FC3GZ+o1cHgEy0jK/YV3P+KZ7qyNV40BlaQVQbGAbrm/7sgzxxR6oLv7+EvvCcJdvTmyn2K9wXfo
HoLX2w46rmd/YyfNuL+/eUm1nbfc0kPewwFQwVWT558z+8bT4FhwF5ghabrHm5cxqThYYTdYe6t6
L1XjMTFTQwTwprxEYqgL8IBTZ/5sISreA8yIBwUmxSPeEcggOR3z7PafoIluQ36N0EQlRTi9NQfp
8tYRyXFzGGpfzkXzUhzh8rW5YarA/OLMbx6BIja+kSsnJt+gl7JZx6IsQ9xmCh5aR6PZNiUjpkE9
IuKUldyQpCLY78sudoqxcbDlMHieDzurdf4/62w4fRkyEavFxUyRof5pqG4PiInbDKxA+FQyNmWO
QXIa7bxwmluU5FFdnTDr8O0gZdKS0Rbyp1VkvcNf+gLH9xIFw1uGgmlMK89PqtV7MBciN06mY2E2
e5cuw0wm5+SDU9CNDTSuRAPC9d+grA/hMztO8HlHYPFflfivziw3nI85pJUBBQaq4eObH5+msvoT
Wo7WpMm5g5p821Qm0UU7KevXdI7JMQSZS5z0XNKfUen/EOgXXAH5/6TGG5GORrZqyMzm+Ag69E0T
VX/inn4wYPdhLOO3RL7LCCc5BCTAzhbTgEM5K9grLwgce/MZ2wpKt5GdezjIzjSZrcv7GTWM7gGh
1TfkteHN+HdxRJqXU4Q3kDs06yKZ+1y+R6aUnMEFkY/xO3TLCXiDnYhTZLmE37J8JIMdC6nYCD3n
qyUICdQsCbjh2678f8dFPzH18bL8F83pUhfkSWwFCGXFUP2/hX+wMiXyCxB14Tnnutmqipk1xuMj
QtNzeN3On+h5zD54UaC91u+SuEYCFZux5f0ew6iBw5LLbVANEtJlQ/36fW/d7wd1VWxFFxKuQGEQ
gKDPljed8ISh+ElhtZdgvpU/UahlLQ/rf9r/pMvUxJXEo8OQGrlRfCoRTf13/hT54tZy6oEyBzgC
45ODGI3jpApEJWZB7AIwSZBA8W9q6jmOZAQr/oxopEzo+5kzb2FRVRlrXPZ39irZADXXbSHI901C
2Pi6R4MHwxT9MzYp4JB6r3+QxM7bSA/CDm1+mq7p5ISEQKRimUHzZZ/R9q0KBYbyGiIhFvgwTbB0
m99J/HUwL4qAGjV3SxO5jAhgMe8eCL9wjZMHy87wLuBdoNH6t3Y1nxe45hGiJjyWWec19dFQNizZ
nLlx4eNxOZgYDpgyoVG6lfbaUJkGL70IiBVyxB2Hn7Nb9jCQmyLq9429DfE6B4ZEmbw0sZU03zvo
S3LUcJ02vS0xzyKa0KAVBZAFuzlBKdYCEQA2kUgcUSlBhrm+gGeFIyu2b3aGGvIiWlQl7keyFO68
Tg/FStrQ6TMwh+QZePSgpr5qTccw1AN92Oa9o9sbp2AAt5hxWsUQbpjyVQC9qdKq/8hAXMSv0jlt
L1VZZfp+/J9PSD70AGRYMKbBG2NvPtISEQ5ewoXNY7i7XJrQ6gh/c9hd1ghwDL1xQikcifpLgU52
g93E9YSSu93Fuo85oyMxg3PH33lPuW4TBmQ45WogNPkawvq56mm0KNMkOjB56jcEKOoB36YC5Llt
j0GkU+5CbA8Aua5Pw/OmbhOcxZeKmBd4iRtGKgfmirKiZPjsHDsdOtYXxZvhJmzdB5W4WPSgUhwD
7In7ueffzW3gpv+XvVeO/F7fNDq7ggXbaRbCMhASxSyfcJCLr3tdq0HzL436QAzonG50xlCvUS3K
z6vXSLQbkso2+dagcyB5dBqHyhcNYVZULxirf9XEJK/4+azcfDohZiIP3EkucZ95e7H6Xf+7CWQ6
IgiTkFTmqJTOulvXL/GGqlLrscoudASyUgeHmhVndEH20pfzY77vFReOHBDuPHUL/lT9B+MOUeUY
SgTqsRvQgei7xuiKwUyPQtWSc8+tr5bR8ihgRYcUx7iDe6YD5agkn80T0+LA0VsUEc+PhRL76oJg
oNk2oPXJnxDiKBe5IuG+SCbDW+mdXAI6mY2bOsVsRQMlNowN0QWPAO9aLMg/Ntf/W2WhFM6Uy0zE
4yy/l8eQXTtZzQ3KBXlyC2YFPS67mUSc1UmS6bc9Az6tfwuhyf+sShfRY9NpnQxOnnHq5Azy193t
l+6YvKlv1wLDu9ytPBw9cB+j2dKktFO+U90DM2ZNptEf6rXHXNXVlzBwWedE98J71bwTZ+tIJHxA
zkBV7ujrEQlA6mQPNthLV1DoSPjp1ydOpL4ubxnjZyGiCexAXraj6i/ke8KnPpBDMaKmcINE78KA
MYorDpWZGdrJ1O1QwtmA7HCjNUUzr2/9z/etqisb9pvygP8xQP9DxgKefx9sm/3LE6Dzn0V+dtnx
4KNbclFrwVRKGsaDv2DXonVwmf2Lb8hI36PkEByranRIDLRpj2chpGZ2vaev++HlTV8BhtTdWWgs
3ARZ1GddIyx5kP4Lcq/xPD81Z3xtaEP2Onj/rdhuDXWp0YOD6HdmVSURWl/CyXvDMf+L0rvokuZC
+7wDhJwhxX7EbnAUrZzCyw4NjsBbpqxJMc4ZVpergbignyBjicDkTHQ2rPa2/1VU6kJKs0Zpfngo
ayJ3UvIPS9+Qew/Fn02be+8/Xd2JCOl26MoqvbX2E+li5tCJu/T+nMhxDbtRYPbjGxtcKRH/wHyd
3oUHZxbhB6nEQ9zh2Y6padL53819RJmbEzUMk92VDHpAmU66ASDg0jIW0Ih+GOGs/9z1IBJPArqG
atVmdYlre5e2PYNFu3vyW5XJU+1qp53tCep4dZq2yeehKSyH+tIZwh6fQLmpkksCYb6C/jFBR8zt
pE0e/Jb/uUJ7kJgJwaAEUw1XHfRBDjDMnCDJC47pq1q1dehzQpGB64flcJP0MHzbaPsF0hpPtWEj
Kq1P+HUfGrLz0QQcNhdv/57EWpeCLZYhmihzl3HFn4BzXyMag5Xsf2lRiUZl0o2K9ribs4XoGD+W
8h1Bo8jyi2p9F+1cEUJKU4BHVhnCPygnLnNuVfQGR9pAcSpdlfRtgucpR1Tn/B4p9qYnpSG/Fyhv
1f3yDIUZrDmqTm2vWr25rnZ9fVJLvm7y13R55Ny6lsgE1vEQfTrvEm5Qp/H2JeDtgBLFLC5hOt80
D6hXMBYAuDfXyiXEqK4ev2ZLsN5jHwNmQpKjP/GYKQ3H7GEC8qZys5R7r8IPSJ//WugLL3siCv33
3GZ77PgDng2BryHeVo6NWgFsh8cYi14nbJF1VrysALuwHjjlBY04812xkL7jPMFIGfNIlZeEs0ok
+VBTl2pqqmIl0Y7J2ENq1n5zQwheLDUxVVnmvQXU6SX5wUUMUWUNuKf8pL6jn5hT0VHacVdsJJIw
wQgf35Vlu+CRiLxaYs+xCeBRpf39nqDQOiz7jA7zpQXPj+xNosyGXpEpfB4U0x2xccbXXZ/6MZJc
p5jqXssZ2Llx/tZGo9P1Yj4Bs8nfW0SysXZ77pqiI71Il2gJ7JbqpAydNzuSbrHcrAy/1mb1Hpgx
svbd+l7w1aiueoQNeg/XBvYTHdX1gnNIUNoAulCyf9qRk0ZX5f6MhvNgZa9EXVJ+uevVkkkxwMOk
Kl7AqREO0sNp4yw0ZBV6nFzPDwJ1kbWAS6KuPRAWB/oOiouW5z+WGBjxTrrqBYdxAkbtZnhGhGvA
bXcdFij8Glpj2ZvmItkiGttVLB/xNqRsCJmprTPDYcqkWN/LV8fxRBDHABrkQXCCV+6vlNuhQNEh
/V7BxM3p2BwHTARoXVIMFrjCL9DEdL+7mePxjKaDwEZbW09HRZjep3SOhXgUooVkXDpv0u+Lbhpn
hbJ7aQmV9J6xrJ71Re/c13oaosbZUKfprx4mE234aRPN7Xpi6a8fGoe9m8X+BQ0VdCSl9kmGiuMW
VgUQLgmrqX/cJ9/ZXfxCYFC4WbpIyxVNNx605XdbbBbThGgPqrPsITFRjHjtrMQe8vmuKYlNlm8t
BdJEAB3EwSCZUXokcISYJW2bxQ1rPT/ybXl3/RGYM++kOxW0+vuL9AITJJjJnI9z/RGKqNO7Unqv
13nFbSi+jOh6ruuFX9cd9jWFd0hNkWhU2fcTP2BROtp9OtGwrNVocHolBSSGRZi/0itpt/4MPboF
8uc4Ro0tFZHti6L1px2M+YDxiVnl0SCn2B8NAWpgAdcsw43xlbdu+AS0lUiJSpcYmZAIcmikluOs
J7VlQ8D36hpin8AYtWVNp76MAbX+gbs+Jxb/NpgGx31LVglU1RGs6FJs+zsX6V8NyMFntvnDFnuW
UcpQUrHT5bKHVbbgrLiBtodM1QErrsCzPgP4xYVJJO5RwMnPkh5zvcXH5HPVoyOuaqs/AppdRose
7chBj2BxkDxo7jWZ0ZEO4+kTpT/8QTA5WooxOHTpV9Qeap+A921gfUy9XlLzTlYNMcDRgAHpkYHO
kmTDEdsrQ59o6703ZzJPv9OcDcy+n5kSgeS8IqiF+5DcPGbhTXFCH2E8yJGb0Cz3AIA2c5XUytBV
lfkzRm3iuEkdtUe8apXlqgGcD+cZTIA1e9tRLgeb7llUAtKBAQiJ5nyIvnvKcX7xYHDdugAzPINa
Gb+w4g9C0BupSriJWwwYcvk7PjH78Mht9zCbxG5tUPri6+kJ/U5vE1Jw+p9cMgqbRr2y/7xulps0
FlX1ThsbXpvEBcmGdldGXOxU5hKPCSCxXkeP3ZYFjo6NJQ4PgqO2fdnK9HoYv0tr64tMTQDrWROu
DekBKPHctr+PUQS4mCxUL8CZVEpweDht6Bz80kBazASnSitQ2cFfe22Gs1daGRseuL+Ozehen4Up
HPmSPSsCuhZtmOkZuBW2MKxbwSocAhkO7cCMgWJjOQS6XCSFZONJkpFOllslDD5wjG6szBRwRt/m
j9RKYQ/f2dWLDhocwo62I0/cXjULcJRqNqDUK3E+tAzkbOc3OGRJlLOZ0cay9TiuxBRRQjMytFkk
bWxzc/PamGEBB2V2bAAfmYqFGlKRNXqGeb8gK2fSYPEmKI4CcfodqN5JvuZzIgAyiRHlqUkBHzXy
L4sKMW131M787/ZyjgC44dFDbhFFeiNLTTG2dkFMx1YwUQY0MGlLFpQfDKsq0tsN95Q0TexX3LOn
CZtKY/t1Vzoi8YgjsSRXndY7AlZEaanVBcmrYv3YmwY4TVdoojy8VyoKvjBXFsEwzDt+8QDtc8hh
Bj4mNBic4VNbufjvZtzoboon6GP6IVOXj2GRoMGUUu6EifGPJPfbmdH3nbRBCJye9KRLDqr4YN/Z
GxnEiWiPfDRZUgl1HroGmjN57fX6kAg9yu70xhS2DipUFQUTzFZYuEMFEOC8TGuxV8zfy7Zd/F3n
yequ1Z8XgAKUZR5GiL+2Bf6m1KsNn2FxMeVg1yKeD3lrv7PXKybFLgJnMarSe1ZpkmAAM+XMfZ9m
TVPP6xuuMxT08Zvjbl0DYfCjYYdK9OPaVU99dVm/MRvxbAFBiPeM2SfizMI3+jnyjgxEp7C+QepS
k0RUMDzQVIsZygGoEO0OrKdTDE8hXmdchbOqlXSe7HBacLRHejNZW6jYAAQbTItyononBDkT7lhI
hPeFfReF0vCncddPetyMZpxjmQzaBT3kFkUTyNnLAxRBwHG/YWoJzzIzpbnVqyGnMXJdIFJw85h/
DQKn1D46rju/ViPHDLhtJ3OVhL7rB7zlFab02Cv+ahpvGEO7RPD2Edy9PmPNHdHlguvLX+Zy9HBq
AwIkyHi8FL+GEbhxWFw9k7OUwaVIZ2Ep2xo6imuddzBpvydsB32cS14XlyyFH5craoxaCEEjwkQC
bTXTbGwGzBXnjz8WxC8dg8m+SaUnAvnERNt2A5OqHs4aFJHqUUhn3PeqmxbLUleZQXrWd5Z0fBrr
idRvKh2xXmi4dRq9PdwpnVtJtz09j4TYBFakv3CRmuLWrmbLkn2Od3EhLbWSR0rBKhLpL3vSc52f
V2ONiCkmT4r49k0Sx7m51mxIBvaEBGtZz5zFvXNPPEoxz957/n0V2MGwwD1k0cO262MYdvDIkkTk
Byh3r4LvY4CkT/GNu5KhmGXgottxwQOhdmXHlLQg609N7rBgDi+LzGslM/UUTq2+p2jiV5yrFnmb
vhGoC45PnPNatU1tr6JSdmwurcnoaIIH5dMuE2VserNuqDjpDadjP45d/KNg9iRgjCdnrz54Ptva
jOAfVAwLN3xOO9zOsZM3ErCmIBbtvtEpuRqBMV/y8lCPIcDhlvvoKLhymekJCa7NHJYG1+/Xo9FA
SoR1CcCzCdCbwFhenMGGSqzOSSsHdQ8eGdiPHPuiIEnrI8XqrsTrFKZBpPucVPUy0zLcRDbUWQRb
UuZbZbIx67fka2z+N7BGaep4y5J4vngmi6qZx2MuqdUcCIMVA4upm1xjkqjQpAcoNPnN+LCc4Fqm
OZzF3AeSW99rLc080FKGYDEvEiMxKhFkAJTQZa14u3kgidP1NT5d2h1GfvWxqsO9WGWl8stfVq1/
CRC0AwMpwjI64wsVfQ8bAaKLgKmjUWemqGC+aqkzx35kNLT8Yr3fIM1eceXv5Mgd/rH/Fjj+j2QI
MLWVXnt1iuPl38aY9z1e7UdGg6uBUATKZRoJoriMVnXGyaPuqzpCVdMd+KqsnHZIdYQL+d46PlF2
24etHa17GkawKY+cB/2e6mK2q9GGsVAuSxFq6K7s5uYTKD7ermcXlI6eadxzcLEo6kf85hTzDHMS
Faa1+G3lv+ZalpB+Wwh0EoHV7FJOllrP+b3Ve/HenPaY44Leg7nOuVCqPL1Hz6Co+sZyJcNuWHsT
rDjEfuMdF32+l/9lyefiO3I3mAu035cLfhJkW3ceuSMqPHD6rE8b2AGquCbVrUASZivVCV1FvRb9
LAhIM91VsTtDM/zbkr59/BB60FI0fe8t5wm0uc+HPuf8x3+Bw/YVPi+NueBsdjqdVk/NFWMW6Uwf
zlk6FHzsHr1YOEo5TXGgQ07aNfgH6XbSEFELjLfV06RSN0Xp4f8PoWd9sXolg0/o48+4R29YDVg8
x8SV/LHFr5SL4LT2Y6qA9d5Wy7ZkzwU4I9I4CTrO5bHidjv+Ek2BqeFp3wkoWJ45BTIp0FsJymHO
we4RS/TB34HO41s4iaflSJ8jkpSVpb5r1AUViO3/5SZVMKnRPJWZMFha8f8L2DnN2uzoRhh+d/Iq
GA1VbVcbo6vIdKE9VjhfxbXLfyaMicD1a5asfgH1BAKOJRVFyZ2opb9Sz0smy0xUneK3LKQ+bxjo
3Bg4TuGrRqGXoYiF+rscW0XcDo2AiZbOhO7c5YsNvszjlVVvpH76R1ODk4z4phExuP17kBm4Ncem
3s3YfVH2hqwpuGSEmfHdxMlT1WssN4wcDshDfIhQCJg42wGegW+Ozj0lV9zKken5C+ZigyOocgYF
YBjCAByJC3af2cZrAQqe5dsnRckdpIyuu/EfxO0j03vF/zxJljFmqvRFkLg2WvKYPxu1mr1gixZc
Fo1NPyXX2/XljW8owxTYyhxHavLxoSPHqCDdHNxQaJmRQ5Duo2VdNRSp3WAkRO4Hl317yJs1gQAq
IrhmgWlcO8OXYOMwdTiLdmsbzxTkQ/1MWU6GgkBGYa9BTmeKehvoErBHuEPo4UATpe7u/w8F4Sq2
a7mcuU7dQxEVwengpb+n8TuzU13bco8PaqMP/1jZe8VCo65GcTAskleg5mPyBUw3ByMMfDdTxOBs
Z0bi3JfoV7oyUmcGibJ877rPrBpTEOM/yqBG23s60k+YS0H1qGEsFZ+lcB6Tb0L0No2OZ87aj6rx
pE5KPoutSPWQoWtevZPJcI619lspITAB9iFTPvUXZrM+XsFWG1lPRmJGx23/OiYLmSDyj9LOzdKD
U0XBfihzm39BtSpCvw6LlQXewgXhKzI2e41Sfx3GlqQFFMh1Vbl3q8ZDtpg1SRy1DMig17oavgon
hjOL0X1aTkqnpsJFC+Xr4KT4YgHkg2D3ldBNXYk1hkoYFCYZrimpG1c3PQ3q59AMNNk993fJjdGe
1swpaXRQbsVBQyFHuy5IL7g1h2nlz7Il5xxJfRM0b9oj0kiKOPMkeykkzEtIXjYiu5mTI69Is6/G
l0Y7RLvLaqTCo25M2WrjYiy6PIzbITXftfW8Js9BIMWxPG/yaJtAjSRzeOt9lBvBCeMDwwbkuxRk
TM/Y0ZnjrEoyZNGVtNq9gKzujXWQq7CcOkI96/PMBXPgRcQnDGE3f50eRhMjTvjGNPEik+q3y1Fx
zvzBP+kya9WrAVsk9zUMebv860fVLqHs7DpJiPQC5tpppYWdLZKyTiMSuw1VPFCGwuRozlYFdLjz
2fiWbDIauyt4PBdl4j65+kn7049k/WKBMh9brhQo2nuCjjr8ZpDMRIzwQN0W5OeXNUthAqWMzZM5
juyDk2IGhx+owdiz28My/96THSOAMUEmhw6je47klBWBbJw5dpO+0+Ix4G9xDXivryYtuG9E/pbv
Lx6KmQRVUB4l223AKG8lhb/Z41xb/ejlAp1SCJ0s7BiavvnKqfalBY3qMuCwWtKPGScIcCcV25On
mMGMNgILCxqmjCKBqPIDPLY5lMknFEcvYrn1xIhL/yDTcN7kuRASV4vficb5ewq9DfDQBeW2HkOn
eyrE5ud6ZKN6bulk0APDpVsSOM9+w4aKjUbCnDNyAHetFWaSh45HwOlLX85wPX8UKH22St751JLF
8/VbCI8+aaAd8syiYBv9B4VmkPQV3s2yREqR4OkNdlULqkTOqwL78ZI7/K2QBoECbKThkwHv2mPE
bB6BbmBk2lC2DJN2gdXizIjcOexA1EkvjRJcYEAoaig6DzhKH9COwZuTAq6v3wtX/IhbywZuyLT8
YeqxWf1bZadqwmxff1sCh/WYbFQSe4EP/C2rLWc4Yh0n4qxJzKgOunRUwafBrlMRA0QOFKa8FAmd
VULybB7rnEjPPtHWOJX8ldNzzyEsfQorxBLxWlUrAgVRmhXdUTGMuZEoY4AuI5q8TQelKymJh+/v
Ni4kN1vUBSKPAEhIIBY1jKxpKlBa0qxBHByh6brhnT6wHSmOb93y55DuWBZ7U/05t1MKdu/L93IU
7vVQUmZ+SzGk7Dh8MhOKmZA+lZjW0cLdi4oZlTheJZgeyZu05Q5r7iwtszzRxY/+STUbktlEjVlu
Vr7SBQqkYNCoCcB7g5LEW3grSJA4ek7NW+811yYSTx+LpCksXrgIrJUTu0xhK5QntWGwT69Pf9Sx
QPneWp3W88Qmp0dvtaD2iwlZTKDfCmUYMOw/g2b7AKfw3YnEVPisdle9za47x9PeYt/wBQ0baVYD
Qtn/M6+5Rnwr2delYbhTOeFPzFkJIHguBUx0ZZeG1WlzFv5Lyk+shdNFLAx0lMV/rm+gFBSA8uYM
LEo6Be/5LmeyRsh6gJopfcbLIHYSq4nZkLXBvZu8pjCn/inJAszeQuT/FeMpKQsaybr4HVwVxUBn
BCOifUhzQ9BYTiS1iAa5N+VcSlsiHHyDFlKME5J911Lj/YtYjvTW6Tl0jw0RabKVfF7aRRv7ii8C
bnULeFxfKAI8jWmWO9UGjsEngi5G/Nh+KAfqeyGylHSqIeMMHvjgkdoTsHj0Nw5A2d1Jb6MOZZaN
T5obxKyJQQR/RgH/MbG7uFQeI4QpvLtW060vnkmjnZOmwS8s7uFEz98suh6wdl5fMvNT09gfVcrr
AWaZgqq2jdX9dAyJ6jFKpwavGtPInK3+CVF4HUDUogpjcv9UEMS9nOlJ0NXfIXecOnEjxcusjHNf
QOwqxbhp9rQrI9F9wBaEPtiXRUt1bsxq+uan3vImivspvGmQjIrTv81bCfAlQf5HJRFPFGYw5cIQ
FqYP5SPhDyt1uHVItzLM/H46l3XaApK+aCTGmtSMfo0PLt8jryeZTGWlHeNVaLLZD1RkPlTHCebA
X6cJ6PYtPoBXlC0ZouN6gnyv/r3kWArORfUqoLYfjqJq7WkPSybo9JNPSf/ee1rbHOPfccKIjUHQ
JRsx4+hzrAf/7xY4P9YOFQvMeqqQZMhJyT8an6pp+P/WbOGyAL5wijYA5w8BtrTGauPdBCAWx9tA
tkjvoSjn8K04mocNRXSL2GYh5qcOiHFFmqTnIbnpRfECT3yGeAMpCAm8DiaYbKLpW1zMu9b9dG9v
eJWJ8hEXgnTHKnAZtiqc1lrB0vWZCHWotHQKDkLEPHdCQG+crh9v+0Ik7p336cJEFIWo1MmjQkc3
BqGx6OAGileHWT2D0y2vL8zJAbAvpsveHIeDNxR7WOpR1JFWOuwSlMqGDX6QL2lAR3FzeoJarqlG
ciaSJ2kvhQjaz68VvXpohG1Vv+jKB+TutNR0QXxVovsFAzwH3ifxweMMb4AcogpjLsuPE2FS2oF7
VpsU0Lwz2fYTrLRFw8ioPnpHlh39vQJaWy/SgE+UCo3Gi2UjTJFIgQadVN1v+42fgAQEFDUJ7BSE
ETLRtQbhdrUipYjuTvO2XKU+ESsO+NpME2kVq+ZFzaH4Rm+f8tpTYuCNkvdzmVeMzH+/xYwoKb61
ToDC+wqN7qPVEsaKSJr1AbZL3oY3G/AWuuJlIg3lXftmPpu/FEnMYoUR9jlzqgvZuArBNEctVF7T
tyywORWp+8zJQZUi42Z3ScNTRgXIe4HCmJHYT+19W85SuDvzwgAJCvA2JOy7ds3kDViI2M5ZQY8S
HctCCVBPMAJ9pT0z4b/RumxuiBUp/HsQco9GVn6Tp1cdYSGcCTDJFzzFahYr95jcTW9J3I2FRPyi
pVVwLCXBtm+xxUYswDtbviUaBOSWuNaS2jfz2XlMKvM2Iud/fTTeFPM6bbgW2kbCU1Gcxe3UnHs6
kSgxfBCy1LQpk61U/5Fkc5GTB/+RjP50rlH/vGAyzSmq0XRyteg8lBPNRNYxQdW72N6YuyDD+9oz
yprykXzdkhT3ZCaa9Sr3LqFG8WiPyiRPcqHfGGi11ms5IDSXZeUUONsZ1Dvp3O8Oen+he3h7GSjT
IyRin09ms75WhBlBq8WttYehUtW8tDo7VtMTmnBl0jxpnPPSBru/jrr2nbWjfIAlJZEMfuDaKUT9
6oJOWINGQJPdjcwUBO23a4Omf7BeYkieZ5Bp69nanS8wYmp6TNImLvbiLR5hMXb7QOLiQ9zeQ0Y6
+HHE/ZbpQQ4N0w8WLYopBvATWQj7ya3yEeNH3XNz/9cAOa8RCMWhP4xTJ7x2keITdyQEvHFTqwW4
W2yBkKbD52sXHkrLkgI9YK51lyUWTnhSYQwOYL1UA//c/puNbUStSsjAS6VBuj1oanvRYRtkEb2W
mWUkIDSZ6a3DC/KV02EDYfYZnhq+dvo4dyDrx6REB+EPna/j49GgCT4YHvELF0bflywzOlT9STpH
NJVFZCtKynQdxh67ofceIbnq8m/xRQXKrk2jmHIeje1muQA5aWKMICqD/c4bQV3Nyv/nkGJINHe/
+QWAD2zYPORouPVP0a0OO2fA+PI0p14oYcC5F0mc361uGi0ryNsw73iEMSrJyd41ASZJYgLirnlI
TmipWYB/yLQmOL7z4GI7nji4Oed2tvDoKl7hRvxeAyR18o8axNQ+VFVQ/eJrUE5VmNRr+rl1NRv/
89wj6s5DzBJh83dGzZA7kJHd4s0g6CCG0vZbuNjtsNKQ6vpSMdBTr53qq/hycceik1qZrZ8Qyt/C
23+lukygEeCBKedmpp5C7/oOfIjV0cVx0Ck59Yi4LOi9MvAtTLY77QULV36kCwq1WakB0f2zKU0u
7Hx+7NFd1yQ44b22LLuR0OL0WiFKDFEaQARyecm/1qAtrcXVgEyp+oDJ+fx4YwvUPNK0rWZzBXgc
NtUFJiwW3zP/v6Xg+4Wp2vrHb6TzaNBTVxz2UZ1PYU7/1Ptdh9SgS5GQE2r7mL5uYv9K17LJTPg0
7LCdv0A3d11AKVfJZY2vbmj9h3G3n1lFoRSrGsA13+yKHO3aKzmVMgOBF5xLIfsqwLbo8JJIx52p
Czblut5cmBKes4dfeB0OI0iFsHeiKVUtK+U+UMIF96knouKnvzRELawrkkXNUigwJHtm0FQRNnQ9
G7bFEVdyZYqZVXOQ1mti750tNd4rLwVfDaLJ0x9yobuIUJIgUHid8LRXgon+ljRN+nXa697mwC2r
f1+/ip7AanBjucbr++j64C4V5u6cJK7DZ1DHS39bqW/ZuA3DD6xReO/b+Urb/URBY/UaIo2iGSd1
HG2PypNZW6J4rKrzVemBVzJUsBHmQwda4UJ4+mffiUINLi99RDcLRqj19QhexgxX6muYu71OTdH9
RAwKZQMqUVwGOUmVvVIbho6tKrqV3t+6LDu1WrP7Tt7kGQdjsD+7SBFBK62pv3ymf9K8oSCqjS6l
Qkpp0nz4PVmK1AW98XnEYU4mm6MWo76UFQ4LDNVw3IqKpTRwCknI3l6OfwooIwrOOitoaRWY9nKm
/WG5XOrh84BlUogBiOOT9S1fftPDTDB7fxg+MFmRMQOKfWr4NCJdkHMEVt09g0HAcSFObnsbHZDG
x5temjP3Boi5o6jg1CCQfJZzxQN4mTncNJA/zlJd6ZLicbzAbxZXDkDzZJl5uO04RDI3rFuMcNRe
AWJKXq71qr/McI0FaW6l30awrrxMxJ2q2Pcay4OB0uxEPMQqEiHnhtDooaCEpOE6zt9wZ7H67Bql
TNvCn8pwF9T5oHp/uWTv4lBqMfSEhNTHa1swIdAilS6hORfC0SvIoO2OTd1zifzggYtJyZ8jGOHk
X/+ww3/KVKDCjwHMOWJTR+JDZNWXkrJAa/kyMvygqcrQJVCKtz3AjDMk1khv2hWiOKNU5WPp5Htt
Ob478wQBgNogjlMa9MEcB08QVdG7Ih3GFRkkBdTtRXNJvQDbM7Uvlk8ayZ48HowXUvZtOe6wVXC/
OOHv0HM6wJNKBeDJskT00hZUGwQIKTiB59KWHIHJYnDYXtEcoATWEjC50Kr8sBsVHb5HslBXw1fy
ky81FH6T3bayrgfCf6qGSYtKkOXQ616z0HbN3nK5Lfl+TVXc51U+Ckyb1HFXZRRveaARTdIU28JM
Qvx5TARQbnygZZyLTQOctbsHq3OAt9ptQLLFro9T9uwWGfDWwQnVGKnuugxyrQQmuRJqpMDTu5HM
Zn3jH/n5YIGzbJZVS+FoEBZTl4QvUVObqqZRk5qpi3UW7gjvx3SJF6tdYsjPiHLRifkSSsbeHmH0
TLmmOWqag7KPetG5KpeG7fTSTFQ0N5S7nhdbGyOcmXRcMDpd/ZPepYEdOIYE5YJSf01FVAsOVuDC
JQ8o6dVuSrqHPWNaAsrUEJtexPIAYVAFsOFoFA48hTYl32FU11jcEyQH4lMrwuPseJaOkALzUtTV
5gIVIxCtdpa2hE5T4ldh+Yk4XXwRG/vxgXEdWPDnGTSsZVgB+7qwvypsNQzhHz6Bc5qnLjbn+kO0
0r8meFC1r2+q0c/PXudV6NpPXXu2ZkS6NflbePZvejdtv5RduJ3TngyzdMSF/U1wr3P8NIDmCFeq
TGi+Fu9f5tAyZvcioT4ju05HIO76DxGcNsanK9FZqlPKPaqj6zC/CHyAI1OZI6H+UjcSJ+JIFBgy
gec8LI6CMC/qw3lpwTXFgeNf8Mz7lgdmCkkKYA8578XrWmnbeXVK4Lx6mwoTJfapxTcyQulc68RJ
yxjBPkoAozYKB3e/C1ofkqerQp8f6j6BQbQPubv0iH4andPWSHq8W5G4Fo6ZvIPYAEIPUCMBZQbP
Yo/UuRp+0PRQNOxdgzEq20MxoogBYJ5rDb5cvq84h2f6siFw2YJ/tcYcEhJdnDpOwklYiKvoO9x4
K2p6OAtKPMRU712Qf8sZ8g9sBYynqZ/hJBLpLdKsdZUmZMbBQPcCK2qGBJql48u0SO0G1M+z0ukk
Wcev6T9ZveM+xDnrE4+dsClafwtiXPeYkjzGJOIUy5jCvLEB6lqx1TzrYcSO8T2t2aL2Ndzb8jxB
VfWHncnv6v5O4lM1b9jkPnPeoX6HOnxv3Ss1SL1MeDW2AhW1M1xtkNK1fv0Oe+O0WWhZmyP0n69l
z4idF3PAJKP5iW42NbCVNY2/e4bpuTxLecn4kcHuNhY6JYKxmoIQIGAzMJ0/rbgcyOA2TOg3O8wY
Ug03BuWnI+kwUg/1DzY7LYEMjNGKNSD4XG3Ud48hKp68cGjXRcQIqU5tymMDS/I+V8vBWw2XK90N
+XgoAewtVw0wyyYC+icFurrjaHqGy+8HFHrv1t8ReYl4Gkp5iL9yVtNIRTUL2q1fazdcxUtRc3L4
KH34kZWrVpbKCzbCQxpCQwj0bcotEyip7xaacGc76Llm/8Ajve65ia+J3zq9uCRY/N0213tawO7D
shmp28NcfAjqTy93JsLc5Qhm/C+4G6rSWe4I83RTQnVrYqhF/97bulS0utwBrfYsgI2doX9NC4tN
/IAYpv0+xzN3d/VGTg8+C7mZtvzOqem5GhyTZy5Aw9AYnQwtaK1fYFHQekFZjW3iDfrWojkv2vIp
i1gLjL2QM7auVoKXh17eMtAudSP1TdGiLqMrE3Tcyzst1qLTm9qGFlHiALL+4zEysbYDpOOs5o7w
lVfRsy0vDPKW6YLJHHLywIYNqMZoHXInEmCBqBBmxzaHQRRaWy54OoGRcKXIyB22lmQbB2No/bat
J5XRmh1/yj/N6qh+9RkUiv1LDn5gbSw2p5x/dGEIoyR9XdfdsWrE6GCNDeHDTpOEgzm4HZb96kjT
zGXLb37l6gpL/DI+5dz1aFBoFUrzCC+3HykNgB1fT3SlWfZLJAFNaBGnPa+AZwIw2M4pZxs8JhBN
zgGgS4rVycDJXBx+NuegMeMx1XOUsTPXMcJT1NzSE/Nuy2VB40mksgOoCPRyGSk78V4kS3ldFOmy
LvSN5lbgSC2vBdg5M2qDYTGl+0BS5rQFq3nUPOtl6HHs2eA24mJX53GAjMxXsgE5vv7ZhXmEFl1W
aPCtaAuecbkvZRFcMThufyony3D5GZKGWNRWEWpwkME0+81/178gUPu+DnPjnvAtA6jE62LGDHa5
Ks7dAcOH3a5b3YMUMZMU7RB2mZO2UDiCGbl04xJCFje+1Zfc++r0qEVNn17+LzmN2pfjk+eiH5f7
0/qdk6s6sR5KihD5E9+HDGgpJUNPIGDPZdXE53jPHNrm+vi1ZKBEWJo55PlhFD5/LTOTznQFkUlR
E5JAb35Bt+nKN1JsLhb1usdueKIaa4ndAFQnHkcEvKAGwhXMTvHYPRIBvT+X+UJXnuLg0CqLVWHQ
sVe5ZXkhcQiKN85g9z0XOaXpTC8D5qyRL+xcA6HXvh7NnpmnNXJglgujLxxTa+z5pgDyaJAge75N
0KNSbMEQHv7hd92+l6yPIDG8qbQ1RNRvP04C/n+4DiOIT1t+KvfLtYgj0258nJg8S03zzPNQkHzM
CgqTh/+zZEgA0xG3JUJNQobRmCoOF90Dmj3T87HLoigF3p5kfgm2vriPMZFUaGCS6om/ZxePw3O2
JmHfSSNR2HQiTq7OcSYobxcY1OCUDmYf38Do/n/b7IjzN54t+KgpFucmQ77ZozgqJcjlArtWfcqu
NSM22iSWZ752rPp8gyJDpSBNzX1A/jux5DsXhroo6cT3Y7H13/cWZcMN0DH2EHp78IXf3J8r59P8
L00syY1EGlYvRT+mxTj1S0H9qnUPmG3ogZxUH5u5X5xiZrUlTuPwMQNsqtbFQGa3BQiyZvaSeuX+
5MzU/S5PbqSO0nxcpGPzO05cNyPpC3eeNupymJWgdJNY8QqlhG+/Cikir05+qpO3+XvFDv9nPxSE
gN/UMbjIQyC1U8NsweNq1LOVDyzkGeDrvwg7jgsudkr6Geyj+Pr1pqmNf3CJDEp7fT9TT3WbNvBx
AZnKcYGNH0B5nrHi68AbTZhYg2SOjTIwb4eng6ojEHI23O/2PrUUsP5eFTBPdsLikjJcnbuUfOOC
hf1RyBi+AyfkLdVefVoKqLphtuKgsI74JGQSMtJyXywE7tdVJQ8hkr1xdX8ZZgpvz0V9TqB8aOy4
7EbcVR51e/OqQ65nJ2FEKX01CW/GFyxm9fPU6r6HXnH1psK6zRjl34DribNR3rfnbiYHv0Cu+uAN
AO8Onnn7C2CtrJyzvGxdhxNhdHMt8vNZTW7LXst9ONg4hWlxwIDTVaI+EZy5HHrMOhix8i/cTvpw
8ZJLegbMECvuK0xCjbt3AzL4uqIKn1akDJSA7KUKnqkSP23JwKoXAupWLbssZX9esZam+yg0Fa0f
SO5W9v9CyQbh6QtrVkjW7MIzgi2yVyXevXWOEj6rVAfU6A7CC2R1BF8hNyQzBFjQGeXlWdM1ot4A
+o6u03VMkkszA25SbH81QTOwiyPzsNJhPg5iEJejLCdz/JYQ5nq3HrAz00qSL9MWIkouAiQHCcNx
9KHKaBlGZxQ/FUztdOl1ZN6cVYZv1nb5BNZ+D0HOVNGU7oZqG5LPozKtp9B4ykTam5zfhfTTiorS
UH85B5U1QDfHfE6onjY2QnAZJIUbCIKgxtEh5OlXQwTUM0oYAgnzW6yNWWbDu4FTi4Napc9mcKTX
tm5edyTm85rWCUmJnhyhDLzEmE6wwVJCd6DJQUTIeIb9FYKcjBLTfkOfbZVrkZC7+2LZkTdNJFCL
JFKH09umrPNn90tWLilNQkqd20yO91bnnxGfwU2T9QMo2sPMDF2N1EvPPuw4dVVN8hxdmqiScxvO
MU7TZ/9tMwSZxRek4ynFSun2+agF7tNLieXjq+JwtqBhd8HyDNK6LycUQSbkroTk94ELNyGJMbuN
6Y2T3v2d0G2bVD82DQUoIseEYYiNKkF7ZFmJ37DA1EMgTMlCC5mDEDZ/t+bsAx7PzxdDwIdRdSLB
o8U8VoSmJXP8RsxuEKJMHGJON8hYj2hTCPt+mKJ88p3SNdaa1F/dW/f44QAijqeUzUuYQO4zisoB
/4q03VMaF8p6Y9mALkG2LszIBRVERPBffsG5oZckNNBxZrm1hVQ9VgM77NNYxq9iqDDTqXNEu8gA
Woym3Vcm/5B0lLfU2tvoDuw9CoWuwWr8xnsn/dieBA9Dc+xjziXR0c/z2SOhdulU3Onm0wcDwTSx
5v7f8PC/0Pjjf67g1yBnwwR0eTMWH7zIiljeTHJVkwZrU0y6kjXs+2EufCwf+59wSryvsSXc6FLQ
u7+EovfQCiXcEPS3qb16lKu4uPgpo4hAitD5DvrCB3xVfRkC5TVbVA0EKk9trSnaBuDBbiC4a0Sf
95elF+3sl2es0UXwibKgqO23GxeCdgIw+RjLDRELMRs2zprq4mMeCkWm/btdngOBF2Bc9YiTiYMJ
J0Gp4BJrGZPhQtm/ljN08jKkpYyJ+4kFeEOr03759hxZ+vGM/qsmWiAaxLDgIzd0A1pTC+ujBYi8
C/lNC9I9/H38+9PJ/OYScVUbmWahL5B2fUBV1gNdFCL0RRhu11HVZn+Ehy3dYljGy7TRnWWNkY32
Ilp1znMLGEEGKGfd8IIExGVeBybglI65/KV5PnDi7m3+QI59c5Pzv9FSLW02xVxCSLYQXSgK6Y3z
PfI0sYT4/WDOw94Qo7Aww6Lia+XeL3WyDOW6DQRvdDEfbIL1MNQISEelTWNDX+BsPDlBFx61+veF
vdUTt84wFWIpmP2gKID7WWJC5JMbR85F6ynzKzUwWmSB69JLeKKA424L8u3FMcQiWd9PfQ1pScu/
hDOGXvaNtxOauuPi+Ft/xxCxT1IuC5pdsLYuPc6gaUvKP/QCH3CLT40SVDIqVnWA12GJTA5tWfvz
C7ZASylex4eZxKFIgcUW+7owY+hXGuQTZey7oSwpBBlCZnPGTEh/OUzJW5QI0/oddyIbAnavd9gu
QiVBBSgmTktN6Jrqsl4mhgeslDYzYe+Khpkq6qqr/GPoouiBrhmNRCzGeg+Pc3ET2HM4rMEnaZb8
3YjjzqxM7+rmlZcsn8ykiaXSNfk9OiFshbBcFqQLZpMx8OCILQzqPoB2VxKIq0JXCZb7rmDqMxrp
2Pckmv92UgpwiKA1HifzGG4o8zOx3Ssn2neBlTcr7aJ5G6ehI++KDBnpShB8jt9YTFVtBn3igLb5
2VR2Y0hXsUp/HXphQo5+eH0/nkKN9a91gkHvlBnIy/KafSpy3SF4aObTvxSMg3Gvp/421xI1cELW
uYkPw90giuJRvS0Ei8OxApsdvo94k0tCUL2yMKULSFJU/2a7sNOZ40078srul/tP4FcEuFEHFXOV
SmAUnc/DM5p+ey1oZUgZEAzme75IOlbmZeV0qWAdRufeKqTtTfvmdyKz27VT9k7+/fOP4GWxVSJX
E9toTQVT8IEiT6WnoUwTlMmU8SXh6FyqtBdv3WH7lszTzUj5Bo28jZcjoOAPr/CQZbuESqnG2O2h
gsp2Ccby9kek6GvbbsRYSVqIbbO2WzDVb2rEnp8o0RuWX2jlSjP7moseVqvyCHxlhe6q9rItAooA
6UVGfOmQw2+aRc8zHIw0gdNcgSmyIqXmEIzJfqUOQohOyE2pkqLih+JHG/If2Ulip7ol4uQE98L/
DLix9FiV/Udr+RyOFfCenrAqELwm2Ma2VTpidvKvoaCP17e1ZFUL72OfQVIpP8OxBOl1Ujoicu9N
UMCysd/li4lE+lcKUewkV+bh9Td/74s62g/RPILjNQ11cd8Xm2ytyX4/JAjnVHe31DZLh6Jmt6jz
IgJv+G/RlUfHSDNHX/VwIVEoH2rKDsrj5GtZCJthrsmdDLNuvl74Ln/Q4Vi6qSHdh0kE+bfHtIm4
YYuqocF304+qCAG2NSxHzWvIRf4EWKswSvtADceOafXl2yrIaEsrPeanMOXmbXAmEk8uENQx/BhL
6gu3MWYlehFSmh7x+YPKPmYQUL0sAdFZ8vfmN2YJ2OMWUzqIgxNMdXKBI+mYJvy5xEhOgmqJhurh
j1hy+JAKIWfxCO7Iwte3fpmWlSFHHqacvHkfULnjgqT8xqynBAlmOCSnaLuowOsbFZtYjDbuNi0+
R63BQ7cIQKneKG6JO8DUjU3fOlAZteU/g2IKqfxN2gv/uB8URqL7vGOS50dXNmR+whsXdGIOeu3J
zqTwbCf9ooTcr8lxdsKicEUADUTqXgeRkoWL0675ODDPZejA4FsOrgi7H3HaeHGqSXIPp6qMP/Df
YuftJwlsXQGiUTBGj3pbibreqAlnoRdhlulH8Fiu85bhjSPo2eNxf+gguy2acKrefsHuqijjMk2I
Fo4XQ0bItmdIHGebIKk88ES1FkhfTYTy4K3N2D4gy5NIIz6Wa2Ng+ykRxsQBmrJRSsFoWkkzilf4
XYRfcI1wZA11SwfI/IPTzU+f06+tQUfCP9bT1ejWZ6ltGZiHSSfz9Wwe3lTlzeWbN2lmmRZlJg5h
lsAdpkSBq8YlZO35oTLUU0/bWMg5mLFRJpAxO8R82SmqCK3qMe6A/tgRFR4svcKZJuHS4evTFOVy
cIguSzyGxAZNBwcuGZpZOUcg0H+aGas8BsIqW2fTqf1A8CkP/hAepHYPAShUTzTYJ2re5MR3VGkV
sXRBujITcdXD6mbqzRW/1oUrt0RbBOSV95PE8zWP1itfG+TkiZoqaD6YBJbp/xi2o982WgakuEzr
SJoVAFkwj/TQIOX8ShlwEVQb0qvd4zOGQ3imrqOKNtD164UDseLiF56p+CTMpzpesjMcC4vUjCVn
qFg+dX2PAYghY2EUfrXAKPR3mjyKIfyxdc7lVLCBWXbEvytLJpO9KkO7x/jcIQac2z/hoEA42Wdi
sZfKkiXn6Pf/eMc/6OPgrUfAznqM/ayOodVb1k8bZATRX/e7HGQQjXdi9IxT8ebrEaLIBTwz833g
op8+UFmDEkhYIxwEjeSmy4HW9TdVuJ0dTz/UMm7mL8xv44HAm8y2rgJ2H7JXulDHp50IbVBDYWR7
O5awp610yadaGTjD3//0X+Avk1vxjWAsOQKAhDevw8xGDgZRpkyT8BPyaL81N0e5fbvlZchL69nK
CONp3SwdMmVIDn0olDVa83RsJQA3TkQHmtDVk4sLXmvpGJ3CDridGq9j5JCswzp9nFx1NVSxcBWW
IXZWnEo6rQmtaPsWZHPyZ+HAmto9BsR+k0K4YP0sP3R7QMfchuF0zxRhAsBd5bOOAboh9vFdkr0e
AwalGQ8PWFgIti7DCyhYqNMdxTKchCT523ID78OygHozEDWROmdikWxWimU/GJZ4MWk3qBiwrWZq
Dcm/SaZ/ubI1hEOXDtli6EpBaixrwYDhkiHpngYzGIW6YF61iuIBNiOVVm8el0CUJHzpayQsJx6C
VW2LsmtF+MXM8X+MPJel+VQPPuG0U24J1qKjYoWzFXUttFx2Qu3Z+rfxQtVRYGTgJj47abbufHBJ
YWFI4LecMC0gumWucirKTpeI3S9q/JMk3nkdrHDzzWexcfA8IxjB3X3CEIlwhekTJgwBjYxbY9e5
UMC0Jy4LoX0Wagpg7QnlewdtOh/93Palkg6sM6SOl8JMW9BgpJzyvisHKyjRN+89lptGEeJIjiCl
6s/5AFN2wtyADTfFvDqrwNMaS4s69ZGDwL3i0oifj4YGouAw3H7fapgQr9OHXsTdLKC3O46sNDlJ
OO/1LhR38rfDlJyxM7atHXOeEqN4IR1MFJlI5NrtCVwUg9qqWiyZ0JA8OMSyhAANVuy/xYfVBczy
7xb29JtaXo9JyUxNiHZJYVXHy+6Q7OoP5G7zL3Msh1WzDjEM0yGPKsn+YTdRy8e2FsImTX+SqKMZ
ex6YezHH55JKwhmzp1XG2iwV9b/3p0TYZBQMvd3AqtH8Lr5lR/zRLtj8njgTYBpCgsDIW0wGUloa
Ee3j/If7mTWjMyI8NKgr2i++KlwTHtt7zSUTSof7/NYhFi/SzKDIlLQpPmE8Mbm6TJXHDgiHVLSc
KuxSnQuWu5kkAQoFrumN8gQM1YMMHzaLpQ3BrcbSo6s3NQdySTidAcdrPjTO56D52wXOdXQSlEpR
trzbz3B9SCkk7aabmmHp5Fvier2Hfwpij/qUpCkGngycr+ibz9zxXQF6rMp0Z56P+YLaYkFVb7sB
v1dNiIMp/fIpzFZY4V/3Oq6B3dFshGv7ZzPO9C09xQQe4f5k20hF/zE8K4kx+qaL2LVh1opH3lGn
MXY/8/qbThnVG784e+WfoYGTfuZhaju0KpI3tPrv8HP8gqGD7aI+l4dARFtTN2jvkBtiey4HEVhN
DBi977sVvQQgW0fjeQLOO3eAA44llGOu/TgKQzFJ2VDXVDCLr46mLLz1NGdU+VjBCfKmovpVOiUJ
1jCm7NOM+VDmISKJaaXpZil69+YV6n2ZiSwQVbUBVlN8ZzMFI3VuzGzWo3WwW47MqtJwm1o5hlhB
HWBbYkYskqMqrWns4I3SdK8FQ8DKs/LZY44nbuctLv4y080PGd2hO2pxZWnVbhxsHozKxWG0j/Rf
4c/SmNezolTFXPm+uBxNQOeYU8/1FhHd6GOwmZ/QTBAoM3ncBeyevbF/FJMXPPZLMKweQizvaFxW
xOjhH+9xko7OGd1QPB1wrHfA6IVG7HIkhkL/TQjPjEmFUs9w2VE+S15VwPd19ve7x7/kGL1hcWBw
PBp6ivBdO544O76VfDHYsqohoMlU/VSx/tTdtjh93JgBPg2ZY37i2SHiMi9fIDYbZ379/lZ0yVqD
UaQtrSGYC9kMG7X1gvrwIH+5+mUxT9Xl3XJn/5pHS6IMIdySk8H+b3zXDd/0ahxZcjZiIvA5LD+Y
CIjWHDb3U2F5FoU35TvbDCDP0Gup4FEKnEbf3NkmsbmE8yj51v2XvyiMND98hKhtsZhsURLGcbCu
sx8IQIKzMhHjoQyMZMb09k2+DCJZT9RpaalU0b3iNHYKb4XFIZemqJDMEkdJCSrz5tXT5VyB6zOT
dkjIob34lF7uO5sXApwQPK4WQt5xYTJqKKELW0+rUbTPyNlyU8vjWfkCnHnPOXBJ1J3sqxDVLOX+
yZ3Vhltnv4B+8/IZMb2ENaYFOJyscbEMzNXrh2PoKmt/Cz75xGKf3crzA6+dnX1hj8TIPP3UqMWB
+CFep994ZnCqOiDyxMcSTV6CfzbELbcK6rND7BqdyZG4G991Q/cqNHWZOkCsu9nr802HU1AabYDw
yClnBwTI34R4j6V/rzMLa/NVNZ5lisFNpGRGa7mh9oYqZvrtZRwH/LMoccFMgUUqsmX77Xyh04NK
zu73MLEniqtZxu+Vtv2QJ1HicuxjtGHip52SlReR54KiQNF84wa+3/ztYGS0yKc1OHjIDv0ewlA1
caRIw7Px6a1mZJxZDw9u7tlwTazKeR3jRCQdPR+WvlBqjDDldqpywkwx0O2//7PEV5hZt7oqCIe3
N0CwGWfEdYeiVvY7LbRKa9iUDIP2R228O3JwIJeSDISJ3hCIjCMbHpLzJUWIi4WrpFr4nKzKrU8Y
FCqscXfsJBrBNL50Gpi1S5/UxAFJTJnLJ2dDf0aCIcLUXqT5vFZHEsR1+5o7awtdsQKbARzhOIng
Kr4bDV7yNoV3cunLlNPgz+25O53NBpLVI8+bPfeUUb5wCb9P8XMuERuxbD3DWrqHbT+ssKpSfUR/
fw8Yo2CCsCLKCRthBxIP18GTWImqf5+koV9JN1Tn6Of72hMxkwS0q6mWXwDSQPWjjl5MZkF3cv14
lWDGRCr2fC2ULE5iNHjRMY0OSJe5XMBlQVWLZuSvW5fewGnY1Ipo2br44hx76RC5WlGnRCCMsXzn
1wUtzxbj4f7TZc3n3oyOS1xLO9JT1iUR1edJpkSYw1hO3Ub+i32B34WyCGOIIFtxf+ueMCzNvx0v
ryZ+RRuLmak/yPTpMNijHz+neJd5hNW/nWzwLX0+u1IByacD0moQQnivKDRfh1HAz0CUEqDttcnR
ZUuEld9Eikb04QUp2ySWneQUyEg7liaI6XI6Zo9vIVD/ZNNWMQwyCiZZsIbGSph4cIAPkKaQOpE/
+moyvcb8V7Dbg3hYxMtVcSaDwy/20A25ipq3guO72XZF6YlneKrf5dgE4FWAG+rpoHzusoP/LAy+
398j4yyKVJcXk98VmfD1/8g6ETrnUQ6E3D855RHILa5hkftXvtRbuweqpHv1ZHmoTaHF3yU84pT6
sUHjTYY0QQDoTkMujPhqJ5hE+5lDzsXyhwrTVBTiAoWJT142XmIj0XW58Zy8JMgPQzfxfwib0Snp
C4jdKj2/zOjjjz3PHWfzefu+5Y7e12+3zaZAusdjCue+owWP+VXzeJb69Z9PRNOsfoPzLuTMMXu2
0lZ5G4B3/0k3qcUb2ad+gqc3AiFLFgWcX7+UjR0c///417WEprWR/oLcFgODmeSZWG+wEv8f2ZQ7
pVyFUtxCAflRzRWgEdQhlvgzeTuG56s6zMN1mEn04wjteCXrkoUa1n3xvFQjlqs64QcsXmr8m7k7
WbqLNTJe2uAiYO826AK7cOwqOnxEa+4Cfvt6a59Df5ZcQvSqBXRSQAqbXgSgjHNHkK8yMnF0gQCW
pdKmHwDw73ObZwQ2CdnltlIN2I5v/OAwDIKtTeaKjXSeVfugSjbrSbksm7pN7211g1mh2UGjCDcg
lM6LSTPo+w2Mv1u1T4a0AUtK8GN8Vfdkc3Cvpb8apr91nzgjlD6t5EuuecwxxV4KqOQIHvZMv3rD
S8ZvOYZNIZs8+DZrnwJEdz/XrhtEuWgmWaizPuMEYc05cWyU7DQCo8vYd9aYqUKFeBAfaNOXQbO7
h+l4dS+G3DiFNJuizyDR139yVt2rn5uzk8KVG4QBcO/SMKnKxBWA68oy395xMWTvUciPnj34e8oi
zbXvxIfWSj9VdaJcOt0Hp/BUJHKCh85OSBqToCSu7B2Kd0j0TPmwhinSvLl6MRnyKNNJV7/ZK7xT
ryTOL0UAbbZw/DAa1RO0kHFla3Cr7BxLKep1it/gR6HRAt6hka8oHOh/pRaBa1/00WFznnJ16mKg
1Vk++LvPycfYPVNYGcO5t9kP7Td+WL7fc5wyVOShKPPuyJU0RV87jgHtU0Uue48a8JPCjgrB8K2W
5r2qg95AMWzwzdPtqASrEEjCIcZaysTgSR0G0HaO1VHZkpAVHLGk898SXYtQLo5Sj/uHljp7yY9I
SMi5I7AEiL3Grlt6WO7BKrsd2Rm+5k+jK+HaRFYcMJP4YtG1JWwUvDZfCizZEG9yQHfdsR/FVpjd
2X41mItlCkRUy4X8flzltHZgYLrguaBdwBBTtWOpcWisBu0XP0bb7G5Fc7L8lHKtj2Z5rDQiU3qi
mJaT79suUKxCdksA7kJ1oOI/4iVKMH19S2l415XEyzSN2u4gl4eDmfg43boRSbmja/Vm1CelkVQB
gWjISSEyuzj5a4WyXMVBFnC5Jusrr2vC5xMJhGFEsayroyv3CBk7Yr2SC9/yzauMwGfaKaRvnfv2
w0unv5SHlcdCvLfZiBejpvKNkI7WXvqd/4gmsZc51eCRGBiFogXDEJcXQ+eYehFOA6AW0q3VppsN
7nIRfKdGusMktZI2TCxJ2Um/2jvDJVKwwC6depHrG563dSKev2SCxnKTlmfiS08Wn2cYPgub0BFy
KtDU+GzFD2wimkVaZ8wtXmsjgonOkc1MPDxVDu4xRzOodj5C4Oa4hDVh2ZEAevqWvQawtAKlylvD
x9cbZnODXFq2hj+t1tpap8UehMyXXnorHxYrWYLiW+D4EOt6r+ntWcr9aoQZUqxFJxQo29dkJlg0
9IlGgBgrkqyZ5N3Y4aOgSmoo6IorB6JmsLiLrH9zhhdq9sT9czj8AZitXxS3qM3JTkxiAXR0Fq5b
le9+WjheL4sxGh587+9dQ63KEZYTCOcLWw7FlAdD+qKSBn+Jevpn2Vds5Ki8q78u567X1mHXpF9L
wyGeA31a/B+m6i5b0OG2OzDM6boZSyoqfATeOkbHaX73L20LC3qyCc8ZIJywroHFdg8gw4QUdl4G
Jx0bDM5+HHcptvf6u56NWgMLFJdQAv8M3E6zbCGnIsQXqmnQi/X3XRPAyVBBGUmD1KP1pFJrZbYo
wGk1RA5sSK6Qk9WArXCn4TAQ9OOtoLRiLTy+KAnl1xm+pshSKGFYcSmh1/F55xiINu1mhTlg3jvJ
iGJZHCbUVoBdA4F7N3LPxx+84itrFac562J8yxVZfXp9/+src/SGiZZSSxfEGg4YtMH+DBXzFvJi
pCAwHedJlE0YsOFvaYBBVHAWWUrmnde9unHAARKkZ0WdjGhEeHuIESDSadBJYR+IT796udkhmy6h
WalC8SmvG9E+oOTEtIJCTUHJ1KzXeirNhnOhXGNGVKUqMkmps3n8TOgdNjlIHmeFlV+BmVvuLOBC
5Ja35xz4DBvxxO+MwFtCVfNFRig+0jLP+4zKzS+yaqXcmFL7Aw9eXjZW2XK87+7VvvTgTx6qFf/Y
43Q1fjxY/RqZCC64CCEhnbu6+Wn2Gnz2Vqs+mHAyksO4FCmjgrFElYelR+eOWaKBLvuWOeN6/w31
caLjTPcRM+p/qqOACaC2MuFkB/4nTL+kv2sPbgSYBYMcQVeZ14SFZrnvgEind+Eh8Z3mkwkRCCHo
HDJEt5Imcmd4BTb4XvEBnZcH9pls5PiMj6KPypLRG+3djLSBCfIbwPyCEEWWbiL2tt3xkyayFB7N
+nWw7651HXnfp8GroQKTrjjlnqX9D0UOZMTdCp2oHL85QlXFNquPj9QcMFzkzMLP6nyW4wcQVT1G
yneNrcy0Ck2qjr0gKt1gE0773YqRpcqA1qGOGy71x1xsLcBxZ0Fo4dj+qYcyOloUs0kQ4FITE8ME
GDgNiAF0Imq0G3JZ+U9YlkIERY52OTrwdxrQkbM0ZItpaSFX1gPnRPVioYzgis8gpAoZUt9SjIMx
tODeFDlLehrp+3pFv+DYemPpVKHw6fz7j9aeB7m7KLMn1Hd8ZTq6hhvcRD22y3q+BVk2JAXoi6FY
fehouJTPSbLOR0EVhrTeK1zc13YLLC3brCYtAya3Xs6icxYsufg4I3tCzzFvApqs0k+pEPJQLkkK
4DUsfSzo9Cz1wr+ZaojGC/IxVCCsJnnzPHhii+np3Yu2+WiFbs+9JeSqX7MYQxWhpxi/FGD2RIel
fuzWbbpEb5xLjddI1BU+4spBKVDxxtVKVFc3SY43bX2jDQt8Xk1YFh0OxTW+PTZYchijEU0j3c7U
4RgGbDMGc5owgvox++7YNz6zgLiNLqW8dqKC1Nst4uuCobIwy0dTDWZN1y7MoOI6eljmRem6YGCy
dx1J3xXgF2l3wJhIVqeFp/VsJqWDZVOqcJrTdZutxCItl+GCtlKBcY0Ph5Mtnfp3yyI7RaUevKYQ
k68VgFOdp78a6I2JiTbmwS4oxUTK3ebRbv8MbCSqE3pasmjLQ5pS2BOl9DpaT7laU5ArI5KjmlHE
c8UVUaUZ1dxegMcaA4CXfReo46d/SAISR1HdbyN0k43EC1aVBzW5j47wylbKrAFaTcymvuUlzE/7
Zc7hCposUe83Kd14AJH+T+dOQ3MlJByqO6XefueWOJswa1dzrJmXZMM+9jeSm4YGDsb9I2ZYCp8H
CzkQ0BQszAkfguLIbJKkdx8uBUHq2QSxsVWpTDy3YMgdT7IlornYpsyOTUF7uv6ExIFOiZI+DXsC
9esbUji/mMRsswd60wWQlAUYGI9lhEFMa5ojOgvtw7U36X4htKo2vdmG/Oz+kO3u379phVyGXDkQ
/NvkRWw8J+QiPCNP6sK68dvJm8a8Xa6Nein08OKrGf7rZ0zVYGHbfBF6caIVB2+OzXxEOk/Ojtlm
NPb9MK3TMuYxotvrjC43nom3qIqobsYJw34Gb08JnMqHM/57Ah4YCaqLU4AGyqJJZHWTyCZ1ATfN
jr4VYGU4l9tLgW1jgDgLtK2LPsy7REqeHLC+UPcHT0r2HyOLIblSfDnl1G3PGmdTjvyfaHAdSQuS
T/jZ6qqJpCcoiFL819+XFfLrut88kSfHdEA9K+s4WjfjbmhkxPbFRSddOeEXk99kxKJJtDrLuaQQ
giZBig5UhGb44oZLHecpA0KO+oltdiqPbv0RfXj7i30+Wm5AN8HLx29rntkR0MCjFn4cyMV7cNpR
HyvGe6KZJm3SwB5IbiejpBZzBeqXbpafcBf8oo/NAG/BqCxlWDypYol5NQbjgAagmuH1kmuQIsAh
1JLd/bbzJa2mrAScCEuM9PNsaGTqMxOvd7EXuNHcqW9d1MZSh9M6hg80InMmTuBWTUht0W9ay81Y
mYw4JhiHUZkWRMlI7t+GIcrFrVG5bAWJ9gqza8jKxpdV1pk4hny9KV/0Vvp7YUUrqW74MCrvHZXx
JVuiazijw6jNdxXdyxdE6WltV6e8mXhn1GKeonD8m17kh8fWmVagZx+3XlDPjn+IX9mbI6vcmTMd
7asHWkOc25N8d03T5EdUW9xJBxuTcb4FE7Vx+VfSlG27inSAbBZ7wMe+GYYrEndYxEMieRjQPqmV
v62NzCmxIUtrn105JaB2NgieyjumiAksT6/XXvfhIu0Is8ZO3Ur7/5CL4Frxc1DkHMh5ypBO4IfH
tsF9t5c9iwOIdz4dxeVP+FaZfyiDemijfOYBz5oOdDuSXvelavdWZpPndhbrKzMYLxX38BZs5wfq
WbfUgxQD0+moXFj7AgcLV9ASrLDzDIJWi7/Jr2rI0Pz1h7cqkWiGr4nEQn/4y3mRAjnlmTWjWVnY
lN13SgWXIv0VwlPXvxfmjCFWPB1JOGCuasGvhIFrtMzp/xAFQzUH8iKfun9JZzQFvhWljL/4hj+6
fyupAhsF3o0sR9QlCf9HeG6TRGFdz0E49OeoSzWQsyrXHr0qy9pZUpLTNv4NzdFYZDA8H5t+AJc8
0KcXM/GFvhGV6CmNH1DxhSKPAyWmbJKy5QewE04JxlJ+5CiIbpQSdEUnjdoqvHt08YggcF63jWlE
d/rH5GNuHJdcaUK7gbJIYdy1kqwJtzgpd1r85eNcep92EcSIKf0eYYgd25LLuTXvRyLqH5xM8Hc5
R3ZE3jBrNQh3YY7LG2QLviS9KRNmeYLMyxAKv9yhPYdlzDTKjZBPLyyQvpBEijhphxRPzSzOyBCL
KRrQ4ZyTYdO/IiTjs0zCKN2Vv3ygueBPuq4gXTFcKZLqn8fNi+DnfJVHtVrO57eKeRfTPNFkp/Xb
fbDU8A72MaRbefLsBNGHQ376rzGlCrkdZwRF1lT9ZgGGrITK0dyVPGPexpkk16AJosI4NMCLyPlH
3xY12lIZc140eciE1PcsTxsEhQShTmAv33171LRJw78bQlYz4h5WLx2pCqR454h9Xawq1cuKrOKT
0Pex+OcX++L7tbV8eTijKhH054+o+ZsgHGRN6N+6/QfE/dmmfgHx3cbxHKLN2Q68eMD17iKM4Zk0
5/24zpKfJ0nDg8cfbSlUDna3lVoA7f1IFvrnSaFB4wQ7WM0sKRvBCHze7W8HNFpJNfCkhJD6OzId
X1QPwZxsRdvmNvRu8h35ewrhQYnE/dPPUuNKv2M/g1BU1iPUBapVS2ntWgum6VLJPlqhhXnpEdmQ
ZKT3rrNKfGolohpJGGNEuGSIZzBZM7+Kg7tJqfiXXghZZi/LmHainMmUvkvCcDETx3dWiHq5yD7c
j05puDisZi5J/p3vBDY0vO54BXjRDP3D9wyvrQ29GetrYwQ/M3Wdyiadf7L8LtzMVhKh4nwaN2oH
Xig24j7jHERUamdZxAObnQmU0a88wN7f8QotzNa6xjSwuwMLyy6OnVzJYtDCuz0Yp6bJ32l6JhQF
FAEOm9fyy49MwrP2vDYjyF5sGbV4ODKJKB5xCDTifjCOvxgAE26pqQt9I/tHjNDWP83gMhnNsqha
R1LAJUkqNPPsQKkvFTy4PFO2C7ie2klzsnRMJmoly5avAeUPIhC09puJQzy+YtnwMTSGpGLv+Bya
Y1skkv18/sVVfBoTM66GoCrlhwrRmPezuBxLTPq11p/2/9OpybgxO4usDB3c0d1B8tGy+1N7IJcx
u3RuOqvzE6zp50RJM+FfJ5G5rwO5qKRqoAnI2tJqG8KfcFEI59plktdiTedU8n+FqGC57fP2O2w1
NJJjIa9WkKvty9b8lIW34oy4axaqr66KtN6W8LGlV7txcltHmoPMLv+MR0x30SR3SWJyVrE/qusS
EZY3O52f2uVeInnkS9IX11PBkgwq2Ofw26UuSX/zKZkraa2CkMy/QAgLMRUb2Fxc1E4/V5e7ZuPG
xzN0NrgxiXo3HVeSq+SmsjeyQoKwO5aN6ovd9idMuWEDlExcv+1+qYP7IUGjLuRZI1TUDm4VpoCG
48HFCBFPZkGgYSATgeIMG88krvFTKvOGpOrqjXfspOXv5wtLwyCuOd9AmrzQAnx/lmqjnhNKz+Nl
YN9v6HKjDbAb2qCE2Chz2/20lXMw9OCf6IcvBHyP2zU0vmj8rj+JwDIRk9TM9SYfqOt4ZuUFqQAI
I0KeOIa5AMUipi1LSjE0+pm9blyDTxYIXOzc/lZCJQtOS56IPnTR7zZNxX/ol9qW39VOvKfz+WYa
EgEtTUxZXdQSuCFWFR3sT+QP7s0PS3bxPkGD3VkNjMDWSzjVCYX6GtHRZcDI2RmveBpC2aNviRxh
FM3fDmVQR2kXHwHqDUvTysVgGznmFEB0DFgq/YLIR7vorJA2syCPu7oh3pf6JebJRvqGklVVtCbu
PxlhxFCi/oWh/IkY2txdT18PCqLEYuIyxBBh79v96V01MiWhKtL/kyn0q9PIzqsTQ0TxarGH4lYU
ZUPwHnjpG4LJKdYLEhfA4aUB55L201FXbRUdw8z4xK1USR3FtWRnKoddkbjKB3SADz9Tjj9qs1eE
7LYG2K/YJdxAIxGp2mtNlbWEDRpfiwBCp9jwDddKv9iVJSrx3ZVjFBoyY9u8Q13xXVhgzt60lOI1
7Uct4ynklIfDZ2hE8QmO0QDyBaugkjo3Iyh/QccfWwwTpbInpcOx12RnYgkIlqHxCkGvrI2Fzour
EevLmtBw+g/zfAkF2wsj60kyZw1vLnWFpgMVq6ZCLjptHxQuK98Dua8Lb78/YUYNl7SXjTwj/7iv
x8PvxbKVGs3uu0WorEd97twuD6hRo8STePBro9wZ9mLQwOdQb/Gfp6+QM6CV43vLddiyqCeRLZo+
Q+XO1WopAu8IEWFzGY0NXBuUDHF1MAuVgTiwyZSdXKJcFnqosbXXBaKkwZ084cEtN8uGI0TdbDcB
/CQYePbj2v4swo+MmhSOAQcZnpuXYgkRnCWdnWJ8jXzcQcURT/ZdSMLnMdQVM0lSZgAY8B6fn5LE
PUhBCrzGATyzMBB+ARe0JZ3nG5+0nh535DnnYg+CUFWryIIUj5E8tSbyWRrtxEKVHi1ISGT1+Gg+
lN3A+ntOMECcPYO8yEx+h1rYfaCpQYQ67T3SvDUBqy4+t5V6QIYPRM8N3aC6ek+R2xtWgWvC18sw
aLFrdaqx8ndvNX0cOSuLhbh52FftKXTDSg/4HwtCkHoWdXx6eKM3Az039Nn2j2R2hVrsroZbTjO7
2rE0EWCRnJibHUu3CeuAvkZL8+wM4OO/7jIGpovmH13bx0S1G4n+ZRTzsz/ZdTb0X4y8e1Tp/4X9
+YeK4V3wJzbWrHaopc9sOEHPrJf8uJ5XhaFA1nk1sSIQiU4q3yyc4eC/iMIQ10F8vpsMYXWbJGcG
lcjX/NlAvAS1MgqLeSCfnqdGd8qSYnOUnbHb2zs+WWUjPCNPOHMtrnZkUbOHaS2ccrbqHLBlqoIl
1cu1CaanyXImplt+JFdRgXGin9cbb5Ol1j/R8AxYYwgdbBwsrj08rnkEWYklhvX6s0hmi7PHSSAj
dEgeEAm1sNfKBurzNW9xJeFJdMzwIolS/FNqmd6SEz7JeTi5yJ8r+QP/EpdM6c2FDyWcweiVq4dG
/pFthRPAQrnhikHX1GSrMGf6RSWZt6FfZzctFz0C39lbGm0X+3Ipn+MpG5ErkQNwfqXh6on1klYm
X1sb8ed8VPUEN9N9m7JbpLS8UjJTO8fsYYLxH1hQPZMT12oFc+ZMqabRS5w0tAylsPfYhNrTFiE9
LJYRo61QpOOmYjssXIIiNhWJOhQ+LPJ3qwBik1DyB91y5KXMGgvhL9KCE8JdhnQRU9eaEnj8bM7q
LleEsByZRXS38Wwj9jiHAvrZUNPxuqKa/BNcfqdgGIw2w2pcsvBOVHohOmqOABFx2HdH2c+nBxHQ
9bKoq4sFonuWZP7UQYzhgcdTQ+/0pu5fidZH5QywsdKaH8VfhwMr6R/us3Spk7MbrhRLVSRnwbkz
FUMfo4Qe4qd4PD4JBxB3lsdOKi+QmqMuaFtK/IjCiJMin7y54MKKUjIIAIual1QA0jS9Wve1J8bU
gEsgQ8MhFkVUPyTsxj5g7dKFhmD0lJkUT5B1a2RcVghNIuT/NhbwcU7Vd+DVHt49idx7L5eqlnjt
5gW4z7UwpyX938khldmey09dXP7GPP3vXFK+U7xuuh29ZT3q2Bh16vtl40P4i0QGxZdw6r+Q6TRl
Vst/+FZb0eS3b0QTcPnYv/XB8nF//myeJvDYFox0j/S1QbWjAUpxFe2CHzFwOu+9HXbKWRxwmSzg
GHxbasFhXpWMytVbJ3Shxz+Uz55xSO92GINKBuIS2SydzDnrOYA1urCbHnyG6NpUlThLkHo36Wpl
HgBLbHQDie33ENHsA4ghn09clslUbrVmmKnMC9y9DVGPt+IKHPpgPjDqf6ZI6OZZC3bZuaGQHuD1
f5UYKw6Za5grYc7CLV+gRkZgzX4dc0RV3yHnBGOv7yhjhn153f+hb1Avi4dBTjfJf+2s5pMC0jyQ
soIqLpVubyu6gCOobRaMreBSmZQRx7D1iaILJI3THcbVQ/da47fhH4d9Kl/+WU0ASSUWPMLD9Ul2
hYn2YNNczUChYHcDDe11tvvwqTebV5Hf1476HqPX1arOC8YmHxN/Qkq3YtuW0ZUi9C3KhhZkjUXc
lOPliryALhXLB7JUswVnquK6ucqZptE3Vz2fhAMB9ADGfetZ4CpL6oGnO4AQCWupoGX0FoK4kI3K
Wjb1sQ0cbPpHaqBA4hHd/lGsDfsHO1cbWoKd22G+1Ya59X6g57NdRqzIDlpoMGkXozY0aD4TLyvd
Ppz0CJHReA3cqXqkMoJtvnttYNqBSWOrHkLt3c2CZP4HBoI3Pc54R77BaQ8wW9D6JEN7pf40PJAZ
ktWGQxZv/B5Sr/8BB4NdwIyrEMhQTUYu/2kVT20Usq57+eqRF/4aGhDVfhmuHsjYOmO9/0WYzXqM
70AjMY3+qwOEOheY+iqASSNmoEd3PfWTR9zNNNS+fGxXWyFC07k+1yMRXEa5tSE4ev4J0pbQJY22
BIqvm+9SusHURaeOwgwj6oGu0bsWYxTJ296lCip6/a5YqtHsZvi6mgzm+DJaL7fuWp3+Vx2BbBeZ
FoCqHTVdmPRD+sEskqoepRk0j23p9znfwnQNNqx2So1l6iQSdhmkXO65aIYxFni0LOtg5UrhK6Ys
5Sz3cVBFTYQAErusVn6xU62I56f6XQnM6xe9Km+4AnmRGZaHwUkHnjwQQZMkyBZKytj0KitrQVQO
UlTh9N1TW18Qhbl77JVSEb+GUIqEFWmt2QwC+oTFEWsVuGdtqP6OWIQe+wDE6XKS2416EIi/aZRn
MkRiROrtBj/0iXuZsfxW4qhjwMIKn0wHVz0eRrRuYfWi/V2HM1nIW3Bn2Ly8vAECxAJ0lf48v+8j
D9KRgivrjj03FjGu35Gd0S8x9inPVdF81OEoXHgJFGpdzE5oJITRgWWL1al9IoIypSGlbmqdIT+i
tqfcZnLOSj2EeMuu5dd7IT6JVD9j7jWpHpo7jh/d0tDp/zv5yxDBYHyvj02GxFVN339hB6co7lpz
6PcMKBbd7Fuvl1+rC/eNXvwN5reTME9QOmHAWIc7nrroDoCl5tPp7SdGAqam0yuGgQopKgaQ3ZMa
XrWZK1neRhx8TVb++XbczM67rRZu1UZzh8QkQGh1Gs5wKSRI6iFblOnV9gmO+wX0nrnxD51wmZLI
gAoGQDFBQ5BXL090CVybi4pdACj3etUx+A2lbGyAYMPpvepxh7OAQir6xWXadrQ99BMqFFRPyMK4
HMv+x5DswY44iCShN/rTjG+ZkU/K1wtDkcyuG1XYygdlcH/hKrT1swPqY/+aXju/zpHtkAi9aJb8
A6Z0vKlw5Rv1kPi6wcbyfmEYmFLEgwz/YczYaqbNtF1Z9Od/02Qusko+19yLXtplGg/OhzflnHVk
aU8HIlAcfSyh0KxFymlUavWDi7qDhs+O14wP3abMUR9LK4hzmWgctuDZTEUcgT59yS1a0RIOaaoU
Efs4QRbzqtJfXxzFAN1MNRwEQ/Bc2dlLB1g56A/j4D9q1pCpd+4nz26f7NUR64mgg+Qiw90Ecrp8
uHhfh45nTsGBaJotkURLjB+kHGbbx3WkbLI1cRGBPU+Shqg/o2lbVLUq1ErjeLVe8cSAuYPpDM8/
q+LkxU+GF7Mq+I+GzYxz9iwonpjEj6Z0l0djjebINgNnOtwYPJ8DfEXklC47aSkLu1sx6cevPCSq
V2utYXr0HfxdVr6RcxS46JWwAl5OizT93Q9SsPmOCYD7ymiDjAZ1LGKo/TIZxCRomrHGND1989DA
prWPPpzozqYZ9FRFdq9Ca1m3H81bUzzmWIqzfKrEDAzSPltmsDPD5+YefWN/nECiaLJ9RBc/uQr1
k+0TI93ELLmbpJqyCgOftFF8Wai3qKdjpud2kCNKOtsIfKWdNgVeNaNSSuNmy9Y0um/sgOMR2J4W
9aYlf1TV8QkALwK8DhMVRJFuNcFVakcvyUU1WPnUSEzpImNInmmQFzrkokutaMUFiI2QqFdcMDVr
0A1NkXnc6rGvY9QKGMsyyUbE3RrWdYXBfA9+fHK2HZXt5fYHw5cXtclOINoXvvisEFtmmfhYvVMF
2ZAJGWR89OKxLtLRYYOYvxTsGzTlqfowaxs39qMM4P/qu3JflfkVAvWirW/cJjh3Pyr7/diCpFN3
g7hVK1vxhoQCmXNSwuLvwnEbxbnu7pIjJsRxDEwM1wROke7tf+yDjXmHopoN9Rys1STTaE0m2et/
QjBsMY3LHgg8liRRbafbzQ6xPgHllMbrOOgKPvtT13k396ZCTuxb+LiviglWbQH2cIt+rsWtU4+J
fRYxZzpX4U1cChL91Ced8iX5cqGZlr8RzVJ+kRhuVsGpovAkf+9dRtWvO/6ty/cACyUKzAJX7xIL
dUuN/j5rRQ9ne0EnZmBil16WLaZkrGikBuR3+cN3QI70ZNOEt1YIE4bVmbCyh/CMhDEVg7AIOEwg
5zzKZrJMgO0GnhlDI1S9uebFmZvQK2tjsXBELEVmsmmd0nCrMs/TInbA4XUyvHCZYoWMI+ff5UOj
qfXmMWn9Mull/TT1Dhv4ZJ/262f51qwBTErtfN846w1/J8OFVgLnCUlyqoTLiSwReupGjArwDF47
LjEFZwHrzOGML5UNONc3IS0g1cSDh/+ExX8TxYn7U9Ts/ZvydU+eYaXq1LqAP5bI0ZHuJBM8pggL
/IOGyUso0mk6ReKXSDaDzRD3wogvgsWVHM+xOmm+s9dz1EMVdZNrvfw0e00pzOZqWzcp8jTsNSLx
OK/0TOyleW205oF/oGbVcKjpVVh8q6AhV71uS0HAoqufAE1jnRTrTHKM15mBqthwByAzxZJTqK0F
KCmV7HtcsQrinRP90SJMk1xdwPVwzo1cO9kwSveZXCFHbv2nZPMCa+H0l2D9IeV7S4mN/HYb8XMp
HXAqFfFpBjdV7drE1IfhxrK+VUnJrpfUedOmarhGVNs2dYm2fdnVru+6QIBSClxy5YevPRsjU8sp
0wJFE5P9OO6tds+/NnEncD084wo7QFIkxiQbsZS+GxPH2FAUNJj5FVIU/lV9ZIu3O0BNZPuO1FXZ
mWgxw+UILDDxnxvu5c7IXiejo1E5UawyWHo1s2wu33M+HJZnWliQYZjIIv6YdlSCYVrKmuauZLLc
Hu8a7szQpQikFU4C7+8DgZiIg0Rfq2dfay5FmPfB96WHlDaJMfbktSEEHI2Hk+4AvDudqK3pi2kU
BzHSrCC4whu0sw5po/WPkgaqUL3SRQYDivOrtjK+XP465yhqbPpp9gKYZMc7BFeZDRRDOSoZn/iI
yuUWtO+ipHRtP9OjVBGzMAbnKyTuUz4NccP+kVjPMe5rBsRgcL5zdTEUUbbxhQQ4lClg4geNRkPM
wi/8ccWo1pQOha3j5i487wb65kLgZxlDTf4o/VzW0qk3uOHahjCzyUSx5QNPUtMHjDyU5cnQ3E0z
KHbHfOm7Wp1SRXlbfCf6GteBrYlrWYmyWNCuncdxphjhG9pcebdotgnLxlPyx9JLSG2ntNs6fmjb
3uTuIa/DPl+2mqXz7Bzqtwnqo+Z4+WIAC8c+l7oje3+rEggQf+bQU9lSgkx7ndKJy2hSQ9I0Kll3
9esXnPVhAbjjlWm6e1/wDrq12W5WQpvOlIXSPf54abi54Q+b0UMJKa069/k22dYDZ1yXYh/qt9sX
ehjU2kY4+scMyVBJ/TtS1xNJph65Eb/fUm7+Ge9aT+YcihpGU0BHJ+8FswFV+sP05eXgQ9M/KzFm
XAVHvQ3U0mmRpHvV7/MstJqGvdvTG3Z07CzwC9/z+rvomiqKT5rk0LNKCSuOkQ0BIFFkl+vP/1V0
HR1p2nc30oGq7Gt6cAii8asCxIN6p6kpM5kaq03o1l8BtZeyL+INgVJxB6PPpYcBPLXV5DanZT+I
A05HSh+T3JR6qb199yiznipFSyxffcRjvODsd6zS5exgo3HnT/6pLd7hAnBzHV/r7SBPgtrAN1O4
SEay728djSwSSLD38EX+0CVlJnXPjs8VIouuBqjCc1efLPByKInKQMYAOMztF6v2kw1fAH9L17Bq
16CpnH5yV4W6pUDi5PaSBVLDlzKlK1kRYJrYvDd5kazWKHGLoTDAGh3DD2JqsDn0UgLPwxrNt4iN
yI/4IBDj1bVaRLBnY/vkxzbCBwy1We/v0vnW3XkxSMMsPekDkCp3TQqlGYrp2ZE33o0HiCLlr81a
t+gwywr/CMRMK9x3MFtJCV7zkdrCqjaMIagFutljALDGwQomUFTXAN7kICQhGdGutdFcOcZ3bt5l
tuFMQpGfaMh9EivGJ8R8swb0CIZ0erqB+P0ADk0JgmQvBiEqIAWaUwFoCGQBu4wtjQhsNJPy0FKQ
8csTxHuIvLGMX7hYeK0mbM5p1ysPWfNKZgIOujgfRw8JKrX8vMs9/5GV/36sS/ATTIqGpWMwJ4+I
MYtX5ajkecdl+oMqgS9bozH0aveW27LArs1OhJbuMwS2htmaZUgohWbs35ZuZcsqXEl+CTY8eS0E
HKq2znCi1me1XqbtLTjDNmpVF5S5wBjC4HPdoKNNMwKMf5oGEqvG9kE6Y857ifzWOhNSYtAnomZK
aB40630yhO8c3cwRfjZv3um5IH0+phHLKjiVbLd0zBxZL4R0XXXFFBAZwvFKbf9z7HMlKXs6B6ZK
flmcS4jOW+J5K34JbITX+KsHsMRZXyb0NGyfINJuW9boMNApE4XsHqMbrzrZ/VXxFtwjIKGlXJ4o
UtPgUlXNEetwQsh3yyIdOKR8bsO7kB3Oc2Pt33UbUOZnSynpmm6WXQ8RYPJbA56xCN0SMo9HaWt7
8PLFBtXB3Y6PEZUWpmamwTLf/hZEi4/BNZu6EAL/Ir4RvD1+uNyLkdK1IuQDubrz2sOnicl6Dciu
nUHBWTfeLRyaybnwHNhb/is2lpe9Hm+wcKog3W7ahfAhtfse/m8WbT0S4wThRP3oPWQjBITTSIzV
ETgvN5Um6g/J3RmXWDw5ikbsdp2hN/qbVr9fnQcYH3lYvxLJDkz1gIPYjst62imprVUvG2d6c8xF
EJgpsSDq4VdN6vqXfOhWD++XpOXI1sgFdnOftcX4sHNU61IogmWylKBZqtlBUuPU1fVDsg4h9dVh
x32yClp36IrMOBzjdZr/eMeDlGb0WlGAbxBPrELGhuVyy7xO8ZHl61pTdFE7flmsHz4moQGw+Ozo
WTa0hcX+eQySP4rC80rP9lFuGUAtx/ZtoxDe5Fyf83MRGOtpRSy7g5R/5JZsMQAEhtqpIrcTXWO5
eUapMt1LhZJT+1sFIhySZhQD/Tgl99K/xZ5fAXaCK2ecKyZtgg6A4Ts7VPH2k3BWRHWhrTawLq81
9+fRyxip8RMbrCQmFuMOnV/VqMxy6PAkTJf2WQSk8A413/0lOQluyrmPKG0JoKAmtURVIeYrvBPz
7cyoI0xtJpJK0oXTg0WUc7cZTwo5mSz/67h4JL24XtW6S9ejImtFpLpijv44GpLCP8653oh2l5LR
6+iP8/jz8tvvTcy7WxNcvZ0/24MmqNj6ilsSdnybAin2jYJ5Vr1ekJxuhWdKd0h8yYeb/8tdD79o
cgdaAvnMBaZE75ucST8MndPZocMjBd6blFANBeGscvvLPszqk4MYyU24FQsgis9mz9U7uiDjuX03
LotYi63rVjFesT09b5ZCjNNbzYJrTe2W4LIpZ+d9xWzKq6f/ACvgHN7R+43zPcep5EveRhNO1CIU
F5GzvpP05lRzOom03mLf9g0KllROJsv/r5+zwMcEg8RxP9gfZYylksnyU4027oMEd9wA3N+kbJCN
eqiG+ZRdDbdYxupxeKS6D1PH+6PcAI9nXLwz6ueTUmabrmlWZkljzgdDp0Py0QEFm1zbFL92+mcb
VjcaaxJtraaXUdtNYrbu/IzcAziAU4pxkTMajjb/t0zyDwMcVgyo6m+mLIvUomFi3cftbV+pqWNn
t6RmSbtJHlwEonvrviLKejUfRlJlhY1pfwQ2d9GC2jCU5JNfMg8j4n0aOaT13PjvxKInhkI8f4uh
zWeN6l7lW7HlZerfoXvecrbo9J4i54Uy6tiCHovKdVE2OysG9e/ETljJQENr7oPx6gG8zhyMpH5P
zdY0WcNcuV3HaVfVpzsuNZ1v4Ddk8+AKsAOMJNDiYuY8FkYDGQ4PMb97peDZUNWvXOvmFqv6hsxC
lFu4Nnw5qZGT8xT/KqD61kPdgp1uvVNEKLLy93Pd9+2VJfeaXVl0yOGaDios5hs7R0sEhgmT7zVP
N+ool/u8rvKw/mLXSKmeVcngPOE+YIVjfR8zg/34U0hqG+L/hKxEcsrUF1LGhHNtUzP8aNFwcbK2
UbO1alVQScanjF7O/ekTDzKCyXWVQ1Mns5M0LTP0eT4oAFyDeiyFTVKz/KJIDGzOzYWH4WW05+Bk
a6Q2T8/oQALMnoWl0i/ObupuHF1ctkDQOJ21e/xYYDOe19NEtrBnuWdEbHOG8Bfm95lR7amcYBuq
KNtzc40Rohtf6ykaq7vy9t0LoX3Gh9N9fO1tsrSOuPek1w1sJ9Jcx3VV5IiaEviugj3u0SX8goBq
vUXue+/40h63XaLnT4OywgaVdXI6CMV6H3DG+0FyQWihExcmPd2OZTPN0u+9OlzALXApFEqBGy3u
tnXX1eSFkBt96/KpjO7GZayuh+38PSc17bYMK/fw/8wJb/djE4+G0lpvoxOdpj11owKf5R5crsAQ
3KKitM/dY6J3HOqptBd+S5Y5OVlwP1LgfFddCgAolvjl2+05ngWXyaXETsBAvtdBHYJf8Xhi9lIN
BPmVoVpX4SK/pB4PNheXNW/SF93HcYggFY4Nh8sO4GqXWfd2xlY9iKUVz0gjaYxfDc5GwVGyVFRQ
BSZrmvymV6HfJEULFRJYNxPEz4Dlev2/SD7Q/rHzu9zkBuAYYDNWciSxajKcP1+blr/35J1ulT5d
aDMUvT+PE15SJShDhA1F0Lg0QBcX9YIx3kPNE0Fwt9aYxl0O9CTBmKN/Oo0kjoIn9CMHfgyGKn8a
Ju0kHqUAd0AjmV44VJ74bw3TpMfd+hPKpO3ATIrtDafxJFqyJqB++2TY2XYXbOHX1BjZHMdGD5VS
9AguPHnaiqtqTe67eklbbWv6dosvnw81lGqUJy6hPHsF2iK/Bva2+VpNgRIwoUpVPcJkWHtLWnDn
NPQdvzDXM8IcHqGHtNlPMazgzMqtxoLIg6Cu24+iChPp4NqW2JjR7rmTeduX4SRw+ruWDvEOVpGI
mFnVlYnV0HYi7/KmCnFuRVyj+U88BtIpqGlrReS73mFFufXFGzJu5LDbbclW9+PBphzFeywiU4Qe
nrAnJPDnR2yT/RJDcPwP86sz26VoGiEfLFlUaLEldirt4nEKN4RDoHaUQoj7cOeIaUMDxNx0pBWZ
MX0rGyOyeID5buFo+OCLmHBLJGtxhnn8RQpIhaunO0ytU4E9WVIdIa/WMgmDa2NHJRi/21x949Re
upvxrPvjoaxTGChkhbqxNCnYILz8lbYi27hmEh8LDKLK2QcqoRbmQxXkY8KBlOUx0UN/9YMzW7In
X4or54osnfYsdLzNnaVp9tdX0Bm66QCF1RLgKry7INqo4JN9KGTiA4xYii1gTGbLIn8Z9goL5VY+
Lx2H2oqRzb7t/k6NvS5gzrQtjPQ4rPO+PoW9pdR64ftqxjRGCd61fUHFwYiAeeTe7N0aOc38Gh5b
hvVpAZ/y3ZcaeVa8UuhJLwVPZUiY8gqIOwUEDk9ilArm19klQeLmxZrnyMX1ZazZnT8SLFC9LJW5
5pAQsdhmmRBfe5jgpaXDW16kxHnWcwcPzidAiwkd2PAS4LHdQrBEb2Fz663IjUg7TRE9XZfk2Z07
KIx6FcMuW1p8WssF3dFtrBWFT3gDJGScyBX7rBtblJcK9dfTicT99DU02dvQtwFUfle3j5clP1yh
hOu2WHM8NXamYvSFbWdWrbvtDpvjw16nxMy5AciSwrBwTaRSSpgWh4rYuSwe9r/zTeSAg4NQ/LhT
wL9EdI9dfFfbSrBG6eFzqHw1Nasaq6ZBHDNwd4qx2hiZACoS1MQHslkrQRqyjFfW3+/4CxkQyA3O
21udxhZrtoW589tbTpl2OUKzfbjObxn/Dfy59EhAG+VXtI3gYTlzHumOd/pPHaSeZtdptOPz6RLa
3frSsBgwHFGrFV3d9Q/YYkTNHVUMrb1TC7djk8GocxtlbvZRHGloXgZ+intfaRrDxqmedB5biaem
AocMC/jRI5E6VuHLhZv9M+Kq/moZtLqZdhZbM9VbzT7h1A5mu6X1HXXSHeM+yHneNBpT47CHKHAi
JlKtic7wd6OjIAbIimGztwf0Vwc8kdBVGfG1j/IROO7fTHnb+SkPEaGPG9zBpbxgfXbWOjEZI71m
UzZzXKvwCfn5qMyHpAzdoecInGjoicH5ICgNBOSwi9S8aU2UYuLOpEVy3zRCanC3JUCHW+4KwUq0
++9ZmTix5dMoKBb7EhwLUbAWIRQFuGuqlg43VSpwHPe7XLDQCSlg7oLkE48Fo8U1dTJBb6vEyxoX
5g7zPa9da8c5KB+5sCZqOpvhKKImM5enJ/GS8CSc/ad2R0ziGOWg+vvB2OhLOQTNOsymrIRsTqnW
sCGE3g87Q2SPIGEeFBthHXJQnIVze3zmicc6JAYAtvMI0xCMpamFnX0MnYlr5vENQ/K8TRLcm55U
WiDKxmXyNZo4kMEELa9R88w27kizQqJQkB5mht8qCFyOfNG3R3nBeqxj0tscAbP2o14SsaOEQwzl
yBHgLzWlFpHtDy1AWYLLHRNWi07+Hixu1eOiSsZDtyfhwX5NdcIXh/LDDpOd5o/ga6jXlYcstsG3
dZgoBKy3z02Izcv3s2llgx4V3r9k9DD3j/jr+VU5p7ImvEbEwHWkfhOyKMVev1NVrsbf03JQYZJZ
DNJVhalzsMCqRZ5JDo+PGXdygL4aOLXYvo8N7ANnH7/7kfdeRJYhBBBNznqAeR7FQxlpGG0But45
K02TnDWudLR5AjwE3uXqd8M79IngUaVTuAiMwPnM3B1diU0Phb3BW34o31PPhoTF3Tv7buzp/6GV
bE7Q+kaGa72lw0E4RI4ChZ4hpLERkMF6+6mkxuHa1UaRZcN1Pk6uuLZZzskYRsvNS0m76EXtAMbn
CPPQ7FrhxAVGP+sLCLmhIF4UTSIlfZ5s+HcRI27Rwty9dtQ2BEYYPSXqMrWX/hqmHoACnCn6jQGd
C/a7Fu9J5XhRTBnsKj0aoIM703lv3JfrLwHstNIY4yZ6pFstO9wGYyfiMYOB2wPtzK+XwAIu3hS3
3x/KDfLFpDD9o6jtDPKx40xA8AAM7yZNYrSueQw5IR2h9JS1KMhgtjkpTO+h0Cr5Y+tqxyouNusd
zOfRjChwWoC9ROi2Zw8McigkmJRtJErr6WOkWt6rnc184htZxbYCBKE2ToqWlRldFHkmRPR4GPlm
EUuKrZNjL4AS3O8go3y9+B6WDzwQzzoj72DgpQmIIhQHn0nznMG3kdV2aZw6GK/nOY/rTFM0U2kk
0gKP43l7KouCXHNhjM/rczDuApeNh7+PhbcG/bZozG/ttEa5qazVMK1KAM6rDZwd4sU0YGqz5Ppv
l2YnogzD7L8uHAEPl2jnfpT5gsajaetkIJrqewR/zY0lYamI2HhHw9/UfLzfuSKVTAFttrRZSty1
sViuDiy9S7ZHICROlpMtMsXQxPMtU8rx6pfzL07NPXMYcN/eSybcnts2zMrofrr0wzMatOatoqOU
HnuDmXVRtPHScFMbQy0SI44kfwuZh0Q4B9jMyWzvSTtmCQfmHMbmTTC0iz8viF8pQRXcj/gLonOG
Vbd5/5H0S08wkeU6Gl9YRa9vpkhwAd43NqCv0pxvPP2A3fKFHdNiRQK4kWtlu/NR6jyu2dLu0ylY
PgfuPq9KJ5DtEVj2jKeqAs9T9wXsoQUYCCwGSFER7ywQkcVu6COipikL7eACbYiL1Gkm53ik1+10
bE20JUL5UGE0pilJguuDxDVYbIvB0AnPIUZqsOXCibq+iasShm129mSaBSGiZuyglkJPd/YilnHW
1rl5tB0tEqd8QVerVSufTUJJhcT8gPTPCUd1fyheQs1/2sXjRRE5TZVt1qeh9PSOtxONI1q8DNhE
9yVsux6wcr1jhwlWHyBeGmUgcOoeZuXJyA9syGLtz21eWLKfTaXXpTlO2rNnA8tLiYH2SAJ8shNq
7N4A4nr1iKjfQJ0Yk8nfS8/5AhTE1zaYbLn6O8LTfup3OTfpcKqq9fjhRBPPq5JbsYWWwYoVE+0N
69RDct7ICEJqMofucnbk+LzQCLSwk83YtOEAfUf99FMaS4nHxa3GmowVdItUH9jTaKXtwSxDsmjE
a2hD/farA8wr3aJUMwVGJ75nkfNMWyUnSfuMPdvZq2OxTMvXePK67g2KkLxxwYJ0XCpqjhGnpj1o
59L2euzlmkr5REbhiwzuD14TjmvUeN6J7ZY33VI965GuuCHmrBSaJqiq/r3sMtvjxsZ1846K3kFM
y11keXVbj/vUVMbfPd8fS/+2JpRROv8aVSylHFdj7l1oJ+52WqGjHX7lZVFLDeJ4xdH3GJYpYoak
8f2y9cuOj3yul1YTuhc/lK/dnotvRrKtCzQt0PXYNCMfhMNT4bvgZ504iyZdnY3YVyz58W92FxeB
9SIRiNBhBP6K6oE+iTcInXRjWL1jLcp1IVXd1zyOGhtwaETt3An/oJ73RAnaD1EUiUIi2Z0xYQBx
X9YhiODR8Ycq/JQmbk6qa5LdsWy4V0aOUlJg6yMlgWecVdsIRDby8dD7u0U+xHBK0TAHK/hmO3Gq
HnNHAlL51Gm02Pb+Di1o0gN+SW6l2nyUhmIr3zvfRCCATZJZOMPxodxsejbYFnKRNayDMVDpwLfk
fwjlLYB1BH3jM+okjNpQaAn8g3/qQJsGrHCcm0YAI9q0XCks9RSMt7DDHbdns9Ceurp03IfnxFLq
LnO0v3tgo/HjzQKLxu0abU0g9OPUE5qnxTwW3/PJJZSzyTvLWiH8XsiXKW4L+I8SprXLzmiCn7mT
WzIR4znRMiNqb4jAo5G/+FVJL40SFKb18yqVp9DTBHBiJZyV7/iJ+haOFvG0OFNvOlTUa5eqiHnk
qaiMYdT/KccZAPdlGzVnCQC9+wwGzUYGQMwTplMpiQQyzkYfiaHyAvpQPdd4szOr55V8PETQznF0
BQ/y810zHlg09G2H1xuY5uz7FGsDvf7eCuBKjG+agdMNxwYa/08LeMxIidNEx/LfBmdN4gZh9bBX
2xm4esIvBiNoXAdsxLzxrp0fjgdlUV9HGXNlD8gxYOTsN3RJ66Dvm4rmgM+StduG8LYt5rt0UIal
1lQ5k+7SGi2CZA8XjmI8h8KF9oHMR83dHTcETCRJAAtkNQaex9sWbvuc/clLbWlwEnETOTd2+IS7
BR4RjoKmtscl0sTvfD9b7orYYofiT3KEgfJl10opFEYZFIb8YdPpFFNzlksHqtetqMMQNBmg/LvX
GWk1TRws3/cWJc9XYAqRhpfUQHmqOvHDpoeXA+h5cORUMcVdHCVCTdmcnN/5h51r1IDaXRpdk3Ea
PsoBNYxP+xtyQaenBRNE1FoeH3+3N1BQhP6hcAuPbbpkHbaTUR5zKNjIQixhkPsUpU0MsUE+pwx9
K3PrmpcUMqy1DxkoSUsjLzU+Tfq0dRDW/l9ZN9KALQ0Eqf2EhO0rHnLhYHbl5C5IoVaMX1QGJXXO
yrMa9i/sSTWVH2uOcoSSLFyMpX9x4L53ff1STQGIBIMZoAGIEVzWDK3CWraMm8oI/mrCQC7MR8el
fLBbzYhnEgpmPW53Gcj/Tu931HIf7++zqk9+ADVvROUW+a2dgcyfvwomBkZ5SdbZbQiioWKKYL9y
GWgpt1S1rkRtbgvQTXyrEiSp9YdYtDo0vjRPEZOgOvilymyC9AwEhu4BJnFwHbdra0F+331CzkPW
g5dZB9N5WCK9qkcFBBF6PKX1RBbIh+1nNHLyROQ21jje0BAUjKEzzmRj1Oq5pP33i5JPJ6QO51xE
jOVJA/v02jW25SwRsUI0iyWKvuak/OzL8M0Pr4sXZaGsCtUyAuiSIuf9rChS635BUG0dgnUxUu9Q
JE3iWxQvGiL0i2DUZD5M0WRO7Rnknqd0/JWUB4FAXqqqQCjKakFrI7Nl85bh9TPltHJdOtJjVWY6
2eFDj66DfldrOhSaBc3Qkp0rkE+zrFSnAr5MXzW2xtZuL5s5OlcBcoevr04e1WGeK3qkE4HAr9/j
i0kHafM474Vsc0q8sOqjuZsfFPZjtbizsRDKp/FNzvnJrAj+TW+oT/t/jDfRY+Zt/lcZ47UT2Q8W
J8Jddn22wIJjyjqb80jCWfEkxFBGmpRCphh/LOMlJnVjNLIG8bx6jBxNA91EPfhcY/ZxHgH7Knfj
tcssqh+B/k/v6u9ruQp9JOLoYN2kC0th247B17qdXGuM/jO9K5YD1W4fovMsj0bc9bXVAMKfP4rD
PDN7CvOq0dzgkCFROg5BBL9p79OB7w8Ku9hlMLiH9TNrw8zciCC33XYql4kqEew0L1ANy6shC8p8
uHOSIiQD6TVElIeIsnQXUDPRm54B6VRqzRSV6EPd3fNrQghK8DLXiXEJ94aP1s6VtZs+p1/48Mvp
RF+8ioJwoQdj+Cc8WI43Nq/ZkJy8YWiphOZI+F8lK5IQcUeMnJhrPEhbKAWb3apHMQD4xRAfnAFz
7arR1RGgfxafOG6Pi5mKqWVHTumiCW4SsT7dXR/2uDPBwoS/pTxT/s6sp1zKjZknos/aAl8bQB1V
ePAoyxe8AbR2CeBMsyLZ2uqGMa97B+NDJXl139DpYHPO0oUWuuw8HXfU+Ub9TduSIPTVc2Nc3Xfl
XPMOYXG7O0tLqkusPTDhoOmOrWf9j1+Us84tNOWGcxRZU1tdrzfOOSCopNQHOLRVA+hI/H227p8w
Ay6H0CCnDnob2WYURLn7PFoTOA1gUkA44O5WRHgy2hh8AssuRm2HnacHvvDxo1EiqdFQKRof/nHD
3ewMRprsnAR78t4fH8OMAonPpDVQq5mFySsyOJP8qkFOR7JbRwfzCDDrqXWEEzEFXGT/4+DVXqOR
0HyBpD2kfVG7N/YeGVLi3tOzSd9RiH2UwDkackZ/moPmkTo30X+flq+0NpCCpsd49b+crbqjogxo
R52roUYNPcVfxEQ09FHbu5Nal0JQ620kkHiTI/hYrxnnn5ItXaYlDUmNcnMyDqXvFbIvcDCaZZqG
Fh8xGQmqZwCQYjnS6WWzJcRHe5SDbX1jm9MbGzqgIcMrPWYZoZHK/8nJcovDoRthYaQMoCKq8s0C
Ezk5C5OEzIMy8Kf2JTwQjPSN6ZK38ERvlICGwH+3xKGXpzLLum/8nJAJh3spErQFC9uJJnp4vujb
xmMCUiT5st+8fG8TMp/wJ79m5GlNlxqg6cMh5OdDejITqsqQD1jGvbjiQQMVYKCah8ZwBoT+cVxp
lEhukjsA3fPR/Ph+3CqS/pdjYkV+1l1QmcR07l/YwCTcijJFTbOgep2p4Po3/zGhB7GNWAiwYpCH
2eoXR0SUzXzbX+Q2wVSaJHXDMlnx6EvWa0baiqCn1rg5ZJjr4T6GPqpLvh9ADSG4ueYt+/87sGeG
jJJh98sr30kwQaSTcIvLqoCJOdAKgb02uCWQ50ji3CUBofYyhLoddOLnclza0j+o1PC0TjPJOfVG
iyoqa4wTZpJG7LCJossPNV1dobaVM+V1kpqAQuQmudoQ2QJz/Ugl6PAGPZHloSJ//UcXpM5bQTFq
jYJVOcHG6Ujr7K7yq2hXytpeOGtbmbK5LRn4FBGJLX7Ko0ImKDJ1h0Io/xrDjQRrFOCwL18b21Fx
96zVcs12t1KCDsb0IWfyXCoKqhlDHfvgJbeiYrhgc2zYMqoAdcIlXDNTGRQrFTN1MP6x3IReChPM
/Bb9MWDuRLhC5fU9G9M3IJoE78jrv2qklhPZteMdEANkxkfNWPxz1etH+ZlzBfJb0D+bBNFQUJ5J
77agy0peLdVWVvKhxaeN2Og8GsL4A4D98XUvsA43YYwzpCJMLIhPMFZkEGEtM04ptNVocJhzPe+j
GyrI9zgemAz8OnsDn3kipS2AdLXuzBPY46kKViFxEQq/I2Ae2iG1kvIBnqB/4jg4lSl9PI5NbtXh
VJcxf1JQxMlgNNAteFfnsq7JtfOJgBik0NE9zsBOJT8rN0TQY/9LZT6lOqHonTmJX383/LwW5Qpb
8ay9j8QdSrVXZ3t9mdQ0PRShd8DNZAFu7jZe4CwFNO2/FPQhQ+0bPl5IBCrTAEF08Oj8sTH98tUj
+1QAKwYNxH4vsli1wuo5VkEe5WcpIl6rwOKltyKqiiDM3giVke31iUv2DHkJPhTcte06vce3KgYE
DERxgLfM2435nqmkAguThDy+nP5qD0qIHSnz3lnZUhCjFSU6jXetcq83Ti0KEm84BTUmSOc1fCUM
kCs+EuWwf8t6wQvnjPXnP22no7hYw368BXFcT1afPz3aeBb2hRIviOE2ZVUzpjRFYPuqXgCl3gIL
BS3t3UYzSr2fOfJP1FBKpiEw7b2djFQ0v8WVQM9QefW5lQbwaMhSNdr6pcdgr30jqWnMdamtkKWG
PpbbbT96eDn1cv7ydBh9bznzEcjk6cSAgCzPEqQFIH45TLbpZ5Fu12cj1Kj7jqc5FlKKSym3MFbJ
BYVRPln9UYWY9+a75Pmo/xAcAFTqbARWr/ZlIs29sIhFIoSBzW5liC9dQ0BCJqQ6iCRmLi99uDEB
Q8OkSvzHMlfT+sKGchzYk2OD1KoUzlVuzxHD9dGpJoIL12jrDK+XQBrZsU6v+VQN0pD2qSsq5R+Y
PY7kWCCKB8nCribI9tVINeWnWVAjlolzqZycQdCTQbcNJjYjwdqhEfFnTXAgtFViY4vSmP38wqx/
Q7b9RRItrVKj/vrh5wIvmVpet60RdBwkI5ijxGUkZUVjwrZbtJWzwi9PRuLCV+tBwZw9i4e0tkT+
dgnAG1aU11K7VWMINGjbxWB3Kc8Ii3j3JKiA40w4Qc9CSkPrL9NFyjDs9DVwuZnbb+m+KJXxmxwS
KoZCImh6JVbBTGbXTsql4loAGZJy+sLydz9bz2R81Gx612Fg9qtI+QpcIs0D9bWvABMtzU+5wZXf
2cgT0BIRekSknqMOTCRW7X3y5L4n1S/HlCmzyIgG30ygIciKplStAJ8rAHoWIq5GRlay13WVqAXT
XQFqHLv34Tptb92yQ//j/bar6+zw3t/AETZDIJm/8JnvHlRtYXia/bsqp7hsqhd4BPKWd6B/UnaL
uN3i6XXv9qLdAyx3YdDiQ+21I0wPaZ9db+8QWa9u82z12Mg+9AUCYXyCurHHQhCgDX1cjYyVnnG6
lhenEg7ZtVRq8wMZRDeu9oXXyXR5Xu+NV4H9YVOsqfxGhCS4OGT10SLsM6mfwb5HcLOgQk6jecTe
nwmizmDAEtyb4u4mN0YFne2izHs/GYjUedEx17WG1v+Sskk1cc84rMwmdvNE513hA1vBoaKC6EvX
RAyck2EH6bfyqWgFMo+wJsl0JrmrMHIoB/d4V/H41mWIGRRykGXfdcRyJc2UXc4A+L6TcLpPoZSd
woTJpv4u5pquukESgLirHxsADvS1Mc/qCg7y8p5AbjDg8lhTADASWNDpfDFaoVMPGMdYSYJePnPl
5aO4l2bPdwGKnqVj2XzsD2br1/vzcYd5x9hBYpnY6d/wOT4a5R+sh7gjrkjMEN1JRewWsyxVO10e
9OEu51DhOxLL+vrTvqnXBsoG8FzOCbOxwWJi8/Vch5hgrnO6DWXOM9IHw2619LJ4ptOhybGexV8x
Wgv3Lqn9zaoeHJocpr3snRbqrgK4ZD5L6i9rWepzaGrzDsWBjsVWMPPQ6wR4qQ0toUYhgDri1ebZ
9k5vQlRf4EnvJ0iVU1wbs1sdoSfhggpka07pJOqLPn52iqeWxfWSi1vszWRVOOa8RqZypQ8F7A2S
QFZYpfWlLCCUJDn4IHnViGInKdE5LZZXqItTjkJFY0NhA4eYsMGgo5qETXT0XU0yyZLKs88HQvkF
lIhuMvj9Qio05GBauNjiiWGT/3hy9mK/CpKjRbskVT3kQgH9flIM1fhQbAV9CbgnJ4DgaLUBlcyp
eMueSsWbgky7+Nw69obiVYFonxKhPovRnXzKr/ub68cZtkllLYAothLzlrV9IU1vk3EVMT3pth/v
CaoTOx3tQL9+wN7HazIuFROVRhemWGrd/emcLrtXKohOTNwRoPnlLwgwiGzKfhY2Nql+LMMS5Oes
P1gQ74LKKOdfjTaar73xYapNVeIrE4fWPax6on5Elf+dKpwZA1A+0CpMDXP4hDA9Ek4s1opzX+/I
Trl9nZiGIWBvXqPO/AuqPOcaqKjUCteWqTejwvLsVmAIw/6JSGq0nhWnnxwnluzCdTAUF5idiWmE
NUgVE2/5zcH2xlVfMkrhR4H4xchNgYzIOXZ5RU+9wkasjBf+KtA2wXU8UjFClI7pFQIRNEGpcpc1
yuzzfrJHEl2r2YW/Vpe1kIk1yx0PIobQSXQaNYoTjkBPOl7slwfStWRo+gk6TGmtFZbb6Y7MTC/p
/0NP8JbJUUeWJVnCTRmR/xgsQgOwU0qTMxxlRv4MfJ18Ky7i1cpZeglyxEMxNUeLOvPZqZL85JYT
6FMsxivtgONB1AXEH9A/9TV7wITAQJGW7Vqiil83LAshoh5EkCQnbpzFkipx1FtL+7nUiS5ij0+R
fLPwTgvy/YNsIEQ1H92A5ebBMU9MxcpO0iQ5SjgKYSPKGo7kQnTBRilcCluuGTLbHQfYU05PrF2R
QJLNV9owwnikzM3ukXuVIxago7stleximIV3zDzSy91yuF/XAg5gnBOW/iFoHKIi1pC4HDM/XBue
vyyjzlgdsIqZIBS0yBgFLr6QxY0EPTLCts+AC0gTPW6oVevAfIMXJRqf/iXGwper33JwrvjeOPpj
HYTisUthPHA/nPFJWiU67wJ+VJ0vXc5XKienbMbK/v8HppNqzqXXzbkHIK1o+4qc5ahXuk0+8YLb
WWnxQBcHB5QeXdxEOnVUpgb//3yu4hhmAvmLzRO1cXmQdargjG8dkeloR4tFHKIk7ydzw04JF7JX
Ja8wCI1eUv+YPYP8cx9z4Q6LSsW7x98hh9EFcvMkqLxYTlEBeuMACCHH/2D8O5hNcSkF2HUm8aXG
VkrjxNpvhFKXayCW6J1mVHNrVu1M9O4vk4dG+prmn9D09SKqlEjxeLT9X9YxHboE0MNVKXmqwYgK
tbdsb4oK6wYPnKkW3SQxYtYIGqj9keY7xq8j9HmjCuGYwrY5qRC/z/LroYNPiIZBpVex/6sv3zgZ
jGs2MUZAZngUFnaRDHZ80nvHZonfm2tKu82E050ZtZNwHG0YwgXNh3EP01uOcShlpnzizNNf62Vm
Iw2XFTs09xVU3mUnzpHjr0Z+rPzKDj2l8ZvPf6b072E6lj9CzWDOdKZ+eX/Ek9u/GyWBX/DECCTx
FLpv/q4a+OiFAZtosyXvdV6bj5StG8JsFp+IbgPm6JGDosjIhjXma5gMtURDIY6m9mWewafeAgCp
nRUj/I0vDJTJtUS5coObIb2Ib/aREY+g1Tk2g8D2K7PlPlNRcpX/v3NHRz+9YM/3QXnamAugjBpu
DXHW12c40hedySg08V6Xw9Hk1Dtw0vOW4wUqgKNZY/QzhGhceSLMWKZzmNORzZMr07opUmyHjC9p
lpFBldyRwgbR9JgOA5gP2xF/2C9lZD2y4PxXRU4jNNXP91Rq1+sK7t5hBI0jZvYz5n1ycfVWslCj
e3W4TsyO7dLUXJZit/D8SbLLhIFnnymyAnJGWZ6fNXKAMyrrVbxY9llUKpDF7CGAip9jxiS0QsHp
uXTkuhypujFxa3BkiqvCohDDmJeDwzH7NjHwCq8igNiZcwFV5eiIgdBNnudhEb12R0vAR0/Zzby4
aCNTfv5rQk8Zb+JlUmv32yuotedb/QdYYOp533iK0WELCg3A7/iYPG7Z50W6aCecTFC7+AbNJzqA
dZK/DXOyLTF2szPHU4eIvq2oOUGY73oZYyvhCttI1cf4y3mTz1Ep1IB8msMKWcg/7MFVoAbCFx9m
VtEx6sGJqNNEgGAM5oY+6T83+CaWJTf+DxVfg699jx2DyCLWQv1dnqNzgQShbuOrcpIIP+Dw0iou
TpqgizqMHPv1t4j/Q5MTd6HkExMIJxJ2ub8QHvWutUUKeURQOvkMcEFhPOcQK+muiXf1ybKFm3LJ
GwiT/JwNr9QKlgjvw4bVGPbZAmnJ1WL8XjfbWTLbi28cav6V+UrgQ57QkCo3nmY5dDOb8ltajvCo
w1PK62V1+IF4kNExaqnqvnPMjVfhaEvP8Clj7foBjHNcT7v7Vmplck4T+H/2pbIceKt5GRTVwGje
3lKnka32veQjawnrcvKMd/RSGSjfcVBSGYtmdAunZPfj4jBPyE9CWqI+WNgFwE/ZLME3cX7ggjmM
BuzHhKuy/Du8fRz1B8jC1ZCcod9pZmmowM7dvv+c4v7OI+1sx4Y8ijjr2HlNVeys52dkckurOsTq
WR59giezfpMRN8OyI4j9TFnwXFj/bn2VohiaVtHr4cwsjs7m88mJA6Oz9fcv6wIsrO9Yc5TVynY2
tnCv7CyuEQWIBVDjO1avxrMRa/c0MXx/867z98u6Aal/z+vHTasfK+sUneVBpm2TNXh3QefK+Ygl
nA6z1138heh0PLXrGhfln7QnPsIYkxIUEA0LqeG09nJIlgUE9J5OYScxEohxfExhVx5kFZkdDTya
ShSalSNrGu9EYSQ5RtwdCHiLEjsAyR7lwfv3IlMOUb4I/mcxKv2dIjU37ZYgJxlXqf+RZ1IpR7QF
owYwPUVmC1iTeW1yIovjJbcciTN7Ks1uW36Zan3Grif9nhnOXFYoLG8jyfemyYyYvvOtM3aSlHNE
cIfk/qLTDqJ1bKbhXqket/MVbBo7Pd2AmgOr0G9N5ZofNcrbag9Em84RBrvYfDA8x8DxfBFK0Ux4
fyMERjI9uRxJycN6TmyhFh5W33dU/6MCL2GYDy+Ezsr28zw4U8Gh85Yl2o3BskgQmMBmU93cnhKf
GkNrxOoh7PKd8Bl6I4KfvEGkRyXVWXkaSaCeC35x0E8r2e7+aoXUIiks6nQHg1lPMoa+D6VH5plp
6QYGwF3nW293+HWLyyHnUS1hPaXY6HEYBIhvtc0kicE2RHLpT491VXrHE3SJgLVE7ltNaTBHCoND
2+9UMPRSjkzleeYk0ZDPZM/XiZnaxVvZQQZ8CMxu3kbgS2pJbIJhJjyb16ubHg4SdZUMbCthlo3a
CzjUAmd4+2CuuO4CF7WV2XRMu2VX55Y7rmvTnmQm3n5PZ4/2p8gBBajB2jCQS6dKwNTVHxEAEEVM
bnlHLQYlCBeqh8RvJp0QIlGiGXNhbZZqqQDOC2R5xqB1GpH/lNktsQjs7xVFHXO999iPor514hOy
jifgBS+2FqpNelRB3Cw4Pu1yZT7r9P253ks8N3GeQhtdGGq3TPUWJVP1AumS28OcIveDAXJBrIks
RpWMdcPt26emLE2VrsJy28TADf7ytb8Uquh42KzQ6QGx/N7tTWh2WVQsKL2/oJ8pPxfpl0uMtwwO
3I7hSg/md6BVUGL5rBYynfpELiDWIzz5Id8Jfhz4fQi8X33KD3OyKsFAchNraIZLLS+CuE3k7dv/
mLz8cHKDuYPFdBTHzzBtU414dL8vaTgzdmdY7EE/qot3SVbLWnKlRVakVWIBYVYG+4dBAhxGxYne
r8a8SBxVzfza7Q77zsA+NMEnLQQ2+d6pn9iGr+MxE7orXyzv+eF8VKpJZ9HB6PYm3MTxuhYcc3i7
6Nt/X1648wRDUAT+6UcnEisgXCGGr0s+CQaMNHKbSKL5mlhjlhozYYGiIffJn762zemGcP6ucaAT
YfguV61rVzNRzLXrpwEIkkewq3JdugcxU+hGHiJ5UI9sQ9zZ7mOPZp8KB2cRDEnFnoL2uSdRw8GR
L8sbRL2YBxa17CgrUotwCS6VWrS6tZH3I9TNE3KoT81y0yD5GPKTRXT/Gp78QyEH5wv1O3AnxqbY
ffQqp5spjQJKsRL7YIZUHNguvKT7IEfrbhoOTXXCJlWMnVYFJZZbpzP0UwaGVACNZiTiddDj8KPw
lVqhhEwCNZA/vO8keHgoZ63NQu3BuqwqRIndcrRDKUub+nyyhk2a/3GVVVR++lugr/YYzSNn6tFI
H2ibFZojSnLWfSkRpLUrIGpTREvNdnlT6Oyrobv1gXMhrIgeQLCjDFCuB95wF1LEnZC+PYwbjuuG
ckLQiKkon/Q8sCR9AY5uxbsr6cH5T+ws79mcz7TQ6zCd83XZ6GzUP4XE8D9RluGyH9c0Lq/jX4UR
BeWjgsrmgu1bhn1L8CpMn3upwrFB4ScftZ7BMsZruNVbvGmaujwurswKVtL3qkIFJAN72wWtf2fv
ObFppcpU5vKXiXcQkaIv3FJK5zDQDDYPCsqBrsP46SKLx2CGAM1GEqVrkxiLuP3FRJY7/wyTICJf
lqxT11IeQ9kGLuHf0HIOR6Pb0oaZB9Xzb9rZsrMGBtToiqMGChFvMtM/Ogu76Hk+fWS8VcSH+ZsC
jNMVk/bI/mEMJhX4pux5FLabWoODFBudPRbil/b8LPtMcJMIHtHwL1bDuZ+PuTJTQFMLcEJtCSWt
Ee55PekdQOeHmDr6NclMZx+COboCPoaDWyOuBGqFbC8kmmyok+MJdjSCJ1E0q1DO5vO6T4wcF4SP
r+5XAUHChBWGNnT4aZe2ufzSbYTcdi6rD1TRW11FyYyxY5u2Nc9PmhmAfr6lWcjumi55ezQpO7UW
6AtACSNSJ+lKAnENlHCmIlCKMN7W675A5Ng8IisBHhMem4Xf7FC9eJ+Hk78GBavs9Eoji9G/3g+o
5SjfWnNGuTlkPQjckBAO8h1LEU3U+nNn0/XV8ZQLPEqc2B6ysCdWNmiyQiQULgkxwR7svH3bYyB8
jZAc2zJyy0hoXW+vTETeQssKQw38LDQNqQCQB3xiObj2YuBdDOg+53WHXlojdjM5fhLcmLvJkvc+
XWFeoOlPc4D47ALlhN33XaN26y2jJSRKE3++p1whUZ1RCwQ3cvmatpeqVqyYUo0TumYiOkEgeZRp
I+qTSByZBxFdvGIOre68sXtAHTxIAbtnrUJsfms+ivCQHYkS90hpOhR36O63AKIMtkZAbz5OJHe6
qN47pZjlrR1E5nNRkhajsG+P+6veETekqcXdf5tKDBDuglgP+e/G0yMBhydlsHKLp6wksSJSneD8
7mjcqVIkEMEjJI81FFt3/HdJLagsly9egtyHOE4lNFCrfDfNdQthyM3qVv8pJOE1E931Luy4H9xn
b5KMdKJctXD62Bq3JD+DG2GmDeSEs4o1Pw3Zrp1+NtWl5QETV4hefHx5pX3c1j5P+RGRU3A/7eiT
JqSJMzykYUqdKDMxu7PKeIrYvB5Pz1YRNJB25MxEvDDQRK/KYA9TOImUF4wnFjPO7551aDO1cHIR
aIMz0+ePdiwz00efMiLRYTezkP8XNv1eKHeQT1emgvkjy+xIsaMmgeXQmw/9CzRtBoXStrV8bJz1
lDRQ4JlA4eCqTns3n4PYLqipYmPSWA/lozRe6lVRSkG8IynHM7sjVOfKN+AeiGTi3P/YeBlUr4Vu
xMnkT0sz3Uv3eoB77d4roTQee3ym8IArzMUmqSXIJK4EdH+w10cuZb7dtzB64Bz92OwJvNvxhxex
D5o9g0eHquH9frHTec61VN8MkqVnu7+3efVnYkx4yFkHdIe4qqh0b7/Tlj1zAYBnoqkqQnD6/6Y7
pTsy6zCRAiotPwP44BhCU1d0ToD75/LdCD8JsMD4N4FykUNbx19Ouz4pvKGo0EvcHNFrLKqT1Ads
2sTXTkNaPtVbj9w7IYn0OcouQzCUfYuq+KMzKD8vm53APd6QmcXWWaRi7nyEFKvmZoMAwNnrzMsn
dBYRmrZQ/zT4j2Ah2Qk899I1rAveX9urNFakRUgkO+DEDA7++4l6HAnDzS8yMyRB7kCRqrcVixk/
3jMjo/c9RA6mdqhJuHQpy7OPfpJnlBDWOr/3niO+rOpaV2LELW0wwHEOS/CV04Od+2+s67nJ6lxo
R6sKcla72+ZoXGA3H3CZW8dZ6vVN/vXtXyoaq0joyG8xRpD8o+wBDuUXk5MHlh4UQLGvB715a0Tl
02BIWlfou02bUJpcl7y/lL7nvLzW3A55EPtIVlTTlu28FmPp0c2DEr7PatfuMopioIEXWu2X+S1+
qPqWJ685FpbuNeXB/SAw2/8nK4pCDG9Dg0v6rpk6HiK68C2Mp0EdOpz2ngoxncdEiet+qy41YpTB
Lb3Ftci5U9V3w1B/mHVSfRjiqqVSI8wbNSXajigvqH/+bf2xmMtIZg1U/pOu4x9zu2PVh9GpeTyo
vwzONBQ9BtC6+GX00XraC/3gQ0Ntb2XWTRiJx5XnBAIjgZgWwRKSSP7sbTzPZPIPHApjb2HYbjxb
tD1MXlGDk8wvlZkEYuvVEa6OrO2H21UQ1eYA3BVK+NR6zx2CkJ2B6/pD0nitvPNjRewFTrW92/Dg
wYd8i7E84wbJd/zTaZTwLlK0GJbo4sOn41EaZAn6axvkl8NSJFybWBxP3r/Y11kfWP7xpFB8KLeX
GdJdiu5NYjHnlV42KkoEZCJBtkcTNnGa701viM89+P2AtT+Y78nIIFhUT44aWiUfsiOhfJebFxVA
j1CWZ1fBl8EDdSUkhIlEvPu4Z18PqeUqHm84WTeqQ/uHPm3Xo3ndmw1vEyfCecGBza2InfQLaVPF
FyYW2eAurDWtDyV5ENd29jqAVhArevDPD136yd5i89R+C6t0Ly6mA5Tk7rvhkbJSnZePZicYxtyY
hv69wOZLnDFkmRnTzcRFu27+G71hRe1IaVZ6M1AyQKLLlASm2jN5ssN7BQCb/VGQrJT6fow9wGeO
qAnPOniv6zlzGWIbxLYy8GkgGb0B2pavOUp92DRXCHAeL075NwL1SH/xC5P6jER57nB+Sq0jtjfO
/f7K4ukmMj3WpFYyyy+WHqVgUVXbBZFQXGA+tbS3v7eaVAnH/dccd+7rH1MMoT7LODFIYpMz9j8d
lcpx3n3SO0FOzdgWeVwfx4IXHu9huT/87wtEiSuOGhf/kCRCO718BeKc+Q9V1dv3SCPXp94EbO87
syzRDiCSFb2BMYicfUh1pFtUCxNQO0Bk8UHGeGN2VVZY/c3r87esORWKAEAqnQJJt3l5ut+SI75F
2zQCrZ7IoiQdZNfPVP/IY433l+fmfJ8dJD4A52DCq2owX5AzsqB7jXf0GxR/N/X/AHXy8bNfrJ/K
904/7I4/ib8jG6TqIYFOZWpQeFXPKgX63I3xq8TEFgyQz4k3TlFekRuUjdPtT/dy1gVxG8A0D9PH
0UucxLPqQlk72aLpR7yBsgksgg6zj5RBwhCLyyZWq7P7XZf9nsKf5FjcchSX7pl8dLyIfRbvlJCR
iTvd2vAzY7FBb2Byiw9bp7isJW1j9b/7ffA0ufjIvB584S7l/qeyAVL5ht5MjnTnZVmjWGYwHdU5
nCr/FFtKGwV1H6Yi9H1rUSa7nNywBgpEBcwNMvwhXeBEZTTwt1S0TThWHS/nivOrEeCIiB5l93ML
C3LZsQBwB1O1vkOEoPHDic/xK6t50u+dNS1KwyK7I/cvTNhFij+sayWWRdt/sYwJmG90Rik4kpYE
AC1s+FgrVeOopQfvhmS0FrwRovHYj5pFWtXGmpKTcOOYd2NILhomzJ+BbFDpcu7GrtB3Yhb5csUa
VGzYNEc7lZqI7kD85Y9BGNNpxp5CCIIC/ePBHOXEjKMrZ3lI0Cx0T9WBl60VDC1aTRjLG8ofbPL2
YpVLBBv1vOBYEIPPNNL6KYnmyhfy/n1iGqS3oizhVZffhcRuUcwo0qV0X4f0eDBVJorlxvWm2Y88
kVXpPSoYCZ75KIyrmxVh2hv64xEqym3ds+vhI5+lpCwpZBuFLGke3FZbW+Y0sy9KkVDFr2d6dKkh
2J2U0wQTZJGbzshX5BygQm4maWywKtBmCK/bNJKCPHNxmSG6C/LBePx5/3Risrzpqoqfjsg+l/qk
vM+12OLgwL9oAlmeftrK6sRS3zxWpVdGi+MmeI1rAYXqmdcq8fe3DHQXv4VCw1Te/tLnCUEDgrUK
wIvw+zqrK+hBqe880BdFveFzUbBH1eqTAO2SUACywIdsGKRA7tMrVnlzXriFban/obSxcP6q7tUd
OhVgBUemXIm83PIT+bf5fQoOPsKX3vp8MJEiwe73vKhOryp02KLcwvs9mKBR7+B9hxglcUvBzuty
OW21TjqagiO+395oi5lZqQPAq70xhTxmmw0gDwxV0NdKkpaCar3zaqbHS+ObINkWsH3y1e7PF/xU
iqVdvB/jV4fsF/JnapHhtJVXxcbY1XQUtE36+YIlcPxU0jZ0+ineR91XRxDd2mpoT6XEwLt7ncHF
Yno4pZo6LQn1IAg1eDLqI/sMP58hkbl+T0Qpm9NSBkv07QKRdcaFD1DecEtGAqYPURIMBQ3JDJtf
/cu8f6/E2uWLI1lifsZzASjeOATNbSif7yNvXH3HBUR1ETtcS3gIrVUa693Kwg0xDMPi5vzzwEFv
dNir+qpRXhLDameDB1uRH38uYnXNIWdB6e0Vu9q3J+EzxkZrasSZlL4PpfQagKY1e6TuTgRttx//
FBAOldHjfYiFTN+9NPs3wMJilv1GuFEDr7xTILw+8bHSFIEAySRMJRtT0JMyRE4NY7cxGrcxcjs5
UP0hfgKlYUQs/Js3OnagwZz6kcGTDuI4lFvyW0x6ZpOC7P9aFtOWwImmMjaAHzWAZFBxYTtARZ7Y
LK44NbdJAN6RJ3fP7YqWGSl3YC04S/Hcv8DxFjYVd7gC29WisykYsLiKkMWr9/C4zJpFZpdtuGv5
n07cRtpDYF9Cseknkh/UMhboki0La0NjYf/yiQKBUY+VBFR3gQUBcHMRaIon/DYWmj15Q4yncv6J
mU2ffLtxpy7nepO3s/wF9wzl3rg4HG7gO5tM5UxlpAUvhbHeQzMJ/+vH4KEwh837HD//+7mkfT8n
F8D4Q3qOVc11KDiaARnpKQ0MA8PX3CWFMxLeErQHIi10D65EZ8qGmk+qn+C/0ikCAomrwMU+e/N/
woZ3VItYKcEm4t7Za7i24zZZkueoEBY7j0ygXCRPHEY0Hd9LEhLrvyclSTKvMk/1AtY6bjwC5i29
DVOaacmhLBXvso1JcaVOezg69R8kHr+69Yg7bwkPORtB/8Z5qdAaK5GtHymXJ/gZ+NSmZuYbPWYC
go/dAX74WRAXTAEFkNR7hXV3sHP1B+o8ke6QQ3OiFeyskeB/3Db1r0UD759EG18091G7zGAq9QD5
WwgwWt8r6RMF/trexdjJ91mQvDyo/k7ONrcyn4JAKULxmbkbKwPvnCoD5mT77PjLOOAMkUYQ+B57
OGhDpsicDls6qD7Rc8KdZuqcMFoaHS94oXVZaBPxDd96OLlROZFuAtj3QEclQdPB6DmkgiJBhCsi
HHNFMSFXewGwUMQp/ED7Ftprq0htN2/Qsp4TyES0yg1sihK2Wi6gEH2iEEIyrIlDyv8OJKEkcO1c
SJfuhlUaKaPTx+sRNrQlH2jt87bkXgUdCO6E1izFjss0GRF09X0F2HOeheoB8bVGu1DKIWNVeczA
ab/bFbJhdqX1gErXbTU7bsdtGuSvfe9zBEBDVaORiLU0MOMFsYSxzyYIoNVPnVeuAsQCBqOoWUKN
dqrqXR4/T5jdr20o3YiaFf8sSu9o9jUeGrIJ6RwklZY9Y9j1NgsBx8PvYyGDkjE8Tp9vCr3p3JYY
T54nriICRqbs1Es8vxSBVyMQu/4kUTEJRQ8zV76zdpgdZmh8GzjNH+KsIP1n3M9Zz3ZK4mwtE3Sd
7x73MupSZjaJv06AgzK4iobjBodUE1nDE+DVf3RHv38XlKRIN2z7xTOCL1M7hlH9N/ZrTKcpWM0+
SlFPda+KNILNZz274ywkzIZCVR0GVhsxZrq5FUzVthhpQZ5wsyN5Akx+NV2kmki02Dw0Dac6peAM
3hmk0V9NXkoWqUX225cYJOAzthp4R1mDur1RVy2ELSJohBiySLBoFQqK/Um1ufboWTa3ZX+CSN4E
7oseRjSVU14wK0bQujvQIWE0ya+3cLCKXmlm5jzVR2VxrUiGfwVW0XR3JjUSay7kr/R20IZN8Qwa
XFhI9Z0DZLgIQY7GSRW3klno5ffMmgn29LslmLNxx2h576NzC0B0yncyhGqcCLZD6iMbhnqJtdCq
k6wXEIAs8sKdTdFtzh9g+C6b9RNf/ecguHfMFTTCGHGHotdEz/ekpQmq+59z92lKjm0W8Lmt7EF6
gvzgY+LHOTHwXFSCxVNwDwsb6PiniKtgVrpFBK0Kls+vnU+3Cz6jYX9IR4c0hrpIh52QdHofZ2pI
h/Yrubt3waA4wgxztMBz8IMMd0G7B1d1LcNe49nfWfMQ7gIGuRx4n6X/aZgrFpWoXAwHVtcsQy5a
GihKJ0YzjC1L3i67ARhNEMZgoiXv9ieUOmyh/85d9MMNxjPuNYJc4msilhGyo4Nnk6OJ8B4YV97b
eW/QHkliL4sqmDE5gdRAjadfQV06BFhCyJGAiw0phiYSD0Gd8bXnHnww7LK4GWsMan3IbQFDX7Rs
8e9kVz452wgFWcsvOiQRir2mZ/hWflMIXEOnbJJ3nbXkG+v1ydtRNbz85Q1UQez/DDWueYttEbyR
XOHFkOUrV0jvZoWUqiIwok3B+21GjATJ5ihhNwioIaU1zzv1TGOOWFH6szZLDqzFbbjtT0QEKhUR
SQmv0bDbOE/9iVoYSxD/rdv2F6+53PNRS5JKnwCAo4UJIIyXdKHfU+wldHHpsDJex8L/9dzasA32
GvsE3mKE7IYjwcgOjpHG6/WeMA2dmNtFESUVRIq3GKedsLv9v2khEZghfRvF1PP7j1/UzF4Xoj5v
WzhWvW7mEnBqqVwxDT18eHj7hmIonrw5w+Zh+wAYYLyCh/ooGCscziAUMzIimsU2gCkazPmIc6Vm
CBU6bvW4NTFY5StlTqcbh7uhcMvkdZV7MLpozvU9mpa6rFqVf5zB1Qxb3t5HSOOTg0Ob3vMGuEYj
lIV1Q8A1kfzAxfRXGsLQ6WK07B/fDwNt83bGtGGHFixRIEtlLIEt8z3/fK6/cAQLJ/PuQhsR981v
1pUFCmiM46o4I9P0R5WpXRD01B6cGu9tB7w9hfnsDVFGfOIUvE2zuuS+wrwO6ZkqTv3yu9ZEv981
EDDCiuxnIJhgn1cGKunel8RQRqHFkPC9+HlhY3v+qzryGTL192lQB0jSoKK4S5ShPNXXuiwoFXAj
IOLxBJDyf6BcnWosPV/JZF6Fj9iF2EoTp9gaycFtYa1FcBOpc3OWsGM44Z8dxWgBaE6yj2ky+EWe
t5BdnLEjm+r52o2nbRDcNsKrB1OVKrxsPzcEGoeG0W6unuAXHurcUNRx8kKtFkcmfvsHlNLzmjb1
f521UvchPqzB5OSOJcU2Jw/8zcohR3bYaKnxSC9VlSfCXJErrG8F3YCmVwwjcgAAisNBHY7CdKAu
g3qnIZ90WZml+w2NF3XbsWQ5UAv7J2KqY4t/FXBdKOt4ZCkco7F9Ej4VFEIr9UN6BJIHtZXm/UDP
rIw8oxrsabB8hQZrilTprHcJul120yltf/MHmwAqrTR8B1blIlPgFTw8JcBd4MFZutbCfA/RycEi
VZQB4QbGuWjjesWUMS+SjRfnJcgcDSgv4TTKeEOK8FMH+3rENhScKSbwHA+Yqy8zYvCL4YU5wgGw
JCIie4DcRylEiz8xH+qUCv20sLHMjcq8BHMu0Eci8iPRecG/30bh7VztzWQS2NI2Bn89LwDofMeQ
9qjntFNm/crk2JDSeFVJudTgkyq8+qHplc2nUbWBEQKGOSQp6qJP7HZ/62DZjcgAp3BDXpl8RNXW
VCgm0PjevLW2O8IxLXymXEGCp+RTWge2noqX0oRjiCbFzdeBZfovqeepWedAqVEbrHWRXcihHMha
KsBU1BumBBbxE+1QiED3O9GKzBrgPySWVuceTOdCnb7iRiNWt+3OThvX8ioVxusn0tgq9MvhoxUw
ynUqzlyIxNzcmcnGzeXMeOrB/Qd0eAhaHIazCZ0r2L6DKnq8ly5YHGGXikGfOVkikM89DIUwf7tP
tClzIDfqhq7JN8w47wScbQIiCueMkCZMgKE5HyrPO7Q1AyLXKdbHpURF/iPol1/2CLzNRO74Bt6e
tbTYlohDBTLKK6rEABlafdQZqj1EqJhVyApkSHo+eKA7pKVIGbI4jdjN9p6fJEpgd/cIca22BU8p
q6S7zzvFm0iz4OtdWh3suswa9ukKboYMblwtwIcb0FkzDcCCFWimYI8hufNU7XNV7oT+dfhQSR7v
3oolF7HBMDkOoAwPLdzDU8p0ICILwfSnzq67HZQeqX4uDyQbcsrnR3mExQh8wHBxMKs7X3IjUMzr
zdmP9zlD2h+13Q339qvfFwQpwGZqsWOe9SHLzEHQKFEbfVEbVtwgVjVYeuJY5w+vKJlzzJb/gngg
gUnFzfRuxyXWerzJc6sSrXZhhF1cD1NlnzdjBnFOppCXYivxwpKbW/iRSuxSB8KP8P7RlIb1UeXF
tDWiX2v2K+Zi/ZbueuDv/HXU5KB2XTLLqY2YPvQjjY5BxIQ1LcUvhf9LmgdQWxL+Ld7ODQaAoFGU
Uvs1hj1WnuI3QudJKJ4LMVoUCQacCdZGekr3NRcl3X2cMoKaHdSjpHzezaLW5EIF6HBWCjWjh/xT
4voxpz76eVlAbF15a02ofjLMefSbi8kWg9+j7rSXYhOuzL3nH3cHl7i295AYRreh5+nqEmP7CdUt
ZMV0wwIzLvKzu7Ot1K+W3xN9uOv67t+tt366qO07BQAzJ5aDEf1+BRzV4c24B3W8aewHjIeeZ2Ac
1E/D0JQj+SPArtHB0vyWAmxMhzdR/QOPqEMn08aprvH4zCEeDw6WR8pKupVnZN2BuH3KBZIXWPfs
fwo6/Cx/sdnguAoPwz8MnOXa3g8QI1yaN0ZVQ16iP/URAZJYno/+uPdtUazi7yuSx8PClynx2sIr
OYaiTQCY1P12wAMbrWY4hdreiBFIVbdsA0lnyFcA4dt4obF+8n5qFdmaX6PXOySZWWvEQWV3xkX0
P/wKLvsv/5NAjFelcZrdyIcQIBQA/+ml7CiFjQnLqu4uq3eUEs9PY1+TVZX+Zb/K9bHcgqfarV6r
TnsqQqR0Fj3Fldw1g/ZrXR2Gv8O4+X/kcdfwaGY2OGIiB+xcNzr40EiOuj3PRAnM3mYdy2juXyQk
/ljcwRmsd0bzHKBtlw+7RiDroK/b/5EKxHq1wJKI/W31vy1y92jW7f+3aYkI8Vub4ANWJ+JkRYzi
FxA6g1mRpxMUoykv8mthD/S9bJ35J+jqSUdPwbWXfD7wdn6xjsRGJ6fbjw66XyruGgkCt8SAUSuB
oVOBkRy+OoidUiLvtfBLciKFCubC0+YHz+D1hNAL75pG3YoFag5BL024ZZSbVNN3WabOa//iBEik
cw8OLgqFtLhoTBhw91r+nXgljsO8apyzts617VE0BWkyfucOsmdkecMun1R4MQBBRA5KnYdCB8IY
0fZaTOH0sLW+CjI0DbViaYPd5ml+ZMBh/jTru0PtcI9mC5Nms2RJF9jGpunII5hiIjoMVIcqttkP
eMHT0jMMfDc2LzAH8/S5PK/npdeI//8b6oGI+cvh0z8E+9pwIlR+LoxuCvzVkbuH8uqV+RbrqG+/
noVVD1PP5maNvTYlqfizY/KdaLBZM0NTEY4qlTD57iSDaS35Hmrh0J6Y2aY/3G+ofOKFLjy/QE0F
vxsvwiT7TW7kfE5kcH+74SzhyRpiEQRf7Pp5TCZEuoQ8L9Xk/ucIS2A7zGlrmi0OYYNX1KmG6Axw
pnObe5Gth1bnUH2siChlIsWZATysE6QaqAO2U5oIqAC++LAdcJux3w4bwEm7n8d+eCVA5g3BLaAt
A2Q1rEBhX7mEkdgD/0Xe5Is1MvBDJ8qUnpVy7sGIJwJnLNCcTe3pxFIH61VXjQSMeOVW88SKjgqC
Iq8Yc6xhngQB4FsY7cJ0/XVwo3TG4duj1yHoRFGWHbsd9hRpVNRG1TmOQ8+hULhqL3Tpgxoghkyr
sMmLJ0TnNmXXfyhLk1ZR89CUXMa4o5tuAXBhgERdfkqAdSp7TJEilFm1JO1QraoOsYL/xth9Zyrg
heNdArQ8QmmX6Qa7vLvfQr+zYHIxj9yhyqNA7aZrvh4/G8wK0BI9JlNytCDZAkAj/zDBOhmSLYN2
m4i5+LwUN1f23O9mUUVRRHhqIB1u8k9zQ6PLh7TdKLQtUxOZwnPpX3FIxcXKt/QEhMGkheC6erw+
XYA/Kxal9hCgBKGSvNoS5IrotP3Q5HCYM/HcpbzUSIg3FHJPrypR/9jTvjW162qLd4LUJwfZ/GrY
Wlkbfzx7lpnFOeqJaSnsGT30TD65hZxkrpr7x0XlICw7ISxyExup2Wgrw8L6fgMVrt+U/RWOO80E
mlUka+zkHt1qwfEYKQbLrB/bCzffiTNmK+nXJjQdUv8TnZ8wW6808pHa1GepQkkA5bVE9mvsqT+n
vZh2nKaSbCbniLWbnoauMjmRk7bvx5HFLYXWhAKSelPZUlr0oELszaE0bS6TFwqKSJdLHGCFNzPO
Y8wu8wLmQKibyjbrC64L3VfzV4Q7knBEILwOMyjJWBdgrwwwoE5tB2IgZ8HGi+aVXLDfGo4Ohrsq
ORahhVnA8m2Na23a7AjjbIslWgie4XhE0C6unCpnznJ8RYFVgNNSJwV9X0RgCNzGs4TA4L0xA6nT
jc9Kg0K1useK3Xa0UKCv906axgJWXH+PGduuPJhs3A39K9STiSzhYSpcsjsEU1KbHXByWjH8JsJg
TKInIuq5oIepowEACNDuaWDBdND1ScNxn50w+s1CRjfdC0Ma4FH08i7FGpMepARUJa1ZBh8ly1dZ
oFXSeJWGEYp+O5ma7s7rzCGkvnpZ5hZloenooGgTfM6g3CR4Y4WgDqowJ6JPZ1NJfZ9V/iOP0I3x
s1cY5UjnNlwIF2Q9q/iWXjB07eBH3ATkjtKxLCm3IfnZ/zBmwNnilPeMh8bak5j6rrG7bo+uwtOJ
QfyIG8c8/SDGEjEJQ7J+ulj7hMdRnBnXF8A3/uMy+C0v9mDfBBCz1TrXq2O+YveQnQYnoEEvj5gz
BDzr7s8J4X5uzzQBKciwqeWqLhVevW2ye5W2TeTRSgcx2Vt4M3mNstnwp/iXeX2/aNpljePLbSeq
tX9WV17UjvJb6Ry0eD2bUByH3qO8SlDN8FCEIRgqLnKt/f2D64ZL2bq/nYII+A6zebQJ++PXXEjV
blRXax09fBKr7MX1iA0vkWKMGtrSI4GYhNegAs6xUineemY/rBHAaHIVir4IjAD8V/+R4HWZOgdS
+54dtfHvZUVPa1/G4wArSWDRDmiERMu/RdqKjORs33zVr4Xt3uzXWN/qSsrUa+okS7TXILsXJIIr
Ss8+1mQZ8rUAp06rVdMXTg2c27nsvFynw5w5ju1PgknmVUrFlsTFa8DoU5FZRHZIJ/MpniXD6t5S
n+z+GMDM5nzVMDQf2TocB0tOT8NxR7069X4mmW1i4PoOcg+SCk4hOHm9j1uI9McoOB6ACUdQJhns
U76atcFTBxGe7bSa/EB9pDvn/B+tpW+iFdbAiq9++Bnjmm2f/nL9OV3spg5Tjd8PB49lHX5C7PrE
JvZdpsXvBc5SDiMPwbXfPPWGqqTJUau9Fn8wtTKv977iq7XtXB6xnBhHCiC4v3Fr42QXbdLtas4h
5F+jYJ4nbV+p0AWNq77KWe695VyGBv7E4uDeVMvcRFogZYv3+qZ4IlwCAKdD09KEUniz23WNH+Jw
k+596dMeGKhO2pZQL1GaPqg2s7zRBKN6VRiGf2LE/sPkgi6DpKdqNNmNbANiZPkIdh+dfA9b1+az
pYFR2PTXSfEJMzxmhePLKgFu7e1QfRu/fozlsihyyMXF71Y2ehblxdqaX2acPD+VQxo5iJETbZsL
iaHWSkfdreM+lHILTHBw+rLyiFcnJTSy0lYmAWFGxFH9dqeLzRlhTk+P0hQt6RxrR+S6h29wkDqO
+emOf4w/60MBFB1Ufa9l7Yx2053VVi9PFy9WbR9CKVRCvd/qp1RA6eA+z223f+ct4zbdqQ8m0DzS
CxPR2MlcpvSj9nI8V9e7MgE2/8U+QVDLn1Yun0tIqTKhYP2HhekU0Ac5mjcv5Rw33Kqyxtpx8TZ6
PscakG4wTvkJGUFpHW2UWArVrqIE/oiF4LlP2ENml/JXuXijCfpoXk42hYsDRx3Qqz8lJIfRLPXU
wxuqCS9YtZwLlspgG2XJ5RQvG66JYVuWqu7n4M9hI46aDFKAOM6X7QHfw5daR2d09nO4a/kSW5FW
QQhbhxfgYlsQkJFsUAtInrnJpxiwmP+9PRJdcQQJsu7LboKFQEJQmf0PMdgvOBE/rsnD6+/2zjvE
lFDcWvUp4JuCDGsmpitddOn5HLodNaXSIRVFpVQQi31OdQZsVLfN7n7duF6C49iqHBFsF3+dlcS3
Sd5xLs3Z37Uux+/jTmRL/ueEnfab4Uy1lvOtdD1yxar9ZMPISqTcSf4vzPgr3zcrYRF1pFDAQSmB
41ZcJlqvU7dpbiUx9raBANN8V60TSaMc/EWQYs5956mHyC/OnrYmovvBQ7WTwVlAoSiE2bxef+6F
8Nugp1IP5PwxvNSMOtdqveNb3/WhqR0dNcJ6cLDBMu/CsUKtU5CJaxMOjs3HpnOofkD2x1fPQ0dQ
5xMRTCb7Mt2vd77OZy3hlZBWDyK1W2LeDnXiB6w6w3te4rxoPJ37c1k/K0mc7/vXt4i2s3sNLftJ
ybJHSJkYF8rBW4xJc9K7IjrXz6H9i4/6x6qh1UnLlZINOhySia+tOa2qWWSIYlcAfqyAlBvPjWZH
N9jTq4ZZgsnIpJvpucEjdLp69uTQk8FUPQWf0PpvWyp6n7rjsIkD3meDfCp/aTjTn9n6RRFc7h0n
cgiOU9IbQ7+YRjVc0BClH9KrBvDDpz3jadZciMCp5VCZM7d7+DJc618ZVL9mGsgF6Bir0xErLKsE
vKDA6WneiRn0LbXE3QM+8nnewfVVjmtllHXVWPGknR4NYQvmYELTJzs2S6n1dKnzUn9H/bYjXpcc
JTvTCFcSQjWgw9jDU5lp14HJd+1KIBB4bNSCKPYpv76leVkGdTzN5fFRcxytJm/Mmrs5aj0oimeq
3byMBtg/2vqWcIHUoKhep9XtggytnJpWjAlHpFDCrnw7sk6GD6eOIG+EvWZXXiyj1zWiQTjapBcZ
mmFo28Uu3AHno/ZHFWqpH/T6lGOJCiT01ST+TO8AmMXAWivpE3YUXbnMUvKNjWLd3aQQfPl26FmM
oDA/lfWwZTzX9v+g8wHwEnG5o5FW4RfuXm7RU3oljSkFNWTkdE++7KZSS33j7TtZvZXzmnlApIgr
9PyUsgMliB63dM8J0LFV+t4HR2E1e9PHti+msdsbOu/ubNQJ64ehKMe6DuXzu0eBrf7HDCHfmUSx
yVttD6GrIpWUrKytBfpuOqp9Loa0s/9Kbhc+gI9kPOb63703mF5/6cbgBORXO4NP4e5i/sdik75N
NfV80Ixvz10BajxUVlSKYwgnVh9x4zuiNGukwROS8/udex5HCzhgO9Ap7taCBhEYmpBs3lu3eGM6
NqT5EPiiu4prCPMyf27u3MjTG6hTc78V7eUEerhSe3Qy8epuo/ARV1tKFrdv6mJiDBwKDENT2fN4
f9kKwtHX/EqIXWrRVcRO75t7A/J08Tvzkpp5N8edvOpuzzOE19/4elI244GbnS2aC6G7M5UMwMgG
rJ/EKq4OW0IJ5pNet56yhUKoH/TcIGb5UDcRvj7PKoGe8nvf0tE9oiycVS32GwjkBlC7q6qmWd7j
e23rgST0O8JFHq/xQLbTjl+tDn5OsQogCjDB034DSV7ginlAnWALxtGLSH1ZpbHBsG5prMT18fdH
Wb7oFtocmbrccXIGTtTYGnTOO2aW3yrs1amo7Yu8WPw8TqPqBwGAE5ZM+2jPtr1Q93vdAJNiqNoe
eGxfX0rE9yFZpS4h1xBLV6MfNqTWzCpwZrUGETLnT2sre7w52FkKuCNsoUBObfYOtltA2NuGzJJm
xNY0uBk/g49scm3xi1Hw+/ZDLetaC5aBn1nQyFBALbUsGb/0YFynDhXQuzdV6VGB8hTfOVsnATUw
KQCqDY8ofEOADpyc+N1i33FA/VLHubgEaAWWcIngb0A4qVLuZlRQUs9zki+KQSnJEx6GkheZQz4C
0dRJ4r/1kyuzjB8RZN2XCP2qyYBIWj2Elum0t58Vd9gjeH6kHRzNStu+soJU8RNwu3hQgQrsSaqg
Z3FSwvKt9j+KQAwNFYbrIev/ANhpZa6tvOgnQHxzNtQNjR/bMcmbX2qFRkNdCIYDytdcrB+SQVwr
R1OF88lNNWMmEudz2lfW3ul9CZIuR/WJurku30EnHynn0FuNqBIskdt81IRo/g6sPyGm6/NlDlWp
Ovp4VA6Ysk8MZTz0ftpB8uDZ6Zp5rAdEds/9ltz15etr8xIIM3YMU/VLqWVKCvEwZSx5sb1dXzWh
BcB7GUR1pVVBWxEBvx7bEvJlQahUXp8p9vS3Z3HIpAkHRrXt4oku5miCt/SeG0jIaislPm4L2ppE
LMPusOzTEcTxsKw7OeWhxgIHgUNkelT5ZZdt6yhAxwqoHwrwvVky96E6LHu6aZUKvXoM10bgLJIO
otJxw/3gSOsXXCGkHwYXVSWLrGlVrB3farbXQh8/9ducYY//0sbYYOvSN2HmCowxLMHLUhGzWy0A
SSBS2JaQbM2R+u8u7KQZADfVhyrhVmDLSU2EJ2UgOp5CvE3R5st1UvxMo+qr1ziuJZS6tre14SxA
V8eBddgQrdzXe2KrvINcFKTJm5PQFb0Qmfl67UjsjnszGDcBvDXPaEO3xpYtB/CpAOmIDgMo56rq
ZQaLnfoQBRp/pCbUcj+zAseuIEatFvEYxF81a3hOCztlAGrZsZcJFcECri3XgGbZz2FSz/Mb7ixN
yqZS/URShsc/1Jb6fSO4UOjJkxZCszpW4u4OTbvDB8h+Ups5ia0vujYRE1BFQ6BM/cRZZs/xSb9M
FncN4D8xJz/4fEeJBFb6DAfyPbfKd+Py6xqVyRSqW6LP5IylKsLyw4xlApKvz4NWesB0utZzdbCo
goLcEji4ZrP716oL4H7mMtqXbOJrT7u4++rsbQwzRKaLB7+b+sJCsc+Oz7phq8ZS71pksnFvjJmj
/Lq+p5IzmjbxjjDxzUQr+Ffuu4vhO9ZWbmrPE7tL51PAaCqT916bz4OWNfCIvXpRMq/N3mCd0/V4
nVYFwblrQgegoSJYW5POWG7konLLDULcncqkGUivvSKQxUFBanu6N/2BAF/eNFKaxXZI22APjnNU
8uLeTLoEfqsqEcYg+YbuRISJaVhIL0oufZ6VP7xVUvqN/08zxcDnEWVeXeCP+sbE7hz+bv1NlGGc
qQ16kGZ1zXpP8yOrjBS5jfsiFWiLdJX6RAV1jfIcz4Sl01uhwjOp9CIdaTuvdCcwmu06JDtQwSJt
CCcqSE7OaeRhH5sMLSApfvtxHDDMslc86LOZ8cw13k1OJH069YCTvtEjxzybjIzOjtDi5L5OnG40
FpgfY6BODfST6rvgHwF38VVlzEFOHqN6pIfGAeGHZFcgCoNc82D/LSNHNX2QMOF1vrnKtpE1AIDa
mlvyC+tmpCgq30BoI0W6SMxFZlgGjjyz6U0/kGKURIuBx7yYYxyGTBnoW2DWYTKo1BHwy6JWlJrC
kYjN3XYDm3yc6AruAdKlRBQeiZiOwmEzf2C9dvUhYRPhUDeSoHImy6jNVdBqd1Us6b4TGbHJplo+
FOKXn9WpLaFodM0xbaQHsUt0Hq4WHZMRhSX/VUoGUfjpa3d4uDZ+yKtQO/cK3OoR9ihenuZE3FMl
ggbRjW8iesuNBFhdKHBlKTJowLdgpvNm5m9aT/5XOgf8jOqQBSSBdbpeGG0dQoNpz6LX+zf50EL3
hAIiyCmabYPf/EmcvJIE0HhNM1MpSvUpZ0AdnQX3OURUxwCywq5p/HLzEZuKfVCheH7T+BrfOMlZ
BN/8xI8k9MQnUr50Ufm+VIFv1R6rqdIGuj/3Sh5wtmcbooSmi8iBEkh8dIMVOjEgOuGc3q8jphqG
SLVahzCVHU4yrYsN4BZcx5UdvYmEvvzLmTo66WH3odMU+0rsCw8MMqrmq5rDDlXZ8krPDl3R+6CI
92nBnOBt4ZgmBdtIt0xpf5PuEfMCIcdGmlm+zWxiUzbWMft9tEdEf1W5gkMlt83Mq+2EMpNucIRr
ar7hYcR6HiPmw3YgL1214Dq+GNXT2HIu1eqc5rds+YgMPwa8QbZdL+101RToNg+ArOhb7CjCEr9W
UeUSkxbFbc4YFeHqvQkcbTYwysxPatQK6+cE+6LkT7zpTaLUh9SY8kwuLt2GCtyhoxuk/ARRp5Tp
yZBY2HHsZCyHOTY69CUoshuuTDb/oO7Qua1auGU99zY/zb1CJN3BM480vYqd6l0SUKR7zQjbBvXW
4qvMROIkAZMai070G+TL/bHhDEBLWeYts3fsINLiUhPjyaGMjFnAqSmoOnvh8FZuP5CIHUUlPcSR
Zf4MMYQ0fccd8Zqmwav9ySQymSaDZrx70hU8XGRtS0ACwb0voMeHKsyi6UtRgexTh2+qqM60VoyN
Ukb1i8977/BFn/AifOACwBwhpj5xuR0DWJOZiXbhEAa8Cm/XmlG+wAteySHHmC5kYuLFtSxX20uM
VZIZ3QiqtguI26+cwYpPbg1Rkf78k+36GBdH7Ob0rdns99l1aF1c1dieE6vbzZD7tzO9JWaEyWH6
JjOPPveJmzQd0otS0H4JtNe7G65kmNnOS0YWhv1TA1LgMZjItiZ4Bp/G9OfaK4uImQJl1wz8KExI
h+CJ3Pa8O7cGn+g4kMSwvIsc34CVtkWThNeXpACK2iCOnJcDe3PCPDqQDQ+gJjLaxNs2LjPZfGq1
z5N4W5l76wmxXsYyipNV+T8yhIaGyYHD23Of2uT7uho1S1OqlbbqRk4sDCj3LjA9OFBYLRfWGo2K
D0+JJyl/2YFmpbtFpxdgtn+uVYsvURPNIE/9rS+Wm0hHIulfKTCq+KC56qHct/ZgRzOfcuIpboqa
y2Z21n5cviMw15BGV02w8Qe8yVlj8ir2wT9Wrdfd/BMudzWvLtuEGAqj9+5WM0cKKEHwW+n5Yn+s
6gwOJhHM/QOC/ShEC1fwatFILrspKluNs0x6oFCA251ltx4FutDzaqWf4JhFBeZ6GvFjPfBbRe8S
rYPMozHknJYzOPHhO8Cd3lZS6j2SL3Is/Abf6k1JC8/gBrScyja/lTN83LrGfCeBHgLGgG57bHLO
K3E+rGWDFFCCEL5Cnyina6T3qQUxGBkDvKQOkKNxsYKRhhnwji5NEv+L58RE58P28GtC7zb805hp
Ij/eeQnMr6229emxBzMv2vx2eSznnLTU0pwYGG98jxBZEguVdyNJ09DoCiZxXitR+QtZQBxjpc4h
6k8OA/iF+l8IiKYPp3WGSNJ9ojo3RLdZuBLFZRRgkGv9mIRBbhJ++mE+hazh5Fulip7epJ87um4K
/o4TUJvHauvZLach7oy/YAqnoWoZBlfPjjabHyoVBoYpeAedfQeJAVScPjIYqWC3FeOPTXv8Cdke
1vEwtA1IUumeUrnnyIDxur1QcKHZ7vLlmoeHGXG7RHoqEzX8tV9VmL57pr2x/eH/V2CD7npxn1ZT
nab+qnK6IdePY5qfXrKC8sH4RDJivEmysXq/VZlZj+D+EMI33vG5j7FKK0BsJP3arXnz3/GdwLj4
hp6pAB8iHY/+0/TTByezguOY6pWlzeFpa3oamUFnynrXqlrOP2an+6luYKnlCpMpC6r2VNFjcfqY
yalnLtJ2aGIz1xCBL9sVYyBgLLGXSYEMdy3V29BgYydL2P7+JcbDK2pZwCuxPe2rD9HEhckPkGHb
zKzg5NPdTk7/VMYYBS7kFodgwOq7ZiR8D93uvrQFLOS3GUiLH+A/tZsgXa83BPaKWQHEFF9nF6lt
hNbzWjXla5IVSk41HJqbv+Yin/ai+SDuXviJYxBYiiJDdY/tSwt9Bg5l09/8IBzY+ba6j4bKuZ+3
hvRtvCKOfXqhf7HQmzSZ6VuB5h0TjjhiC1Ts1Rpmk/b0j6teWZMM5GSPremmCvhph3lDCx+cBb9b
tbhOrj3/Pr0h6G0GK3fqREXUQ34WgD6BxRtP01pqr42VX9EozGfY/sfp0x/2NFTdVXdxcXmr7Kjq
SAs4/rtquFptST9OBcIqVmVU8CT3TqTds0ky6+0KeVvxL/+FXgKBs6iL5TYBSqYttbvA9A1y7iPV
YnV2Jq3YNbkduDSC/RmDSdjpTmPUzZpQUFg2ihktKp2i+BFGVC3tkOcJwKG/QqQ0wGcanPgeMTpu
TBw44NzoISmUlQspRT8lwjr5RMmTBkSNj7lEka1Aq3SXwCqCsu1U/tP/hxIBDjvNuvEMuuLPR/Ng
u0S1c6jh5RbEecOIF9IZWn4EdtP+zHgS1wrpEFB/Aal9y/ddF1SyP4NPqO6QN6exNG+Zqpcwcrry
lSUNhbgl0w9ptb+LzXl2jIvSJ54mR5oXhBkeLSRwaH3ZaudqSKGZgVUxT0Ar0KiVGZTnCw8Keh3j
JqUKHAm1ShXUJ2fJof9/sSTc+NkoBIRccLqtV0oZSa0S8alVuIK2+WYpCanxlulhCeNTr8jk9DkI
RHURABaTvNVEhLgZnNxLJohFF3O3wkb24gGB7IHy2NiEzJDJ2IOqBhN50iu+8yVpGr8FecwDHUH0
MotUSHGKBtaNJbs2DnWZvRgsy13rCGvCPPld4FMdblQi7oDOhp1H539uEybEaxxXVFA/k/cZIIPz
5wjpfK4LnhWcc15EFXFytXwD60xNN+hw8XRK49xPM2ORaAmC3roTTslKYUkP51uE+jn+6QWOwFgq
tUY1HDVBdJpZkuJ5wbxTorB/M5DttE1yWEZipR8huO3uKrliQgkAKs7zcW10dij+3tgxMkLhwAqB
rzxaVoFDqXkIS21TRI5ibrfv4WieKUQJpFMHEJ94TCEsGMzujkoDWxzIMP2hhKjBpHYbG6wbckXl
jPLmnKN/MwnMv77zYXnQThxUe5jvJCLmKtYvKC7qKLCS5FlOo/geq9s0mgsvTE58z5agZdsrKYik
Mnbkeui6sH9pfYFY2MjsDOsPDVAL40Sp/9FFN7xgwFCWnvyapOIOPb6lkU+TMLR9SJzPXhA/tIbU
IN9ipXk8z+J8XAk1SKaL/ElSdOrBV/CB6dhY1rUJiVTpNnBKLqkolDW6aXnghz3cB2knmuGqocPT
vOjo9f8JQWQ/ls8niE7jNPcgU1JW4GEiD75ojSzBm3i7ceI3XTfbXuN6tgFKiDRU0jacuDUy6UvW
aERXIP8viTTkxYLLXBsc9aSGDYGDodLjvk8HR1XSoEEsK42SAWP8w2LpT4zAe5ezLK47q5vMA2/T
LDyTLR+jLpvVEVekfjN24c0aSo/1BbkpXZvnv6aDhWfGMS8wwcLz+lYLQeFdH0EPyUnKcbvLjwd/
ufUh4r//CYlpoWTtE6+g7+Ajq/Lcy5DAbb6fUnfVb5664MpYrqU4N5a9m0ln8h+iU337D6/fcLDX
rFmrxhXmQ+oMYZQwOGdC58rXdAKA5VTL01U14335kpmtTaE0brFedoYGF87yLizUuoxRg+BLVIVb
Vq0lRn2/oURqLUR+xhHNt1OT5kuthAcZSs3q359gjmr44rb/vtuTZGur5nwdk+N1wL6J75wTlR21
QDd3iuqGQsQjuYVDIY+Rwtj1erER0fxGcRYAm23x+kDKZQcjsHzARdir7pDwf9jKZ+vWXSG1l4YX
XogbAy4WukshtIvLudP+6HkJghtDjo5HsfN6qgfnGaSc0zWZhl/o2+3m07SKXB9gctL3XNUi1sp+
eZmP95lzF4M8RSX0oKfyaEsz5KLlibGDLZctfGMi/Gp/zvwu5fB/KVq+SA81ZWubnHlqqTtMBJ9L
xDE8upmL5atmEUmn3wuECBHudGollyswupQGdEViqVgtxhrDkBtIq8MeQ+semt82iMW2E7byP6hf
AQYW54uN6ENhKnjr0bWlNkcmxeG7NEel2Q2fqkk4yaL1TTHdfsA2E33Z7g7W4AtyKn2ATrSQ2jZP
R9578c0GyrCobU5eIrLNprYZixbAg6mJeF6A9CUBCi7ro9TcNFm4p9Y6VOhq4iMtFdFZsWqnhLz9
EpsA5hPflk0NVeM/4HKqq/mxWkAB4bwlsMjM0+TWtVLjBzSfaliod0tWxxeTeakFm449LsinTg3P
thsalajBVnl0z0/mnjq8QwhpA3AYWr+x7uPx57R9jzI4sXc243uwOa0RvToIOHNBgQl9fBHwahCW
/qjhtpatZZ6TZ6Xh/6mhhx5+556AtxqwxnrD+tpIxgHpT5+an1nGy1eOlNqk0i7dd7UVMbLR+Hj6
C8Ir2g/LsEfapOx8YjMhL8Pg+5IN4zX24XyHlL2ubMcHE6hZGTX/0g/K1jnTm4040L1+P0GNSEIe
OkGOGkwAsp3RL9RKjA+lVwTJZhWOh22rexRCpuSV5vg5FTwMYxSGXPpx5PoLFgtWhruCgctckcIY
KedSsbRJA6S01r8ZAqdji5ZN1goCOo5MHXQ/jcizLKHd0i8vbVrt3wtrgf1EFLoTJlyJ9r+6wXTi
s5prnNfoA5KFvSHJj/J182SH/Ytr50MhuzI/Rzg6332pZ2dKKh4eEKiaggvvT0UTqEaF07nWfYvf
5utOQYkPeGTYkY5GhzYPcJABIAgE36XjAXuQf4/YZVc72XzvGBEuzXrEmTPWteSPMza/lmZN0+Re
lpsAA2mRfhQIzbiWbtBqr/lBcINOdM5++i4JyoEmPU+BNqqD+0OX6r2dGb9LFuki5lpupNXf3Aze
Fs1xn/SqVdIzeK3kM9hUpxVQU2025fcoFBoNYIeeEJYQJzqaLhtC9pwmCxIucvHaEy+BYxJsqvyc
kqVDTqwylEWbmeUd2DwPQ5Ortb8EiboHcR1Tmqnyn71jn1HAt5I4cnYK48lhhdwgKXUtRmGCfMDB
W5EOZ5Tvo+5rFBkVCC6pc0TM8WcRPCfx2lOjVIycLuQTg4k6zuQZh+H1vmK+U9dEaYu2LSOdTzYP
18W1E9LBaVApRlN/sBF89bhFCdt3ULMrvoSJ3fw9y7rVqfHoSlPNHxB9jrP+z4L6uhw05JjuCQRg
M7JbGAZLk5rx50ggvZRGmRvnRN0SuXwLqhKJtFjbW6ljejKAjW/bOUvjPwrT3W2xELxzGTkSCstf
SBJX3B5SxjnoMIPEUAq6sxHrXBxUL3DlqO6XcSWNcb+rMPcvJSFgK3Eq5eetsR9Ys1l1Hytt9Ylw
Oim6CPvzfOBawNQiPOVVaqmiV7r3VmO+yNoh2NStdbLOUWFIwCI9xwumt3dncGa/YisgncxjucaF
lqmRgys+kh4W6m55pq7/nWK+V6dDmmgjkEh027HoRlNWr5FhNwMYPUzxzwxKrcShCKkm57SxHYZV
muK5d8KTmSETqHZSLbskn9PkOOuJy5amxGSwzgzStybcnW5n550/76HiB3xx1F5X+noqKm4Dz5hZ
N51but0NH95068nzZgH4YMLnwOoRmNgVYzrfTd/9tGZFzVsBFQ0wPa6XVYhuLwJY9qWuzvFRF7nv
jab4idbD+vxZG6KDL4Ftw67beH+ja69+p7qcSVcMi4WC6/yD54qsvX23u6UcrbDg/XT1nW9sYoDG
XESiOjlsnxEpSu3KuwPgmTIEgMSWGp7TZlf4cFZehdP/XkDtkOwGJsFwKt3Rl01VOlHjXJRGVIBz
AY50tSN1JEPXnC0Zdijgoobz/5g1N4zkHkyMuDJrJ7tYwc7pNXaq5cpshjqFgAWL4IILo4tC1od5
7WGhj4krSs/N4A7lmbHHC5WPwQxTuYiRx0+GaQTVBOFGcKn/xLdMebfZ3guXtggo6/Znbu+SmHdr
PnXpK7olozRDzeeb77NLFis7elT6NWZ8tE/VY75HslFZ8kHBw5/9AWaZO+1muY5D5lvfFTIzehHV
eZRg9q5bUxjyUBqappJ6yQjXwJJX5IWICktnNYG8H8z/CYQhvJHLq8uiRWLt7gP956uki4olkLw8
W6PhyU3+sJ/dSavp85rV4yhNMJ95l1TcBgLi3milcr5dXv5WrEGZd8nm1bN8/Vp7iFhX07HfySAt
2NyUcpBLGnh7Imul/aFXX9J25Fb3xi9s419mGrLcGKtezhvsYLEBQ5yMFmYt26uJbY+P/U2Jq9SR
9tO/lMOh6Qttv672xnLgU7aqfkGSmCZBLVo3QqM59EujaDvl+j9s8LUIMJOWQ1f79BMQPRgHS5XF
BF1VPns0PAdkdNwm7uYVA/ks9K+IKV3y2Mho/2G7VXo63Ag1GZwOszmYY4cw5+JE6a4yApp9+6oB
kR2KURl8L01gYdZb7s2bKfv7mDJ+qNRTTjp3fM9Sytl8NiaqaogEDmreWRRK4AnbiRlBSoT9TmfE
ecL2kVc0B3FDMh2iPqfpzi+zr9D2c+93KwdWf2WkzPVdovPqEUyqUi/mqIcbra4njlw5ZonojQUL
0Nh/OF9O2ecLzoGftorDnbKecjbw/9JOnJt2f5xCxt0v1e8h6kW+muCHRsBtzdea2DlcmpjKQuBt
g3hi6iCzG3vGM2RQgZi3iDp5voaYm3V0DyJJfrt7mf6kxk0TMbRxm2H5UqJorQOwZrt++gdzmoyV
55mvclD6Dm+rBV1prWNLGeepH6yqPj1EMRgjakaVGDb/k1rbNZHdIggrxcyAGR4RhqiIuH+TVDOK
2j+NWAlZaIGbofRxhzE0OK18u+7BORqqPlh20A9kizouSeZbw45EuRqJbtBUcJg5zHLAhPp3Nofl
YA2uUsU2RoOlF+aW/r0Y2oCqLQ9+OSWVEJgelxvat7R7Bm/ZbFb2hDmXBD6G+ph3DK+JsJWoFcDE
7TSFGX701U6K1OBE8ix+HapO6h6xR4AOS4MhjxJhvEYFUDhphBXTP2/L+SXadCpVAnwdb+AARG58
Fm2V25q9qHFcuNzwiGgnVGltF1VdJB8zlE+Lm3P8sXrA/WVeeDm6XNLkm4uXEKCJeGEX+Zcez0q2
Q9ZL6M/I3le4oS1fXUlJ50EKfCaV8c0DLfIIgkBFwHoIwh6k1Q23WFcr9ye2ccLEB8ey5J5lf7zx
Xcouqh+Vbyqi6gRdJWDpxD+uJnrh7R+AI6dfomeNVWTjMTdD1I1jtL/MXitLWdBI/U+Gkx/uNhE/
MO3cYxLbq/K6xIkJoy3/9kRay6FZNwgULwdgiSREzghPsCoO9VgAIxvhQUZ22nj/KBCUwuXC85c1
mdkuWKL8aWe1g5M1bsk6eTNez+m8+ptcrmlyAZJfDz0a0bDEDpb/g+tWLtdoOs630YkFtaeCQzEb
djO05H11g/Vdj9UvFQCI/pMbP9jne6iHMmaYJUXwH9hi+ltSnMppk3kqniP0TZhWrZ6/ZEBusJmE
C3S4RXykmNm6PyFcoE2U7WwrDtBf5yMgoiXXS60axzesKhK+W5T3SVWtQoR2bN3cSTWMOZs90EpJ
dnu2zo2XAeCez1IUJ0GYRnRxjUUcBn6276wXn0s/3tHyZzYaEqgu0L0XYwDsO+RM9rJ813yVuiq2
IVBR2eq81ObcwTyqfSDDI6dBY6xq+zB1FWK1iyjwNVWuoUHVJfLkshnd8X9ss50MsL7VvI4FI2PN
gTe+WtifQha8BGU89SIEZBEmwz3Z4+dgO97vx6LNK3I4533Ti/0r1G5d7fIEyVaM14ImK468AUVA
0AHa6ggu4iyAavAy9TnzQGP7QB6qSIzRc2k/76Mc3Qs5YE/uh4aJNausuBegQ4sRCYaa1JBECGYw
asjnsNXWfKBnBu7QqefzRQJdFUNdgUwU0Ci1di0uqej7LQR73OL6kLPfzWosFaUdZXXx41X4e6/4
6DJ/32nJfLSZAJ1/+7SayolO2k0p40shyXhfOALL31FY49aYTa27XdefbMVsUYzpGknxAc0SEe26
TtUonm3/+OBlpyuQvDJlD2bwA3/ZSE/cYDS7wg6unBpmJbymdI/AVNSm/93DcT2R7s8ggodsiq5M
YRJD5+o5ihvW6HRyjFeDN/3VKXw7Iv7PoR92bL9nE376/b2KbrU6dNoLYVqmQJ1AuLKqKgr7OgLm
tPFUQiG8UQSxu1ZCNg8Ckb5WoWqVKWAYk6bWyxySJeZCK1DGysNH88Dq+9b8soSDftdfX+eJUH/B
gn2KSS1cYSDAfCE4enVbammcNp26HRJp2lHU8vMjPEIjLl0vhBv9grpwA2NzhATJTNp0vsqcjPc2
Jecon7no0PwzxtuebMuxLkoSvemNZ6DUJsjPC2XmCWil6lZOeK3PfNOHnd2iUjVycST6ajAClmHF
8fA7F98ANvxhyyEuGEt5LHBRLdqzyrmILkLgbJbMRMLcLZ65DNBbxklFegUMI+Q1pdh5vaLSJN+E
L/HaaZHeCViYqePEUT+ixf34LHjGMZvZBQ+avR94MP7YEcJwwBSIRmcleNsTBdj6UnxsgL0yuRW1
VG/SbviAO7LgZvdobYhnbRZnVv5faLUvLD4woWAtsBLKrx1JqBzOQWeTo+rvfcrWLASB1/4x0q/4
CNfwUks5Cu2yfsG0lhaQMv9P6irCa929TdOGnAx85r0Dz46SOvtmMd0eth3JXXwZAiL2cMSMpBQK
v1YVgcvzeRHGQAttrpMb1LLUCu3Nyrk0uaRrE4uc/QjwDj5rp4KxHKHIeIEQu86xN3dK4cjBW5RY
U7vkSsyMh/tWdL/edogOaiX1Ts4dZKGvNrMAOkm19g+RfYafRvVsF7YeMlnXEhP1jVGRxswtnsUT
92qXoDPVulUg9pK4RmfFoRC91KqnGJMRJZb574O86SfGH8O3ZwKfbyEyxWQIANU5kXN2H9sbdyRI
3Z+kA0Gr5O1jJ5C71V9qrNYDf69SWTiC9IbPNa67ODIks6SzSCtXr99232xvPvhwPNFKvzltqFsi
1zYCbYSzy7clpJKElsZ/lYi+s0ys29sW0twTSYMlLXN9YiOwP1PLN81BdXdbpvzldrswCpajHHZ3
zWX8fT+jhPweBeo13L0Dczfpt4a/ll2wqQGmwC3k/nwbLtm6pY1weeyGc9q2xYo6QbaUHpNRTkND
ghXixaJCHX7bLw/BVWfie1jBKOUb/QKXC8HS4yVjAChbok+QcK4wx6zX4D5I31kQRNPxFy7eOVFO
b8cv9Csx94xfAAwG5wwcAwpd+Am4+T3rHQxXD9nZsVMIULuRXEPMI99Wvy7lmCa0SDasHBvRk9CS
FbP4DRbiikLGOBjxnC4wQAtokIMvvZoGIH1yCuBAU8dcV1ElvxU+gxFZhlUGzF+CXmWmjVsIZyDI
cbDs44YvuBT6OWWAuC9wxESTr/I3C0r6TgqgtjMQKhF6mcTAdHAzowBjPTlIh0H36P2+s+rx+wZ2
4vEl/LGNsiwVWcYY2Qtqd2HVIKkVP9w/s7a83gVl+2D+AOZE+HdWbfqPmtvmt1gDiZ0O0NmBPmCn
YTMfFNf4CSuaeDcEd3YdtMe3B7ZcA6dVBGVMeUrJcIfpOsSfvWPGb+nKSZwa63qFcsscTAO1ZwXL
0kp35zmJIb1QkHszn5lBiqhHKbnq4eHTP9e8OhZVB9tLStpi88sCTlxe6cM+nafaswFNEeW062Ng
qUnSIZeNB6C643MR9yi+s5Z6mhkBw9YFm5+n32PqBHmuspF4LhQjDXV24CbBU8RPnucLtEf+OKgS
rvvZhTF8/ZhnwREu0gwgTIJ1hbMnMnbU15c2SR/RDbQguG/720mxKHqUd6NKK4uVrDKqOBDCpqs9
34a4kgAzDmPSIeCt8kNH93VpUbO8g3e4K7OGlbiRWiAYWcnFCNuihRKYM/35E8dM8k/h8ovQqGR1
EDf5+XM+O+Q1PR4se/xQvsNnYkTwugywxjjQTNMXgQHRC6ls+Hi1vY4kbOQtZKV+iMwZw1oeThsw
7ofcnFmURuxIGX/25KmDSBnWLzCMzERLFY4kyNajXwzz7PaZ5+SvhNefl5DvamUs6sRGV0JdtPpo
WMN5XEg6TiVTX4m4TZFDFgsHILvUF6ziW2QPMLc6khOhaWOuQmuAOC0SAOAkDvVidpMmMaQOQDr2
YTNrHa1qfXBW2UrO+oUgertO3CI92a9Eo8Eus1M1SDHPCukwE7MgLdrLqcSxFsfXsb0Ln1aJd0Ii
vzElzqNgGPErF4LO5hacthNHBpX793qIksLjvrVATk3YQNWNwtVktqoxziKH4J5hj+XgpUkjG9SO
2GpLrlns3eRyuqv/5A2Wk5+z3X2JvaJR5bwYzod5XY95z7yXiWu2r/KuT3zsBmNqgTJ/dAPLUsNA
MpSvGsBxV8fiLM5YGq5OmFPAY4BWBsD5GNSbFzZqanEbS3ZS9djq3/4I10iHzGufbT7de5VJMsOZ
PNEY9PVxXQYYRDOFVVhATkXBs1Z+Y/t9P+EH3XFHogW/GCXVMoHEs1xuN4qIEr2sqt0tgFjKr2Qp
p/SkF+4ocxDWgVVM7n751y8xXJE8p3q7ZMOeb48crHVhAeKk+MeAhOgA1d9DRmobuIiCXkTsFwgK
CvdfV+6qbT4KaRDyw+JgOL9o3EAti4+PsRbI4gDzqQFTXoIE4jges2FyilVSi1OVAtgBLOp9RyfZ
vd9n/bG4WpZtbfw24FAPFV6uRPM1KTue2t/U8YrLhdBDSoPba3UTFtvwTYP0SWAmksAyQ6rvmFrD
XJ7RqSLK+gkZDrIFjVjOblKlVrwGOca1DPAnliMGoblmavByNvpR6mDPI7uTtx0fGJHk5G28lxOc
fyvCXZi4LJ4W2GD9IlqF88FosOJq0I8OGIWdYc/OjKwzpG07gCDCDbiH77vCmul6PNyBnWPc3/2B
N2qMT3Z4D7Fn8NUUqN/iFAV3uXiRx7WMn6aUcowYWbuwfhXVtwjRiTqdtjgpyzjLkqPWPdj+Tw4H
3TrSP2Fm9AloeW36fkMt38ctXXgvFBZVF470sot6kRedJXrbFjMDY84AQJg10sR4AKztbLOHRoML
KYY8flvWAB7B+RXNLIwMWHHA8QgCxbtMDfIfoy1FvW3sipeQRpZbvVhJoYOYIz9pCvkfg+c0brUI
sIU5WGmWP0LnDG1Es+vYECsVeqOCajYNjZ/iQQUpaC1RHnS6DaydzgGgfvCj/UbW9CC1QBYIcUPD
1oYr9Brsjj4NUe0MPeCaJqlyCgOZQmXA9Tk74sKW2QokbvdpXtDfOIZorvtE5g80cSR/Zo7KARI5
tKokjssbH69rR3xEav8a0OhSlexbIqzpewueoARRenIXx5Nei9iunoFunfp+/BAvVy/BMjq8ihsd
Tw8+NEmGieC3h6vEmFWtrlcT+afBPca+zkHFzQVR6711RxjwsfnKlP57aNMkZh4lYgOBNkyRb1VS
fRtHCRWrPdXHd/6K0sEmGxKUlA9D6KjnbPyZxNUzKQ+F1bqRKmyKyBhzMC+wHtp8VizEKWwKCibP
CWWmbZAYV8JMvecSAXYk7PEQQTEdtLMJreJALtmqC006LoJWODHVE7bR17KI4Gzf5ITwn0Bc9njI
nS2c12GkomndlMNUiQ6NCgEiCNBcVkUrafw1cQEa0E0gNFRN8ouWNaDpM+YNN18WjycFrmVmZLaL
tEzKs1bBweM7rLmR6fHR7gsbvJvuBFqZuLD7alxhiMxCtjzIYdvnSSuX7B5lJVkhWg6acgQzzbii
2aA4lWVC7vDcwqRGtRtba/E7H7hQgGfMEK3kz4gLNuGIRS/8Mj1u1ZEGVCJhE00zrXlMHm6Qhd3D
z6xW9e7FWE40MYD7kXbHynLtHqPdBAPni3SPz7LuSjc+7RWMw+ZsxWfOlPV6gXl8sko1pe5NqAZL
I6sJTKpTiRPoND0hbAo+DMMnJ2+O1jCMhFFjHByVe4/zxARA3Trqbdkb2AJEqyAw7BLR8ZPQCA8g
LFYodmXgJXuEIvU08CRW0pQAK99stPC5r7Pn5+MWLVgSKN9kjA/yzMXg2B0abQte2KVV37sRtF0X
5ZWoVrYkCRQhQ0/E/w+e8gMdBlSNKcD8sHCBPOKZfqIoLius5FgmcTr/j9VF+w2klU40fT0Zo3Sj
zkTRFmik7uMB3WpuQp8e1v4NbNw0h8m2iPlFYqK1PJfT3B7m3CtcSukNCTFtQTYhE2DZo+OKsrKa
sDQynED1jRdZQspjZi6xddxFY6rrAXTMfxyBo6RQjs0ftINSPqNAz7E3zEgFW62qjKXp5CFgsjiT
EQmP3v71dAwS5bw5ecsy9Vf3VQB9gwC8eUJ4HdvLLwFyzKV97zumP+sZd5tGQCXwjNs+UOOwgTTP
GBAFz1XKz1iBT0Luu2Bk/gU/1eXwKvTaJVM4zaUYkG0PFKvgIreIDE65fBiZa75gsyRDA4Q+nmem
8fzOjIggMAsBEDR4F7oXonbN4GnaIZa0nmMxVOAFnx8Qb/mhqL5Qyl3FCHPcXrU76hxvjEMs4hvA
/iMrsuJ3wLiFD9p+VQfh6M8+LFolS1Suq53N/Is343tOxm6ntd+B79d2NTF+H+2hO8dQUQggSVoV
o4q4RsOxB/2WRZTB4cOpJC2b3XOoL13pZ6kbHkJisDEwoljJTSJ3jT5M6jroC0bkCANDWIMnyR+D
kwIXY06XvZRFtIS3qnpv3Ypy+tjr7n8MjxY4JD0wJF38CADm3GhzmuDn+PoxS/PZ54Fxa3WLNWYl
OcsHVeVbQkq9+GLL8SjTMQwJZkaIcZgVK1kn/OWzFVh8tH9lxVilgV2xatfBDREZcMte3x56X9jR
LNZ3k2579pQm8DTFaP/f4OR9GqXC2LuZdthRhF3X8ArxoDQ0WBJ20UH1WkKytM3V3SPhFnJZ2OVQ
Gd5Pu6NyApcDZ/6wBrajkM1BanU6w15QHEbold9rkp+1SiuwV5tbVm+hxbP5q2av5cKJApQZ1aep
AjUnjavXPg64VGrFKzhyb5sALSghNvcUcsd1ahUD3CDWPuYZZzSVGPniALW3s4BtoLdsz9dwH4v3
JwKGjdrPU0laDdPA1MUTowj0Y4xz/jsuilIelLGEJsOYKIA5ouU0snP9YRa4bNSdpJrWrZFET9M3
8DPq1tvityph4vgfCvxJppqekLsItgXQue2PReXpK1iIJaFDQs/K8CvGq7Xv6a1O4Z7dcw5H8ZkD
TnI3JVkOQY7LFGLYH9yfoQyFiRRpR8n4IEzmsabP6BQf2rxC+D2LSHid/yB7LYpJGSv06yTs/wYr
z+9wxvTvWMGE3GfcVv46zuR7sNE1j0BqiOJF/dPMYFY3uDeD0NI4jK+rI4YDt5sMXwB7qmHP0mTp
DpvTn/n0Uc9x85oWaewpV8hubZ/RWQypPSDRV1tbFxh7T8Toy1E8ioViksnvDrNODmCNz3EqQmad
GkqWjrDz0TE/Upjs6wYlV89FHwujRRdb1E509NxXgt6TGC8mKsRIQ/NJ+2mhyBWiLzjTSVblmUMS
AzRP+8jyxU3MnncNR/s68FScFUpXH/l5LzwKgmdyuMIAdHtIiDwFPeCbSy90rnDSnkqkGVd/PxXG
8CaOJ8OFRUHcx93gYxT78x2Uq3BiQXkV93rZ34mEvF4U5d5LK6T2I05pPQLfsDAaDsJ/stHN5DKn
eebHQSaP4sXDIddmqsweBsi15evbUQqEfViYwCAF7/MBG+LymAdqJnZVvI8ihHPLG8UvvEjv84QU
Ofk3gJUpwmz/fe6kwFvme9nCdfHTpDgZaLt0yncwMK0NdUt6r/7GEHSm9BrYu+5QbrudGr3U4yWM
MlXHlKkb7V+xJIwqruvRryb0EvwNNzNhpNbacK22p0OyX+zfK3N6U+YZW5+TXjCvl6E8Tf+nYKvF
NVDqIgMBXMwG3dtZb0owm5dzJWpZszby35bX+znRghHs6OOeYb4tifdjOiXOEbBGRguQx3gBn2x3
1zuB2IbiF+UkjE3mrgODXNeIg7I+iyqkArTiahAMY6a1w+u/glD/Si/0koBeGrBIZ/hJhhsw9xro
eqiuWE8JljejIiWK0ZWgQ7b+QGjXo7AiFzAGERhJMIpmj9XGSHAR7gUwc7L1+sHG8Ftr4v3ehiwL
lbMsVOy6MT67p3s1IIPzPm7rOEtxv35qYHfc+YB472A4IyikMzAqCQhuJc5uT48e2sHwE8OBHAnB
e3jjzgkaFN0A92gLLJ4hIBth9/KnMy3QB9SrIgmn/FGu/KAZOYzmQC/SVQ179+e2kQbQWnW+uA+d
dBnEt+rYSl2Z2JZbYKaPpHtc0/3I6AOebT22OZjDYhob5HwdKyGod9zkdSxCr1o7QgiAMChdEE+m
29gh/irFaJt9WT7/iR3Bo8Fr8Egaeofj3Zv319rjXL+Q1gEyNI0Ln9diRuWIWgERaOjtBVhGTs4p
EegLCu7IX3TDD4bZneFGqCHIW1wC7F33LkpOoF9ZC0au5N9jLFuEtvnujF+aZKN9CdK+UNp4E2V6
wMc36dsxU2YDNV/hti1Ybd4Pvi/CcAmDM8JbTal9HWdK+oLJYCk1HkiYeBCKxijB1M20Fm+dwIp6
KWrJlXxDTUh7sNH66GZbMzySc76AEOd2ld2Zu4ox3ALx5Gmyz6HzBeakIkwjXmVD9KPyPtMVSB0U
n+5zjv5zZtKZtmIx86WpoRZfobF3zbQwv6gNJ92xrYhsO8L5zwJLtGMxhDUwaFuJnJRVQZVT2Fr2
jKWtiBxxL/ca4TMa+aLRRKQMzQEarG0CoG0G7QT7tPYXV41XNuCTo66SqxDyLNJAluDzO1AwLHM4
ON+gRQCGdWJJhysyTSxVY+OZ+Iwy90Oz+rKX874YdQpaEl/SYphO5kAvdNjgqj2cpv8hBSGDUZO5
C+bT9WoO02jOVq4/B0L1EJA7v/NTaMyLAZJf4QruKXihoqinYgQ79muYU+loQJZGb4bUXJCdBPuo
SydCKhgmR0EWpVFv7qu63Wz5v4Bvlipa2Vt8WpppGVgcw55DQUV+qCtwf3y4ugQ2awQ5s7jxgjHy
yqWI9t8ekuGK6CItbqOWG2wPR8l1UWbEiGENGUIIHZXrzcxwWuLI5/T9aX66JOzObQ/RaOUzBopO
easvY/4/hA+O9oCjhvYVcm1ornnYbOMpGaH1WYX++q4PC/Ft2G7iMYNVj/X3Ln/XydkI45Js2s0n
TSkVg2HuV3/6pIsge1Y5KNBqAwZuTcjLh60Knbtu0AscdPjpT6OK6RfUG+Bmb4/sAdpakXhj0adG
8QoPTBnbhfajqAGfnwenjti2J8XPqB2gDx13DKeMODGoZQB2mhau67s4XQjxOdtK+/9nz5D3O587
P8ddjkNkvJW1YcCDqr+0Y5mzWR/XPDCa2JasiH+Yi29zIpDjZAwaQsWxvicXRjGdWmIUR1atuxTb
K9g2O3cxzjmCFrDFcRoSJB0oW4jcHwyljA9YmtFK9FEP3Knub5p/f1ZLVo69ob2yp+q6sc3NTXi0
4tVky6o1cD7bXZCN2x5Amr/RGlMuOsMM3pJGPeltiQAUjozZcd6dY0hk9eDgcPThl2z47ubUvVDN
jXIjzYTxrLx9nkk0WjAXlDQAb4z2Kz5j2wNdz6+NAocXVxzfiQpGgLu2xuI41hdOyxx1Wct0Vp86
ozizQInubJf/bJoxNlOW4ufPAkitiUPe6KK60JfcAH261sM5J4QllNHYDRsxAPrbpvfi3dJYACSs
hvuzyWdwyTYwZHNeFsPjz1vPNApPAy8E19QQvuEpF8aHIeR7ch2mkdOmHur6iSsE5JONTIvDi/Ts
XnNuK8uFj4qvnYNZdmKxoQdePjmyqMNpwCZBtr6kVEeMsYsVa1hHPPzFkILlWnOtC2kE1iBZwqch
uWJx7cv6C55HdfSwNhn5OL1SNjSb/QSQv2ofjj0F2aEG3LjxTZId05Uhl4jBjxrrC5Ql2ecj+WDn
iK6kzu8+WXLohP36Vn/gh9gvFpBQ0B3dZebXhl24AlEL+vQ6uWf9QrHy0bgvepk6lM9X+A7RgAzb
HczQZ3ILwOQcDEfdv0cSrigpJkrKF+DHU43pk34H8/6Jp7nA+Xg0GUjthdzDjOPCyF9tmUrvliFW
rNeNqGCfYNoKivcT/egKvJkQZYkaqPuN6fvQ+F6bazMz2PvyGn7EhR8IjPTEjZVJgl3v1tDcwnlb
sTN9dWoKmfwzMXF3uWa/T1V8IMJmtLCZZIzhzIlmFa6vNoStitMZftb2nb9s2itZPYxKPzY0UOwe
CgiFGA9f4ClH3TICkA22r3U61jec+LWuTHhuXMoZxRFYU89bxyc6Og0XZFeMCjN34+albzchaix+
Ah33/EQyqdQ1lDzVy7R2LVtOLiM9xMWQONOQz9W+h2iL5eTlOOx8sUDACj6rlz+z4VwveCP7zmKR
yEc86k+uTpj2t/o93ChqLQ5B+XVwUEdoGTnORYpS3ARWrddW/UdMB5SXCRGqiMt3x/aVlZdhZrZC
14KLw5p5ze88fYSpPLzMGgRRMsXoqVkwynOWV87yfl8OwafVaRZMYkGemIS/tP8cNmlRJkmneyYW
nQFy6QR0A/n+BQxqlzHSPnvpFC8FVVrps7udVzhi67byGvaHKygeme8Ygk9obzwoEBi9acZO2BEb
/7GHRmaWs+FL2jOcUxu3M3dPWfVofrCLJdRLl+KthB/8cCYtbZliqERg1bQT0ANvjHmEXfZ29sVI
vmWxfL19g7iGGT4kq6tZjDzYlq1YVQkkGt01G5bSOz8UUn9neFmc3nREhISCG+QbFMZlzQ9mh1hU
QHtaVvukfRotpz2UyiO+ur17bQzOuYNUKedTeJnkdQ/nZPP2FUjhwjZljedvxl+TshGQZ1w7L099
NuW8u/bTPuwLVPK8cExsMTcqfTVGPkd1ge2TidQzHHTDHEw+LD98Q2UZfjASotYm1cHJI3cBDGBJ
fWsohoKTDwMrpVCnO7Ds4A3uUArXO2+9fsazQ//rsXl2ZEEe4t0KIXfUzoiiKivYt7mdrTwzLy0r
5Mh94pqQIouohHiUF8zbk6n0V7flUVzJoTi2eiF9Emga3PUwS6t2SnVQJLoCO1L/erpX8hkqBdYI
7CSt9vEbZk1S8STgPYoh5ydmDv1mete9JEA1/KwhDu41fzSo3NsHGOVYg95ElX241A3XsZCLh7P7
FUxi/z8WtRBf21W78zuwaoypdH7LcrHMUS5oiTUaiqLzbaFZ8n+6Gvb2yHs1+jTVrIqRp6JfdHcl
qv/NQ+afvV+6V69FGYapwRBnP1lge//7EcKe9P2Yy79iuKBCU1XYGiMLC7WhvGX6zwibiJEfbb4f
zVmnxkejFtRktvNOSadevcynKpzO5c9vFbpycyd6PA8hO7RiVld1aTyLBXNITWDaD5TnP7Y1gydI
H0X8CLCJiBVy5ewS3O8t1bcarO2PveX/Xo3m2WXslwCG5mJGa9nmOcHAFqKr2GPbeDks9l65IXNv
oaEBpZz1fGiF9apOyNbKVO2RjcyXCUJSgeuVfz5PV1Cqw62S3HJv+Kts96fbWqbNYO4gtXPo6Tyh
O5uvlrzdds19/O8zcCdnjCTJQgLMt1Pdzhy60puOuBOG6/G4XtsWUEbIiGi5JQhOW4Nt0ikOUiaQ
xW4eHKtG2/uyECV8yC5vaUVWzrB3WUkEt/NT+6maMtAgxukh+Rtni5zDb+hDXxz2SqZPRQDXhQ3u
AQ3AP0jmfT1rMpJVDxNZvgXUiP8kaOGgFUpDpL5wEbp60ETTnSZi4Ibzvs0IaZUyMS7Mf5rgRTmh
EgL+qmPQZx6zi4BRdyfyLo+qeE/EFO9DdjVkUw7o3IXgZZR7513nAUcszQUN2H+QA2+f7vCq1lg/
qa/AW4AOdmzefMFMKYftK5dEeIYUa+H5wLNRBy18rxGXCGQhJ2YQD8U1HXNHW7W/HCdnnqSVzHww
W5ntdXrFF58YuhCa5aq2nu88F2UotQew/U2kGLx9o6mkOK4/ZG5MYupkdvcYzrFpMls9nW7ResTA
r2rGui/7uHgqVwmTCG2XvYheOkigEUm/u/RfoH/5j8haUBfemb2S3hF3zy4soTeV6GWv67FtFOnw
XcBPw1q6zpWFolZuikcc5YptnAd8engH4xfFKkgLcDp6mhFBlTavQ9e4sjMetN6rg/q6WHboBXX8
uVg8U4180+Hyh552Je0Av3kvK1XPTmfOxcwBm/yLArgXvkywBOIxJzumhm8bF4UEvv7GwIH19bZY
lNAPwxOmp3K5OVaZ/b1SBGQL2etOvHQYaBvxxNcbeSLPcJ7mkSSJ7herRrhBU+sGksWVuUKyRhmc
diZEi13GWDQtvCCpRa+HMV42rGgETN5zW7ESWPQXExk5HfAapx9Mvj1falza3kqNtkkYTu137raU
cZa5a/VEGwCRBSUAL07at3dq7MUHpcU6a/GUawHA7q2YHrS/hbUfDFD1sMMC5q2qk9i/w+bScBr0
3Qenkdiax94bE3kbQ0Uz6Qv2qaJHB7GfyQRs4kWaUYyEQO+6rdFhZGqT0Gmj7bXS93ae9eI6tpmS
ppCm/djE8Bp6uD9a1Pff/70BO+zASjtjyTSQMJ/FQMHi23KayCTZhGVXA+y7ltbWcFsXXMZaDg68
na6/4EzPpOZ2DxoiRz6Kzt2Ye+5ntuJAzYaSJ3ep75mRHOplHnPcR85K1MPBhf2yeXmgs1PmIBOh
w1CMd/CkV/Ev71S5+0SnDC6mXv09n5Wyg3nKXIPoDk/7p/9qCkKVz1yza3oxdbuyxLEa4sa+kn7X
/zQoSU5ekQ3bMWQzOXCQH2mGnc/CPjOFyJSS6uv6ukv2vzB0V7N78gfxVo8n15S+DaKl09LDBIx/
KZmGiml/VaAdFfNDQ1VHpnGyfrLGQ9B6tv3dq4MVkpZXkB7DmCi2MKxAm12LHynQFn4pEP9qNoI8
7vURn4b2Kp5t2uFNAhGRtYYV032mrBAATlOUFNZvFua/JEM6BNKj/KASNakTh/mZtv6KqgzwEzvw
wdNCgrvbRZf/ZigZOUOFjnz0RHEAJCErEl05NkmZ4KK9noImJ00xJOMwIB0ti0vVpPLs/p5jvy7D
yHuQcVP8wjk8lEmQXNcBr8USJKCaBvLiifs/bp6tV6/irrmx4lM+mpXhkTjSVicqCClz7/JpcatP
kunQitkN+jBfTVT+YXIdf1uUfUYMk50ytCvUbNS6v6uvruJKxVbH9fp3dceWQkKIMLIyFj28lyCq
n98e2t+54bwBAg2btMFftvlb2xJpBpYHa4XU0OhqzqXORHLH2h7gpbZ4PbO/rXklBjLM4OD8OWjB
MLzbo0DsODv10YNTXFnPipWfsz0tz5UcFEg5advEeGxtmNHHoX5PNbC5fy7e7VcqjXpA+xR4uNR5
o3WaK1lQqk9VO7fTSXRZ7vCJHTzOW+2akmBpg/IFoWrRXIbpQSvKW8GRUpBIDRYs6Tpt4fCWv0ui
fz5NGqCdQqXDDOlLlDd1TaMPXgTNszypkzdpLX1yyGrHC3dbpMG1C0Wihz3neIXPXvxxicrSUX6+
tJeEY1XGVXUPdJ6LVAoQeBAf4CuDW05t6REawLP7Wht5v0NKSSQUFzWBP2N4CIWL6TXG9a+EZ6qM
3gSudS+oNBv+no3Nfh6cyvjTev22LZhahjUqbDoizoJ9FlzknmgsTDoXzyritz/Z0iWLtQJ9CEb0
3CFhRRX/tOqhWNcnl/pswSomh8JeOn9wBDTt2PkYGV0Satg3fo7y1lC6SG+QFtTICaVWsOzz9tLL
lfebd+i2Y6NzAKnjrGwMP8VYP0MrO8Kg7Ct1yPiJtMMTI1LWEh8f8PbcxMwJLSUPTsHkriH6Tox0
akZLvrNudLND2wcTbQAvGDRMnffQZF9GrcH9ySY7sB8bAJj9Ar5x/YAihUZXaoXmtS4ER2uAptvt
k6lr8ABpHBgSMiXAl8a2gOJPJqdZpFJincH+/B0budnZIUBS3DRMwcPuE3ZWI2Tmiq+YmY9T+T7m
IxAEMxva/L1x5aOt57FII3yg2mlO2IKw64EzO6ZF4XX49R58nsJho2zmwi5WuJUtBFMCxFA7KbHM
tTdi+RNElVjxOlwWZLQzdPWhMmjFxDflDXLCZF+FKVDEZgzp60xj+NXujt/Kgcw/+iPLMzUBlbFo
+kmrJHDeejxvY9IsyLXksCAqVJf0GK1qMDfxWwM8dGydGrJyyzUt5+0dNRIo4xwbJco6QdXCEnqT
43TCIlb/KUVRhLh5GchlzWPg8LUtu3rGYiFaazpvfTmTIMyNZjCaodBJ0MXjYLy9w8uimIPzZwGe
5r7dfOg3jC6HrBlrjAqA2G9RF/wbk1iR6tOniXsUDwQ0/0bDlGGlOqiVc/ESM7lW7SVtxygS3UK2
tiN+DaEXzW7YrUdehubr5nkn/h62w+UkxBUmxodc/F8OzF7S8D/J2QkBliY292MgOaxJ9qV1EEcI
ePrXlYI/4RXKb1F6MZc7G4kwsnfjPqLGAEnWGpD/c99hRb+Hcqrs3vPYhFObGLm626XwI3/Fqk49
k59gxMES3BeGPLMNA+Wq7PnPgGVfbrDU15cYPK/BHrz7+yhnWed1hz1aXC7ltujH6TuhPJ+z9oug
sL+U6ybH3AFxqzULs2djSMtPS+7GrhiDWRPhI7DLKFKvjf4PbhypVAhh8vAqBEtEX3cYDaQDBCOI
J1bud1beW9LOJFdAqAKa1yHVEns3OGYZ/GCVeVZxpIG5ecu8SJqD07wQpjUHgpJNUczLn6lgE7/g
rK9QlmaNzOeK/z0aQK6eBaGHqRmjdohXPWbmm3B1anbmv6UoWkTcK9PGdHq9XF9RG088YyDzYh5s
3e2F+nxEUyMvvK0VLtUuTpP4mmJ99cAHFwK8mQXYKt91xhQOmVDIXPjlZCEPeqemx2aVNoR54Hj3
eMRIeyTWA74Qady0QpDuRXMW98ZYdVKnZ4gC/lb5cxBmUolOWFjNNmzwy8v5RJiy0t2ZDTl46YsJ
gprx5DvRwVAL1jIvbSdZELJHUVsNcKsLX0Rn2Pc0r5vv75aeeX1CvoRoHhXD4bZtu/6tapchw9c8
gJbfSkbBl5kUyKhEcx3lS/66VIR9yzyvzMwk3N3wPQyQoBepqJP5i8gbTUgZgUSlqgxZOegFD35h
qbKBIGJ5mt8BwEymlasukabUZZXFIp84W3RorKdwxDgauqGznjAlPGdhqeSLW25UamnDo51Zby7n
kfWr1j0MJuchdP0SWO5Q/HUaV/oP9A9T6RnPBqhqISWMQL1Qz21FjuR4SWuW2I17p0b19BFLEoKK
O/Ozd6YfyA0TdchR2TQOyg3C4MWPjl4GNXP5epAFrX2SPPTO9rCe1ryRfwHkj5O3gR034L7oq2y+
ImDwyKC8T90qQfMxYa0pUCctrTjSEQ2XFGmHU8ePpwvnVqWBgVdgYjNfUJ2L6H8XoGF3Nmv+OhBz
h6397FhixpMYXzAOKycqlS3QpSsALsa0oZei2ErjGEH2O7a5/y6q+wfKoQ5ifwpEusxbiPVCNfPQ
H1NWenb/ElPfpbvWnOfkpJ3PgZyeLZo/nAMIDonc5XE8BIKtrmcwDHl1InDRZKQIr7ixpVjdvvog
J3AS/7qGEh4gnrAbETT2JXbAstAxA60dTleUhiug+yyoynZ6mIOxTpVJIdOOt6JFhMp70zWexKTZ
ArSB2iuWvOAb+1X9jCDokfVbHDMIrcukyD3+/x9OrSAFbHdLBVBbiywGFRNh84V/PxAC3gB5PwQV
W01/CbKisIy5K7c5M9kRBXpVmNHFk4xIXC/lIan0ZY2vP3Pl0dG1esvpF6Z2/BxtbUzbuSvU+C/Q
i7RVZz4OeE9CGQI3wwmpo4w4yY4XAhSBX4jzUR6a5fF1ei8iZpjLcPkeuCmCcI1IgjlAMaad7igI
a8ga8v/OIJ3u7z9s1VwDi5L02H8JkWLFdEF2qXd0WwyJh09lpwFww+h1UH1We//CFSdtHRFh6u0o
KcVb33IUDHlp6VPCgMnRAq96h3mvyjKdE1XyA9eRWSZZemLHrCW/aKHF7W8uSr5ETueWl4eV90lf
877Pn9tTyIagp925ngQTnl2/dR3cFu5DvWOvG9UmxsJJHiu2E8P4S7Clu9RWdO01yYFoLLjbgKah
B0iWLOZ1zMwu+PocgxrDUWWJXQLvOpHleN6YBvM5AKiIhkNjgwXnOFUPEvDM7Rb29anwa5/vbi24
sbDD6813585eK96CJIqSUeJSBGqNSCxpr+tP0QDLCxKZD23l1hUc1RpXb4RejhpAlqMYIT80+1ek
HbWJ1/BxKuAZmk4iRv+0ZRRPftO9/LXRBmRorr3VpVoVUOU1P04JZjK8JjBnraitG8ifJ4ew4GzK
5KEV7wT7/sdX6Gh0FN0E4w2V9yUhAlqYX22Af3PN1UB+Ud4WeADauL8gHvdeQVHhv80uuAbZKaQS
1GOYDNiqYSRsTEAcAM+ShEx+jD0M0hFtgdIs+EH1Avb2hy2ibMgHib1Zpem4sU2ZTm1JLa1cMJEb
X+haoXAS3OFIRhGZX/MnU5NLZlo6ngOJSmAzinoz/08dwnzonbALnROqLez84fOBAOG9QkfOUAnk
okmCHFcG6jHU6iPSbYZrwM6YJr0U4tNVyNE8FTaygtTzLBm1KJbpfPiMfhp/eW7kYioqdSC/9Oq8
NNpTutnYQ6SE2s3OTT5T12RLEZEFp2XSHJu22xTzvR023gZVrBaBL0Tsg4CHCTXWrGYx24xT+9oV
Myf4jDWYUfd5xJiddUMAei5RgmKw7aFzPP9ecumG3kP9uGMXnU+8MrC9gKUZPxw2sOChFylZfyPe
bwmvEyMM5Dtw9VAObRkQq6a4lTKTnYpWYSMcTZKt7ZXbTRDN7J7jUC+0SXd+B4V27gtbfaZF3LCR
WpzCEKn60Veg6XN6utWOXnwXGb2TEZvXGmUco3hUcJY5jRe+CFBKRVXoE0pClSQLZAnQseWV3mph
/DiX7GXuNSM/JbkW08EmJpLuJ2jQsGIjdwPVfi5LW/I//Sfipp5OXpCJQDUwXxuhm2yNtBdbzmkq
SOcwuJNYRaAmScem4VJ69+GlWDUClyN2TonkvEOycnCsnjOem4yTdaZvBKW1mtMaAMfx2wkyIqjr
fWMCfBWJOBu1wIHcdHTgpL4eZslEe9sanxOPPjC/T8sXEWssF7FEvno+V3V3pQwIkTW870UmrVMd
hkQ7rJnyuk8RLoi3pHnpijggs59yrHsxV6BoD+1kkvLfVuru9c5E/udqgcOe92LxNJvtz9MaUUBI
WKc8raDzlmA3d82RZ3FLwxla+eDd9l0/rFbjpYhSTpNDENw8l6ybR4lygyFcdvbzoyRlG9qP6czn
YLKdKItcaV65VnyR8QWR3BnbQ+vgIPRGMtjOLyzmquzdT2PolveTTk8o6VTrce8Fp7iIvks41Br1
CXT4FV4PvRPArpot2mLb6Zb3qGLaxdgljduTV6gtIHH3zACL8ooYGBpREiRyD4Y57PW1Cn051nrj
IrEDbfz+r/0CRHEd+Ixll3DPOyKrkED1mi3pGMv+Szp7f9WLtvwgN3CqdHuzNNNTW8dHjVRVvWK7
iXpP05qLKUX32OVVzLpNmXcYTi/QlxBV0sSLErTZrP91YpIydgI7ofo4dc9GzHm/IMmGNNCPoRjR
WkdU1YgG79gkB+RvG6t6XCq4Fi+voWG+wVrjjNSEEIDuPDQMXYxKhp66cMJuHLDWQLlLU+Sssc1K
YPQsk5ArWMrGmfBOdPM8L6KaXxT56MPo9U0C+ZeJcs0oWaKUbguJytBX+FxNARzEVR9LDmazcbHZ
GpOg5dNCyfD/Uo0cAKopybQGzgWr48TvNwUGRL+P53bsGo8tDI+PNT5LBzsDpmOM/1gb8O6irnp3
lw7IRjR00QXa4wDBslqMG32zlQWhHHqvJkzVieT9zVTGhYnrMIsLvorI44Qd5ZXaIY+9rRznR2Yb
OMqPJJQKNk/6SGxPR8hVvjLvyKvQm94xFcfTrAKYcd7IKLbSM4Kh94PUnr+oVlR1zX4IusqAnj7W
rOqetBhJvIcXMkZE1gevffoHysQ8jBLgrB7hHRkRdE7oEkTK4dLKTvCerM66rTWkORvHBZDts14r
DXiVLVDTlPOX06MApMkKF8NqXNjwD4wq/2/CePjQdTe0GuFjB6jqqJ1ewToTO4CR8JUGBJ9rPWSZ
9fqYI2RZQmP8/v7CgtTm313x/lATOHPOnIxwEihJ6pzHV9Mut2ncFuPL9+TpJ0ev7nhHE+rAxaQo
bRle2cddRv1QD4yyNH2aENK1l+d3bpSbyDkEtuE3k/uLmgQ1F9ETfmeq83R/DUr9iy4HJal9sYLs
X6WQi1M/pvIsLYZHqtUHW+vXzMgmgUOA1tBZPJobtFalc7XKkSX5HETWUjliAcbfI0W5qs8AKODm
lV+XcL4HMy3b6E2Bcszjvwqai9q+rKEcjr1dcgKEVKnuEKLIG2KA1fad7NujbTevfs0ofVgoQvfP
2cJ9yfQJ4j+EWsErVJwb87weCcwnldNuIpQWy64vF5dt/8M+l82Z3G5I4plqtsEeyWsBuWfqh7kJ
UmjegO17kYp3tuSSO3OjKAAvQSapEB7xYtTZVRdDNnCaf3OSg5LrYloBgpF50swv3bBYjpNWU5Nf
VReHeJxsO/34KkIXEK5qYS7lwwF5CkvJf4Vp47VPErRjetHgNf2jyJYnbkweaAGwSY2cD4kqapW7
i/T7f3/eC+NXNgHvrBggPc/aUisQUtj3+B58hixqVC4M9+xsnO8HK09kuviI47CINgXAB9mmaoz9
qDUj7ZdKpQSJP9vDjJ5OvUNY98yCluUlBrIRPImh2Tc1mztXv8eWIkd9SVZAzqFd4JZV68qVAHOU
Iw4eZqvsElUhUOs56YlsKhWtSBGJzSnVjBUzXN+uWCVBVNAaPMLTnmOi2ZcdM8nLSBtxrGyp0f4v
VnGvKr+B/Tc8HvLUrt0SC2NsCsFzLfEi/fPbb6M9oIpDn6eLGRAHijbcSpjbII7Dm0nxnlgFk3gZ
pkK96eCfqFa3eHX52TrHFQnpQmoJNPXsJkf1WQ1zhrcFG5iRyISS/VSVR4hj3tmG1k3mQM7K8Jrq
AK5f1/v78FcuYir5nrcNtciKHXynmjjgcv6QEdVyfhxCrxEtwJmx1DuG5KzhMjhl8697qG6rYxfE
LUBhZu16UghRU3cpChdNYGhAVy4tie+ERtatUgK4+YxgbQh0SdcgttVVraJUAwHAgw/TW35VdShr
VVFhx8vx3ntDlkB2f2zPXOHqckd2oY482pe6eO6pvbjBu5T9VVObjW+8EU/M02DQR/OCA0eWyBWw
M6ARU6r1EaigiIyKpfH0e5XDRXhdDRsa2eBOc++lM6/vi79cb55fZMV3G/M03ViUdMJpJgqdCOAS
6l2/90wP1Reg/cWQx5jFQywI4XyFscNm9ATLKrezTS1MZH9PUlbARXeImHfVi7tmpNCygwbvxb1D
MlSCucEFzgdkhckJdgSm06wSG8GGKVHQV2YxLTyFkA6MyLC61hkjFUBsHJCC8yxaNGj6jFTAEph3
uNzASa1Zzbd4s6T21e+94ppO2jMdq4pWdQZPj4GMaK7cu2ymkwkFVbn73hamSSsqSvI8+LegVqpk
xSjYTjWzkWw1mOvZoaa7cweW4andN7vyjExPkaCPocSDJTT9C5h8r9e8CFFH2C7QX5PbKr71nfuC
LNOHOUDODXhddm64OTYk7h3OV8Ui0si6MTMv7iDPyftUW0Xz6fsqpCY+2F2/PTyTsKYBZCnUQd7b
OxCMUpw+Tb6zK2Sp5bUn2CcP6XgZPK8ZmdwncmoOa6vD5C6oNimqRnYNwIw2u+HZQxSlY0pzMHzN
+uFk9Gtdic5kM6qoSBQ/rz2khyRIYxHVdWeBKTNIrXbQDmc5It/+pxh1PNicQtuX5RbKI5ilC/Tr
Ps0dLJZj0t6v0WNanFvpTeDp5eVGrIIbzs+c9k/iwKXGxRwTtwCZ4b1nC6OCaM88aV0vnWVX6Fsd
BCpMpL7OQrdjg52h5gk4IEmn96Ovw19B8JnrOax5tnNqwZm9HStEIA6bqDZcamr9H+0qdFl8/Ir+
NfVGP8u4fKB2WOoXRKdxSq5tROjHg2hsQTAFLkmmDXj2rkzEZklYRBDqlpNa3UahaSQYgUQSyGmP
oi1s17S8GI42musQHjWkGkgYSrbUnGV64FpRN8omUcb/fge7XyQWIjNiAk3lFs1a+HQfniL/VK9c
lqVfKvtAqyMBpSythSzNkj8KA6e63Jo7WpVXeCk81VoNsRj+VEIFdqmX8gB2xwD/BC+Ckv+2OBA3
1PtJl3bDG47ewNBX9ZYx8enogjNQJHCWDhl4shA2rz3IprNE5C/z5+KXgYokqHfWkS4Acit+hQ/C
MgDTNNhJZMCss0t/M2NeAvQdn4raodxcrBBXRSosOS9gvaENR/iEr/BnpsqKnUcGhgHVbjYRQNBs
+0f9cW7xjFtAufkKT5nCr7KbNTuXZoBvxketwJ7eymlwnY12Npsn4bLH5StMprdqP3V0FIwv3kJQ
Jk6FxX+YRwr7MTF4himeuqVhKg5uj8w+r4gVksoJxAzv/LL8vIFMH3ViRTG0QN8I9HBEG1AwvMYi
G/XUEgxekUywm0xSf2JjmcGIkw4Q8LFEbebW7biiymVuRxgL003h5h+gS7QO8cTO6EpV/He/Vwwt
rp1+O2YZRAEwdbii1Jc+n/sj59Tjwsl6Pshrmw8Ob22ulK94L1tpDrerl/WyhP3h7c/gRNCnJOaA
o3YYmrDDtLB3lIsDLyDwNJ6EOeDu23pjZvJCfNXq2qtNRGJkWtb2Cg35/XXKLqQ9tCvb/Vv0qpd9
CyhWEnObL1QPbFeF3JLYZ8uPZOs0vOKzGXq4zZ/OECFy8MJNCmvfQCAO4vfCeAKZL1ahI2cHKUF5
ACrKiJxQ/mlzWzgdVzGc+4qWVAuadsLmHRIUttEHiSwbuvXfZkmbSR3DrUxYqnTYgWIy++xf0o/k
bjbDfDzG79c+0fT/SkaZK6vkwxX/7/x9Q4oJXVMOElWaz2FGb8r2S5WvcAUBNz42RuQVAZtDXfy6
TnrxHUA/WWLV2nTtoqV29maPVQDsOCD8GO5+fJz2JZ38HeYv2Y6XB51JFui2OHhWcltI+CoRX1Gb
Lfq5DybMtx/wSTpPbSiJalRhDReXEndZV6SImHZzcMx838aWfV/L/4lxIS34uCdUXa3e6akuHhUc
Jz1mR3Hu3G+oicfZuxloKtik6xs6kAoTz0PSRLstHw2tT9yYRNDZaBTeT+Bu0Q1HNGRHgqlPkjC9
EjqC9GRe5PmT21xUSiOc0mjLeDQGlQgbIyStxWvYQbVmxt7JrrICKEEF5L3fRUhnMd0UdPid7F4g
sCnbI1wrOw21uQfhmAAETUmV5IjIHz25IQ3b24IT+5LShqc4QsxhnIlon/oaXteEHSPMi5rDuOu7
KiwASbfdQB/wo7u+ILvyH2tNcOusFCudnyUo/Ok2MubTkmAwXz4RflJWh3CJBalKrpaKxUGRf4Gs
akmQ27XKe7WqJS0EUYIngRcc6dFj0wQSN5J2pbKd2XqHhPfx20/oPwCMeIMx93bVZ/528SF5Gvmz
bINSynTfZdkuFGKGIUIYPBl0gTt99l6d0ll9ZJhFJs1nmEyBCCIOsfQipFPJnl9t8KhiveVhSxPM
x68bCkp//Jo6a4dGWT2jin6C5C+UhX/RCrzpZaYkrepcHt41bNfoqdBOfq+q3Oza9XUau76LBWwH
GxS2GU0TDr/qyR9FTTjwLF204g9n3/A5wWnxklghhqCxglcHBOnTMr0ZQxRnGnHifiTT92fiqKA3
DOzZzB+mUwGpLx2d434x34fdenNKldAdQxhqbAziUb53Mlt88Zw2uUIZcpgXdZ1UQYwOPrj2RAnj
KgXvYRAxHDU4Hw4aa4YI1UvTTyDZro1oSDKkOLUF328hS5Yj5NiNcpBkbE4/3CpvpQfE2O96h7bZ
XYrZBBcO9ucnYRe/lc0g4+MIM7gcvO9yFpkHJlUUJLPC2W+pmH/sH57uGQOwT+bIcXop6Yte7K+g
wD7FVg2NVn6FL6R2ZwR+Cb4IDBYaS17ckFFzpF/buumt4vkPoGhTASo+nUYqfSbiV1+1FQUyOvVI
abKpjbWA/GuABmV59Twjeat3Bsy7IUr+5hWsSMUoBDwLm8KUYPzM+kvb90a+Y5JYxgEyvI5RCIKZ
uXxloeZW3fMSk+fXMtUDFTy2eLKz5RRnUcio95zDjdI4EYGwi9zGxEZFneegBagYyuTI8Ve3+UOM
7RgweCqBV8qZ5NdPawbh+lF4WeydgclQozmtdG4GqmtXk2koNZm2HlOXBxXf0SRA9J2hbS6ZtgTd
8jwItkQhpw7lEMMCyDaTz3lWlwp2wZRtzHWzR4l2xjaH3Nt9jfqeJ9TkfCQ3Z9t8rU+0qjPy0lpe
ehHhJpAt0arWOjaTo14NgohfKvk2Q4oBfS1Wq9/yjFV99Rw6YWY8wKoPlGmhEIkvHqqX5CG4FvHz
Kvn/EWArjxVTJeOUYYcV90ggae3jpJSdh6F/JTVnhX2Yr3yMF+xc+2Vuw56F66h/oTviOIr/IS9+
Tbjw8Z/7Sde2y65PXksPNBVPBo6pSxjPux/7czaeE85mZdN3/scc6MDiAUyf4mfJuXYtYu1oF+qj
OPO1jhpHaj/d4DXoInTdBf24oQNUcHLsxhyuiqJNB++/Oap37uk3l5DGAXLzAELf7DE4vfv8MGlr
uKf426RCnQnLMdxdqivkOOQM4CfyzML5eRC388x+8X0zX7dRnK8FZ1mhNwIUMkezHxW7+wyUzeX9
izil+I6rFd54fSfrEjTMTf9liKiB5gh75xt6jX4QbA1OTYWRF7Anek4EcJOZ4R1AKECzcYCHzqdB
2mQdMU4Hoh+QdQIEtTzYavCjFIOIQKin6IYOhiu+A/VQG0RQDzJVrt0R+qi5pBLB9YvCqk4sMAiI
ewkt8CQ3URojYbiMy4vYmnCSLQeS/ll4oyyJLa91jgNe5FF20LslbpnzhRLZ5zNb9R0ClCe6wEuK
Y2vmUYcvgzdbpHuh6hrwfyvj+pHsUlbf7qgb/VFFwUjUXlesIe21NBStZTn2BBwJV9KU8Ir618Mo
jCR6d04sHo/ZOfxlS1OP7NN9I7a49blzLZlq1+2Ps0Ot0cgBrW0OcQfEYVzI9PeDB3mqsqUf4sia
+t9s7TieatiRheLyhiWw/zJrcW1ZyyviW1JDOsWAbiXYduLWOnvjIkMJGQ6ZKEWJW8do0Z8zWcG1
Jaz3ZXWqpOd6myfEjd3ZxHwhVd71J7aqp/kqiF93tCHo0DNS72466vRKLJ36S+0KPDeGat80MFDB
/TOYvWIHpEgCXNledpr57/+NU7P170TNpJ+1V0VFC/gy9g0rVzae3PcMkwU2hnGV9E3sBv45o0TQ
3A81/Im4K/RpEjYmOTDf1mIdNrVX7If7ZIgFi74CHxlTjBzUAKzgqIqZ9HpCeCQAQn0cHVLA8KhT
2Jak4I9HawQW1rorgL2NqsGmovBWStO6+EllqbXMpHRPitTb/Q7ehHidi8ScC41sgVtrq6g7SMY/
9Tlw68iDtlox2Zb6CSCuoYAKq5R4me15KdJWTnIJIQikNHv3x4+9c7w7cRzQITdmgn7u1UGSJMBH
dCfaurcjMSC8EEiruPf2KZI7+c1chGimPQLhUuP+58cND8RYAxbZ3fFhfsqxUols60XaLvTbIyUM
pxEQ9OiK7BPpiupa82ygDFq1+4+4cW1VysopD4rfusEP9+YP99K7MPv3Lutc2Pn2YdsthGO0TiNf
CJ4fesLUI/gaaYOdG9qtOS8FRn34GlxCeXFf9y8NDO0+D0AHbGd0QTdYY0v2aHP20Qu8QnM/Ignj
waTvscJJcojpFixlUQwzfJNUy8zOc5WzljT7iCIIxrpbKX3ZbINi1sNHxlSuzYWYIv79y8+/GokI
0dl7zAln1LMm5sLst2+JMfGAv4npYUYauFpfBG/F4knjn+0TH74n56sg3d57o0isiUwBZL1kNvM6
mWek/6FZJRHeYZAM1uuFIWVy5XF8OnZQOQvNBpTDEP8J/NWoWvDNtB7dc8rPfhNt+pCeGzLV/WMR
PIhRSUO+e7p2yQUL5Y5lbEJduoHdKVbO/iHsuAUpz2TlLBoAZWEJDyWtq+4bS0vdr6BtiQY6z6LA
C9JjqKOPVtMPN1MrcjP81PVK4nzIpwY3MBZXnIok9XPIQGya/4q6xUEJHrGMIrd5E2CO9MgEncyd
NvDwUWrUMw840BN+muTiVTsWoxtuMOA9p+Iqp+sULaLjrfqrkQs2fh7Q1oxt+phaCOjvp+BCYkg/
XOd1LNFc9w4j3ByCxXJO331L/B7cQ2LGIRqZKd0d2euB/lL0EOhotJaVOfbUFIq3debSH7JovivN
ynie2bVeex0Wn/faNQPu8/EoJRztxSB4/ajHmXxcDaiMukdQo4J+RjXSz30ERehNYqQCWmimncll
5I+4B+AEi2oC+5UqjGXrEYfyMfcU2qwfIm4LR+Z79Dns/2oEcdYXXttzOjHxbIeg2x9K8CoJ1dmX
6f5s0ceLf++sWmulQs6bcOc2rynYN9oVNYCk0j/zS4+GvGr1/7nsW1Rl+RzdLRONL3ulb9ZYYZeH
OK64MKjEZBxGHIRCbb9dzH73no5zY8UoPb1BQHCKyFe4WRP+IjFiyGLkFZTEw7ovwA7kExt8FxfO
XUs3pARmJD1X5PuUAlPQFYm1CWkmzW00jRzAL0C1DbJrXAuRVGWwDxZ5hSMfWqB9bVjR4gHoOklk
N8DqDwmSkd5zEs4tWDjx+t8gPVKmXD+pzJlIzUIZw7oIR7qzIv5Oe1dGpeU85wduznpAA+LGyNi8
7otrX7qp6Cvi3T6oIEvzHoPS+d6nQ4xpAUSBv3OnRgNCfC1wU7tADzSlfYp4t8qx3LZFgQPRK9GU
Bzrxp9DhnE3l0k8hUs7e15TPRn9hM8UuA5PErzy6TWdkO1Au0GpuSOOWor1IAN4Xc0IH7VWoIRXr
9s4UPj081lU2Hqs4RkQNAW4P23UMe+ejss6aW33bFt7LVnw8kteuN0GfgotSVZyAQPL5S8e+7rR/
DRI/qQXmJqatV95qLZU1VdbqyxKb9D6wB8r8R3snWIH43fTMpvd4PwiIylrGTF/y6/RJLtwHDCat
O5z434eTtVPey3GjU/u59vg/WtOsxc7qj1AVKTzi/qU6V1pY7jlbQ88iKbRsB4hAbnpnzCqQRN1M
zagS7EaXwZ5ej7mSy4Myoruu27g6FJglrasZjleaPRXMvC/Sqd3OxueqK+c8nQ6s8qrX+Tfve7t4
Be9D09SXpBjiJWC4p1Xw3vqcSHbWN6T4E30lRclA7VwHMmFL1ViNSEQLCgc3BpCF3J2Gi3dLxt+w
fk4QJSmcsZyjnIAtbRupjSF8vzaR3IN4+Ensfe/ZU8nZx8WrUyN+IhT84WNh9hOA0xn0niCuIusa
dlQGDvA2y0wWjP65glcPq9JJxJAr5paws/OMybbgVvuoufq1NZzn405VKMSCieInauywefZUvGlR
dm3IXxb6aMFMZPGsl+otJVhXiYw7uZcAUVJJbhOvjJ1RIdhn5GEyNzGlQPP3YJJv0QvbIp0RMzY+
KWxDqfYs9N04B7sJuDuM7+GwiTaFgi06v+H3YA4NJaIJ3BwUcyr9Ot430u6THHQhhge8dSg6pcvQ
0Gph1eGA85MY2Dn8QNWkeGJWJzVfeEYizsq2xNyxH8bmTFXu+M0xEy+x8DBLud00lGicKlMzpKDA
mJEoED829Z5lSIyvvoZvBRdo4m3rH2A5NupRw+oRaHn6Q3iJq0pmOeMxQClEPPJxI6ITmut/oQYd
C/P1X38xyQV1r3e0rWErstRzBwL4D91o7MKnNx1bFBeQyeMJnATasMpi0m2pTLiaSsATS6hsfI+k
UQeLEtwbohwzpRHFDuJWt+mSHvpIibmvswljRARz5DW5FlsresoTMRImpQs+cKOpfAf3ld0od3M+
YafdhUWXuvjIdYegl1norfNi2mIjBv8XmpNkqcEc53Zm5CIxQgXMCQNwPKOUxi4e2feL6kb9gn2S
NrAqw0YzOoljgG3/YrKru2AUctIV6BY/LHZLxDxi9TYhtdIPQvhZfDFOidvBqiVmjhgPuLSKbDI/
PXEAveU4DyPXeHjEHeK2RnI5r0KsNx9JKWr68bDUg7nhBxrlsPO80YvYo3QfISAH5wJyEwMvjCHQ
0vcq4u+Z7xgOgJPg2A7PAmJAJoXfkOhUjn/C5+zofeu56tAhHJ5MoLKj0INTiPEZLMknFxdY7y4C
XbV+X/X840MvVEDNThFBzJMRtEH2atXVgl7a9lBx4LA+9J28vFFrp9G/TXkdPfrJx/ZKxNQzq+8K
goltHAE3uaTehDynjqXW4J86GuHSueG5dmx/n2mQj7sjsBxjqATR7O/7ZZMsb7mYH4KYE+xsl2B0
xEWxyru5SFhwL4JEGf3gAOiKtQnCUBEMGMwi/0hLeeHX7QICOHbvxndhC1Fm7KHubrGvbqwYndoM
7G9NpPC2bXdwtQY+qW6UwyQp+GnBm72cFWBvPpHElLcp4+7KSYyafTH3nErRBizAJq3aHZomXLDh
wraTRry8sLQRVirpxC0Jwob99UQHLb3VI1j1AseeubxpWlokr/L8SkZyghkPr9qLDO//iU79UUtU
TgpwsVAzCbRWiEgEedqjk0GUug4ZgAY8Oc7zHGWDPLPPU3WrAuW80vjODrSFXbw73kTnhu1J6UTh
FB5sZb3XZNy99RG/QLZZlYBAN1J2XR5OvyshJREFHjeTe61/0LUUGWorw95lcCmNYl99Nw1AHPej
Jc6v8nTl0l++mBUqPwlEpDsIHNWhn/ZPjQMwW51xZavn0oxaopUTaNT3yBdi/Y0xz+s67zPQeH8X
xA4o6CS/UBtfUYCdTAhPf3G/esXCDIznOlUntVkzxRpokBznzNFEjysWKELYoMXg3ddBO1OrIdYn
dcTetmqHaeM1lRuXZiffuvpDiMKvSWwx3GPu/KT3BU5EhrCYgVJ5bFxhcbcMaXMyxr4tI3uRTO1E
Bl/FcEXI+DFMTAHUicq1iUwswvJh72CbAKJ+RZaPCs418HkrYLTyjbrZAkSr/Bp0MuMhkefymF19
gX31nPbwZd7ZR49zwShexen1Q79leNaOqvfOnydCvlTwc0BkpztVCRR4Q92MumJM5qy/o/qMAOxS
TfWyEqsxNPoTzuRyytjXQhAsTagSDxIMwp6a5XGqCNi8JFZOSqJtEwIdkQP6OWzCT110dc7d/LVk
l7wDNe9Tz+MJChYQdY7OA/kLdTa0AzaPddn3whezG6qx04e+mdpftMBFFmU4UWerb4OkdZM+2aX/
pajMtg4n8rUjpfWk5mqocJrpshWC0Fuk7famdfa7fwVOOaH+Nt4p3Y3OOs2kC3eZVWZn8I5kgr/S
FueKLoOWQClevOmmUlYNAFuZock1nHYbHAEkzcXSwOSySMZ3At3U2z4u0gW1XUpzL7/0z4M5G6Xi
I6Q6dLVpt0B+X1gPHEJ9higyx7UHmgUN5rWVD53Q71dLbEHW178mhB3gTMrvTfZcaLZPr8COH2RU
LbTirpJGDuNdLI60LzRYqlaeeG8wuy4OCqzcmKI8c3FDtDfdygcos0deUkQOikRE1bJWyiDwC5kO
gnnQ/S7kxVeBpqCpdvH0tMXaLWRHLoQ9vwH3NIukqSnAK1kP8rCKgannp7pL1KkOhhY2sqLU+tX+
p+ZX5rMw8a+xbWBtxuTXj9iFjgMUbdQ4c+owQ85/edJ6y/BHH5+HytAPaD5BhKN/nHhhuQxls+hB
X+GqxB+Zt4s00yizvG5pqVPUbkympG+a1Hl9VNU7X3lRV7UPFy1rofSPW4X+gQiL1pAj85hViAvg
IuK1GVMsX9MrYBNRFrUD9A28cKO3cIa+3mjnIEWWb8Zj+iox2JysE+UddtnCG++ZXfssi3c+fRE5
VdS5r5MBFXVAxcgwOTjl2fYXClVp7MrwyvtJEX2TVRYrukV0MYInP1EE9G/RRBAOKC+0bhTVwOob
5nSpyk6xH4zsb6J0m2xav7h6PAH8DUir391qRJT2Blf32X8d/H0YuxkdanW1xD047r4JMXug6UR3
3AK8fhTmku22XSSt+++woOyiJqY9OjK95tCtiduZUj67vYwAe/tE9opUOt2q/zJLWNwKvKUmAMp5
xRdUDNZG3PkptqZMkRpczq6DzHZAneOLC1ZuHAyne7y2EokXBr0CQU33B0j1S7sLPpK92Tk11Nkh
3yr6YPY/zF8vIs/BP5HHRHzIm3mFpXjBjMqeh3pnxCRgtRXXSP+Z5s4y2JjbRElwhmrBWRt87Ohx
01FKljc5DcOw+Jow76h+y4lIWC5KQoRDRzFcY3KtQRYbKXNxyii5nAwqpsZpH20UMWgIqN8OkTqp
ehRJWw2L7zBvNNLD6loFf3MXGJf+YznMztgBFAaZtw/8t8fwUaK7PWmC3K5CRLaXLYBGBz7aSGKI
Mkzge4cvaxAanI8inDj4br009axyaepIe2sO5VsajOG9jgyxf+m6URNGK13Xp7wtacoVN7BNuOQs
Qsa6K2oti4gQxQZljRO45tgPDM5IyzmqVcyss6aDSxXqDvwt3T/0mYMc/stuzWtxh0Zwke0qNMdr
tfT5gns8Ucoiomf2uTfjniWtZP197ztQGAKl9tBaxCIofI00vTFu2OI2Ita6jrclka4HvjUOO6Vs
+6m5qwSPL5k4MRYoT+bWgPnwZh6qy7dAf0MDkO4BWNzEPLlNGJI+rYtsG6ViZ8Iv0yWuacxJDOyR
6OWMWfvQ6+MYaFf+VwqtbyjQKiivQM7A41AROJvuIwpMtsWHYV+iCZCJdDrO4ZWwH261JMMvPb9u
Rnm2Jx0ixw3KN0Zl8MtnVpC3Ong979P0gWpFUgw+tyttcGApj+B0Bo+d/oO1c1LITNq2jPr48GXC
iUkzF7xceT6F5/2RsEMaAngKZQ039VuhAoTM71BK6KGS3Sx+bCaDaGOCv47/mZqsNQfbgAH0HgyS
FbK9pZ0L8TTz3qwoh9l4o+N6KS6fnG37EbQoQe3FU8zV749FblZcz60eA83hzmVovgVrljfwZJOQ
l9OrBIT03vCjTwrKA3fBkdFDZkJeyxFYkdjqvYgbadn9An3OSIRjoE9F5X+4zMJFSqWkcfDgUUmO
dR2omX21IlnlkVI+R0GgwEI4Nv15bC2GzWMrJmXJB8aN1FkavaG2jyLHZfSoW9teR8UBcH7VjqsS
UEJPhplP1jZzsARkVt7DU83KDmhv6uPcYYZwYHirlPArZrxWwZSZS3VgWM0LxV9qOdmVIo1kVEsu
DbSW6L8J4sstWaSdpPbuNjIhRjbjs+tbwmUeuSZsNap8v0FwZJ3R1RsnTqeYKox0J4OTw95i/poG
35thNPC6K+2W2t5eA+rtq1lioEEyZXdF7MUaOdbDfcq8VHBTuY/cdlcDbGofZAfg+whhqWV3f4Qe
iKI8rywrlC/r4FqV9+xlMHsWO8vIf5a2ewal1XJ3UrvKA5Kifh8LFP2mC8XMI49vnFghKW6LIqlD
MWQY00hUZkEvA0Gr8pkXIIz581VIc40IYno2F5LijuUQc3BR2gTX0CB+9KdHak6qOdxB0CGnRGxS
/NQvj3PypoCZ+I11L9ea3rWAFJV4EfD2+1/rdjs6X0n/TztkxM1f5PJve7tA2nFA2qb2rduWcvSK
7yrCrl4BjGDkxOpSNa9P6MsxLvMnIYlHJjVoJK/CHDLjOdSWtj+MHBdoWud/+DJ3S8Vx6MpOLUr/
RUgSYBOhtMRLtNGr0GpeUHLfxxIseI62Kbb9jJ5+XeTDLyws0hMZOtn5Gpk9MbLASzfiOgo3Wq5t
fTbrEfXoqhLUJq0LZdfMzpCOKZUzJXYCajVaDJutUQ3sYK7+n/Hj1fhCKv0ETtJQyip3kg1OAXeV
PSHBphgztYnH+m/dWBzPIRl3m8+OEep/0AZT3y8S4cYo9ZhM15SrPY66rm1FNbYo5sxRXPSbiR03
au74o2e5t+SCwlSgUHnvp8HSVWtuO7tSSDtFdwh2a70hJHuTyw+uDScLVvFuC3o1nlmyTzC0GwvK
sqEhizi1pDw2EPE6Blj5liXkvgi5M4GBnVKFv5yNWrHkXGT1S6qP/INwctEElsGFEXTgd3f3splP
OHbyJw1KzVuP+L7WSqSpM2V1D1O3Pr0tB0G2MZR+0PFSvxaO/xTXD31MixbAnaaILhT7QfOX+kMk
V0/mOoulQQCwIuT3/F7ePKwU1REdyzZaSaEo717qHQk0g7dv9ifmNlNnpSjuTF8667A0bYjrjHST
IqVWlu1qs7kn9ZFu+UbfYO1B+w/BFTgOzOTYt/KwuiH53mj0z7f5BnTwK2Hc7WbHCKMRNkzt/iEZ
ziG7SmfVSgQ6puaPZtib8IQlEUIx5TYlRss9O1IRkJ3q0cAFnCW4vhp51/6yAAAMav97/ldaWFI2
SPWQOlNN+pobVelI6Z3ooSgkHSIxT31glut2x8oRTsLtAxaSFPodISx6Yz2llZ/iQxIBk+5QG3QB
c4bII5N77hSJFV288wVPH5cFM6a6nYCCErlZmN3okYZDU8LMo2lcM7AEDgduxuq08UhNSFV/QT97
ATfEExq5jY+x+9WaZ4jgoToSPY+gR1h3ca79NRY37rAB8gk88Z+xxnv+xCl63bB2TyTgbRl6p/jh
V2QGRGezpU4nz4rMKveYJHotpcC6ZD6iH4ZJmjlHU4YTbp7cnUEujhbbYLXycdv+hYDDynVa54lx
L6JNHeEGTft6Em1Md8ppgjJ9m2tCNZ7QwghiQyh8//bMfkntz1MrqWL0Xf58+EMg0YetSaAW9QAY
ODkufR9UvUOl/Ill89iVTQAP/pfkLYWznKSCAhSAeo6JZB/toXvtB3154pHV/3vjYB0sRxlQM0X2
xXGdBVeJv2DHNUFeVmv//0bFRLA4JT03+OVSq49xnvoM3hL3Ov+r07xeMYaUa4omPONMED3OLN/g
I2bbWC91VdQbxCopHXaPf5scN4okScE1a64Ow/7/xSGuSCkZLLBVvjpJcdUjrT4NqgPF4y3nvWLk
j1IE92nRpf02dMEshDNF/ZQYFDINV5oQhBuHsV+ld9wHFEcaQB5GJTpgBB4ED1B7WAhvThoxP0Gr
4pe5sol6r9LpvLunt4rO60eHXDHM01wKQqOyNTJVrxuo6gXTR5OwMX1oTIXFQ0XO6IonHSIdvnXr
6hPAgCqVcoudYOLeYk5610BXj945c8l0bDpTCS8o6PPsjXbIKGNz5yyb0RI2iHV0qkIvQlaIFnyy
4OIA0rnfqnr31ir1C4r2zt6+EHyB2AmMOn5GuXWO0Be/LgH+TruFpPWPkpW8ZE1myRSkRXr4P1zo
ztl9pujhlCyF09Lg0D0ia4M7CVqJ7rHNz+OSdmfug/gPpRY+v/DJw0w6IbeJEYL7KIWNRXKxmOSz
wl7+Ey7tjMNFcBM7xfdCX3q0MpK8ZJhqmgDLgV3YD/4ydxJuaer0v5YcrVH+t7UFb15tWDcDPglg
8LZPvJcVBwt6ERo3FPRgR+WMM8uvZ+533mF9++VCY8YKAdkrs3fU2eh+jjsKEB91gQd0kqUrrLdy
coF9Pvk4Akhfs7zlOCy+xpVB6VBbUNC62ZFhZgyHLkINRG1x5xN19FNkAOtPKG8sYvtWgkbdJfbv
YJhSENLDZ+dMbkY+y8l6IdcbaW3oe3mkQ50vCuhO5AijOJZrRwvkp3en7Axx09tpBgdkx85FMRBY
aJSQZyJDlh0McFFd032dkl9u+MUuekSKf62jUB55Fgz2vZpmERzYCAIyrOIuxdNQe1hzKr8Ctebs
O34fpxOo4l+KGjhn2YVTjTPjB3ZS9dFD30SdVboh3tQTo9RrmN0kxB9yTkW3S89yTNgLbJkrwlVu
rfTEG2DxxeSCiykRXWka4FSqbpAtPz3AOYeE5/sS0RvDZw1Xo2dTwMuZo0Btrd4bNUZHF4VhPI8v
S+GwSSU+/S/RBUgCi2Ejihvi0CQs+3e4T2pYfckfvQ0oWAhyVdakxX06rXOed7bc8DnPk9Pc9bOn
K9V3m8cNExa8knw1xZp5TtllCSbXSGLTZ2nSbog6yBhBGBMWEbpkbUMifiXorjhwQtDDldTX26cu
/hOuf/olZ2KgXHQ1NXZsC5eB4uSAWgWqhC3XZLrjVxQoO0r7JA7l1Vpn4od3YFfFx2g+Z6CRnUQN
TmuNX3aUn/64jRAxBKuzclLudjC/J1mlAwKKNCJYG/UXYdNxZ6BhdVFQbZZX69VSkRAU0nlJRdTf
ro761K7pExLawwQg2TE/WyjV7jZW6MTrnn/qYlScT0oK7FQXiyNhSGoqXJEHhzSQr4rPWmQMwRD6
lqStTfwWoFd15ikMUY9W7nu1h7qMIZdB3ml1CM6rrWenFbH+pXTr1v5jfkFJSF2lUu5lLP40owlY
VJjhh49gRn//fWMzARDuC3PApT7ENlKlc9pbFM38uFO4knBaN6IL6U9dulV5MQZ8JkOsy/2JHY+B
W61Dw7+oLxpS+fRNUu7aGPq8Uzq+31yGXhchZhVHgL/f5v9wzE7IgF8iuyRtzgHzEHNYTEy6fnye
MzK4obRHB4v2/nmhoPikJNpuvPk9uZG0rLmveDDJfCuc2wGsBtpjlyiKmsdGWjj6Qf/xwblCs4gu
A+e5Gn1x6H126V+sxLepNCJwMHVluJMk26X7sGcNp5BCOFalSwaamWE1D8rDm6lNGEJmfmRkv3df
sertQvbXeOnJ88imK9qhIZvYxjPGQK/wF9AGzvdDYMp+hSHDOcT9hRslmkvCvfexIcMh5a2/hPXW
+uNE93A44YKiDfpRIBF1RpIoXbLx22vYvtqYhZ6BXQx47BScogrhNqNnXZyp+/4VrBdUvsLXd8+H
aT6sBARxlF3JvMwl9ukyBhKSIFDfDTG5gfgUEB0OmdrxMjAfiVRCUiddoIdcVL12pFKd/TyaADPP
rqkKzN4zGOuNDyHsS3pqDaVGBJAlS21PW/aJknhsB8E9hMjJ2bFCuwLNhbV9ARWw4oIHpuRIygJG
P+2XWa+gpMuFgOzmDm17uncze1BosPznjpwHCHn3igZ5wKia+EjcxH3QDinEnlQOXWTnBPsRvHch
mw1QI1gDYoZkMM2tYBjt70FXZzmr3m306dPL7Wt1YmR95mVJtWMwNht0tzkZkdjev1+9fAU5QDfc
BPaZn+3ryQKXROxUQScM99FggLBcNO5SJsfmAoC+GssqI4g8XpyIJm9QJpltW3mXx9O0aoM383Lt
3BVhUNEXKmCu03Tnd+PV2APxG7A3JH2BwZx2Ana1T8VH17pO4zDj2q6uhr+jmmuZiG8cSdBO2yIh
pdgu9ZceXJ/yf1L4o2i/8t4Zh7Pw9Im/v/Q5q+hVNbo1DpJh2nsq7lJmni5IIbe3PcP4MZTag/K3
J0/IA6V4FloqborC+9h5aPQ+T7jvfQK0GWmnrSQgf/aJE8JiV8lQae89kBp/7szYMtpO7mdRr5+w
v2N8TH3bBYHFHZA4X4TOdeoyjJ+tYKgjwh4hq2yrZW4VubtywroRLf0Jv+F33MNaIQ5JjPrBfF5B
7XkAGt4gedxJm4Mv2LAXc2sRx743aImd0/XppRKjgV/O7qMPgE36dcVF849lYoAuv1BH49bbLE2q
q1xrN2rvGGxTYsPc+kgnvqL4pJSYjBoaKk1qRhpbHllSEYrS+JqOwwTWv9Kdd9vhJv82eCNyQ1+O
whohUvPAPFRjTiLr53nKukeUUgQ938Xq7jf1xLmf2xzkQ+RVtx2vuUziyB/2sdvm3Xtxc5EnwI6Z
TrPo3Jsb8E5tf4L/R8wBb6Z3cLHebRkL1VB2Jgq5ad5Qr48I/8OMalVQDx5VMq4W3Sf8ya++/RG+
xtH5QTdEakCvNYjIY6sjZzVIWIvJ6+geRqUKqeJ2518Z1UiHWcW4lghnyMcQZj+18Mj27njtbEyH
iQ3es/mOO665Kqbj8ty51Yd1jhoTS40CWmpXrWTZV/SilaRYS+uUWZNtg1gNeph+G+Aatiy1Duko
SkWcjU+L3jggDfyILOAvJhq4vUIVUL9eHRfIb+z1XKTR/lYrcaAUWpJyQw0ulV76bcSTEps7Rvos
CbNO/gSsymPU3fsQ4SST/94Jf4MD+8VqZ3rRRp33tVzEDnldcV452jzZPi5w+AYOJ9Qnqg+c6Lcv
EQ3DM7Jyq9oT1ec/AY9xHxvOkxD2WvsioRzXr5Sk+IZ3KxfId1d4Ce2Dt3yit7sufHCm1jl/wqcp
ccpxhsJ8UjoRtkrW2JVFGqXkZ3SmB05xjGIWmDyOsY3yWrU70BH9na/Dc46JxAwwZrxi3xCiVZrj
6PzI/HkPfgdZE+4oXzq2kjNLVJUAisBLphxXHtIUECr+34j+B5U89+7yaLhml/xofO4pXwpITCSM
9DB9wo5mjX/udd0Gp2+9GcyNut7NkWkFM/5j/DcoT0KUfrEYm52cOuOB2Ysq900TmNVLmYQvvGNm
mWyfFKM7KoAO95UjB7fiG8pmxWkcF+dkU0fwkK334uCM9KjKSihlMWSpPNCq5+rIie14c7Rw2jEh
C4lVAhV5X/NzOiqXq3rgodw5gel0iXAMpTMw4Zs0vxYWlhFBmnOBfmnxRzDdpjOZGEpl67GWw56H
yuWs33kkzF9mWNr0NTYTruAMxqdnaySYQHlpSmr2fQ14I6ViR5pFGiRoLdP3zqxzFE/IH8FfTYWj
aNcxjZvL5qWhA5CdAsFbn3KOYUCXL+OqA40EJvkXxcBMGw2eWLSGjbrQ81sIkRX+ywG1o5P8mse0
gCKuSAetBEnSaVQy/i3w7fYrE7bLvSJ6x4uhE/HZoNM8vCK2CrGopB3ZHCX5K9orSYXgV+F1vPPb
0WN4kX7Jjrt+2gp7hmenMq1lYHuR4bN342hFIKc5aeTLJ6q8F3VTnvUXrrq2a7Qx/hC94Z9Y43aW
HkV8lZaFwZPKmPEbOXkDx9olvgLOJwGht2VlXF4SScjGCTTB0k62OZecYjYCbZ7Z4gJJSbEQy2je
71KxjOVWE5MbcqBU3owz9uBPY5IpW+rpu3bd3i4xfkpBxJ5S/vu4LIAY3AdWnDzAIGmHDSKOXClh
ReW9dHjVk46rA2ZaoW1SUdjJCFqlIdXIfXDHypMxxduKHlFJu0cU+Q38H/C3IyPpPBRAXsZ5eoT4
04CVBnmXnFWIrX44udhRkn7TpBTIg7nvEfz45NsWhImT8vWLbwKX3IigMHWZS+yi82Q8q/OSpBvV
kJa+M2BWuTW6+3HbzLoX58F4JT6/1AZvIuqLvRqhrSQptS8QswErn0HGCpt8iegNvH0X29zufu/W
D/EUEYQu8wjHIf9YbSIRnxsVk3X1H0emBHgfmo/E6nOiKAtTqLCjWwOlWtsuxMrEruyYcmOMpXcj
2dqS6oYCjiUyjwIcsUbCzl7F80UErEi6GZkx6Xhy5YATBIFTdBbzpscNEIzPOWcZdZR6O/drhkSG
BsPqtJLLxtlMWw9zwBAyGFNUXbzBko60NM804TdzQ/VlEYvVNXnoABYCcx/VT5otSj95c9Wd6ETl
znv0WcZQXZU5FP+y9SR4/5PPORl6NTmDEtyJqRKdJ6JBcIGEmY/UYp0/XqDrK2IwgZtxCZclLBNi
XQ2wutweYGj+qKh77grc+43ua4beWbEDCfZ3UlE+T5U91IR2aEHyLqCMpUuIlSyRB1EvsqW+cX7R
0l3Ujm6cDFrLY0AgaB0/aMx8xUFinlaJJk6t7uXJ1vFCGYMq/6sqDWU7sFGZXxtKFu4eA53vZBWh
3/jLr8olk0IA3VM1eh2tjD0MNl0DH4FTKK3xfoatpX5EhS974UagnZ7pE940k3COOvelGWk9GpwU
UJZpWDTEuOoifjDMT095BvOQx81wCuTpjttJBAM45mucbRW6xm6DK68LQS1E04frYg2c5iNugYJ2
6WJUG9DyvwKPBeExjKmmF/vjzepZV0PoDDYDjibPq5d2QxxSoYK9mqXutWm3CXY1l/Cyo1dOcvRb
yJ0+MLuJzgww44yNB1SztHbDZkVtf/VEEibAf4VEzKttVf3VvJgwbCC+V2vJ7GssuKUJ0MMc9yo9
nH6nRE8Mpg6OFqwo5bhpM+zgUoNjZfesIp2yiNZQcYjo+M7/T6WxVjUcG3VqJgmSSMst0Zr3Yj77
Z4dc2OA5uBGi8AVd3h7QGdnjssBpgW2mrMUkInD3D2UIlyUWMUtu7nkcafNZJ3Yo6LO1ls3CYeDb
P9ODbS8xTR/QKOu/X1m01ltDk39Cptp7utJwRve6MAElON16+sXLLOa2hCFTp/3F8+xQh7c7EZTb
9GO1g8O8sXqi7XIejyOlDCsyA7oOkZsFTh5TGvxb3hWXUbsLU79f+dqig9CCgic0W+HCfiIJytD2
OLIysqJxm7rh3iHLi1kBHbOQ61BqIQNm1GIz8F6SyoAomyuXI4Vc9rofQXucz8dyNuFP8p2KEJt2
LexdNSLjuTaVsDHSv4ZRcg2SVf4eN1KJnpMxFKpNA+W8pRe4zNEyR9RZFo3o9d+xmMn7vVCjaNvX
O6Xu+wxkoyDLbrfDY33jPGD36ZqMWNARAbcmfgksbSdidp98RVMujQW+ReTBO+YfQ6K3aigh95KE
YJF6LpTSpG6DVfcSHNhqIDBkNEPOmSDXUndBcfYixavhNye5kdqeaS/lx8KuCDH4bQ4YdoeHOMVI
ImOigPiYd+vVse48XGVIx9ICloNL1uhbJbgjzSAFpQgsvXeibDJ4OGqOfjGy4xyKZXHAGjG4uESV
6yWfva2SlK0YElVB6Hglk3xKdJ6FZiAbyIhbqUG72Df7g9NJEShjC+QAt/uVXOsPpcGyvfn53avD
qdHcm/UoQbysVnlNCgs6qXNxKllLr+BTHM+TvjI6KR/nnCFijdSqZa8AdC+AXDmMCSdYeV0U8hMM
iV2ZEQZQPmfDK/a9V0uGsBio1qBOqzBTGfq/zECBomhV4Q5RvlHTH1PbJbOsEJjVbO+lY1dlZLEG
6x35svQ6acS6WcNk+Hsw8z6nzTUaNqcsQNvd/jKa8HJfbsl4waxaaMR8VZ0v/jepnD/JlbZj+gXc
hkXGjuzCfeYYgchj4P5UnlRRBhAaWV4nauenAiygSdn7tvk0R0fw53uTyrwMKWzAygNVx6vbEekB
XNqpQFTigV1hYNSs9uKmVU6Y9ZwTah3nywEd+HA2M1bHm/6NqQYbekid9FJwrszWieL64E2i6r5n
UlGyzhbsfJq8xYpIFcwLXEN/K/TXfJh07E+EobyPqaaA18d9FmjhnP3OGYbc/cXJMeCBMm6I1NvL
3iHAV2FwtcQxSK2oTDZfZ4XnzAIYLzREAhExjyof7yUgC/AR7lnlfNwS2+Y0IFQJS/YCBhpHU/td
7yURclchoVQdYKJX7vH295udJQ5iBY5tRNkf9Lg7PlfIGgk6B/j1UTPlodXl8rrOnGrrX57ikVPJ
iwW5Vx9RyGxgXE5CPKxQ5foqInXikvv2a1EJutlqWbM34HOKayHCpB5eEFN3jOKcYJ1rwr12vkM5
cxRkzzeppW6TifOqTbS6Y/VcUsHWXLSRwPhttGy61EX3F4XsbUGyjagANlMxOiBvHMozwyLjvJvD
MEkFudyOAwIcHSRsAM30lzm4CPC7qzceULBXd6GK/n0SK2EektEXY8+sM0DbNymLblbWzl/Qd5am
QozlXDw3czS30WHSsONQI0XWJ/7KR37/UfYg1ZJ3/Ygf09qNAVpAVfsZs+pC8+tEQS02uEI09zVM
0QcLLN8dqvtCyWoOlKSPE7NRYupzIlT02UwrXkrt3JwWmNMi1wRLhLu3VEL/43f2rje8QCSLQw4K
nwszy4NnDqW9Yt3BwwVzNAaA/1DmlfqMlrtRCNA8Pud8zzPIYvZYrnGp3rjk/0GUCWEDaF6NiutZ
d1z2QQmdTQsUcgCaXitXj8oOUi+QRN8VNvdBZXZK4/tebmXsyA4fJv6tJgNLvPk+6UPbRxXz2a+K
ltUHTQ7ppMolyLo0t6li/ubblq4RMhaQLFTcaYp2XqfOsbxTGGCMpf+t0hyoPqtTgRFCf5mYlmQ/
QkUDNAqF5bpFC9IACcJaZ9EOx4d1/QE/j6QUZnV1as1G6dSe6HOqKICBhVjN5pq9D/dM3iooor+N
3UzmKfw+Cgt9oSNQnXy4MYeyL4BoVzLUd8MkbxT62ZWoMjksPy13UioWT0P3n4T8SSP/vs5teMEF
bkX1sMEIzu3GfSbyd2Qh3g7ekKWCB+kyAsR3W8W2r09n8W0JIiPndS5pd9tAi+1EkJOlwkZIcF8w
RgA8k26vIJpOI98gSAmYbsMVucVmuVjloNpmAoqPYKpleWBff8oXDFBO+6UAhR1F6MK/Cjtopjxj
3ew0EYXqkWxNn/sH04gBnEZDC9oRYLoWNLOEog9f8B4ZuklWpFN2bnmBFeku1vF+Hiekevj1QL+O
ctCtUG+w9ipH7dtGnDGqsyqqMayMJqnY6H9vadDdTDXgN8vLFkGeREDgxt8FqG3DCgeCUONogejZ
5wmkNsSa6NsYdAXoYSpbFdIj4jEJ0GXdg+jmSiJkJD1DsAHth1v+PuSQxI62sPLyappARm8FQ4+R
O1UlDqfaJdSk/avf/7inoBwco6eIH+0RiwtGSMUA3wxL/rfUZP9oTLiKhLkt6rXgrTuH0X+gdQSQ
1+DsrANGfYrs3pLqX6oswvmBqXkTM5yu2TpvfNVy5VjIEFTXZH5hPdFOziGh1D+tuqG/iLLPNKHI
lFr0Rq3gelLMSwJzCu7oDQuZbUW+uLghjuX1ogXz/pDc30tY9D0I3TWD2KN6/KpTRuRDuHtDayQv
5FmSv2CM8G9s2dc+UfGAvqdmiv7Bl4t1oRgXni8BLWtBgJFEWbRg6s33uQuT0JyiKkJ5KcUyFn7f
uDjy2LkdMRM3WZVUkAipG5Bh9leOuiDhhKKDjNe/ssKBFJ5dodJxCMEaZVEka2sshNk9pZ6iIZgK
EAy5+hRCcXxcFY8CHe/vZhDFAnAzv5n/wOKp7pCjEp8W6c3VP6btSmtkKRqp8wlFm1eLzxN44Dm9
YLgTWTMbbsmxDxT+mpYEeFprQDJQ06ULJ5khPV7reg4vZrRLDoBdQQNTaPN2JypcZE7Bj5VHsJrz
4XBhibwrQUqtJm54BOakhkShnnWCT29CihEEbKv6YApaz4K/dLjVQnMzi40Kmw0nNn+4gGH0UAPQ
ExPBJbQSzpij37lcsR3lATy1MwxL96OauILpgMgkfEr645lb4DmNT5AM6ROVoQgTdMJD1yX+CXSI
N0cF8upojH5U4J4/XPYKqvrcxrCUBzTy1V6PNQzYvk0+Y2Ps8w4o+Bv6NaZVcChW9IyepRqwZZRF
gBhcqKGhE5MYJSFqcBbHNPC2tx//gqrCGqC5pn9XxSWPm+6KtNkCJwK+W+sK776CZmKocjr0W/lb
8GZg+lXNxgHw1P8Y6exKiPodmAFm7vDRAf+SZQ0BS8IYIc2yG5+Xi4odWujyPHVgs1y1ndJ/RTvs
o2kg6mwMW8Qg7ThyQi+PQdsgQwF3sB8hB0ZfokMU14aHM+fS6UV8UAglaP2tSVi0kQy6H5OY3fhO
HCV+8gCzcHO3zgrxB6JN6gHDrNv76QNmNLYumsRND7gvGuqBeuJCzeJlTTrpdj7v7Hq1EdtP3IQo
a928UghL28GVx06cax6BMGc7ZmnMqRcnCNm8VyEytrDBjVOsix5hnJNVUN+DpHya0+fNqfwxMFs4
36TPQ5h0vJDR68ApkphPJuu3MjeyGTprJZIkDABagVgHBFqmRrJKt6Y+y4546nFDIFPyvUsiOoM/
D4NFOoatpv8nN0ygG2dQFut9ACI8ByKZXUxlPwK9Ri0ynKIXvYh0dJMbjDwdonfEKy+PBaTsDrvc
1nVwUCB7ic/AZB8k1O0HJMcGxxyNBnkldUyvS9WLdFojZYYFK1/2iWw25ptxK/gXV6FeS6y71fsW
2cRRAqlhAIzzbD/P0/GUvuv8Z0B+Seil6XlIQkiTPeSpZjErNp3f3PuPjP41GjfpHowaS8Lvs/2L
VnJNZLev05gaW0zLHz4Aeit5KFpuL1GrpVO7AkwVVxOlxnQ3xUzz4aXzrBcmj4cGip/gjjQ5pkEP
th3IELaL5eJYonsizfDormQregwqJ7M3rmTB66Gl+5CHZlpGdTF8XgcNk2skFShIAggltKMLLAaM
13/pf9jOh0MRF4v2jGOUE81ZYJdGOgqrrqQ6a1E1EryAhvCZF+KUbKuv59lR5o+GAp8WX8O+d6Zg
h787oZT7JrnAhnQYwRQsRgPhsRGj6SdtELE1ASk/ak4GnS6ls5E+m3cGJ5dmb4fBi9CGtZBeWcjJ
Aooq+9Pra/+RedPKJCh1MmU4vQZ+L82NkwpjpFSxVohssj3n7zsokQWLvMhBI2bBpVWZUlnYkZkD
d3EkwF2gFL/02vT9aLKemo6F8F9xV9Vg+o6aihueAvbH6KstmwJUL8N1zpG5MPcyI5hb6kQX63U8
lekA9beatb4f9nWbfxOYBXupkfAhom6xrWLXerE0uXRTvEa4YQmpVy7hbSWTi8SEOjG4T621aJTj
O9C4ZzHhuD/2ja8CQ8mBVHSZs3k79WNKQenEDLSSioruNOaY9dIoVMzC6OC+V51ib1EdazJ7tGxB
QUb042qcVh0SPrL16Sgzl+z2B7EnOxo2HoJkSR1cVhI3Yiz34zDbvKB8qpu/qiG4TP9VVRh668Iu
vbiQYCv8JHQmC9gRpw5w+NneNWw1PT74jNvoXMsb17alqZ6ObJ7p4FuMM3U3yvfkTD+kYO4H/yT8
r3THBY8iPcxiKKyJBeyR+ei5+G0eyW0j8ODw+R8f4OP5GYb19Y3ulhiYMmHqWPmahv1dWjfaQpPV
uoqhv7gXBt6uREEetYd1TujzcfSd2CuJ90BnLL+SDLVHPpwZPAhAkQp687cWK2kFHDLxWPPoxuom
1yxTzuQjDV6CsaJnO6tACaU9jRV+E0yx2kxrX+v4kBtYSZM1+rQ79p/F+a9Kwfpj+sBcRpo8wiOp
9BmeYtiAYLT7nIPWgfXQfop1RJVDYI5eczbjm0cLFZtynJrvgawTIlPOrMoCRMA+3PnTNhVqq9YM
AKRDiqwc1OKQzfDE4G8jlHoA0DSnq3bbn3O04khjHntWGrkB+1zXG/fNAS1QFX5wZ1n2mk0rJ7r3
opttIeuJIwFlHP7VKMhIrgaFEzqT0paqVr7BnUR3QgOxX9/6d8k6d76O6P6ZkcLp1WRi5fBVOWge
cLeG3g5fl18bbeVOVtVRmyCX/k90Rvoejuwc+GkJmkSMBPuqkLbf2Xo9+/preH0Dljl4ibFw8GyH
5qV9qfr9+SUJZkcCFdNxbxG41rZXqTEwCduyHKLUr5Fjg7vtfPa3JMNsh0Waagj9s6XH8783QLeF
SFzn51tsYz86HRro/8qw096XbO8dgYUvx2AbZg/JoTzd/KBRjR6wwLQaezjQSlyy2hBkEVPIR+su
MrDPzBYSTP61AZN1F2Y+z28c4Yr9mQ6vMTuifkmiP2t6gFinjyRq5gFKBU4vjTjKrf/H/hTZHUYH
WZYgA9ehQhjELEBGikyUCnJaQBXL0vr6Ofy7MLG6im46PmghHhNC4XPJYHua1jBt0vgVH0qVRe6g
RfgZF0QTj55AXz+VPljWPCKiit6D/pJiA/h8s2zpHP1uHtxMzO8z3uYUA0Krkp5q1CEkEXsyS4NX
XX1ojdhu+i9JdMNjWFM0YsHmKPj2zIMzg8IQ1xf7Gxfyro2ozWsrVhsQsLCAwob0sVTtqp2Weapy
f8GZw7DA2IHkYKX3xfqkWCjzbcwgDnkX2f5pv7rmZqe+ChNNJYIgpYjhkCLZ1wc78hJDGL1pept7
1597jvJ+oN3NXKlomZOLIYDgX4uGvAHPmgSgq1MdQY10NwUgx1iJ6PfmhbGzBvaZl17aqyJdS9aV
Cqxk7r3Q0a0oPrs57tBHeGDOaZuNVesDaSAwdJCozcHfH4u5auseEX8qwtO77McnObse/pf5b1xR
DmVBR19I9AWW2G7xtnr86Iol4/31vwiLJm6Egvq9s7ouLQKMxpWdPUAg0ZOhea5lM4knXVuB8Nwh
D+47QN1Sutw66sFKRmfkp+emFozYvOkw5ity3+deQN69E4OBC+i5Q8abCx0CGV48//fnuutNqfPU
JKhefwHSjt+eMYgzN4nHFyNOS5wLVoS5oa6Nco7fn+1i/a+7Kabw7HDjJQxnqpOLlhlQn24RU+EX
Gy9n1q9uLR4i9v1f/LsIeBsCyX3DCposu/JV4gDdngd1Q41Ioi/TlyDE4iKJVzz5J8qO3gfFo2ma
8MSBVyqYL+1nTLw1r4bYbzX6+coH95H7Vc/AwFhEAS4Rv3lxedy5WFE7i6heiS6FjGdDSncGpfGs
XfSL/uQ/94u80QP1dcNKtIsVkTISEyKvG7ozP5UKKHX/xaE19S5ecp97kORBwxUhVTtyQeRiancr
dmwnd720cOAQuWqJVWrblEHsa1JykZ9c7NSgSasI6BIzmQyJy5ISQmIlkbXnQ6hPYeIjp/oBNRF6
xNYvNzjcXmgbrZP0IT+oJIEXpq7F/qZGquinq70DcVVWZrEcaJh5UxahxLlc9G8eWnW0VL+bLW2f
t8/UafXW5vrVIKIJ9vH1mvBCqFUI1EeHIrjvQ8+i5q1sQ/ieQiw31YG0BPrTVZT5jRGLb5HDIFU5
zDxHJLLdGJ30FKDih+g4wt9KTgwmjOypn4kTipVai4wQaApIdcZq76P/097K4LqxE6qju8iTcQQt
2koSz5uDDvGH8eMjhHV2CH5L+gxm/Jt3yaVW0mgZzNbKXiIr8m7PjXZjzHn4kjyuvCN7p1zafL7I
r+iA9NIkXoTqRGF/zBj5p/NEHdVmwp7Oa/KsWitImeuwQHhs9rd6eHEhj4ARAD+NXSHl0Jaae58H
wSp1HT2Kf9u+mJjWyjgcGIiqcNGcoxrS+0V486BWjvqsbuzzYsDjGmNG4WGHKHupRDYGfyNUQ0mj
dRgiUAmwy5m8lo+rZ2nGuD6rR9MgULJHW+To5xJYO0ogz1gDz+JgqIoyi1UJiQV5uqTVYC/tD49M
wkS22OTwbniXYC1eGpWeChEhFmdKk5+DtJglbvV6Z9nkYEwy1D6eXdAnueZ81ymWBS8//8cvGRk0
YNpmKcAU4lszzAJ7vlwa8XbMHakf0u4IvQwz8Kh/H6dKMBYxj0D2vOxDF/E811oJYxJSZ+ttWVsz
U5wjlwW0ymK1Il5GKgcJ+xLlFaKLxHS7ttrfcViAHRPzd20qLBQKFqFg6ttAclWXb1h5ICxeGhQw
at5sUcP14//9lksnoLsnqXEmDbC6hoBO0QwFDbXtV77gtOkJWXjZgLXV/McBY3UNMgS32+DXoFd0
UrrKbZHYxmKgja4N11UnEPjrY4UPzY5elC/TlhFu2wb5BtjLjFOpPyg0VkU8qafBxQM//ONRMGs0
ioV4vmlkVeZ0XiMAbu5rH5ieg92NCKMo86Z8K++v9EW9qcTGyKgCxfDjUFvYZ0jVbZvX5sQ0oo4Q
OS69yZVTKn+AJxo5gfG2cvmeK4mkKyRCN5EupZrS8JoYWP7lJhE6jO2gtoJE5wvBXalQERVvIsIf
2U2l47PBPg+NGMLxp7pV7ZCn5/W0VMv+9lVypF8blA1vpRXfD6nCAHUk40fVFkL2uRn7LHatl4PP
t9G3VHCRg60QxTax5BpKjNpdJT81RH+99SJtAy/Z9y1HOu89yUJ/JvYy+Jaot3BD0P+cdtxvsBZJ
QcOtsvMU29kiEqGDBuoYW7AMPv7yhlG9EH35AifFHkwEgg6UE90o6HasG9GZRiwwXkQBhFG3F7+I
sccbfUwZfDN5mP4FghNbDhnJHjdD2j9MAHSmO1mf3mQaMS5VvRs8ECbvHNa/7uyuQqjod+6Zr6pD
70QteabDK7HtEqfFWmO+ErSxwqu0wLcZv7dkRfdaFXsV7sBKO31NyrZxtgx4Bw/2LTXRgyui1Ayh
4+ZZKScFcA8SEUibJQJf2eBTZUfs9OMkTqHxaTmbEUjNtW/IdcXiqTGwzen77kCvTu3XGG3jpTik
qMgzLzHxJxzItxAd5XiP4BFlunVYhrDyqn5LN2s+No3/Kg6fUKzRZYP/iVxVyL5U4F/MmBW9fc0K
s/eF3FL7Ipjwn3w822VQveTOAqzfhzaxY/lNOufAObOxmxFT/XCqNH7i3zqPewonKI5VrBgOmKzG
Uyv30U/s5gjCm5NHVu1669d/rFKGd+nQR3SdpeTVMAs5PrteZ9lVGaPd/ygWY25+RnaW/DZOKeBu
+afhpwK26R6PGm10hT5/aMT6AVmxYmwdsskOINZuFA28M6gEHwGx3vBo1amnbBcCoB+7SIDI1V8l
LwcIFwsv/E2TD2avA9Z5uYPSp2W2II9odYtMzcP+Bngz1uLpF7SrDSIRtY2+msCDCR4dI/r9zTbx
R8uxpf/uil648jCpUN8+7LPeXR+rqVJzUymvebOyiY89MZ/0MDPFxDDWzuYPUuPpy5yhTuCzLpMO
8dsmsIzIfZX+uicxKhlMFDuwXZCOZX8l2EKZXTJHsBr2zgQVdnzhNhKXdhvpQCrqaZxhN9SxzPfd
ZUOB8ReUVMYcKvyzccDtbjyugay5q8mUSOJymysiNEGOlyXYJFdYRFKPVhU7lNokr6N7bpUnwiuN
p4LoKXR5LNUAjEx39myk8rWy46s+XFL/RiL7h5Wv0184Q2ALoJB0orUoYZNpecEBPxxcOp4aeicb
fDCDpQSvh5TR2CP1pHeEJFL7IUctssYYk5INWZeCkXNbogBkLBp/BZ9iJaK3co28t0CRCwuTICJP
PGsBdUrzRMNgchjhNKsl+JChIWjhxypm7UzlDdjOYCLM4De/csZlGa/+zCAcanPf0bBwDSARcTLx
+ATrqjX7jDNgd7DaPTrXbzh+WIWCmFCeHGsOUv1i1IXkHKxkEYzIBQiSKS01DhMA1bSKfUY28bMD
mU+oy6BX86evrGqynf4FTzMqeIyNBk3xRQoiHLllu5x17evcQJpUIcRWopc7HWb3GJ6AVIg30+EF
R2HoziDU8AHajfaO6jhue2rG/jaJEUPLshl54pkgZ7dhjiXDtuEjtg/mO1Gat0Mz6YE8C7o7z5SG
8j3W+pR3ic98s5uII4Q9H6SKOzxjZxiQz/2QllxEbgxunfjbnbiuNl7OaSHJCb7gL695DB6IwRa/
UHfh/gkW2MZGIn0874eMRwa5pl+RPwOOg/T/K6jH62CKLUPPAo+butUIgA7GRL3oCchlse0WpPcn
z+WNFgULtT5R4Ra0oZ2N99M9bvfvNcj63STlQwO1S1cBPLrXzfwN9fguSS7ib7Y+j8rDTNRRPRki
xM16+4c+x4Sf+TOrCMRD7neqmO1o5Ibq+y+YfntBep5gpuHmayluRnNfK8Q3x78OTW59mJbToc6K
sQymcb1F04LwH7ehuRxFhL0YRDLR8lw9Fxr6/5SZ8V9ptOGwJvfvtaTQ7NrlbxSWf3QHaosPWoI/
WSVu+LwCXQi67ar2bACbbgFrIem+F/Z2kOgqNjXFS2K19xKZqbltUOQA6qPBJ3lRNF3micWLATPo
IFX4XqkERZCEC9op3R44dcNvyBj8cDukAq0DrgYmrw9PQVjJmIqqhvd76A3NHFuH5dLUFyZ0zvkL
AKJNWWUB7QIv49sYl7Fr3nQnXNwPLMcKoOimZy/dsYVumwwgXpAoo5Ym5o2KMjKhVu3W2wuM1V+q
tCwjVxWNcegNJlwwvRT0CufRZ1j0LzHwkUzBANMTNF1q0r5GfQ6JFqv8f789uyp/zARxVsN9Q9bb
RuJDRtFvmVWevEHARbnzCReWT2h4iMOS1Jw8xQ8QJbHrVZzgFm26AV6FmP/xUHuA5bTBIpZC9iHY
9XdNfodOKziUNWMM4lsowUVDB9JKodD5PoSgu+hsjRGVhPniF/3tnW9hqqL6zAnU1CSiplo50PvD
7LIeXf+fpbjD+GSSWl6dn2/JN2oRBSkATeTLiCnp2m4ySBxRN1erOzGKBw8B01q+xyaX7mJySjMC
qoLKe+yjy3C1zqM5h9X894vn3Wejod6NdC1yGNaPuvat8iUEAB1DsXSswIFDEQvCixRAi2jOLBps
4onFAbHb/pARoeb1k1doKxM+XGtqCIywc+5N2ljplfsXRluk+WmBgeQzOoxrYuCHbtvPEaj0hXzN
HMANpjjJzP2oCMdyJPt9+suExhP6mc/SuSzmL2K0fAjtNX4/TdjIk95fKz+rX5xbB+DjyVd9RUP+
exfgP4ug8MsEd9nQ3kr89KlRpK1adYeK51wFx/x6fIqshCh6/CvhiBWQZortkEU6pZZwXW4RDW32
zzDHClSIXs+9+6Qb8roTgpET2XacaKjvg4cgza3vj+xymQLbhwRFxxrEmfcF/DcbLY5ZTJRngPfq
rGdMVDwi1JNXNdJjCSu8AmQ7JZNhtGPLB3vz9yxbWztMaAtAQURQU8h2IpyZU6cRNnttcn1wi1Fs
AcLsFpZzFtbut2oKghPQ0bij4KlKra/G/aecdk4g8c6MOFAIBC5tQoe8k4oktaKPJpUS8fx/j4Rb
NK8LKLGlnsA5nRB3KSoucA/AoB/A8qzKB7+GCUrfJSgGbq9IA+nixmo1hqhSo39Xm2VRBcq29L3p
tWET8FqfoShESc5EcCQ2Loyl7I2eyyVxURmdq7X2rj8nN41AD+0TkKVFAhckM5QPo1xGG3MI3VIy
bUD6H5+nFYJSz1tA7395+S05l+QKD4dSeVL/7dEeb7DQaQIA2jvJRW4DDl4Q6auqmOeQqtLx1IQ6
hy4eGoae9oe00+c404G+BSf0g/bP1R/B8wW2yMJRr2K4yCOpHrd0BTDGSJEIaeAHzZVPj+hq+d4C
8s5ThW9w9m+Ht2E3gVfQ8WxOrunupZIBE1OFCAySNaUfA1ybuofihZrD0x7ROcDIyrVILQVVJ9uA
ugzVrO5NXenLMlc0jaKTMQ5nOuwsLFafByt+6nDTIi5oFNLT/zmSdswJsZ341PW0urq7TTJn/dfv
FUknfPVpKb/JuaXCJI/AeB430435FlT1v+HUx9J+Lynu99XKyS4cegBbkJQwnMCNyvv3HrLV/wvH
/AIk1UOCw43zN3fqHR83OSj9cOZX5tqkmDvpI+ixpdBlNwHamHdPcGEBuGFpCPfjc+ECLfoLXQzj
QuzXr450lf2Tu+ZBOYeYl9SlqKgq3u2SiV/EthYcew9+H/HY8koiKE1TP2HIYVaIs6CT2c2/hKfg
stk3vBgR7qcXiz+pHaJLw+xNlfpElAanw4GrrCR8a+YKbW/5MvFFIpvkd4ULPdYB53lxpXzkArHn
tbH24nlfJ7GWOnrQ2GdVjPnF1+Cy9VYlCIcndM77m4wkA6DPXjJ4Fg3KvcoF/7YdGa+bNQWeBzrv
VmRbEKp8u6FeXT1ZPtZa1YXpuPlyMuyDwbpqcco482Riw4yPixO32hi3TZtmDUb/cRvQBFxE3RGW
AzooF/ujzmJWga1NrlM9gFQW3RIGd5xFXD8zk6PPB2tUAIcLjP1wKpWUTIt4NZYT1Khj9S7QAlSt
HQhmEYTG3O2MEiXtu/OBog+h3uPmXTTKx9oH4oDipr9wuQ6ITLrTg6x7VjKNxK7N/QwI4ZuAHz6l
75NfB8n3527eQ4JbCsSMjIQQ9oivXmI44uQzBe//n/+/qUzGC73z2S4sv6L3UeqzaXwV1Ov2Ru5h
QVj0CNW7u5DTNJw6OnYZgCS2atqjCQcs8udAyG3FgmadhuZzKGmOxWGwbHXjbQ21ZCGvmYjGfcJU
dPwrCWPK1O4wTfBapdNLDH5FPrLU+5s2qXHdiUqvPC/wfuP3HX7kM3++lKv5wspu8EXayPPa3Oj8
ykP5zdQJjfaY3N58anGTks+aV1lDVEePHSBFXSEUkQHgbRu9/oAZQGM6ybCj1vYkYmBvsw7O5Cwc
ygfGS/L9ZoTXYSm1VoI6sMkLhoz1FBzewMoYI9U31NXsZ3A00FiH6bOHmirmOcOxFuC/+8EZlm+K
ZP8kkiy5SX4CYSIUlOCK3wlynHrfI8Tzw8Uj6RN2bmg8aRWcooTbAUU1NIj93CByHQOhSpvobAqT
sTA6RXPQ5fn4E694rk6HxAwB8Gn3yhCvOu7IQcxD64pYGex3uscvTCxpLPh/nfrSlYP2fiCjPK41
rnUPC8JQyTjBgHeyfq467B3SghBD9mEhR74t3kP//sM+L1dHAMG9/pmPL+1Pn+vuNzJ0UAOuPyqG
iYl9x1Eu1quJsg3VXSScbM0IuRpWuFPLVjjQpxSUtrpFMYmN4gvvt8i7MI96jEd8Zjh9qlH93IqC
hmTikmCtoQWMAkS/RqNqBVticiCspeVoUAAJI/r2EdLAv9kMGQBfoxZj6kXJbVrwEiqiJdPxxNre
amUrDys79XMpdJj5RbwXolo/zpYyIi8lBqbMKKdYgVpt01G4MjoCcw9ma2J80f3nwBy/jIxxUfAE
eWLSc0k17efI6eO/uCH49dJzeDtn0lJgA2q4SJ4aFKnn4SCffca8hiNz+sNFOaReiAVME4IFU2C+
CMOr+4RbtvHZdtebCqBwZbzWzFqhW6KOhPoDyuYr0bmnHQzHTte7ee5nWVA1gtGco5TMRF+lYjfc
VyWjlSFXWw/pDXwtAoJr3v/qcIYAzMQONos/ykbxdn6AqyNwmPHKYN4ZdbCnNJ/uznOFronXv3Mp
1g1EBzS1pYM31iG/5IrJ/xvOiyXanLpO0uE/kmgdbapvNv1kFtOZcMPsoO3SG+v5iHqlrfVzP3Aj
HSfFUQbZLHTT96zOdCf52Y5Ccefm6hvv6a7B9srbBKCxSpMfVuaq/ADV6dzByC5t4TBxV8gbb743
XFHd8U3LvKVOZctTVQPhZhtsLggnavBSOBihx+I+t1Y3u0nNfmIJvrFTYlhi8nKb3B+2iE6VK/zr
3imOZskO09eUVwjGIgD2SSDw1pq/lQhSEkDmq2suwdZvR+6fHR99gPa7TRpu4tkgMDJ7iziHz/rj
i/cvjNq0uW3Cj/1NVW7l9X/llF8iNZ4NDzTSGA9TR6SeRoU9RMtc7lsy1MlcDLs6ql8WLJSQOywn
qK5lZypzyLNjbYj+TqS4OZCy5A57mU4KCdI3D8dP3Jao9anWWKvTKUTTfZpC137xb66G2d0rIU4r
n1oPagE77wr3QH+pqMv9UlNPn1Slzjge9Q6DIb6npZhmXm9IMc4ysB4f1euSzLSb6xqvBbIOU2ZO
g3HdlntBZkwWNRBQzE2ic0midPKRT/PKCR0Bbn5h7Zika4v32Ynn4/RQ/+PdCqXb4u7ZMGvhc+IU
+DwUUpbKVC0YoJW4GdJgfh+uh2jsQB4ypzdzh1wxbGSrCUvpnPE2I0m/e1/Rwf97YkfHfTuBfX5X
LHlXrHZQIJ8Jsirw9OPfNhcEKF5rMZPUm8GHmvAQCQCwjuE1NeNMqYtdr36sE2k1pZgRn4GYujbU
Ks2NL8NddJbGUUfNtRUYY6MQyKd12wrLQRJv6Sh08WwAXPbXqznWn5Ir0AvIVhyimACwNr1kHSzp
OU6KcTuwqC+3x6JPJTlCMUt5Z534mK8v98iBxTQfhhQt9Y+F0YcnxGfwyg9Pby4bZEZUerkneLmG
vMleaMjbc8SQGyLwXZpuh2gUAy7Zisoyo2BghllXQUS8LBXrV72zbPJ9haJwLbvCdHpZ9Ggl3Ton
8HW1K+9iVZNv6JrrfD+p5XBnEF4JrAnc4GYa7PwA1e79pjIaM5wN5wlBNlErBWQCu2EpaWhjiMah
GB9JqDtaotG1AA74UHC+6t7Eyxd90iCDI680SNRkrdQ4aQKBLx9g2ezVNdJMOplSJbSayZo0WN9I
qHRXqgY8TS+DKB37IgVCb0rwOMV0yN5YHKiOTZ9lg5KgNvL0fI+8YOWtTI9PXlQi+Ss4JDCftmK9
vOEVibLkgY+9k+GJB5wUSIDaQ8CnwcxVXFvrnHccWU1gejw5ePxIQYIGSfR/ozx+HLdkho34b5wc
1K9KR9ozgBihf8pAQxrMUbtzVvhyf2sAgzTudB6AjBPEU7jjSnuUPUeBNw5K9GTNmNaE9LZnnWPh
tf8z9Qg2uhBzwqNoeHlDnmR3zd7kpTSML6mHgF3e2DRH1nF3ZnGuY1kDupHw50JIuPTKNoIqZeRj
APQ9HSqJYcCKJVFfltgLy/1BRLywSBGZJ1JjHrsTJmGBnhq6FlSNN4AmLettBTNjw1kgiuqCDlIG
2PNnQ3JwPvBABFc76WEsJEYggWRIk8C1TzV66mF5gBTNgOKpY8YBCvYx+oStvRtPk6r6zd0ScGY2
m9oYH5DdWifZjMQYWUexgly7TULLKTLdyeDWH+4dGMHwP6FL9bi/mDx8zrNz452TUIRrJH4HlrPq
eeleTMPg7qu2hT7gP4YAUZ5O2xYJ6YPxHAeADOu6Q/wDh2OBqbkni58Wi33KSws+2iESP6vXrIFg
gU4/rixI06nM/yWQy/pVifj15/wNPrxUyOwsu21qMhEVrpe9HgacxGmN1uL7lQKZkyXr+kJNDZLG
92VIR6ZgWMgOmkeO3Oi5f/YY0+B9HMInNl8iorw+VSQA1in3GTw/Gth09dDyVn6Hr9DyFtbRzZIC
fRG6nPBXrQVzxhwg1X/A0EYMONqvbArrWMUB7AYNJtg7YOs5K4lBH8ANXXmBVkwy7s0gJ3yZi9Kb
zGL2hnAGkBs3o/Fj428MFWs0sL4cP546D5A9ANbsJDLE74BznwWHAr3Kpfu7Z7DcPI7jLj8RJR35
yBi9tDA7r1VgJSf+LJ5kwy7TGx/+RI7JvTiZNIv0KGlXXoQjMf3y6j6M3h0Ch1PtM1+WeHhuh7U3
fKwTish85UwdABboB2qj4IY5m0gxzVdRcQHgIMOnw2+Ms+1C5NUYjw925s2hXwbPvepd7+oxs1t6
Y0+x/fRGcx3Yn64cEK6oMAkePGIa7xwymNLzm1WtOc8rZ1L9rnykrABdAiE1s/DxeIO6OpjcaGJv
0iHlGquTBx9Tehaatk/OLh+q9sl4hMtb34jzTMfHHZlX/M2Q3c2LW657ezq9mrNlRDUcvJmREKZN
g6IxNAJhlJB9/aYtL0xmMfXrpllqy7jwWYckuLg0yuNY1YxD9Q8P3adzu46A6esqtA0MNuwaoFA2
yV92D7IXZ+JizmLX6f03sm8J5BPoaw9TzKddVSdVSw4IXWsQZ3x/dzovgF47TyZ3bofyCSVef26D
yi4ju4krV1+A+KfnqZ5SNgw5OV2JF2OBGptYmhn3s3QBi+X5x1IGpENHWQk5mRdsGYNCdAHVWA5H
DH9J8higYPCbcgBNdxvv2+qZFvYEuRG6j0Ku01tJAn3vnhZ4G5ZUOJAPmJBjuKAKiwZzUN+AbIxg
ZkaZIz9pEjqL+etC+0JyyHlJn8RVwnumTE734T5VQ5Zr2HnO+K345MnrKF4t5mBfQKjlKhh81Rhr
oKgJ72dztfvtsxw1q026Z/dV4izOngqeegd1A3lZ8dc0mHVp/bB/mlfYp+t6FASV2RGkrg0sFDtM
VHUT7Qfx2EUdoNn0y5QwXrlRYh2LGncnSOPFHoGnnw6nrvWVPtkE5/DVox9ZqMEwHgGfkPEkrLmv
lPUbp/1LTeHv4mpUoC+Gb7EpKghSrdoIcoc/+J6l2kqrlkUP5+n6NK1aCOaypMfeX3hGlpy0HAkG
hAep/aGCP5S5K/AVtGtCnw2HfglT6HgwsznIHzOMlhlzwEbfBGJiTx6c0X01nUQf5LGVmElwv9bT
J9cmdOlPHzrgkGFZ4hYvOGB8WR3MXqbA6l3W5FzMymuEx6Nw4wTOkf7C+5kMeaoGCgcu5ngq1Sh/
yHmsiIknDaO0uOg4CbP+ttGYUZyILL8Cprb5YxagrfoHqF2Usb1664DxKKC6Sp9r6K8qWW36O/5V
tCKW6FyCATq4qtK4+amDReX0T19dN0I95i6dj/b1RcBRTw/WtEIktB46TDEeJMP3E925ajtnOAVg
PojENAmWMcPGLEBMhgDSspVeoP+K3hcU9FcV8LeuLFP2tvJdY/i7FvSgjRnoAzlt7sd6JJMJicoR
nsIq7l0Ptbq0p4qL2IK1XOLHYoc8raJicYXEwoo4KQqTgVNQfyW1Wn/Q/zHcR4AJws9TkyYwjelZ
TltG0UBkznWRi6z9Jk6YgecFyyVXm2k2+dFaxBFPMZAQ/+VMdGPF0+3QJgCoH1+7P9C4KKgWa8C+
/FcSOmpDyct2dq1rpDG27oixU3I/syM14SD2rb5GnW7FEPrbyp94bcHtDx9Jkeclau/D67BgGuBO
T42WQKcQxZf1vGqRK8KzMByN5WMBPYa7gx2c24Vlk5MIczxklS9zUg/B1wZ8YN34OSZEwbd3XlGd
Qrff/i2L88Bv+NXPs6xrZoO/NIoZQcpA56ZK1Q7K61ENSiIQTfiEqwYuFiz5RHKNibVlOn7alLGg
Q2TseHRiKfMGMqUWXopKTbTwAJwArXDFX7qb1gclTPuSdXvIXOucIC/8h1XYoN+H0k6kyNKeNys/
N1Rni5Eva3HQoYjaYaaWwmRewq9BpGxtQpiDcHXqJ9NhY/v0hB7iJe8WcfjFGrea1S5albIS/28n
Rln0FrWeIKrqayRSzfpWD2Cv8ghY8B342ANzfHRasEXYx3oSx++jN2ypZEc2IMejDWFEv+baObKK
edjTeejbKpKRYqAsWa6Q5ZL6QVNCRpwxHy6xcG0YAjCE3/r/dtYw8kX1uxvYEScCNCCU/GPInk62
3VPqTInbzvud+CYmIdaBnHFgt/eCh2AvVocRrJ209Z9gfmLFvrHolqNMSC3t8ZmC2N05dYvHf1Z6
A9v/zc70U6N78R3BX2JotKwwRmI+NHhihu8IwgY8i9eQoNNKy3VMm1alDOF3dmZ04Dw8mZisALqv
/sknOSHL20ZumFdgQpqIEUmHfqo6hZC1T+FS+5HPvqubwsLa1WcKDWzLDSNO8Em/efViUXvC3slY
f2ux1W20l7xmHGV1sWC771Q20GsgSs/OJRUnM4Ukk+BIZVAb+GXYpLwjhaBRwIQ+613X4RHLvy04
XbAv88sZtaqR2XJ+nl7kFCAWO861wZGt0Lp79qLLoHU1czTkxkbqBTY80JcSrxta1DtnDGEhhqA3
6eHniflHFTHDGg4rShvTv8DmT9vp/MTKBRlJ5XsuyX0CuJ36JWtY/8bsACFNx40iQYTyCgLef1If
LhAtyQ710aG8r2hwzDWUzTZQpbVR1hZiX8d7bWmIBXMc9e18bVkGUXn3zS/kLXHM3JyDlg8Sp/Dx
hM4Nb3gNorAA7z/OXAKmnaiF/JjIe/aDMysV5oaMoVdkdM1t9u79w2oYUt4akaWcERrWGVGIhGUG
dZTva3SZLzdG6+/KbGyeUnsf3v0cMs/eSxNq5LPJEeuSDIHFl4mwZx5EGlYAOEf0X2J5SrNXD/oA
xCEtP/RVfOivTW2mLq5KixDELnHbgr/roafdlUjbSju4l9Hiq3SRSrhDplXvF8bYdgV8W64H3lv7
76Ls/7d+ohQ6mUa9RV7mWML/tRpl0cHDvbELh3Xg2/pbXz97h9puOFS5438fUBVJ9BwnAq856NCD
OWH5kbM5EVaL4kRuX5/osCh/E7d6os6CK/i4Vu0oAYhEedPN3cSzE1dkUmNzEZGNHZGP4SPPo/YH
xPSlXMr451Wcnw7mTv7g6KpCXt4hEdWsvb3/We0SnJHcccsWHNpJR67IfvbmAEDzZf1UvLWIHZcW
HtOx+loYPUfdj7+6wjFbmozI0XhQM0gwsY8t72Xe+WqBuIY+Orp5VQ/qq/lBmxnVxCEMV+3/nFef
tCsSh3KAVXdX4k6FobwFGw1p1Tz64nfiyOZKVZ5EV3u1rDxNQla6PT0VTXHe4qm6jwtLl454215/
iNiBEsyWnD2PZtxM2TUSg+5XLdldUr0R5mzTIowcN0lpN7WyXJ84n9duGY8UbF/cIlFYgwZ55pws
7EFT/NHrTFGvdqfzizocxakUgUudnzMCZzJnu+OwGkyscQaA8to+JVv7Wymx2sYelmvjVdBpO3OZ
FuWmHYpA+gtcRbFcU7SmrmuU6z+4brCdrZpFS4//mi8i7jPp2vOQyLJoMKvinQ4PbVzewcdxIeRF
aGRbN6OPcpOkmSdIZJTQekkDtF8PTeXNl8e7L4itf6gzV/8PXCdqyi2HxyQeDK0uwDOjfWW7v2yD
pMLbMoWbnnYcjawwf3nKiWZsM/2EcSr/hHUXRcQr4xz9Lif85Ry3+B2mDIzZbTBdCuYTiGxgQBIx
yoFDIg7bom+hiU44nEf2LS5x7xYYpk4zoPP7WxZ71OHVOB7sZShzgEDPuzJXX4zRw3k/rcqyAS88
/fcWZklTXE/qIBkX2RH5/fVT7gL+G+fJl/0laQ20QZ2FaSse1qfSlsE+mxWI+NNQdPLpJfLw/642
OZIr6upfaJXUbY7P2tV9zMiRwelQnupVUCv9M1zaxPpt7wd6cc0Yh/obwHLfWQ/aCp5KT+OLZR4J
vNuS5dNX5rXwc+DBLBoM2dKT3tehph5Mq/GS0Rx6kU0x3j4lkXGcsDljNoLQyxk0DuODmPdvPW3J
YJAgDzYo9XANZ2vItFMDujjR9RQTb/k6+buEZt46ebTHmVloWiw5EWg4HKExNXHr09vmC99O/CkS
4R1VZA/Vw4c6Ix+dh4r/5GEF4fOl3nHJ2vuxmSSZjAIZAVXrxSktkVHyWEYD0sJQJAJPV5qG4A2x
nTRn5yb/HvoyA8vuB8hi2B6UCKUQDxWtZPiyFluuJ6r2UTRxAVYrEZdWmVxcEGtgoLervyfOb+Tk
7DTJZDS1cEFDRe8/Ze4ibk0MbTmRW7icSWp57q4XMpUH02QbF5/VPQSnjHuFgiZKJ8F+0FNVV5JQ
Vj/bFTzOqqEBEvmIE3UA+w7mliUnR0Q7hgjT2Dzqsj07B6ZQphDQwKwbI5HSaSHm5+ZJMQjAzBTO
5/Jn3OS2aoObhCVHYKn5gW7zmzwFKip5vOCIJpsrUOWMkAozqYn6Ste+LBtSyxvWp9v2w2hcJ4lE
Hjnfn2vJFTlKF70ua70VhQU7v4a+yqjwG3YZiLiVTFjfK37KFHc9h374Jfyc4ow6hDB8wTqaS8D6
Ari2GVCWf0HBrfEkyRl2LO+DdzTWcNFW/BUQWvRAlGTl4wNjOOHcwg7i+/fFabSMNQsrFKD4h7DY
Vi9v6jjij9nTC00fvVEqHDBYfiAOPg5F3mI3AHuW6cZIS4E0Zjh6bm8vImlydLfBlU/ypNZxlkVU
Qevs3vcEe5GSFfLvMAgoGn/T3h119m3i77AsImqTgMh1enBz7SqDsCO736/rmGmx2DlrW7Q/Cj0I
rV4EAxMljrq2m/ZWnJpp8me7HY2zSPNZ3vcabBSLNA8Xm5efq42qMWhPiEwQW4b2AybuYUoGs7yP
CWCx986CkIsgUD1v6fvJZioVxnpPnjUuAKKp2NDMGzzwhAW+SiCsu6Fn8XN8aKVRWC24p0Qjj/5s
YUZO5l8IlBGB5eV7qzPxdevpqRR/7sgJkXk/R+4fwbB4LO0dWbnU3wMPK9dFkRAaiwomSoB2TNnh
8uzPXYyL/s6YsoAshg9oW2rPaVwgvqxLkpTLMhAs4MSPtfKF7raLxYc+Tctdq8bptsYDrjKZp4Iv
di8dYWIzKyVVaI2Q/H0P5hsiMwU6vZhpXnx38K3wOn+PeAuetGM+VdRX0E+dugLHcxvO0hfV6wgf
adqcB2yR1gz5DR0/QYTVMRj/auYoXb0aC/OVpc8DcK7CK7TLnxo6sqSiMqLyDKQCGIbSKlMiSvOc
yGoMDSGPcrBr8vbONjy75pA+DQzhJQ/j227T9D8C6hs5s46yOHid2yn4aUJHKOEy/NtnRs8/xaKG
Nn6nDrJAMbgaD4NRnang412uwXoBBJPlNMp7mDBgVcYm1b95XfaWbn9OOFNOCBoGhBw1lnYbVPcy
fUWNB5kiZkjwbMvet1kHo7aU+DDwjpyiT3L6hYp+lTYVW48SMj/Io6j6Fyj/JQqRxkHgCyhQ+Dmh
k03hY3JA/QV+lCIVzi8AKu8Ve0Br8p0XeXF0kGY8kjyvhZ6nZpg2dt8Pj6L17SDXSRwQnSollNUz
DvICoReJC+cMVRuZGbr1/FjuHcFhhulTm7HdmOE/X9GvR/vjkDwld11cnR8O+Xz0ROmTd1iXTmCF
9BtjI6YU6rMomrnZ2tXj3uOjIwZqzPJKz+BJwYG436fDM6WpQOoblCZ15s6LWttGrHHmm3Cj/62G
uqKwNY0/IfH5NBXCst2w7E8DcGPREBszmXcEWlbbwgkyevP1ZCFCxeJgFAdky5Lprwwz/QaBJK+7
IpCuhp2cw5ylr3PE8U+LwTSuFv6tP5eKYS1+XKMmib9Tm1F6kQiPlu53hDxNXaFwAMAGmjDzYQH6
Ws3bD1rIeAe1Nu8YjmS9MyQNjdFxneIiVVjmx6ynjjFIFZcA2cLKmlo7tQdfNggb6YImDTgthPPy
X2X2P4+LllA5NsO8RWyRRzAlTbbSGqTYPH0kB6hSwer5hXLIN5HPcJjiIi1b6k+4ibWHIzvtx7NF
szFPOSPI/2gPdXw/nGl07JaDef2+DIEX6ARZGSimEphdNpD5bZ64NuC4DhWQpIBsSM0rQODPeV5z
fWWNhLrH7Kpg971bTYzHEbiGY9vFQn9cU9zdUAa2RRAMctHtUhxsTjHP9B0sAUgOg88QaYlKjOWV
0x/+60xxF2ectppyG1IwNtYZfmCL6OLL3rx6UGkIfs35OMPYx8N/BCm2cBJ/vI8iFvbEGQVZrps/
oN97nx8+/a9GhBOWUeGY34px6u8yKlmFwAozFZ7EIrkRVn9w/aa0Y+UMlQnUH7TbtjtjWBVloqVM
ZYfIilbssJ1LKAs1cMRfvtdS8fylEpKs8COChkaXcWesm0oFOLjW794OkQBRyNmCcl3m3Wcb7WNL
uOuMsIHQmarmDaMvDlLSKQD42mf/O/qSitWrftARCsgFmDYhRg1iIAVGHNkmGFojI7Gos330dYTL
7q6c/M/lriMpOpFWCgDHxXq/1CC2+0uacdhFYZeftWgcyZVjoZnk8ywCESy2/d6Ri/3FHthCu77k
7/oZ7M8Ge0femAQRlh1PjOX+rbQcxJEYvIaCznO716ME6Afhs5D2wEMa6ivTNdJzRWI2o8Yqq4LM
dn4oCY0ZnWTUIVDTTHqccgeGs1lO98+YtH/NWkmYTaD9LZKECkoNin7JUuD0Eyx+9HESq5a0Z3dF
XO2qzBEX+y69YGIaHaRVe/aP3tVPseu+Nt8vOM+WhiAV9ofBo1oKYATDw+2+g+nCiLVo4NaFLdpw
+Emf/heu6fkRTG1+FLP2OuUQgDcGuGlPn514lat9zEbQSYRfVSMZi5QnHGNTn73YKDKZfQ5dY13e
qNtM7HomQ/ih9xPtR/UtbeZ8EmsjVXY3olbb8an7bPxlQKC+8o60Jv6JxxjAj+oSn8dxCFb0SL03
eN3/rbRoM9U6btlk65W3RYx7WRbbRQNWh4gWt0E9XuVyoE03AP7Y2nxf1891WITrdWco3q0Olo7N
FzPYJAd8JRcVPXVK+qi8tpVCJVUQJ7J5m5OxCMx2po0v7zmyQ+nxeWia+1kFUffq+iZbm2GtSa3N
0welPTB1GkkChBnUi4pUita+jvwjMG6iv2Xm5viHu6A4v4xi8wZVoEOJJ9xkoh8bq+jpOZ2y1r+1
hgKnC6Yqf2VFiVA/WZGNaJOyitwHdTAz4J5TDTtv7R03SWj8FOMLiYsjF8DhQsVqOUoQdN9WAXyt
Lcqz+PnmqwWrOK1C5UqzyqULuhjLQjO5ZBW9SiDEpYmXdPrunDQK49yI9OrlC6X1Z07GyX+3rbfT
Fj9bYEwC3/OuPgh6TuF+8wDFWVhURXIhPjAxl97FknOT8P4Uet8O8u5Uzes/kBofr+jpCEWrLLiG
ZMHF8bzsRu3tvf7oEnypjIXKhzXtADZqNErXuB0cnFGJXGtA5BnD7CI+ctDnPkIgUWb/0s1vy3E9
dfcDXXy8MD4RedtumL8xEh/Iq7t8fxll0A+rjb03C52us9n9uqLyDjveBNkW8SWMp/W2Fh2girfE
4NKsIgv6jjFQb3U0L6kiXUy353JhfJAKIQwxZaomOSiOKia0zvSBROAHpHZh92nPPJbPCSSPHr26
1Ph9+UIcYtK7ei9S1nvoCEfwLAQW4eveG4LVApUMcVZvWzIoeFZQckw+/oFl5qYY7dDO2ZT3C0qn
nspSGoCpcoEmDIVKraY03uoqh8gOSvRBbdnkg/SQzjanIffLDfGQiAbXoW0sXeulpkSiVNV2RgPb
F2deipeiBVDrecCBac1XHZhDmPIlD2irxUCRTsqwB1u0Wm04jq92RE1gh4n122JoGEiU5rYwIxzk
K4jny5CfGgCRChIvThy66oRjhqdJlSmPM7Mp/1iZYm92HjBW4yBBlrDmef0R3brcMWCbK8skyxB0
KNa+Hmfnb8dFdT5o30+OBjeldHkY77JCEGJtvXEQrpd8eKvTf5Lwo5YP9YGxv5uCJ92iFL8NNCVU
iFA9ebPCcLXU1tBZCU6G2hq2opjVfppCqY9CCcpb39zgRbUI4EHfb6dN0naDXUBJzstF8vqOyGtr
bI9QugTQ+mGjenqbAFkVFNthBzhYB+2hTng2ncgdAGhH8eiKUgkuljjn1IMk9c4VYPueRJy0/rXy
m86Ko08EjIqW5UcUEac7jPdAzOoQFpVpeQoKwhdbZJYkz7L/Dsgm82VMzigj9C0Er9Ecn+AjueUw
nIKyNjAx6Raqw6j2idJLYvrTsAeQ/wTUv5nn2nQUIFQdcA9GEXDwcLrlFH0Qo2yVWOad+xQ5z2uz
V6dizPMSNHJMQw1cAzETLP9751uQRmlkHtqwzsWF3YALmEzbbO8BlsCicduUHShJmveH32qKumHu
MwGVhVqwRzwHyAs8Ra4d5BVgmzRQ5GJ53W1MnQOi/yG0iXZD7B2VxUKHcKgGMwXU4CCvXlOODngo
5srxEQY6lGuTqktxQUeNcTIy+VlQMxle+JY0NEP2m6mYElffLGIPZ15EIt+pa0QsMJYUkQYrX8Bn
EeaQRd6l4S/ZpeW+sKiffYCjiUtgoU69UWWOo+VljTbWeMJe7aQIQmhQYhhqCbHMMcjXEgaf/sfO
GmWsTst0ScB9UWZwjPYAcEfJxsk0ZYfRFib+CgWIS3dflLiJgXz4CwmSr8RbK6aut7Ic/Jl58U8G
+Jw4Mi9LWdLb8pEbm57tLR/azmnoTiTezfzcLWfRIbZusnSTnKpwpdX7JWfZFhNDjv1qstLNGdnD
GmBgj/yh/nGLQry6Gix/BbN1avD9TRKriYnaOifjuT7AZsqyldAfMlRtC74Rk5uoda1WYOftxwds
YmOJlTWx8yLsJSrmY4JlQvrUfq2egJtEvPOzWW+O2WSihImdDMjkxxEaESNoHg85UA6QwoB4tXRi
zN+vaJfviXNt8BbSBefOPM1I/cEJJ4o1mJhKi7jraeZy+lqR/LOd7LmdV5GZLhb5UMgaI7qqp5di
oHFzImwroSrwvV+CNQ+Km9jaFfMxKMED57FDmFNJMdmLuNdPGnED1RsaHbnrPvdNuR0Hckls8zsx
dNZNOUm8qDtBEEYB8A5zUgja16B16m6CaPtMvTRLtFloTNu9g+d3aF28rbAIpt5NH62p6wXxaFvx
vuormfSsd365Aft6sFYs4HubVpxremXKJxBjW1bcZ+KUVUyvMGxKQNgwP9mx4tJXpmQJyfK1gKd8
1PGE4SZ2OEUXj7KBpLuTPp9MG71dBWc/SSkmx/3rsRWv4PP1e/BnPm9pDOK3D8+phVVZ7+TyTwnf
E44wGK6IoSHXx2QIN/TC9G+VDvWcdC2/jIAzV6VZvsoO9IO9Eu24hMG2LtkKi6u5HMEFg5+DNxzM
9or0adU7UWtBOsL3Zf+3cUKAGr5Lwlt1HFxmxWqfhSBkGwS5YqrG5O+NSvfK7JSdG8I4PSVZm1sK
8RSDCgU+7WMQxsdzIbHSIcm7zvVOxkolh46FT9T0sAMFieZo0TuBGwjCZQP0TzL/YrHTcAliA/+V
Wcba11IkMEHesUlYjFqOwp47Tg5Lb5ATWzxo4zS6Hr7VPQ8vYRMLaiawu9NwXekqSHQbQqY7YxI2
kkTQg1LUYISpi5szJYHesOv2cJQyGaC8Ii1sHHshqmEXEwGP7rJDng+e9z8B0i2cFK1lkb9II7+t
0RJad+Cu/VcTpFlKh1mDMP04MuBeVEc6Aj5kz8DtuoOCWKGmi2oq4UK5NKGqrejzLJ5aCfBltu1x
Fkm09ivBzTD7tbjkN52FR232qK8bESfHakAJdUpSf7Wf9MdjhWXHhkl4zMpI2opb+6ooxqxZCNQf
uMWyZjztLZa0upD1nW1iEWvK1kFX0G+UwGA9VEfpjDL+bOhw2tG0sNFfQArRQiUFs1jCbg2dBkYL
EbuY5INafPFAWg1Pj3vQYWvUYbwMJ2hIKwSg7N9Z46tEejNsHKVcHclW7WtuRFvOWWyt74RKKc7i
ruQGR34uqOhUMWS1oAndjWg9wiehjgmFyvwNI4491DqGUv70MMPL42M4R2Jx7vEh2fIrJEuZZiV5
AzZbaqXf42DJFf9D4/wJEGmt2YQ/LXvqjNm8exemnuHNuPPEX6a0VZ9s2dvrwy56QOix8ZbPwraG
+kxxlBz0a3LokmiohiCH+JQ2ingDIDrz8WDdEzw7dYtlIJfmkR6ebcLlkJfeDv6VDWWYLApdlf9B
F1zyIbm/aVjahKsIrCjkgovFnBdZalyqJtznKO5iKcBymi1K+VhAFcWekbuZORGb8J6kjCJYEPZN
VynWoQ/Y20xK/WNSLGgBl/RQlN3U2x2HDSe31PHwyCajHlnQjw6Nf4mUMOv7v3zZMPHB7qAWkKEp
DhhRWcB+TEchu+CxNii5QRpEyeslxDWCPXMVdbm0ZY0BNIUqec+6ctdtuhG0VdjylWHTVvwMR1vB
bU8RgRS10uTe8dGj080tMY374hPDhvEbHPLyWBF7ZjKU/uG53KrNDJpwjG9kAWTnDZdjaXyGDiWX
iUO6jdGJeIbs8dySi07VKz9SkVeE/VKuiaA90NtV4CQhW3ME7cVrhPHDR2ekzH7i46H2B03MkkBG
jX0xp1m0+doc6F4KWKC87dGVMWb4okm+mBcauQB9cneYWlL/3diSL0GXG7fpAQdXJnXfA84T1hvF
r9AE0ZHF5XKBagjEbiOniS6oo+96NNigY174whMNGQJqqetwMw8fIyMiV9IvBv+hjFHlBDRA/Rc7
RWtG45Rmut1aezdZlka+tjqn4EECdn8i3NGVPGRSl59AaFPhedJ+9yUF/NtrI4xDcO5nVFzys0+i
NBzVXoNIzdlzqgR22ukjQgY7/KU0A3ubUekWAZFCr1miIWHD6JaY58KlffwFdN7k6xKipDJq3nSj
1tLdMawXigtp+JALfunfEbaiyuSFx3XX6cP1AOHRgTJtEacP4uQ/xVy3IJN4cP14qNIVLRPwcax/
hp+gLnrQE7IJx9ykpjut6Iu8dCcu8j8lKq1kiuWaPZlrl3Ov5FdDMgM0v65PUrc5Z+cMaZ9sIFfV
tcP5fr9Mcr/yydDHxMbn+AjILpvKyceFjaiKT1EYyUL6em0hlHZK97l+7hVZpuV6tRmDrCz5OHtt
nzREu2atrc2aOX9hFIutzvEE7ZS2J3S+21WtZaiRm2Fy2MwZSrXJvMv89F5Zmve5jMIWIvgEPRHQ
D03GYzCylZPydt9k7F1p26hsswuSCAWBS8/K0uDSIffPbUVlOk68QSrLfCuheHGTulmXS4Mzhnrx
fNu73P8AbEt7NbEFqzWKLZX9+/MtpkxssmlRDFbEYPdXD45m3/eS7PLFIWD5yhaavD5tcL9luony
gWxPUhlADJhqPcoA6k2b+AOWFeT8GTlCCtIgDbV6g4YnKTRrHESFvYW+7pj7j1G7z4xnOREoDc2k
8nX5LBXB8lfTofawZRqYu3eam6O6AjglOQ46CsEaaI0ikXNlVnuMmp1csDrNJZoJiski2DNtfI1d
g+oQFGiiCTk/bf2a/PbLo7tXmRirZ72EFI+bfuKOXkKqiKjb8/F0by2mz1mHFrcEQdbZa+dsLP/h
4za2XDtjVNgnPrX5RcbOkJQFKUNK/tefyWFjDkxUMonQQNVsxkn2zXm2HONRW1FAU477uJXKTlLi
hyMzAygKtO07btXaEhpmYxBFYNPnzHC7n9s45t55wnRBm34byjsU+A3krzH5SzLJYxdHgmFzcvGO
p/rwejxoiq1YV4QdvwQ4tU9DuDFDgfcuUHtBzGFzROcXrMC2CsTzLBM069KSn8K1ixveX8BpVW5q
wv6Gss46oC9g7CdLj7z8nuFxukuou8oMz4Z0p7qe7gTk4PHeASKm8Lha9rATcCJLyh3uvc+lND2I
M16E0aqwvftzyTW1o9SqW+4+MQnR3/tZZA9l18cQKXGnLfRRW/3kbTDqWJBL0fXPmpZKeEZzR5Me
HxylnFPRnEZ+dwQRxrmXntMzJCmhufZLNKLBLvPO+SNc2qVB0cdkkyL+XPtNkTvfC+5OYPNuwbR5
2+HhzQqzSNEJfhTjOo0yoccoT50xk1uEtPwaxYcMD33Cqb4cmAb7NiqRrVv2I6TvJj2ckI0qmNQx
i9aJ8YMG9FTFlESqDpFrBnBeiM5PSikZykwKpOWlW9kVkP+JyUEE7hMr/x0Z2A0aPLT+DTEhAOJS
+zYe4vS/GSBVPZkXu/J+YxpgKPyKYlo4spemFpP74HlKnOps0b3hiITuosOuDrLh1XQChFZXMVDu
h/RrsJesAdBoZFJ/bOEffzNeUOK40+fc3HYyEzQm56HzgsuU/6YL+OVuJO1VDeRTJf65bAWXHttp
VnM2oEwCSuhgst9jcUGtTgMuxbqIlVM3VfnsmLEky/ORBqZgDs421cvBgLLWyktbkQS8QhU9uLwW
tSyGPBDQJJ7cNt5TdyljUtBvhDXavxsdBsXb2bNfwxtFX4/Wps/5V7lI8BxrYEAMF/5zVCMlOcGa
QnztvtXMg7/UZJqa37YvNHV0dGsk9l0XclguNHlovZj3mO9kKv75VabP8c9aVx05/TagepSByLKv
iHWXr4C9DkXscKPBA6l8wjJRJZBF3uekUhE4iCPDExtVH7HMBOwwHe2j2BWZSy0uIDqW0KpHgnjp
YNCztOvFfxaWGnZOrcL1OOiVhmB4UrKE7psVP0dfeuZPM2fNIMrtOn0sFt9A7ea+kdQPvI4AgrB3
TvmNGbT07yzIPdwkKp2rnFRVDSMjQGf4OzD4iW5Ce8ix78agIWIz/RrS5QKpVre2oOJ2C6ou5Tig
vuVTcbegNkpDrZo4AEqWBK2GQkXC4jJs4jbGgp6n1jxvyzAjMUgKmiEEdFoz1doTuqeVfw6P7vlL
bnsCI6zAFKelUo0RSlntky6OsX3bsWx/9yG0kM7fA6tn/5s4JhOq98ykd40zDyK+mcFGXgromgyL
IHR1WsLuqNLEmivtDvGPxBUWLGD8InXYUgEDMgEAyP5k2GJhgIX+3tFVdvp996H0GXbWVM2sUW0e
cMZfnbnOYezJdscZb/Msn1LxsodAxE2cHwxRoH9DLI/DdUd3bBI+Qz6IcqgUFcWTcuQLQoR8X4eX
GDMZjefARtIucjZdChEtISUD+lY/zzfypQojDyarTfCWouTRMq7H+wg3D/OKnarMao/GT23FozyM
SyGtHkNcGjbaUYbloRo6/d44k60aEA5uuguzbwV7LH2TvKSVymQ3TwBWsr9Wk+Nce819GPCLp0LJ
sa48tH1KUogQ7AsKX9u+prKd4idz+R/Ne/00Sm6oHgwVMlemqgENFSjq7Yy1z0T5avrgy9eTqoJ7
ftCMyE2xmYjvqdjTy/MBukZSHTemjyVYFEsM4aYBXwvH91dG3YxdT4MyAjAELgod5wL9tfFM5yLI
WbnFBt1P4NUgVu7c4mQ5J+ukln2E63L+hG6GIJi2Q2FjJQ2g0rbfgwrmPuD9ab742omiVqOY/oEW
Wb239I6fFSutFt5C9bPbsSo8rkSf3opDVq/oUpOg+eNgPg2s76al+c0ceyFhgppn8HMgh29Z2Odf
6htzIWUUitAtAt8vGp1cnIiKH2fVZsuwTSUonpYNYMNHxtq2DzSh1t+yCr5a1bKJL9vItO7rnr6t
MIae+XqDDnoPdWYS1oLXvSwUEmgZGt6NgJyQxI8yqyNV0k0tkL5nkJP/7maq7HiJ3s9v+grnqXfD
BKAuZGN9TgXNaoSunuJiugDUVSJfO9PUDRD4b8/VTxEmNPtmDLJ3ZrT9XLzp4x4WIyml5iqHysV/
18ibnDchFWSwS0OvryMecADyq2b8B1kJ1HryWkkIzOBgDi+PKLfLlnNbc+MwqyOirJnU9CwKuZYo
TJ5ugexWQ1KNdZaYOa3TjtK2708p6Ma2lP6ZXlRQKlWdqSm4AstpJ/bsgxXPMj2DUjOqiayRbQLs
fkGUKS5eAJIF7W9V9gdTh28fNf22UmgKZv+RQOVG2d6faPTZ/bByaBo/kp/nz/tTPb80VjqlSVgQ
FOiKftvYpYOrWI/nD+zWjsp8fLqJNNYyDXuUG5RmYJHBvUzg9t2ZG4Mgu9PUOPjB2b4xct5mBSkc
Eqhb+xTNYe28vEw1GMrLF8K1Z9iv0A0J+pzFdFJAVW9lNS95N7cgPzMRL2llnFHu1unUdhkRurbe
u5NMyfiTuEORnM05X/IY+E0tcQ1oiqezCjqm8xlm+vmP+F4APZg1ULyQHXz22tdq0JlXL7BI3U8C
KALRQQWpx+Cy6AZJM9MiAt4cyZzYebfryQru13L0EuKON3Shp7ue8mUX0gcOQAiGPLgSgOG2pDVY
X5neJ+C72En7mS42RHzF81vz/lbOw9iRDTV7+Wgj06EK7mWRs4FlGGwmmQ4hSMDlaNFK0M68yXIh
qVevEqtQDtFa5iNK5hotGALCj327Wy3Mtr5F9r7JznxEML9JPO1DUmmF/XM0AVkK4gYllHcgFUPx
ouUHegfETBJ01lLjt+kxtCNNhPul/xDQPNSuZ5FzfzFdMKmurxCiCSt5GQps+b7JoVjljepYiMZy
zjoDu4xFqwahLkCjuPNU0Z8kk9cTRNAgk9XurkXMvWx+jN+UmuzNl6XJKjPlr3pGLX3tKfMmd+42
XjyhWsQOzTYBktdKFB6lB+KcRO9bWhGH+8rq1dvNPuFmGeOy2j50ngzx8nCJlQAViA1RWdjzpuOo
olVgk0+OqjsAw1wPGGdN6bC3H5+fU38xr7PSIN31xEXA+Wc8J0hLyaLCO5BelplI/K7X9HNfCZiM
tzxiVgM37H02lDxWkXCCri0mwNLY0j7Nbz8f0hTjN2ZTNoZUkOpOKWXworUGF4JsrRcEOwCyH8ga
GyREQc0t32kg+X06Ichh9rjuiFMxRIpJaEXTG56KsO23RZ5X4O2m6ie8vBoWeiHCzZvdp9LwPiRK
GL+BLwNMY0XY38Eej08fKV+nfVjbEHNj/hWQnMeFMw/FQ9V4437PR1YLixcIDlcjG19DT6O91Lja
hHTa3EWgfhyyXOyT1BTlpp02dom7GvdHBC1nkUoGCtHdR1oBj+C1DXDWEc4CHyRXDoNNXzYr/S2X
1/5jvDltOhNuN0HJIdFzdirWn/SPqwKYA1yFvXkyGdp91FnZLjvZhps8l2h1i4Q9zkQTjrKxiBUK
UHIfYnJhXzvJQh5vju16qxVT0e7WICcKheYyBX4kWf9T2qjBUtH1tFgreiuS8ZglaCBTWHk6q47b
/n0SKicQ+aXji56MejIGSDOjXpx1LRv160a9lOIoY+ZG2qQhHCmfiXcbcgzLRhzprR4wF0gdrP8p
WxOQiHXjGBLKbrmHVT0g9s515zs/sTvo9mEhMq6Hdqegxb/mkNfAAAHcfYialxCElEUB7fk9/QG9
QYMNd59xU20nWpbgn+JPase01hrLDdR55IWWO6S89NW1yMi4tep6YXJBYVsc566qn8fp7flum7/+
a22IKJ4GPfmnPtbujrT5FbOxugkMOhtM3ptqG8GOMzV2ttckd0RaUAMlGM/1J5xbRZ3Z+KfaAjIp
rWn7R3MyQ/R9emxijo5OFu++IxVPsRIeJ51odBAjDvZAiQ7z46dxvWcDXHv6Qx7HFNVGrBKtNry2
D5fp6byOToQmd2763uCJxiEcJzXTy7MVWwDPDUzDxfeOh3oXWjbwHuzpWITvZ2iUqrqTT/Qsgy2M
20YM5Hh5U0UGInK43Ot4renksJV/WxY46R994tLgeWWm6T8Wk7tpEEGEssAiqDpjyWKK/8egc5Xw
PszFoteMQAd1an0Rg4gD7AVi8ullXIUhgKiS0TOsWhByRg3cNWYTEakIj0aWJeiaEwsbVfhX1XXH
s4Wzuq1n3MOOh0UNFeA6CkpmdHbmhGmtN1usECteglMT9/QxRd2el9uR6cc+mvT6icCO9lleybM6
hyU3iyyZU2ruCOcK2gnAHU3cxqm1AOZGivrr6K+ztSY9tmdMu+SlX1Tg2v+8+rRpWbAC0pq1qYfG
fDjDYo4FAMeJcsJt/+9E5471YP3jEgZKM56yOFjSokyXBjwEDHFAdJizIrxdip0toEQBPAKqQDP2
VNtVFDHWCCbJN8BMJrwlSMJkV6+VSlBQg5ThD8a2AETj7ZpYOtx4ZJjP+z0Vs9ZaIqsbmI0d+hFh
Cj9shGacHaHiDHcJGkgb9lm4cF1zclRlMelnG7Zi7f5vpIVNce7OdCD14HkKPFtsQKNkxHBQF3Gs
T5Q7IkAw7skQzcvn1lsnqQMR67bhcyxyiObDMauXWDIgpu1+gObCbl6nZzfrPznxPIWmUftXdPaj
5jZO7kHL7Y+QzGAQbapVwvUxXjGeHXPNS2uRJCL/T4/zNGnQHtG+TAmF+wMgc5cX1gaOFRP32sAS
kUPjdkiqRxKphOa7x/jRtyjyXFYSERXco+QEO+wtFnzvX8EWehXhP/9N5TnirpkQpx6BP0wq2wva
ZXHARKxFVAysoyT3hv1ZDxcNJheQlISW4WbUyV+ZQl84jojUmoKdolYNvusOCv+DBMxaT8l26G/2
V+IqsBJRdfQe0p06NcaT6n3JlhgjHzZcCCp8QnL8zogFWfTiXUkO7CAbJgKZmdbfpwSecB0aWKGJ
A2Qq7tJRiNPj2OfTOHAwqioQRdLyGr4qmW5VxUEdwCKsE+RooDJxYgfZ7Vrno1KU91N+ioVGPXEc
1skqEW2b+9PgYe+JY3V6caVzkrNgLY0gB/paOiLD1Kdm7v1UfFIXdwdIgNXf0vgDeVMt6epQj6NZ
xLZKtwbp2vpCv5nLmc78zxJvZ8A4+LHXoiTb8iSgqzIzjE6mrtqgGOP1+8LQLZyxtM7nmIjHSVeF
DzP3XWRO0KaGQCvVGZquWExCrGtHn3CQpTkJFFz0DqUsnHIcwdKplm/FRJ5icFQ9GsZyoATLFNMi
RSBwReZLHYjH6N0HpdY160R2KmGE4ewautSEkOYEIVIdoruMs01d0cyb+xTuInBBowdk3bbnxx5r
2XPjrL9b4rU0hKkFhsOhYOB/Sv20kkjXTFdJGB3LCcaMjwiqi3ERjCzF0hV79dQYgyImjX3N+Iex
OY7YctT+ZZPhLx8/m6VH+Awv0jNFKZ36ulIvkTS3P+K82327mj7Ay2CCfDr7AsVVgTx4ypMrXrHW
vbWCk7CUb2jS84ZNgRR/cDF7Uexv9NmKqh3i977WfiREB+0BGzGDDRuK2iPRWsR/S5BWpne7bwNm
C7Kp92VyDlmYmjEvhD55BjtlTjx/Qu/rF3935MqgaoUJBT6lvw4X3XUiUkKzLhgiznBX+5LrSpH9
iTgw8JgMD0j0UBe/XT67AqQ5OR716FQwpo8fGYKU3gP93P6kyOZh+QkZh2oGQskWUSfHl/adkcXU
AyC59Kyc0hNzYMl4a9udDx1I4lCiKvQ8OnpYUZBuLVPTqYWD1wUCpFLIJm25wY10Ndd3KWmoqsp+
a1+vC/bp3SobwYBgbsRXbyomud4160tX8i8L6bGzLCyryK77MeoefQQNoRgYsNA5hbp9YBVkI3sH
SA9IAx+LNiw9QETW9D7454khkN1eH47DPGbf4MH4DMsh0gMApNPNAhttuiyESGAEMozxD1IEr7IZ
2surf+YeEXixScqCcD1FftOrtr2e0I3JUab1QcG8JQ5lgTLDkFtQFr3TtZLXEhwcbX7PcgSksfsR
Hu2Jh1BhtVzPz7etQM0SJyQi9/qB+EZG0YDNI9CUsXcocjX0gUloZfRENmQ59ljYsGnhdslK8YjE
U8H8UkbMTTZu0/XZCPmZlDOHHXDpADMAyK3ZGpJ5JHb4Ncf1gC2cG/WtB6wEOAv/1sKmVnudxIrL
QsBc7e7+/74csesEjUReOKHtLYGQGRzRZd84hB9cB4VLy/Gt5CBxLUd6wf4z4b4UGE7Toao3+sb0
lpHwG8wNxj7oNdlnYuTeOP71IBVrQ/FJUH58bZNzQeijCK6AgkHRcdEwZY7p2OfCrclx9Zn7ynDO
ii2oA6d5XkFWRzTE4rUHGbADHwDtRUVU1dtDnZ2YE+yF3lW5LR7bD46n34A9pkPR98+at6uSKNCB
jPdA9nPGiFVetTpXO25YDuAe/2/Gg5rJ4FUTPCQy/gV+0SnI3GSB2Rag8syYwHF4nXFE53U3ctFV
+S8Awamzfja1RilnSW8FlAP0MuKRgnHzOVOY5CGl2gCU3SerPq06vHRVmfp8Y8nyGxrBBqUyuc5D
Aypb+TEhrwMc7t729n1r9xayvesmeMk1wX7AmPvTMCoEuwbazJWXCXk/Tw9cFrDkALazhAnlYN85
xCwY6ZsELxeepcWtzcgUfvxlIXJqPGjA+sS33pOqs8GFTuztq15HI8PzMJmOFReuRLTwRZDJXbO+
go89D8L/wPeZDNCp217AxKyju6Uk5yqytqXAhtjc2iyWKUHG5xq8GHOH/W7ERgTrBNQ4bzCW0UY5
tz8EF6lwkYOQlKdZ5GSo6GGfWA4OFeaMfcZO7CdXd/I8unpjeU4ZNZGapDYkzl6uCU2EjC+up0gT
QLRNwBfIHz+uakDBGmzd01x/66wwdr80w0eeIrkiB/vGcvg4HpRcaK9x2EoCzpn9hqidX6gBG7OU
C2MDEHmxV0wHHFFKUKb8QqPxkbBi48o36sEZ23QUgHAP/JSmt6rLoKbFBcfQkUTjx0e6lYR5CNGg
GvZsCdOh9VIeGViPDDUQCi6wNzgmCVlY6iqdSFRvwCAxAYfS+ZOlNKDD1p+Y7umE2ImaGL+R9Dps
mGhqfn/rmm1DV5F+suNaJVKnIDNjMxob7PDAtnJavmj5wM7z4EMP8SFMdJKWLDbB2NMV9Wl4KzG/
PmH+SsBx53mcho35y/OjX9Y4J/xcJL0r4cpLATdNEX//dRwTjvVwxI4au1Vm/gMWNpTNjtPt7ski
Nh3PYGLe/4oKGP1a2ZBVUHRM3hqEzBom1+YeBb0znS4mNEQLCOgkLryBkmcIVEqu+mIKWCHD00J8
sTIsf9EUAWuTt61u6K6ypac82/IV/z3ID5ht6WCEBsumjoxnXdgLx1apemY8ZWkF0VmLQvFmS/tJ
YC5Q99mVTVyq9lR6YIPlKRjiImB2BW2S26+vklMpAZQ3WS35S5L+JjrvuIcEBtZ1+nDRS9RUmRWD
p42aL2ALWD8ZrIqpkZOwD+N58M4HtVwUxmpNoxVyoEkBekqhK2T6Rw4336ITyuNJcCisQQv+1g/F
qFr5EVwg3d1Pp/NsIEwpzhoA+0emaja2GUoUYDKpCqrgSpgQ9jAGXfPQTrqxfr2f/Uhx2dps8W+h
a9qeUfNAvHWtVlkUpmZQgCriQjUPp5FkFjKLyTJhdiCmWklP3Ok7p4Gj5LRR/oCaX2eGXM3VRtT9
noN7odVh/w2JBX51Myi559vEw+h0rgikFvvg04zX7LV3T09nflzd834A5e1pzuPZj59DCmd3cE11
ADl7cdi1/f036PMAGAkiphvxiTvNmy+6zL8al7Brbau95/Q6h6x7iJiQ3SAysNvieSaWjDuZgJrR
mgwOZVjZpPLhhOOuNCZjogYkA1AGQwzG7YymENgYrGLcTbO++V7oEsb/yoghWcxaQ9WOqgulFvNa
EdUO0C+bg+ncv6eOTC8SI1Cok2dKGEu07wo7dPnVGjOkba3kwy7+54c+3x8kYbwUwUg/r9XKLF3w
rRdiS6vBsn6SjkSCa8togmT7mKfuu7P61duSrgT9hvmtfFoVggY60TICkz2zhf2z7lMO9ssJHzBp
J26yqFU6Hb3cYWy621d09PUYVEQvB3Et+JUxT9jAZw2Q+6RbJ5CL3ip2pSXfF1qjIq5DCdWjHk/P
oQvFdrpIolILCdetKHNsYaSAkHW2Bqzgc41tZ9gatAcfnzSNgU2BlSPUTnEAIGZkNnQyrOVDL5wx
H6pQ5qW6v8N9eauZGIoU0DwP4R7eUOxAmIGk+/xNFx0GwRfe6At8ffwC4Fa9StYCYioku0n0uEN6
BJ2mBDwEoqs/wsBh2Ve1XrwGR/a3XgcTwI2xBgTXIn5OdG/d5GV8iZl0pelX7Kl0c2BoOuL1OOfC
DKxEYnWcKUfoUQs9CfYHwLaPY0yqqf1kzoWq+ZR0T1mNjPP21Wy7cbz8cD6WusBSUIDK7gy+pU1d
8qL1NPgpiJdOnr3OUw25IdgbpiDUfNFi4gaRfKHG3vA440WZGO9kK6ecliNNwKKZxTAJnKmeSqYP
wYGf6RTvXFkjeLEok86dWdY12ghcNp6LbS1DkIAtVcQBqSSy7V04Y5USWIQfIRgxlQpTf995GYna
8wzXMr6Nt2T5ULwmClEGkl3+l1jAInEFmTAncXrOlwsw4eocJsTn4j11gjIAEIbIlT4aGXYLU2Uc
BVpJ1uFtBmktXeJY82DpsbUauetZi4W4tmEi8l8j7kk3/bfEmvMzJ5yFjegspddcMU73vESXODOP
HU1l8AIj3Y4AP8EPlY92Hg/arPCDifqSOWUg83RwpLEm+nFnPaZEh0p+WP+fnwBvLXTAaqkoGx6s
eHH87Y6sPp1nKjroe2FKVy+e/3s6q7Q9vQ9qNaIPGZu9ezWhUmyp3ruyr74cptseUxEWxtmZ/3ZX
HXqADE114sTjdJ35ETteWKVekvyb2jnCnZVAYSHxDbM6EyfuSN7K5DRUJ9L3QP2ZgwNi2qY2j0oP
Y5or1I5NL8vHejvJUYZX7TDpJcE+20njYWhIqzmvLDA03JtyqV9BZCB2dml8L//HmhL5Rh2TWple
VzGx3Y4EZmDKtwxL/6TnkeDS17fCn8Oc/f/BXDem/q7xLwd9OiN2MRCyKMG5Lx8/CR/2g7Eiwo5o
P54pdCFN27aURc87lsf2DeLNrt4kBhfj2BeeYp5f8eMq7z/esuYFYFZha+8Al7rIWnbryr+05mOY
1McGdC0OOP03G/qitcnpcx6wxpQqvt1yVl9eintNpe6UUwGQpXMWcVAFvzlss6Zd93/EwNeo8jla
btZJrlxx9YHjCBNls403oKUGUP1/mdO/i3BdZJdpLp47dyLWqT08SQF5sqnfdBcik+VwtfgbGjhg
KICgPxw1F1twb/ZjlBd5kEXK62c0edFAkAHoFMB3nlKVrcPzQ8iaLEvaWeD7qacqG6FuFIYxv4IX
HSNLNwp6GPo0nmmxo71/tHCx8qCaTmqqSupDPlAskh7X6d9z3uZGKtQMdizJ+0cgK/U2KuBmjQK+
J8fJgaHpQqlBx2hrEWp1A7FgI9Ct9/unevo2GIrByfwSxOEkSlZiipgwjakFMIx1WgZxo3Tqn1Jg
YD5Z8vY4nzRBhT8yAqNe9fkQwzVB4RXhrW2dr1lxY4JmyjPWFl3tiC+oszMVs9njC1Hlyx9bSEcl
iXCsCkfH4I89+JOxqi5OihmDLbA7kEYOeD4IFrfvvIHRSWF56NAt6o8+PPTKi3AK2fEozCs9z/JB
742jqE3cgk8EM2fQFPNCdYXygswVDBF56OEp6QVFFQWQIi/L4JhGRrB94ljczgcQdpTqsgB3DZOW
qMNqRy8667iHvo31VWegR1n9VEpBqnftLNlQAOagJGpx0lk7kFdt1vEi8iQy5Ubt9pkmL0GCtY3E
mzdmolduOhnLHy3xLrQnEjImAHm12gALQzNqsZwC+8I/V//qzUGEQe4CDF0qA28mfivqrYAU8h3M
HhM2I4EvAJmrSQTuHe0GzypKSznHDkXJ9cF3/toH8lTx6NQgfxQG7awj10/ZBqZ/LNVjgvNpy0bc
Wx5c31mP98gsuwotPbpRyZLSXGeKlJsH3WGNGJluI39ZhpXWC5CTAzx43A4pZi6VLoVbKXrKqWEh
8VCiUN3erDojDFh7slOH3CMt3aACSkNjPQCTURw2PIIV/mxPbbMpgsz2aDs5uMopqiIQom5MAgoL
Fxxo2AlGvJYEwocZz/KjBn3PV2F6NOh8iK79K7H/phcoy5iLsTNTgAYfs1pFqziyrnXQx2ID7prC
Y4JaOghk2HkBY6X8Pb0Whj7rKyBf6cz61ewivM2/UfRG3xHmGgbmeZ7PrfnRc6GSvyeoQRRXwZU+
hbCdGoL5lTNtCGE2pDwWVfj4uus2RCXF7DJTJiYgBSz2pMDK2HlZsECjQNsxhV7JSAtICoOmuRcT
9ycco/BBpLPEvXRlQTiSyzd7d/pIIR3kl1f2kMtkqRvEkX0x9r0A1HAlY3GnLoAxQRLIfG/8+sjK
8Qk//n+Y2JkDflBx7BlFq1Gku/mzc4npEpvkFTGm0XJ7tid7AwFqubi7NjcV458fTg3OSXgx7ycn
+l3xNztSF9rEdaqqj1c8PDxcrB9wtOVK88OwD0YQfPoPnbLVjXegi5DxfpqwVgxhbrgeYH0Bqxt7
/Iq3ZrEUXnOz379dQS41pBOBVlv3x9iDwnJ1KYgLRoQf7kDpAtKz4UEJdxCPUt81GgNeT7cMPUS9
Z3Dz6LgESDM7hBqxaq9/438DI5VPB9CqroH051RaTGoH+f9chW6rNlNECe7DG3CXfJBYvca7uOUo
zBdJnLdVXI4UrXqMdVgzAfs6SOdZfMX/o/X5BNw3g59d3yrdtqhahzIxkVLofJZoxfrUds4U1/YS
DRHPr9epOR4+pI8b3sc1BJGKcU6h/gf9ZR7Q+4EVt0HVZpyQiNtazmxmlcp2JVZgq4YZnkOTYCV/
nNBgiSoDngKvWjLiBjikLt0cjZv08AXER+sodlvBsgf+VxyariqpZTNPUnIW1S/Xb3zVzGdFdPzP
6bUQ9WVeVH8eIle1gdLORY1kTVFiIWBsUU1H3aHaszP7dCCU9Y4IJ4I4ZDFhZ/G93l3bgi05022a
HeU0HJfkK7nfKvvmZ74Z3RYYnYb0Gmfue6gkZf4CYDh3UDNUoX7bI03lCNvaJPBJ6yslphymhxho
u11OmgCZS3UTtp1mGUBgijz82G58MPumwfk7i1Ehlfnq5ISZQTUfE0+AuW6A920kNY/8GwRzZqd7
ZxQStDWnADgS3hiBCaa8UNwLmdOYIbkgpcIhEcJpAwdey2ltFxYIiT++5l6azCegnuknYwF5TJMI
jZNL7ToOHvTdCAiB09JP58ruQXBFff1vTUxKB7Z15Xkjom9HGM3sDRF8ie3cH8IZ4K3zaH/rNYz/
6pFOG3pTcqlVVo40yTdrXgh3bkNKFMw2hwXdpm9Sh9r4lBnpRzg4ulLTmEwkS8wEHFlrLCEMP5se
j2Cv9/cmNcSe9sqmOtslCwzSBV9s0WlY5cui7omxGTPlKQmaGsJuG5SngApWGpXzyHRN2vzUsU2b
TyWS2WHlB5APp9GIS8H2jukbXqS7xb3/7BYPu0tQ/Q4bWRp6HxLgnaFZedcauPeiFucSM48SndMB
qd8VvXZkptzLuyPuHc8zaj6GuvbGy2okm6MTy7J7CPZcpCCkW1h4Xeh9pPgM8sphN9sj5q7UDcIv
7PH99+JixLUZtidPfs0rZIfvBvKHq4eyLvhI9HLQRfkur1Xejvr1tfhuCHUUOY8GZjYqHUw8lpFo
J+W/5PKo3Vc2J/ev3krwyaiPYyI7Yu+JiNUWzzNvj7qTOFwNJWI8g6mgDz0AXkZlDyfe3WPa49cY
QyJoPR0jkpmDpvTe24J/mIolEQKjSOYoqXEOVQEQPA1L9BJrHhJqvtrC7dMWRTcBzLqrbcye45m4
KoA8xU9/cfcEzKZFeur2FlCZwhUS1MrMubFIqq7a114jpC1Q+e+gnYmNGm1lhkrXHCLNKJpuxYIg
qNS6zISgKwbztb48/sinZkyE0TbkPfqSPfT55j4tDrv7X93rXMbT/niVchsJxkIVwIodsgHcCNEZ
Xh4vOLt03bDACNiGZ6yolRFatSzlsie/DlOZxrgA66kByNM1qLKqOShBD4d7cDcru5ekdGkhGnsC
ljgE40ZUgubzMMfFE5V62iJbZH+k648US7LXyLYlCYJMWxqJmFszWuCaBYjH8uj3Umfqk6nLmRV2
SzDjDKY8gq/AjrmZSlf9Lcnq6sivN8sOuZ6nClzgV+q6NWRxStDAdmdRjLgdaxuj0VXCl2jGhfCg
s6RrOezBcFh6RgMIuFobbPVtEQBcA4ogEss+oV9Ikai2O7B86XW3fqHrADeWByRvnVMtRXza/Qoq
vENsc3RoGaWlWdmkKI+WTf7SZCT2+NDjwiBdR+Et58LzFnpsG+dKH8qJWNxT/OX+RTULAcBuqCN6
UnbD1M68FtIaezlXgArfTjkpeBfyIH1PfxW9OY1aj0pr//eHOdODY8y5xLRcCJlO3oi7OVQi83cf
sFWT48wsBgtrqixg1Xba64IzkkHDgWVQZlgXByj+7izW+C2dj8jD76ERK+UFoQKYecx4oGFkNTwv
VZOQ/7OwydT6AtVT19QwPaAuzRCzGK0d+UKwJddi+sYdfeDzkb/ifN+DmeJBWVkXm/eGjEeEGv64
OLuJ1MC7shysYWru/grAIrxUsU3ZHB0sk/RsjWu2xdLI2hzOwhkeOt43qkHucEJ7xux8tytRE5bw
J/jR1sy/ciN4Da1Bi6BizDC7i2/+3f9PSrYkrhoIukYbAljP3SrTzuFoGaYmQgLSqWhekQh1NynP
r/HcPnd0L8yGHjhuvjBGQY0McW+f4dvdJUfbkedxES6YgBoeBYB+1PqEcNjMCVHqgAzKGXP97lgu
8KDPq6tbVq7BbM+xHaETprKXdV47kNSPJH++sIT7rUzmGyozU9FzjXrYYcjbwtWzK9F4nktYe60p
s0hy2xen1XLXKRLGv4odtpzxf65HcsU0qdM6NzuB+CquQIPsWNYSlpgY8QgslxzFV9Wx/YYkcUtd
KgYFSeuzEiwBgude3MSdv6ctm6NxIKvrt1mifmfbBhVoK7jYnxAZpJmXsrKkEQiDnOlZbBPRN0E+
HzDhbffjBhZ7kd7ci5Fr9f42c4agHmxXfU7+ezAHzh8xPlNdn7fsV7W2Th9WARRr4m9vBmJkb7Ye
6Lwl0hrLIvFEKdjMm4IOTlFCwyIg3t5QglCLAmvre21mXWyfig4dlUf3PUakiq8lXLB+Ap08YGRq
ajnp3loyKx0E7YaUgfiGUOFFkUin6P1nv/KEdYT6otuKWtl4NDBtPcD6BQ2Zo0uSvdP1JPUtc+6y
aIQw8mm+AVn71LQkI82UmUiVAHMOMpQnKZouvCq4/TFqcwBiYSt/ypPz2//H/SkGQwhtYtWGmwve
EqT9ADBvrzlSo6flqnKu8p2gvAmPmRy6Ci44XswNi34BR+ji0HtNeYJ57+uWEC8obfvvLdKq4JYB
b+2zNAX9rr96CcLLYR0iR+tIytx0dqyNLNhM3gvBYvjU+rVr65AlPNxLFvMLri1AS3CFjYQwdCp4
kk2QsRVVuVGklbDuDmvogKGj3eD1q1nTTqENy5UKnZktd/pfnzU2nNjg0MQ5jds+OYrqUSrk6Pr2
telLmeF1FOHpFQzfgIExSc8mAWX7CR5WpCSBGm2EGkrODne7i4mrxRzeGxTf5zElwN6p2pfrvjaW
zWmrdaKJCOlFe5ReD8vxiOkGUEQsXPGx4XFcT2SDDUtlRFH89G7imNccAP1yhsy9djficus9BPfT
lwixYTipZXiSeCu8E2E0ViaN9LVEaNifVKhqfMjvhh+9YMJC/haMctorUWls99nB1Ya4ZphMsUeT
HCLZQKtVdcfe9h4X2inhEExmecNeIUCnjgreyz++fct/0rRlFZDwEQeKh2HR8lZord5ZR8yEmr4j
LYOrnjeAgdyU4IAA86yuMyXJCQ0sGrH6SoZBJlaFt82p2Fd33vrJ69DOx09pB9rcZ+URNDwWTosm
YGcGaaawVZ1DWTOsTe4y2FR/KA2GkjxVQHH2cZ6lnzFitmMrS04MeYlAOyO9+RIECXFx7lyU1jCY
o/7oBj7dcsJRtYml5jAvkel68YUT9fUn87YuGPc/peDtbIBku9pT1j7Ok4OJqSmRg6nG3w+E2lJs
Kx3toNVakIxByjVhuANUOsFNP3xjTTin93hNb91WtcdZlQNlb6cUFERZUdDsfHTHxeQkZ0F5fvkK
tvneM7+a6Kq/lB2UH3bpdlnhvjqWI+ai/tRl/kX0cdrk3KHI+PRrgafueCwhJ/V+nXyUuJ0Wg62o
TI824U/1b+BD4eZs05L6LaSoyL7rTaVUXaEPSpdjWtRK3PN+WYUFdIlYCOAoSc1/K8IgAiyPvCoZ
4uEtSfi/l8iNkbDM67Tgo/qexbApIi1/DpSLQ2mE9lqT5d8qOOlLbLric8ELq7ORtG5vg0X0IzxS
n6eNmtB0xtDI58kkdojw5FaN2HisOSdz1vNOTQ/bjnbQj4FnIjR9T0AePBm9k218LR3xcjtvIZFq
yxPO1L36kqjuRveQ27+1TpZC8dgAiwfA2cZErkOY5uFdSGZaK253qvKv3wXJQZmlEGBZDkuRyeWq
hKXPXX68VcLXI1x+xY3TPDFSkTibSQf/Sb1w7NUWsH1vF6Dz3QzDdr9GQ3dA3kAkYepSn3TXr4Sh
ysrDn+OLaxN89a1DcH41A9aSBvj6VnwpFYybqgenA2BZBc8T7MqwywTM1gEwjwHsvPMY8M3K3TMb
YBpA0BvRodFuqjeFHBdYzBKOAxpSH3ac+i3X1gy7knRi4vXeyBqun2H84ZXJl21/cA7h+d9+w3ta
Y0PoPr2L8I1FY3wcM8OD8DVydPPxuYAWROGu/VlFllzC8xielRILYTRYinhdmAwBV2bA1gLw8Cll
6F6dh3Xwi2iGQxIrqGaAQOIanV6cLy3ajm4Zc2piNz5Cuft+b/Kwbjgz2c1Ywc7zsEt9m4bGjcwi
zHH/PGjSBi2YSCTuprsIk5HzblEhgvAcP8qo0Wj/z7BIhfQ6dxIr975+Dg6Gp6VshHiuyfNZXcLb
8S5zKkH6hcR6N+4rjCCp4F6QxSwBKILkHnH3I0dK1Vd818ensjCtI8NVjskinNB/I3FAl4N7Qhww
8SPa+knKDXThGTZWPulxT9YnxMHzlSCMXvMHuil/Idv8xZ5Xjbf9k+7+MXMgCMyyc/e6AKP18bWO
lG53ualyWp0G/kbKQhVkuzUDF/FFaJl6BdNiK1Q9uWXC5zhCVUMIYOwDIc16WifivgTpPLtO542g
19FtkT5OXsTijH0uYWuZFx80ky8Nsap1YgjnfqRp5vcHmzwoS9QIUt9sZJiFfO5N8QqOak6lD7L4
9xuAluaARMnNbPg/USbtfTNTozymSwBYXPIqAb3lHHQ0PkPf4JHGLEOpxrly4ZrMPJ4XoJVZ26mU
a7yEIKgf+pSGK55Hw1OM/0b2mUu3oBISMu1obenlG6tZdUCHIBqnBZmqFo7DhbScbMlTRvMKl2Gd
WUCXewAaP96S5hq8O1cTYOOwhFkEbpKk3bxFNd2fFWKSfUhtPYcaKv2N6TWCPaKJ8/TqBR1QhIba
E4Owmx9wPKNWR8XzetNxFvpyEbibjM1bOYj8Em/bzEm+USw59mTjGVWczTrhdQcmeOKfffPBG+Mu
J71uhP9jpBZFubyPd+9psOdNOoOPxtxsRNqEsiEWwQ2CzupaRIxpRdR6QNVt41ERGOIUi2zEQsO8
Lo6hZ/NXgLK0Kklw4KT40U97yclymc5EOYpdHL4WWuJFqSpmgcFwKja1U9B6LC5Fwk6WygyFSwev
dH3w6ioM6IhiYGDmrKnKZUORJnp+XXq7kV7ikqixkxuAenW6y47NIe8u9KdPKFa4h/f+TNQanMli
wztQ44bW8Un8WqqwLyk4fcAiwo0oSXPBrrpZCKvT2lZSiHgeNV56FOW1GVioAncp2ZvFmaejOTo2
SOPUMFxwZxeg8nNbCIW91cKp9jZbJfxdkOcjr864xhuY6QLXvekyJJEz99FxeAyfdEBWqVYoxXUV
4RWl8nRr8UxohOYPWQyW25SZVhx11DpYEIf/Zq0X/T9S5pG1lw4M9M7NgDFc6qQoAPdHXNi98arf
qZQ0y4buILInkYgLu5pYm9MaURWJ6gmxZ9gJECv18/5rxd0FITDE/QifHdsI7yvFzUZ+MWpGcJ/a
JhsP65/3YQfKVH7YX4LQtCqK9KprtJs8EC84OqA4N18atHwNWGsStfzjgK4y1u1RCUuEjLbOPHpK
LCj0Z/uDD8IcRz62b2MdkjgUH36fWfYmtbFumO2tpQXe7LYxRJ2oIiwZi0ThSDxeQnv48Tg9Se71
Bxjp5cqPhYsS3x482ZmTg9MJs9Ytw9g2KNZi6tFQ3/vtvLUzTl2NqBGIyr2duoctxjlrhT6Gnn7Q
2GfHqdln4EXeQCKBOVJ5+r/qfZgoXXHs1nSC9lChA/c390d4lqLK1XvbzKIC1LxkatGXBusWprh9
ZEfVA320r2kosrZp0Ib8SWtw4e5L7TXfQBLTesuSuL0mbs6wsfwm5LBZxTRVwCF8yxyFwqs4YsTm
Wt8XPzJM/c7u72fMHEgcvnBcgdulZwQnDMnHmozWSTBZwB0zaPHzb6ATx+Xt/q69toIEUWNnvZ20
DCDtu0vE7FRrjzJ1kvWSi844/7QlWx39Z1EGNtC3pYU3owFfA/y8ONwBnrqJ3nEN5XcbVfmBXr8z
TNDufWE0x1pWU/1OsN+PLgzk66H6iXBTH3X8cJnIAMBeJDIJMJJGFmeRO75REg2QQn5gKZluWIN1
rvRFKqP1scdYOgUOvqoLnFTtdqap8YhWo1PbkPWLKgxlwsW1Yhs4nfG73lZ8y13Gybg7tULwF48M
AjRFBUCOjcRAeMEfAlPVjJXPbf4/KNknUlZlJ/atyoBWqE4vMW/kd0UZ7TAU45qOmXf1t2gqtV37
8F38oj9MPcpMDq66XhrYgQwmZpNkm2e39lYgkmr+K/gau8uCyhqwFGBmwtCe+Gm4Gwwoybec6eBY
UzH7nrAvedEhG6duWwgJo3t0lEd67H7K3EsFONXmK0zqfwKrn0HSqtb+C2/iChd0vKBWybVfBVsp
j8DaaeUXmTFsAj4sZmn7Hp2ra5K8MqRIGTo4hTr4oAXfHma0kTRtGbkhJQUai75xa79FodUXWeUv
vkyvtW56gry+fwbKfqdY4fngEHCKjj+3FqamU86+LoLisnf4QlPfQ6j6P9vOdyw8yR5bGurB4qxw
fTA2cAmoQ/1QIzpgoSl179EKSTub1m6D6syizSNMgsPzGz+yzViaw8C2OO4gyg2zjqQjaX3sqdCp
RiWWzycRIPM5JPiQDgATStJBnrIKDRzdnVU4aYFymhxBq3MHWbnFsZwtWAW8Upm6x8sUiPqfa1F0
t89PJ8iM49UIx3n76aqd64hQuWTO31vaIEXn91aoxTwapSrJsmTv3dfDN+jjiSJjfDFYKWosF3yO
uho0KldY0j5A7FRm2LC/8Z/mSrwShzLjcWg6W/IgDO0hawD0tQXP27m2LmJP9qv1qmxOs/8cgxDC
0olHljnvbJ1l7US5+oOgZJhI3kMA4USWpJBFum1D1HdPBoXX7rewlTe1BjsHPGBB3DagdfKTEscK
R2Wa7sH7Ye22J+G6QPRGE99o22JGgUq4f03pK8wByzzjRZ3pwoeCbih5+Ao2iJ4B6F6DWybh7ckY
dCEQSlIKrNAijbFZpTVKGZI8zVdw/KLnCGG6nGHeBVoKazKupuaRmdT0MN0zgrEZYGbo5YmBCAEM
59JO7Bpfb1kiJnxDwS1uWQDjM2jkK0ohPeAm66m0HFgfZPTcFAVRQb5+ZxUJQGlDwXcew8dcK0bb
LFWCLrklMDEJw9OCSV3yawkiqwpNV8uwalnF4uyv6VZG9rFoi36bbiv6j6rQze1YG876U2fnfwId
8zeAkC/P1FINCBiinlRKSUYWRa/CEjocG8fE73Sy+Co2ikMOMhRHmgtUecS9KpeGYzlqPcU3lwIr
OKfwSAeeSMwgo6C3sjKNTHkPm2rdoiwylcbYN2RbfRCZ5ZCdnjsbmfv2YabgckuLa1y9e0I+4gRH
kb9VrPBroKlfqnmP87lVgTWgMKkSt3PBe7zyBnmQ+NegucQr4B3w9loW+ecpsirJIp+tAysVGCqj
+ebTOHQ9Cq7dqGMbcyt1RsH6rYyquE5qpmDfpjY/klfPoMP/Fby93V2PxGW6RPhfyNBOHKEsN9Pi
p8eJ6g572Y+6TR8NbZlY6XxiGboYbZl1KvEFoeAgMT6L9+33pV8rjNvJB+6Ja52mJizFrn/VTiqD
i8sPri9M+rQcwj6+bAva8AcE+qek/4a1RtlJ69X1yp4JZ3yfiaItvLulo3uxf6havOk+Mca5kptK
ZrLyj/VvWI9sHmpObf7fbYv7HMo8zvRAqUjRGyLFcs+j07cdPelrXsqEW/p1FOt/R27y0LFkr0I4
PLYqh50bIvx0cohX6Gv4sjz0SzSqrK0BNw3ksuz6jvuzhVuL+KFj0ZMZcsb0kuAEPDewPXlJTLgf
YVN3hA0jHwU2eYjhTUd41O2lUWnRuk03YZBOItsnvB+fmlexzDlD5yvln9piSO7a+NGNlh85aq3m
9Q4Sro6ceT7/sKC1YhJ/DJHanJJnmAazN2d8grBd/wNz+lGXMgp/bBUd2lhbabErqRTpBn85vnpU
ifHdzpMlp+/jog4ISYXkysW7qtAvKMm6KnuXLovMBuv14QN0yVJuagedFiW63hd4XYqw9UtVLHz0
fosTvNLED9S6C2WVQOmvGTO5rxdG9+/IXBZOyUtUApvMwEuZVJGR6ZU4hp4QPDoU8de1pBIZl8hM
lZLIipAZvmCybFVRKO/ob2xjxhnAvIGWl6QyH1FE+vGlDdtQpBCNRdEi823CPCsrZp27koX4LlKH
VQu1qSIiLpxdt5iuwgE3sAZ/Kja8v3C67jxtAA/pFVKcCe6nAnBuEkaqI8txQeALujuSz0YwIuMt
5jhbAVS2ZK5j3W1SY9P34roRW8ZSwNmJ+cElx8K77Muqr4DLgtd+Jbtc4b89MAls6KXOru/1ofU1
WBELk2CdnrWktsWhmUTD290qFasd7kTbKxUQpqDUyra68WeDzIhBXDyUp/ocrhiJSr29+Bsa5ka3
O06KKdYOTWyPWKJrpZqb8FTAfrWpDkfcYrAaxqy55HpaIN2+KkmjS5h9Ptb/1sE4o5WX+AmkdJHy
8J/rpS7DOpHhkbdeqbc+gW45e1vsgjaDSNQGTJeQOqQSeLDPWG2oDo35G+B3Ff+m/rN/rDyUgsxI
G/RQCQuetJq9mkTg2Z0gZq/TdQWO0mqkA3tRh64Ecu3IGJ+kWWkwrkve4gPyvM1vkqty8a2vee6m
/K+i73ufkebxxvZuDvzCgnTZdmTS2TsRVGDbAG4TDZU1phGEza1hgQNKgHXPdmxTYVMmdSHDOc4G
lsR4+BVpZSBnRK0yNPbWvAgMBrSw+nCJz6DmDVetjBzTikavlwiu0veMOpHusn9KWpPaUa4tpnDD
GFMjuSq2mjLvsfra+4D4M+UtLQH8tVDJu1buLkFFDnsLoyonQyJDweYCqycYXz0vHcVypdXJjmhm
ewmvx34izgXqxO4lxEdSt16gk161Sf4Almj0IdGqpxgQd8RLuouLGNWcK6sWH8N7UNdjM8X0csHe
YYM0IpqYO4kUY61u2p/HT1nB8MhNi8elG7ve2M3mscIACCf37q/dkpnGn33BZZZSZ+/dlkzm3+8o
j90qmuBpPSS/qEuwup/opf0yhUSwoNu5fAuHzp9RlixAmbrC0lSByImcOKGscO1PXQLcMb0OBw70
PhBX5CXavZQdsZO1oJdmzoesgp2nbUFh6wNIcHjJbTBQD33ailMfLmInHN/ep+woIZ4sYH78vJHy
5qPamIKnxvL9kXNzN/ehv12mU1QR8Za0TWq/M7d0JqpjvbXokrDFA0i7Hs30b9rpnz1MY4bF6IBu
GWzeoQ66shNwKHsy3srxx+oj5rqn9/rb7aXVWosX8hHqilO723VbtgTIbmwU1eRmpElvRVeQTI5C
TOQhpjZJBliDhpxDlv3no1vL2E26GP9F0Pje6mbpth72W0xROr7mk7GxbYsP8a8IY6p1/pXMW/+u
BV9ubddqaRLq18wsUKhG5U/eMJgd2PFAmpFJ0qea+t8Gh9EkE7pmzPmeWRyxzY5IaW5iXYsYrD2q
k7MPG6s5DtFWHpStxcSiUOmvU+zcMvBHJ2LAPAWlEsK1T64JSt3nD9HdRum2HXeMd0f3K2Cm7jJ1
4dhs4X3Bq+vAHCHz+f0sQWWvyACfPJIZXQ2PXpPCXdi9RnaY/QSDw1CKryU5S3fZdKmoLjH3S6P+
WAi6VoOVCsJQd22F5eScyx44+L6qp7S1fAYycAbnqLWDVoEPO74DQNeIyZt8iK/J/dS2ebt8jKcn
XA2e5pvAXh0qdyOFpWm7LJN3EStEZLVns/e2CmOs7O7QWNesGt1cuBDEyz9nStb2m0vuvF8T0JFc
oPMD5iSd6NAgoUI1vFDKmcMctdCF560TyrSHHUsBm+D8H3DSPd9oaRwoEddyIk2sKUs/z3vF142w
YkypHGO6zJQp/ZyBoRVrNVwfXDMFl3TfkgYsvdpJHbKUda4nTZI1kcGKGcteEXHbH1LfjcCuSUW+
/1cj36csXqS0ENJ0dG7jiMvBXGEdSLtXDw5X0UN2b9dl7dzFBa7MiCT8tAmyb+pBPvLRcWiRHVY8
JUWu1e/L3YNlNrpv/NgQ5q55T4RYTUzkoSYGfxdCwq5bLklgX7Oalvb0vVKaUACUNsCiVh3q9CSM
pogKVWMgJ5YmkRgpse26a8DJCyFlP8q9RdCQdGghhW/gYbxUeUeXc3RFupe84IGmcBGOAMU7s+08
OQbBL6bkWDWPIhnu58ZG261uj9SPPe75mHhyMuFDzaK+wm55cLSGOskmLLxuUqzwzyCmLQohuFx/
wiU6ksCfjBhnzYxAduNTjQsNXgN0xmc73uH99P3wsHY5kTJRNeakonMcUTDOjzrRPJ4CNng/OYGY
98FbRxA/qr/YPDX0lWANLTIs2fxPNxa5jGtQj+iySTKyP4Q4lVtZd7uDGHg0eN6M2JGBFqn2/OCJ
Z7NMuhlvaZlVk4n+JUhLas0oJqFkvfwg6lYs5eZT7p/jvVnpBR/fV6zqUzlbwftGQNnVDERYV7aS
n4dxbTEZrXOuv7IlhrciR7WeU+71/zP29VqlpzrTr2CtQ3b5zUe0VNHttY1aBsQGkZN6vwKDClt7
mClVDun89mbcwSn+SjCyZMbqPWsZWcI4cCf3opeZSpC0frCKZRc/P9nai+lFaXdDrDlNV8jTl9sv
SgA5DU8qvtpOsFglj8ykz5LUQjMxKYqL8cL0GZCfqGZPWD7+QSUcftQKXFtLLZxHvOQ0EPHkficS
cMdAX3X/gO9yndtpPoQ44A26zNvnJupp8DFJIliyQQ50F6/t/DqLvJfrFUzloj+E+jLEEb6FeGII
94xTzQMXOuiOKRcDtaa6IfVRQBK7zxRGSRpIr7mJq9RR0Rzav3354b55ret9S68Tu3KkUW+JOOw3
O75XjcelhWCefnoxFNjmjLwBKcKI4rqH2cMoRyxhVL1UExfg3AlFIwU+9pzLobDZBBog5AzVAtTK
ohUoKZWqMJXfrcbGUw+OQB0OdSUZRY0ZrD7gkQohTUxt6mshWC5HnNiBbQvktdu91W3F6difaobp
1tYzL3Fk5NUnqyLvM9sEgrmkHS/VfOYNR0CY2zc9g8fox1TYAFDuYanzJbSbID00lVsedrmPFR1k
GusI8Ol3m8yfdt3GvS3GehAr4epQtLJ1inAdoruSbXehoMcJt72BQTRGsSGbWZrGARYWP416yun9
eeU0KGMGMmCANGs0IWyLY4XhuAAWTyjkhJqhPsD7lH4ZXE9EC231RGqMrJK6rpYRGJ4FIM+JaumL
cK3HRpWvBTBrbc2mCCitwEaS7/uZ/r0JnnjjW/0uC/BsXG3WPPsCMJC/gQB6QDSmZC6WF1YHBwSv
cnrPjmAfVS/zirCXX5Cwn7F2VAbFUIv0va3oZgTWf3b5VT5Jb3cX1jJhh8Yqg0Li6Gs2/gYs0iHW
UEF266EN7KPcgX394wFLqBpVUb4ijKgYWRr3JqWLcknLlLnjIx70GS0DYy4hPb9IYRwmurYpX83z
65+Sij7dhrAkE/uU/Er0/dgCnw4Kv5QiLxQDQPNQ9XKE8by5KHts0VnLju+u+RGtTFHEbtjm9sxS
rFgW0S+NXWXGicen78iayCWLGIRVp8DWZjPXre/QxAvqtR0jTrK7I35tylG4ZYWZI5kthovFFY/e
7LqHpRs7OKto7/SARXqKjO5Iz8aN3vI/CVpAB/wqJ8oBszH3rkDQepWXAFibk9MDnI+fbIv60sea
uX4Yosdft7PIWDZcFoyEKX5nX0cu+Dex5kw3BAk0vHMUCmTedVlekm83WOR5cywcjNor9R+pVtwA
i9uf6Iu8M78QAPVPHu9deHvePZbZKsJDPMIPaMn34WhqXAk/rpznW5zKBPFytCXBoRLhFL75TJG/
i1sWmoPBD3Mz5L3nxgsX6RY6uJfmzkSvfz1w3Q5nYP5ZXtz0GL8RImZ8Z1WMJACI9BErRdCDXhFz
WiqZrW+88WJoY6CcLKG3TE/WYUH/hXk2uDO+LPjSQZiDz+IeP/wFiKdwKgNphko3iAoFISqk3f1r
RuJlxfJGCQyZCIQg5uknhrSLi5avO7jyK1AIvhuMf6P2+ZevsTmOPnvRp4A7v1wo/x5gcK0Ga6ZR
+HV/6fsk56Tz2YmYemFGU/Du7EfEpugA9Y6JAcOAPcv/0wjhJ2N6ky6wRvrz0mv8N4nfxYIx5S7p
xzkmJlIvd3jJF70BkIMY2kI2FD8Du/MNAglPvUy50EzT9zxmOqTjpKwmYiYCniYWIcEp3mUoJTvf
igxpDL/PUTQGfJJFxA4xkRj8a/IYcmlJuvaQ1wyQKs8RQ1TzYSDgzdGFZiSf4uPBiECIX/QUlyi5
AjaahemEjRCdlh8JkNilWb6Tht1HnqYxzqZSs09jxxjDkDXbqulaAVfH/01lVfICIlRs2lMCEi9u
N5CVloWetAbYn8MgX639VUrgbWNp2xmkdTz9SiTEvFFARjV9SYjKLwI+IvbP7vHNLumfK9kK4e+N
RQHCQ7rnBCGazDTHk9ZxG3o8t6f+cE4vDMZvZhd4QBWG9PZu3LGBAfdrPKqQBdI5jeRl7muvhxnx
46xRNG43cxXY13vGK9WBu3eMyzXnZXbxvNjc173E5hKEB4u44P9Z1+nSCrf7sMvdaHrFs508iaCD
8Sst74cOvQX9QX1oy6po0r93jydqFlztwIRjJKRPmzq8iDnlg75wVpKDjTW50xOGdJgS+ttkV/Ud
Au3y2E57KuACeuc9C+GnesG8EoHnymbqu7jn/H7mxJVdpnDGtF83QeJFTfYZWNEqwxS6S2KEaT/S
q8UZ0oWbM9V6h75XjBgeaSO2Za09l7CueK9ZwI8mVvbv65LMZOGAbPAN3yTOPHXQOTAFibt910MF
4OLC2eEPvgJNj71Qj/gHLoPOFJat01YvhNljuMCQogWkQbf1gYc/Cj7uv5CRTHi23VMf6udCosJC
4bvl27JzFnjRjAIh3tO16KBFwHTebi07yC5HBe0OK4oiCdUEO/M/DACw6HAYkkBqkEYPBnWbbnp2
ZlD1VJ5PkGeGhWNx3P5eoAue/jVdEOc2clnk5RbkHiMuhTsLZDUr+ruHORTYRSBxOY6g2+b02GuF
ch/ZhY44N1yJWk4CXS7bOF8MOzolPYAvrobJy7Oz8vEjronLAFna+2FNnDFA08mZE4aeJwqPK78F
P1H9KakTmRMPk/ISJzHk1hWUn2Vqvjwr/DD6hxg0yfGHzRM6ybBYFE0ZW/tUNYopSpOPDX7RcVOR
nBExO3D/uGfm1c/PkuHMW9YzjXJjI8lRhG/WXlv1nHnUHBfZJxzre7mGWyF5HTbgFvfaWdXkFZVQ
8tAncn+ZV+7ZkHmwY9fwp1TO96ZKDzJnSVJ1FFASaBYKaWntBdxcmXgpZFfsmdm1479eSSO8ikjd
rFGlfAIFLxmSPAVTg01HuA1DhnvhGl+UvzCtHXwrV0e77r4PH2DWCOIub3FwjYkfipLilPQsKNeU
vcm9V3TfPLA5JhDEL2ExFgqBav8WeIUkNIPWLix9xcV9q8TzaRrnv4rOtJu8ZbAQduP7TVlAiQXd
ps2MjTYuMl4OieUV9fGVn3ZRu+dt7r45842EijAfz83LckaM5hi+pR+bsdkc89Bmi88Bdt20Myaj
cTZIZQ6cGGUt1BrWoMzj0NDlpnFPDyKoLMnJVaYU12miUOrAdKn+YGTOMbbYW2TRNJWihA0IYUWK
obYMrlnyjQStQ63Cmz0kzmvvPOyW32Vfs2mkGxtLFDToMI8pjTX7HBd3AVOqsyD2/pgHZfiiLDcu
rY9ANW8kSoDyUC17HLnSKnOuxwRF47GCz+5f5D860FJWWSuVBmeoSDor8Xi7JSloveEOEQteoIEE
J8t+rlb2JyFfB1A7upcow1dEj66E6hNogitgo0BJZtKKCBM/m0ZeVXHuHKpObZvF+w2mn6Pe6Jli
pewIlJrMa1h2DKB4JhLCoKT+ipwcGckolXRQfq1W5O2r4WDoz8L+pfsv7HpN2puytHVhG8Ac3CvN
zjeQZtZRwPeSlh+aZhT6KXEnZ03cucx5NrnboUUqzfRRSxmTCwBFZbGFV1rI/rFwBs+3Z871zPN1
GCumUOVXfDbGaAqSxGAwAtB/P7701U4SX27r//kcUPucnVBUeKTsBvxRW3HKT728dlVfNrDK7/f2
anhvDYJdVjSLtDfYg+kclMrtsQ4cAsNnAOaBvnBj54W5y1dK4A9Yor1Rfts603C1tojsJtZ0qPYf
SffTXHEy2tfp4lWpRJNmlS7Ld8CiZECY1qxzB1/ltyd4pMM+1492k5/lWTRaFEwGh7NsUjpMV0NG
WxPhI9ff5RgaZmQ34DLolU8VoZ7In0uJWnoQ6xzwvG/NmYok7oQqbTRd/M7j3xAvOw4d3QFvsUFm
qq0NQYTpAEYJYFWDOLKOPmMz01rVTnvj30QsGiETOl6FTw997lnxkwLRPjy2N7gfjiJYvqU7coEo
NMyCOIvXpQVbDsw8HosV+TJjWs+pcxgYm7PCeu7kdYsafC6iwxbKIY6EesfJhax0ctn9Tg5ODApv
m8+oNvJllBgpOaxuPVO8POZKMUDJli4mGbfRU6cEtiUe8xBqnCy5SeDgSYBTegZNpfi74T1KBW/B
RAE3Pyi5bAOBcwlFzdCFVKhQSGS4pfArGM+NGWq82sozR7nCdHR2KcgadwpDJEEA+rthj58Wt5wy
Iy+gKrJBOMlkeRR+JYCTBO0RpzTb2RFcHW9GYy0B0sXe4JEDMBFRGTgHaUG1ItbUp5SKZAbKOS/A
4OYbpVST26AkQiClc5BbugSK1f3ktDFf14QXqZq9K5foKzc+jL8wztKaTVberQzJr0ev6v5sc7NO
4TPZ0SBF+To9A1txPDdv+y54fUXyHW1r1O0lxmoYiK3hmQWZR/CzEU3kuKkrVjOFbdF+EbT4SOjK
Nd5jse1cfjAgw68Btw4D+rOUcp4e4AOiKVID4OmSh98ygraqitff2sJL6v64vhv3UZX+PYHnogIk
JR3rAWDj6Y4qGTapaa3KhMlbdxT3yYgOmoTE/b/yhBIV/OVyxYQuS4QXOH+M+x/ylZZzZo7nWBqK
+I1vdFSwRphzUOlMe/4ytCZEfS5kX8dZDr7f9j2T9NjlPFEy+j3ROfbMwistK5zw07Sn1Qc8MZFX
aElaOC3FE8jxcpcgyYg0rCSr/4uiv3b1gvTkeCDgjgpLgoVwOM6iufjwbptpqjTDyNgJZbZJooUu
KudPtLhEUxsl0bscstR2eR2EwBL/8fnY6ZIxdgzf75202sLt/GgmYp4zateEpPQBP7FAuKKHQuaH
FJ4gahS/aT7LGf1JncUwb53quNUy9/J3jcP08O3B0J8Q3OnR9mLznK3uqQw6blhk1fpRfaCPpiEK
PleS6GiDJMV4eyqCobQN3kLnI36Lmjfa9qnvkakDAB4nfgEzDN6Z78P1oGbyuL+RcEc0GnLg8iTQ
3ycFMg/z34rxi9xM+gVylXvgnOIg6jM+bR3QXBGh1RSbF1mmkzQ33ME/DrBDj3zJV9wrskeEHv49
Jt0FDnWUK+Ai4aUsOlSu3Ny1tLUQ5M5rXNWc0IGSJ6K+xARWI1382XREqf4meUXk6aW8v5Hzo1lH
4wBwqlKTynrWLSycGqQ44Zr1cv6t2rxTHndZO9HdZbvVNKgq0idwPreJCCsKNh5X+UGeSJo4hbiR
CAWmxdue03FycTeErTl2C+mzAK1SuN6GqpL2OAahvM8jugfwJsEsrISbkr2lASWqmmt+T3gQLSQR
BSAq72Oqa+kkrlk4S9MljgZ05M+Ayiq8AL0SjbJs6N67Yy2DEKBpy61hiUGA5Q79Dag4im+yl7DD
evQ9KaAtGM65XkCCPvXtCWEGFNhQGkDzFwTmyF9a9BYJ89ykmvfmbHd8G0d7BP+BL1AeNcz9WROr
aK6uQHjTzKrJRnNNwm3AvXviRvY8EaWobKzj9wsId1/FySb1sjg1dakm/WADvcejL9YbWhBUbdNx
Swv9Jb3M/gr/YGszGxxjjEI7YSMp7yZMDL9yicmYm8o6tQx7rQbKBVg099PqH9neLeamqnqzKg3A
lhSqkyKfH3dbRztPDhUzR1ZKoYaauqmfLeGdpOw8a9qNPJNc2FhJlb3hw/18nw+Oq074Gd2Oj1A6
QxLA05MM2V6keHMfZM0sf6tJcQhP1GqeJFykxChp1u7zUAFdAn06MPiTCrS2hyb+gqcheBHL8JDg
PTQytPKXsUIWRucbCUvewwv2M6hQLiyHOHL7EE2+QYiaW4Kah+T34pJyVKBBupkN+Wpqvfy8Qmxa
VRZ0w8miJFgdyRQeeZBOq34K1KE1jG+4CEijTSIR4NO7xXhRzT+xJgt+tiwNWrl29E558UrdDshV
F1u3FLa5p1pmNEtuus44Xs6sB2pUY6uC9Mscqu6qKsKbSQ82G2QXbo0IFIJRoW1LcJD8ygpLXEaN
W7LonNpDsA2xJuz46Hzl5zH8CydYwOGE178HuaNgYTUq1B01WE3ohKVlnJAiFMt2ryYb0POL6zLs
FGpr107LOKZDeJqyHYPbQ+u4TE/7uv7faP8H9xKyRlngnJ3ekZ61L1v1VEVDzZcg4tw+B23kGkI5
JrWBLhzRL4gh8Qq0+kBkfS7S/LP1t21iHCTBfOUaHjPNY+Qa/ujb5jqtQOc1U6E6F5OHfWrSkM3M
knGaLM54pAbCmGOPa+/IZ2ekHpNyXv17wPaw5TKihaey6f3Nk/soYBZOxTt4J4XKkAXL1HUSkrzY
DkQIZIdR9BM5S+YHg1uqZyU59aZpjOUFbKUq22T0hWek+xmkdzJpnJBQvzJLUhmFrQF43zkq7cvU
X8QuIUXK+1MfLY0wdxuf09/u0iZYy/cMcDbG3jF2S0Q/GnU3kgq72kXVgD6qqBp1Wm+AB9s0Mwn8
33u7NeiVb06FIv/ANihBFAou6bEYMtMZ39xd8EOJgwNPuE+JfvqIkonOigOdYKx9Bv5YPbhTsdPJ
xdPsrKnDMx943XbRsqWhRwL9uEyuxRzDWmwUjrp6McRCfzbS2YVluP/gMxGDb/bkuKh9sTX8MVJV
CJBfIH7HJ6jYdRAnx3G8N3aMa++rNpNrLfgaUZIT2ywbOvtHNVciC5Mg4vQ9E+5Vac3WFt4GrtSp
oOch6gxgj0ZkJkh0j8dO5TmCyZH5wZedzBFiECviL7sgRYEbXi9xlfuoy7YWGNQP0PhILFrDRepq
fb64DSU8ndv8bqdn+GTXGQJgLufjsWmeDVGyD2FHm+IZJRRqX0vureBipawwltBTh+gaofzsBU4M
PwoyLq4QPza9S4DfXuU2rLEaWLi64+o1ArBkjzBEhddpN0G8BCm4rSH0yZ5cr4LUKzLrwfsA63ld
jkHnk0DQAKzo8BQ8KJkSy9lJpQeWQIPjdbyTVW3Q88ENoMtA+nGoRG38wwj+k5iypAksFjJtT1Dr
j1N9/nEjN0tzlXZyxqsjW2No0VXLcnEVSvhVNeMXNhagP6Sn4DIjWZ3PypRD1wrQ08rh3yR4tQAj
fce+M/PlCUkUgZkNYb0jR1Igz3PZtLvXLUx7+fJPErYb273/aFUHD9Q26HJXBe9YoszorqigQaio
U5QsqTBfhfvs/iDcRVH+SnSFxTqmMdudh1sgq+u127x16t3259jAHh+FBdSMoowQZcMID9fy0Oht
hLcULGZz5tf+wU8MDAcNe+wBqSD/hpqNwl12X/dNCg1uI34MvAke/LBpS+aXBZNpPuoL3MZW7zXA
3uAO3nXzqMXcwF+atGumKOWdvRxb+Q+TA8QzmGmtTrFR6zy/7yS4HaXj5Vxdujyt+UUI4nOH3SHP
ZrgU0oDpA3equCmFULTjtlMwEwLxfK/SA/hqRHTioZG7VgyfdvhebC2oUX1S8rKLq+UCUWbjMFIL
Db7BhLQwkX4ikxg0EjbmAN5jm562/ZQPzrFoucfrWipYao4HmUtiVQ2rqF7q6L6EXvI2l+6EZf0t
fefU17B3HkNX1OJIhdIYHz4Qpj/6En7oTUY+uZx3McLQQ/hlAeU5VrNTKkmHgku7aK42hmg0fyQz
GcreJJi7s8LjuqkSM9ZYbsrAX0BANzTfwv2FSHpcJ0oPScN5hyLC5JUJJkFulERafswx0sklBb1F
SxkkwNlQVSyFWwTI67OmEL2uKwi/W2yv4JUioqMCjXP1Fun9J6KLYiLZWdZUOw+/YG4Y82dU7Lmj
huXok7LlH8vql4UzGcIxH0xwP71dGP5AeMTBh/poKX6MDZqrjHkRjoDunW+KYonk4plY/4IZKF5j
q+zn92sYL3jBkZE4YBJRHcXY+hbnI6cG2Iedd4K0YKs2bU6SkWTg9+sVVQAJCtcVamKGcerSMoEK
e98R+uepdwpVIw1ikHNe7M9M7LOQhCK5RpMd4oD1rc+YxqkwsRssCGRULMfav8WgPOtRgBoq2FEZ
YVTyCLkDjdZQ/JtnLTf15nQqAYcToPt+RxnI405vPuOwiVgaHdmHOV6qUlqhpnz4DCcSV8/R3awb
sjLJJeVSyoPptKNuZ8fyiMMl4FmqQBXeYyfMwqSTJcj1MA7/VCOu3bJU3yLtolrczmLaLBJQqBbQ
OUiehXV/0DR1X5QQR+0quZpLTatKYFC4QdQ2/vBhYb9I3ipeil+cqZbq+5wpJDprjFRTmeeYBxYq
oM1o5TN70vvw3hgHT+t95ypGDdA0rLeJOW97ys9fa7itQpu9kG8/nAn+zUk0no2q7cTUA+un3Bm/
ymgoXLqW3FZSC3XqnxNwzymRIXxBzOpYD9BSAqW1B9s8PorCbwelrPph76IgliSWbrbKVJhMUPbk
/qvDN7XudkP1wT1pi635elz/T5L9coF76UCWxIdPljjc4AtGpos7sm/lSgB356yJPVyubuY/d1Sa
BM1BEowHKbVJdheGs39/PRcCGT6WPrXATt5OXTuHc86c6mSLshwnWKc6YLA13EuJg6e3We3UOgxK
riOC16mMTl1teqvwGtm01XiE2mKzbXU62jz/IiSr5Lq6dxoGoi5SNejGFSrhPp6QynKvB7k/x8fa
oNt1dEntezVVWku10pB1JDWiypZYVQ9K+fpb7MZmkohgXqZMboAO29Zgjh2zoiaoYaKY5hxdiEZj
ZQeByc1Kv6lJM5jDP6uWqf2DvIrIa6/55LYEc4v4URWNiRhTvA73y8u2pl3qO5rc88+CbVNjNCcl
6xXwlpbZQZmUIXik+WESDRbL0XOOyjQ5f/0/9DlAxdvGBXq7p8QiXcPnimhRW3awXNJHDDJ7h6o4
Koy6lHptH+LUjrrni1BNTmeiIM63BDEACOxWMJalc+D+jB241Z+izouIH3NKLERFeoizemP3Tjjc
W30npcGWNmBYpIN3lravc1dVTkLscvrrvfWToXrV7yopPvckY9GnzINLyGd2jszzBMLI0UNqnKzo
rYrADIlfUntW5BPR084mAf1FAlozIsAM/bbiu4kzy7OFKgbHphaNFO/rNybNs1eOIBtssRp6Qhxf
dJWLVsSW1XCvSIvnz2V62WnnpZERla22eTU6DwUe5I0qyOaSFLTqA37nsvqHgMR8IrLTHt/hEVC+
BEOZV3NySyGb5RXkNS3lDk8bbdTCGR57lcL96PkKCptMZFyWJ9d361QtpYXAkvGIUPOZJXnqLHww
lcDL31rtwA7083Vgnq/nBnqb2sG5sNNdloDr7eetATy42O6/SPH3oHFIR9YaycrHWTAy4c6x6v4I
YSGoxJzjEyYWXeAwB6uP6yCAvGBDpZ7TzZMCLf7XWAwFfDpReDSmX8jno5yh6H+Q/eF9KLHNVHIe
eX1eKviQUGIUW+fui/V5CrO/kVfXgiuKx/vHhupH8c9Sro+u8ozBPMKBRxpfmkglu0xqXd4xypUV
R+2XEuCZ/wF9okJEC8+UL6lt/cdVVmO4LTRzxWQ8wlr4n4r9aoQw+aSyunanH4dydsTax5chZNRm
bmw7rRVT7N8pqALhzti8XtfmIHRU57qrz+ztuUYCI4yGzcNbnKfOGsohvmdSREw8l62mtJJ/Epwo
LWMRzeKLgSE3UkfEE4XztWKyYD4TcV8SWf9W2U2fzknXxVu5HQHmmA+CdyriU2qmeNLy1McCmcH7
b6CjZq0dWtKiGERG3KVEkwlr7iKtOlwQ7rdLf9bNfJQ6DU7brZTA3vMYFFyCjnNE2P83aF0/bmok
2uyFZ+68fnUmeK/SHoM+K7jBe+IDTy0da82uGyg5k0jzgRxFHFOndEywajbVAzuaFtuOVBuWaKnR
JFa5HGhSG7PLX6qCb1mOBHQ+ppoec14ZO2VPeDnHhN0J9ugF389Gr6WlLn2PKoFzB6ehMr7T3siu
qsNUe5BsVNbKpYSc8rkHDGpntUlh1oefXOd1gQL2aomilU/+T4mIQy53qFNUgLA1bknLbnCPSSF6
eUxbxVPS8pw2Ml6P7Gg7JNWQpgbzhRGCfE0nB412qatQXkunmPg1AJDzd+yFd8TYsNRMzANjPoIr
xczUffzxPKoHLW9GGvboCLZXM4UsitNYbgaLNkjEXCq1GZDG3nIxIJD4QG2qPAfax955Z1X4uSQ5
oYh0AQdXv55s5HrfE6lx5OwaasU07RA5itUNKFbQuZ7GonQjm6qvo9Ch8b40FHEOXa+dASAsM03i
rw/hQNzMwE1pDg1Xz1ZFQb/gI1YheXvZFtPKhROqgROJWdYW+yABgcWsZpJtYNSDQj8OaMztVt1g
HBOIPPasJe7EWNsgyig2kQXq+LGZipYD3jnqKw4xXBbVMHc6qy6iwKjTYsfCTnqqtp2/zc3QBbgr
diFRBiuklGqWzl1LFz3ANNaWyDELrHZjAfnAlM4he6tNKtb4XEcIfVb/o9W2w7jsLw6Pa4ZjTi7S
L88sIpvOUlYGkrGUEih7cv0p/PcR3O/dUkC9sg07AsG+VgbV7q764xb4gBmwZD5QJ/OfjthHO50I
xDqaMM2SW+ar4Om8cbp0apUfeQh1Qc1Vfuu70jpx4wUcDkCKDDt+o+yY8vrzKOM5Pbxweq6tOCgc
cIkHTGpC2zsLC2n7k5Ggcx4lzceaFlqNfvAag7FCzRySs0jfWrxkilS+wI5AeuHv8mlN4dT8y9Nd
YKJmjChPi6ohycHYgy5wzf+vXnQdT7MExMJdWTDv3mbCEL5J+3+5cdWF2BwPJRRKnumjNUcHePHQ
ek/wXmPyjMQE/lz3yyY6R12EMJWg5rkl448Nr8gJXXIysp1onyZIjhv8RZRvr4q99NSJnynRJSLB
bfdngFa+zV5s1vr/RCij8yThz31lhAf702glsumgCEFVy/gGeRWk78dyZaFZvLOLdpKONMsjpjLN
+aNmIDyLoiXjjyUBQ0/3SlyHy3DF0Q1pFNOuIDTqc2F2xEFPK2h3GeYhzdQgKf2E3r5s4bC8MzIg
nVd2EWS34FBagQQ0Ax6lWdNwR5mdtiT51PJr3dndLVjM/TWeVt2Kkj9OdTEAc6I74W/SfdpShM6w
lVLmZApHN0XFhHTelKz7I5hV+xCgNLcmEVGI6PVE+DVHFboiiFD7fjKJC9Z/giMnc7v/diF8cm9l
eLCUNEcvAOaDmg4k04SVIx9g43yQzDV+w0JMdaKciYs55aUBeObOSbpKlnjoBc3URaHK8rHQUECV
cOzMv2K4UcmdDsEdZhz2etSd0VTP0c8Db04ALMiCmWIovZHTTsGAp3LLfmgMYqXkdt60CTnmIuGO
2koP5xvuU/wa46+rX+TqhNSihTY/6S9MHuNzpvyUUFSxodsa2pMwWsnoCWxhv9Sh6yTgH0QHvwVz
p6s0u3gOq7cm8gtYQucHuWC6Ebc3dm7rl4MGidhTW6fTlQEMkztdWxbV0dbllVU5BlnzXl8q84JJ
YtjzIH0C5mU0G9jRxkeMJV+Yfng0uJHSyYbIl26kb6eheQA2Y5gjestaUCUBsh+4f0IKAy2fCkyH
0mSKtDxOnlXu22exfVQ/0eSsbs6s4k/gevjZzVdUndCr7y9hJMUXJ0xZgon5Yq69hrmPZ3S6GKpu
7Cl+PykHjpqLEZUsoLsckNt98MjBGs6ZB6oewukNqNaD5bJsLpkfRmFBCI8l+7Uui2eIjLH8v8CN
E5FQl3k3/MRUARU7TG37ltVc3KGvI4BLthnVGK89bFMh1xgnE4ziuTKkhbl7chknSWWkw/kzf5cQ
EH2TOc05O6C169mxMk+VDB20pNkJ1qUOg8qSU79C0DxCsixtrLe29cBD3xCGuEPT5I5aDEPFMz/M
Rc8PZB5LvN7jtI4QZzC1TuMHi7b8Cf7wc6y82dyqtfNq1V/Vvo6xRp1mXc69L/hTxmfi/SeWfVk0
vLJkneL+4V1g9dHetTubby/8jlVzH3YW0cEN+pSkrVFY48r4KUANcz8ub/wjh1gHAPbrfJs0beEA
Zm7UUrH/MQOU+iBb4Y7ETOU6A0o4Ygun03MVfWVJzOumNKEXPZ5CZ/AkNsiLuIc1h6HVYAuC7lfP
LoVQEB/yn0lelscf+8wko0KurA+1PQAcmMApbHX2ltTUeuom2Ym+Ev+dw0nHJQkey/aMg94Z9O40
iscQa2umK56+ySbkXxSeks7CriiHTFdSemgM/U6eFricG5tx0RTWrBj+WY+GQ7hSh4zWe4YrRuq8
GA13UpmbwJcLG5iynMkw7v7YhLAhhat28dMSD2Yfxm9fS54pZVAvq9Kg0EQkZSGFWvxtZ8WX3pGl
xwFw5mYBGp4l6+KPco+MiACSXnUEkQGgELbqNCSeVevTf4EKMaxTyJL/9M7sKZrgs0rY5e9zRMG8
5OirrjVoa5R36ZQTrYkIcmL7gCgRuovQvLogWD7IDIURUBYsjsT/fM5YKh4XWr/iUpETzquZMrEM
iX+uJ5GFbnIaEKj32Njwux5R+Lmts1KNu0ojv1O82BDBll+6qSEslHGUfO+aj6l6nFuj80pC2bUC
rZhPeU0mzf9HaruvYylHJLkmrelu6o+L49qNKgyp8gHCBk/BY10uz2sPntL+2uqr8Kf1QhhGyGI3
kP2lC8GMWyGL2zKABigdwehS5fwTwANQJDaaHZDd2pH7+b8uxE0GD2Yilw2WzO9pdEI2uWug0Nxx
FMUX4zJPhRCjhtYxZzEjaaS28KNgggyLdyo1q+0mZRUNY3Qtv8IIf3LTgadb6lag7usKqbO6h2ew
/G8BPBdWqFBvL2Xmg5Mf8rFDoex6b1b8HHuA+4Hsaoi4qyIj9uLoyLC7/HPmELPBhd45aK9kViaa
njqdvmym9p0Kkz1uR+X2ZDKOicH8UUzgC3K0PdvtwOk+PSilF/WiHHcVue1j2PblCvjhTpWPdHVE
QSYA9vHiy5/WRHkgbE4b1qU2O+SwtIIODfVdWdjEZ0h9nz26OyOhoQ5UzamAOViGDBOhTFUAdKRe
Yc3eSQRNvCHVKVnT94eYC2ABsYvDTa38zyH8177bVsQb20r4xC4fOYP2f5JewRwcGumpIxO+BtZy
xogG/WZvYY83bveb2afagGVAT3TBbxLC+v8Tgx3uIjS4tdP1lfLsmfoNPNXqnkFF/KOXvXYE7RUR
Yu09vepeK4ucuJ21L5oQBDJOUEDQbq/0YeuE5jqT4yNHWL7X6qIULuUyPklqBCufWchM9h9jD32N
1hfY3iqAiF+sLyMP2jdhtbmoMt0srlsP6wZmLtSHg7VcFLnDzEqW0j2Iznab7FBhL+NEsYF6KikR
s6Ukll74r3DiGpqeb899WB7aoRFts8fzVwmqhTEdaxhnbKXSJY0kMe9eGwraZoeUknvBEs/oIHZd
ked26yYvNcfhhCJQlMZuSKX68vnLgn0uOucgY7n6OoXdh4KWOrfO0zWc8GXBYuqVhYvHwqeLt5KE
WhJsHC0gz+Yay0Xh58CE5J4UJ2W2WxUyA2UK6/LkmcJjtDFHo9hUjTxOykmjnqYxRrGkGMuf2lGI
LFb8ed/z9C5lDZ/Xa5RsZqdHWXQ1Z1YLr43pnsQr8xwSPhJv2C7FaHHg6Tz17lC6QCAxF4QnRbti
Q3z+WiixqMnBIJraraTMhtNKelhMcJzJhpfxPNkjCSqdzdEioDBvvLwGJnuwnEtb7u7IGR10FYkV
u6GlmByVPYecM7pU5a/+3titqo/1csu/VDsu7ZDDDRnLqYp7k80EG5CuRFEgIEjMhAAyOaWJqRvj
mN/73rXqrtAn1IS+If4citOaf0iS+leACD7U6nNQ77LIaLjdBbnNmeyfe8kQta3XhrJxcseDYGIE
pbIOap5eVrgGdL51+I5u4VNA1XFonXNi/QE7QLo1uwGC55s6pA2yz57RRkvCMwmdBTMT33vIdedV
WwuU/ZOTYnpvl0vuGU1Hjw5tEov0Kl2WD+k2twe33Z4yX8ERJYKf+hOjtYWSbYuvnFF7aIuZ450d
3TJ65HYwA77fB2WUu7902EZoUQxJGBQTkWsp/Zizuigz33JanIykAaNrt1FSIu2gIT70UslmTH8z
AsF/J550/uNY6QncwoUbbCmBvAsey/XlnTVEQXMJuPwNGLfdDSs8WaoTJcT0/aMOdFPLJ6PRBbeB
JIJ9aNGNzm/BLsy+m3svQyOo0ZRKSKKbL+URXNHO2Cd7wMAmq2SSrkbc0gCmhaIRIcSwmmDyZXv1
xw0yHR35y478MnDxglENJSYedQlU+q1sZpDA3uBmDgiNC0QGdAqX6Sv0o8bwH92Im4hC+O0HtZPh
4+xjwnG51ZqJxv9+IpprDHt3jkbs2IW9MgHSgXmLDKsKzdX1MccKYLcTv/Ggd/Ae6O7iYLiZuJsP
GcAab0nHuT1c2Y0LEmuAf8CbcmBEfVgeL5p0ry2DNTOZg0msDuH6GQTCM6u1ZxbUcpJOqkC2ALdz
SdKFSFlmV4+wetfbtg/iQU3dZd6Ivwut+bICWv86+oGW0BvBfDylnrxdbevkckvmNs9QrX3xixac
64gSAzg//E7ej2Abfx6rVnm7LRWM6qTXhCXOtQd861E5ewwu4bNoX0YDF8sSdrb4kFXSRiEaFnRF
qQXdSrppwYh34K1mYCCmy/gAwk/G42KjXUsZdWUpEdbSE06Q8291/4d01So/Nrci6vDsa1CP1NPb
sbl84Cnnk7vy9Y1Keit6lIMO3FM7DmEnuHFWrrLrksd8ote4lFbyrETq3ZC6x5OlyIzjgHrqKCGM
SatBtWglJyS7e+Bke9LyWpBoKL5h8ZuRrlx+QbLFGi6MpEKPpeyIAXCVohIHMiJpFVs/91ecljZj
7Yt/gq/9bNuBXfuVvmbkvxtMW7qzOwvDQTicbfxlbzL222u0OZadBXcBs96hxvWTJ62VvtxUigwC
lDLl88C9U2auBMVJYVh3htjBHHNsNglw89a4wXR6ptyk/Tze+bS08CQPRQMEAvw7u0HWSqnja2w+
VMJwPdys8Iqmj0z68yWiEdt5YeeOGIyDRJT59DkzE6htxGi4FjOtdK4lh/Ig52KO7iPQ2DaMAQWD
1DLPADFNfTNL1DvBpcnAJB8cTBmbW/2ewfh8VvKQH5YIaBnRZAEFXNg8yD0/gERX4gC/Oxxy/vqZ
cgmjEFxcnth6jBicfZt56tAiZuS0PHSYM9Y/PhxFqVniPiPokG+kK6frOd4za76zuTN5wrqWyDL/
ksP8H69EZs+kQUGEiA4Jxkd5bzzftIWRJPbV1ZfPwoLZnCsJg5NOUb6fFnfkrYQgqVjcqJ9L4N7A
XuX9J/E6zUBeDFhYlSATuHv3pwCPWzzHbwQmsxofGQD4mqRcW7EAu9PdtHpAkrH0Qb6pBkntIpHS
yVWs8fRcpBVBay/oB8bKz+v2ewCiOUWaLgIfw89zTC8/ZHMrOASIOtOmbuzCygq/CMPzGRVVC8r+
UHhPD8fr/QTIgArzw6tFz8E4ATqQzn5+uoBJAFs6OJcZtzRznMqx/wWLavn1OQRdJuBmMEygC+ve
riU2t5sie7qj2ysSSkMU3ih8I0c8SiQjDpCyiRHo5o13tnvqgO8L0JrGoEwHrAdRalXjJRhw5ZzF
1ekIKCMJw8usbLpG/lYsQJ9ulCfa2yHLvNq7XzEkFAWRH737bROqpOouGFd4o2B7JSAcegkRurQ/
bRmpq54aG0711jmql++jkMU89ItG+bAZu1MRMYnx2hOAnGkyag3n249SJ9Z94/9BodL5M1Egy2j8
oYqCQVH1qZHlqDDr0jUS6GCMggE9pJjTG3arsU9376kPlcb2b0YU5xXVHmhl9zg51sdCmaqD3zY4
25X4C/CXN951qQHUXQRdE1YHPIS8stjV6rixSXtB8oov9u8E4IJu5AJh1cpcctuobZRTeglqdA5D
ET/dDHAfCeKN/8ufoqfZysULuxEopEUWdSCNMa6R9+tx2NNIHrkPb2NkT1EMrnm1PnMLw8sdRuRk
ZRFDVfyE8bPN0OtTUNY0TyTZa1UcgTkFHWB4GlIbj/nSJAcmwRMFVeXCz5UtZhyJ6+uxRiRZfJEr
tOdWgZ1GvahLuFku3CHBdciCpLr5JEPJDUc4tGYWD329Uzd1j9x9lvcLoun43xtKlX1NM4dj064R
i2C+eoba3C3C6pK457xaBeIntRIWn4p4uovhjXF3z7CmNx7n+d7PH7fNTQUem09y/IR4Cw2FljhT
voLZUkV9rSmqG1ejX+jooy1YCcO4pwNnwWpQLyhq7eEo8eWHaLMNDwXpKS/J248BD+/AuLs5NWsc
qscTcVNL529xj20uYj0W8tVmVbXUl7pwoe8rIbnb0m+n0ZSsXZPOXpW1rkN/ptSzIrfsuv1BJ7XX
qInr3FuRfWZr9SO4Igz/XWQEXL5hp1BmF8/Ov3hAqB2KG6nQ9qLDtfHcL9xKmra2DMX1JGB1EaU2
VEpe1RT5HfCLvKM9eaJ19H/q8oYk6oh7SrWZRtshrhhth3LUYJ+W/OPg9L9q66Qa97B/c9KQi+v+
vilTm0haAT3WfN5Xyfi5zPFTE2Em5m8exaRJ+LF9Og8e4tPbpRRPnyOIHanWzF3UiltsbCSKZSUX
+zgtY/wp+hz3YR/EOfeNL+arQ+y+4QFcFkjiwizh1QhU0MmRvh5ebiWEgmrlofxJbA3bEKJSkb2g
SG0VZMHI+tLv7F6wLsOExL6R/yi0i+BkdZcMIae9ySY/1l6fCANhjuliyBeDZa3OyW+kcVA+wF7f
DU4+EEaaCBr3jD795e32Cmqoc2H9AfFUfdMcNyQFzbIBMWlwdc6kIqlgL+qzvR+V143r3ocBcz5O
Yw6FbzUpb+Tu/9DAoUAW7ozvYEkZ5/Ou2rxmEkMARUVSb6FBdL8hLiTZIrG5IsHwmsCBlW2/yASf
5GUAlzVMalr19y1FjPxAyd9Jf+WySzYWVr1IhJZX//ws4AdUAtr5eSh7KdnuXh2L+7RdpKdPVtiK
Fr+POVEklg2bZ2naXKK8YA1YUaYVsljuMC+nk+bpKYaZxO93xl3E6m/tD9pjjKwSa1Mgh21X9Q6/
DkVAVO4JsxVmXn64962CCcOAWJjQbwE7xs9Nbr0wrl9GBrGBnnP0FgM5d1CEbTULa8ccN2zn2z3L
0Vm0AJFhjuRKT644T2S6yrvA5FEB3FHrWsHZti4/2mMetzHcJ8npc6+Dpm7+OhojmZKYgyt11GD3
u1rL3k1bmjP99xUQPSAlMLsd7Z//yYcPQdvFmlFeF4IBJcbfKDMYojCLP0dnHwupBPeRJ8HpU3E3
nhSNa/zU/qlTHQ/+v9Gkhw5NM4I3hhCbeEsLO5Vba6BcsQHYOZmfyuR9mJu3wy6SA/ZqaFv/6KD/
a1Z09s5X+VVi9svgKXOmJJH0qj4REkYXUuvya0ZY/r/oVo8a5azUFLI/Mzbv8GggnuFNPm4H0LNc
1QaU2tBYnM2nc3GwAdWaFybp2k50hpFIBt61sQ3humnmuWXK6axLaaWZhLwwXfBbbM8xNZYkZAtZ
gE3F0FYlf+tS2Sl1cE+EgdQ61LiAha6L54g0CdcTLYn8ZFwDDQx7iiOIBN4MqxWEMqGlaIDo3dTD
HgUij6dTKvssGjgvXZjrwgSbV0Ug8Jmbhn7DEIe945LpQxmm4w1YmKGjwKKBGIEyMHlZYnoG6iKI
b/uLd+5G6cuOV8+7VQYEBAkKTQEJA9f5qdt7L4XDGGw69Ev6+ktZEzWYoKpvRHNRnYu2V0cVNnFV
wuwDWWfkqxJ6gLqlCpAJLinWfc2xPCCtEVuB0ZqBVpjZE+NZqBM41IgC8v4X9KvkhH17NeNSJRx4
wYunl/5GgNLgztruJYe+B/sbJgQ0p7o2jUJVLQT6Vr0ZxvNtiOHnHjAXzwKsz6pMdukqXa0kdZIq
scJ/Yz4cpBbZveOrl2zEz6adoFniM6JDihemHAblxw3aZSrTyeg7ZP+xrgw5pTh2s19AqYIT8XBq
g9H3i81iyJ+x07U/eXi12RJty98QG1xTHzZw9AgHtAgVUU8fZoGXDk7bxsZG2/t7Iv9kujChU35/
qB7FbfRJUMTKFgsA/93tK425qhFxlfcWL7NPisNS2Ck9v5tdEhL+mdJFJmSN+XeeeXbRiJCFazih
PfF+5IJ4udrodfRF8YnAgsYsXxF/InlrnC9ipG4g/GVa1F2UwT1PudxPQfhiXyTGYWm/nvsItGy9
k1TLlEzxPAhbpIgXBJFGZuInXK353TNh/szdY915mbZ4XquO+6W1zLlHTTptwLByzNQHHUwjFcJ0
W45Ik08hQZEWqlZFNO5xK9HHyz3Q1GAuok0NYseo58dUxuzv5suNVIX4icDvOcQKA29eKEoTppNS
+KFvEYKAL66Ey0WTyZmkLE6yHr0OYdq1AB4IAp7CNS3p7LW+5Q4wl0JQ1TRZTp2cqe0oBMyKgLel
fCAfP//ygPOeaKG4RlFqRzxVp7SY3jrrRm/XL4LqsMwBnvJPfGugomEMwnuB+1besPncdV/lIvDZ
Z9BBJiNvbd5/zSj6sR9CyxrXg03VNRXSVdR558fcRFe26WMSeGhugnguboOiS3o2FdF5gu+pBGCU
9q3BwOK0zvl9E0oBHFQq5uK41AitsFSF1CgT2KYlFZjJpCMn1CCozMsPi4YFetcGoUPS5YhPyt7b
9M9jw9ZfWySie3c/N1Llr92AY2UucHSPhn8bV4B34fkX6BZSkWTgEbIlM9POqgWftOxl1O0pbnXk
rbELQKi3RCSX4IrC4Dzl1/jPB0ewO56lo05Ai/b4ze8px3IkB0d3wdfS8TZz/xsXhqmjKp4e2NLP
nduADU+HTrlWEqOCDf0KJOnYGJibhJyCUBtsWN5Ad55ooOk/w0XbRK5soLzrXuRnGJ9ExaMrNzNg
IuTLXe6zYa0EmIWo41Kw5dnCeG2UMCSj8pgC+ysy5guK8wgO8zJcuptNinBxoVNmA8rBv9DbwOfa
NLUzT4IRt/PS3foZFEOXR8z/2mtBFr5rLDO4NyjrXXQzYIxerEJiE845IoZYuBZALmk6G3BdaFmo
PStybdbrG2j7TrqQzSCAVXAPqlAxa8q20C0DBjP29fFcivMeRcSyi+m3X1YdNLg/Egz/Q2G8L5Ku
+C1ZEmLTQrABQ8qWhI2mPZ8G6BtDjca8B2Ab87ONjG/czhXOuA4r8r3Odt5cu8WbFdvnkpxXtLC6
ZaqC4Q5Q/axZ3+CQKymwPVyLN3CEqTuZLHTlPwuTlK3fFpqoYxvgJe4oHh9UHfwzu+IVr9KNUxI2
PmCQWlQT68RTC5ETK8b5/N7+FB2cZIhJmg424nWTx7bWYfY+PAMpuaI/QPdnwFldbOB3h6fACBL4
UBup0r3Dsn/GUYSyMj/9ccgckPKz3fHHgBdBrZW4I0k2fHU5WoeZZbIqmWNjG719OjhgAi3a0Cgg
JLxHLPVoiP6/D5ubHR6qS36LUcXgNJ0ICYT/roil9jKQXFZ29RCgNy8oDmP0bje488yhV3Li+vHu
rpLB1+CiXhVmv/a7IFpPUOSaOdwyn6o8OC68JD2KVDD1Cgjz65LvdigrNVvV3Bz3FVy0MwN+N+W8
GkVkAnG4N08s8sSr5i+G5wP1jnZB1qaiIJchvrjYPVu27kHs2KFtjvh6oPmtRC2r1yoK12TDxJRA
Y9iUVzSWYVcqp3ILFUZ0aKebXT+WVLUNY6th01qHCo5o/SJZ15x4d7dlq0Gssphs4f/xiyVG0XUh
R4PFLCb29afc4vpxr+LtczaqS8oS477iuWIKthLQ/8FNczjls0ufKlZzw77nnj7GRViZOgB80K6A
QxL4zGRRr+BIi5jMo1yKhdO7MavUGyevD+oMxm0a3YQQ39iVKIFoHnVTHk/mFpjZGddzbLzet1RF
RY1H8De5tUifR2Paxwqpv6G98Iyb/wUEhyaUg5e9m1q8BboS/ZyvdF+y/y1jQEx0OCezBqxdvFoP
LTi3JnBqjgPHcVkjiCFIp85fUTA1Wy5fqXt7muM4JbxeGITC/NqwO914laY8Afu7EhCKJXZTvGOr
LQ/CH5HuJjbd2cQGCHdy6A5s6HVBqGzgd6AoeMs6lgI5wvwTzfC+TXiqHZh722adPH8HcPPrAtXp
oyzYEV4RXU8H6griIfMXjoPf2rWnCNZ2vU42NiTRIQt7sMXnaIFD484Pe623UowbBuR8e/BLDiVt
LYSUt7DPlVC7tr1YWgKY5InGcGNZeUNvSLI+tM1adc0WCw3Pw2wjKyxFsukYPiwhTwKuiZEExJwV
cLWzzJJK8t6Scl71dBazJcshzFBTSYjpecWqmknb1xZq852kyABG4aq040cvtymLrL3UuOB/EKgk
rLyHiZBqJ9JkH4Ddda/ENuLL0Ap/lrdeh8I2T3URVcbrgAox4s3ijsH+aa+S4xHv9gr8YPYe/gw2
JfSW7oGv3AyBlsAxKoE+5gLMvUsVGNO2xa2v/KiGDDmbeK0/k6cTgA9cEiirRhJyMHSAQKECnKLP
+YC6vvhwSTaI7xYogzC87UHLGsDvlM0AhAigYOCSWwhaBk9x+NwrJARNi8J18Vq5Y2VOBQHBEbS2
oNYnfmFBZOh/HQ7Sb1Qwl9GGCGIpxipDCol80sKCkYXbW++CWpIx+QJwXaaKl/9vQhQZMk7V2tsy
H7OgJSTVKibCDrGwLWZ6WkgZ92ynHIIx/bMxVebVlmCGm50pcsPaxp9fNYWFm4NC9J+FBCbawjXM
HFNbF3aMvFudGmSp8FKepWrHgoWAUD48zQfvtzvHI4UqbfRB7vVqABGn3XdRRIlcv/p4e01o/kbM
G68/JnVKZhMkGqVWH6TR+0+CaTMJn3Zpc7eHja3o9NDcjX57z00pfmZU84S5h9yG/K/vmoebqTG0
ZGIWa6/S3XZOfP3ErLHcxSinRB6WGaKBe9klb4pFHyYPmWyj02h4e91BfGKrccXMKCopU8R471Wu
wx+qqdD3ea9EACFZSoAEgtWqt/6Rpt6w6O2snI2rJdPTJie/TiGhQ2WHwHsPsb80pH4glrep6BVF
uC3co/Ce+5qhMLgZVFfEUJSsMlxE8XonaSYEnQGKn+bo89oOClQk2Jdd9z4kA0VN20M8TzHtgBGk
iRaXH8n3C/2v728zrM8r0rBBO3ZHji9HhrGw5kp09WNvuHlRlSW7rvszwrUlelT+uoLNOh4phF3W
esBk0QgjZEejEO/wqAU86uBXxZgXX46fWsW+UKph4uDQnynl7J1oNYKj26I0iOLDmGQWg6SMBqY/
LOKj7EgViJR6pzktigSmOgukdfkwilgzCipo+5uJZQGr27coDT7WJqt1/OWmoDMJMYwoxGXKynge
krgFqruQUlKg1kTihwwNrS+UbvcDOslPm6IkAogIfX2M28Pla+AD/exKg8RDeyKuwWS0bwnRWI5B
+OBdpMxdtmBfAzTZ/z+9E8lCwrUYIwvFHfRWECzUvAp/GEv8ot5Xg6li7I9ijGzm4kfJMuHyUTJ7
TVOIq7D7hHPFZqX4Ejp6QP/PSc7blhiEuXLXEWI/5gIlLp6z650hHxX76atxPnfXEI8h/gEN0XZR
9sU1x0TlWyX14kHXEy2yGFI7MfWShCcj/kS99tgUZyNd702Xai6XpHKqGK++O7K5GkvakbdEyc6g
Gt+85GE3OsZwYBbOF0LYlY6mANn9mg8IhOFJn1xOd8cdtO1v1UYVsyhEwZnu/TV1Le6wCFNqDm2h
mmmcB8nDx6OAWXxuoteJTZezsXtvzQbBSBkKMF+b249kzV95maBXJ2zoAVxRg25Xbq3vtOQigvu5
dtuAnMImBzCfefDb9R0j6qJBw/lVDaYgR/gNY10pllEcyy00YYFO1t625nIswNRI0qG14xaEfLae
MIBWdaG8gKZnlsXYrFee7GmjG7reKSCb12OOVZ2+7NOhRG6wLAjwPRGHVc20ks5tmoxfLoAvOyA7
UNu2un3sGV1zqCeHGGdjLVa5dQozuXEZViMTpEh0bL6MiuonE/jBlWnrIN5NWcVi9A4fXsyYtFrP
IdqzrrY6xVgNvslD2ah3conTWIF3i7CWqyhZi6eypChh75zZExtnrNVRqHLmvTHW9bRmPg5+vT/q
Q4pnYDWiyFeySUqU/uJ7VC1RhX865w9qkC2nLmdPm0lBAkfhUXJzLm26Rc+0kBPhR7GQaJxuvQBu
nfFLXy5kFTOpHuvrvOTyKs2K19PbpWDoQPXhCULNfq155YkMAL+uZZqnlNvYMOxUQ6XmTiaoVJ4C
/HfhkObQb5Iyk+mVDLN47vnbaL5E+I787YU9RKOhAWrxtdNR6D7qWt1Zvx/CKn9ihk9MWFqk3WDh
+pZGRaljdVKMVCoUDMME9kaWOjxsAQXhtce+f8OCne24Y8dQ8GeFBeKrvWB7bV0STokC945KDXLb
UClUQG3MlTaROM9KclLfqIBoaSlfbWAGhu3VfN7T5QqWqTTrjatv3ogVNCGKu5rIPQ7GXkIEADOO
3sk0jQt3ueJbE88IuvyBGhVQKjCuB3WVHwfC9vt+1DH7qVuQoo0znRsp1gw2FfgpTvAjFZuXTfKH
fXYrUbLf1e0EpteDAdFbyEzbo0WSxsN8jIp1pZL2ohZwaKi9+oy4rFtOl2hORztg4Psio6g3cKDQ
kkcaEni0y/kVnsIyu6dnOnB7PwWeFHcxGolsoydT0SXK9vh6ye4AfOylC8IAzcsUTL0iZ2Svuo7x
k63I4vuwXbq/T0fWOS+ShDBZtLfLRYnNIrBz8QD8Zu1FJEl4HhmoXBMXCe6SWhoMX9ScmS41ETqK
TKKki2JfH7XB9vUpwh4TLf1n+I6BBRTBnkWfYWJV265OZQ4R1T4Hup5cOQ3uODNKo188IWE/z9W0
91TM13JUVw30VMaq5wHi8iIlx5UtU0zBjY24J8fDgT7To5fTIxHGVrmFioGlk9dJ7y5AL06U6kN3
UfUQjLRflqA+JW49hT9Fd/yDu8edIgylTnE0q0Klx37VTWRaa2caVmK/xc8VI3vfa1TdTkHy0K+q
v8sBpghISJcB5roKU+3hViw4y7QWgL+YxUmKJHQjLeP5MiTrGdTzp4MQmZeZ9lakbkps35q4gcZK
v+/29mOdTvCI5eZ45QSQu2/IY4Tk4TyFRSIUimYuTuVLRT8MiQUT8L9lep/l7154AY507kWj5aw7
WQM/GRf/ngrO0Wt6QuN4tD9ho39Jp950m2ePlGjwxPTDMRLLFwKhfteIawspXq5WY+wMkcmE1sGZ
23INnmArDrUAfe/uwLn39SLxFatsSyHNSlFzaJQ4r4J9f5GJ4sx9nUdXYmNnxIjGPaGyYoys8TQ/
hW3asaMekpok8uWuCTr1FTqD/167yU9zibtFfvFuEwMPLyd/2a+3u1ts32qE6WAKlQ/a2HhbjHrT
+ZbpoJfFS4YeimzjKIapV3/wMSbP0OuCHZXuf7TRxIbLOhNJwLTvM+OWN+Z5we80mmpfbKyFE/JK
eK4i0wiuoN/w1JA+E0sGmh54zaDQRgb2J2W5a05HfOcY/wbQfzoeO8aT+vFIjVfiVGi0yfhnktY2
VGpjbWkjOr1mQVdoqwF6xTo76Z0u49o6+uc7Hsg/XtHf/OMaacWwoCPETv+S6iZTGPGySRllJUFn
AT64Runhww+LiC19HtkY5qTX9FW2mVRnkNHyuZO/rVmvKhk40H4I01ox5QFUK8bKJI1VuZ7bavuA
smFje8doSe4YwuQmSl+TWELGfFiR6r3e00zbkgQ1EyA9rDIITEYXRY7qp1oAjagWHsXYu8Bc2kX8
D+cjMjoss1+mvuViYIHrmyjZ4Z5vMjoMsQi4ClquPMIc6aReW+0swzU/c/jborxcyS88qNnVmdy/
dFiOjLVFgA4RkpbzyRZQV8Y+79YNOKBjxQMdcvDLIB7OUVv5g2Uxif6givUwyBeOa/cWLna7x3DK
1ILb2RthkkokCb4OlLvTeu5JTdSC38bd8MJVQa49Inc6B/mLVV8B5HUQBq5tOQkMuTJpruxzE8gs
hY4jhcdaiER1bC8ErUR0jcuMH2IeMzomMcDHrUMScPPYFIdJfDdK1FuRe9d889nwXaeQj44OmR9R
qBNUCFaieofAvDZkjl6/VCEI3bg5KQbHoiRj1A4aLkWpkWNIMMjkJLWqrW5q8pJ/cItyhhNJYwC/
560OrJ0bMmwYIOMln0F2IMRKx74GgI03HuHsCTo9nQNpYNbOqBEyfdeNo5koQNXjnCcHCx8HR/Pu
1CqhszDBBwQH1jL4lmVy8g2RSDsje4Qx8h/bE2xjCMFzesh9scgZjqV94vRNAA2Ithlqf3iQhxEB
Pie0D67Ut2xcbPVWd+pGh6H3fj5MUuzS8gMpmVMLKchxeP1PeSeESwP+TL9GOzVRfwOefbiMRl65
XeDwmVWZ/siYQExaeer5ewWIdCsOlap5/n3GObZ7BiFLzhwmAsCxXjLjwtIOhbfBHj2Ma4YY2fem
6sABxE/TxSUQNchHsYu3/Q7os3IXT8OUwU/izhHAsfwxuJmYqQSVAb5HyB0giHGWCZuDEvcdUVeL
g4VOV9iAYFDN+DlApZTkL/hldtr0mv9skZiHIKD7VscTeEW7mY5uJ9lGkMzGsJjGjDydzVJx1yxJ
dhVOZP4se//A7RimPFg1R1QV52ljP/hB2E/qZOMefemasNjR1cbIdrpttQwT/zzEgj05x/vCISjQ
ZF8+tdZqnPCc6Q0dxVA8NSA/65eh6SG1lN7AU0sazjz4PWc3oCcG6hFYPMdf1P8Izccm7jm8unFa
u2noegwp2QYsulGhdm3Cnq+tPSN6jnDb0ke7SZXvHZMONb22AlYMZXgAnBfX3uYvCUoj6yGdg0MI
bfgccnGDPJQdgpwLjQz8MhhAWeMOoBcnsyii6I9XJqm2Q2lhYPd3wiV0cTJ1ZPWI4VYc2KJJDt3C
9oIJTW0wt+mSRVcbZ6ELh/gdJCnzCwC4EgaYZcKhurmOLyTVX8IE+PZwaCi4rfgXZKChKoMn2DyF
O+fLnOMIR2PUdYteAbzNQIFBLHkDN7wgWIdUwrgcM0XDl0p4uvlK7JrnAxuUjDZLChmZ12XfOPkh
N9zpASgWYDfvKYOF7Y2DybcFEeyMXU5Q0RZUFGlk//ySr9ho0GMYhnYo2RErAgZcC4h4bx6tsdfY
29UbSz5TWeaXD8qf/wQaPCGtDPFDmryGnmBg7oefb8TISU6jddemkziTWkP67GAFHptBIJt1P1XT
XwMXhe8wSXP6paSMXOzYtqHywHXWofxhF7KbB1NUeMjRqx1AL6k++G0p/2zOYZqtW3FLqGh6qw3Y
KKobUkHP9O++eQVQmEjJgVHzXhPYHR9cjmt/O2/dvgKFQXub4hJdOo0uKgaSlZTgo8SnFcYBVoMK
+VlDPXPWe36avxlj254bdlReOZtuFIomPElY2gar0DLNsn/yqj88w4hrs0rUrFmKu5uZzXgGTAF1
huT7vl5kY87UHZ5uGD+cgGjJu3gmx2kafpeSPsU9Plo/5kxLO08GKDBPtzw2cQXczGpU5o9X0dT6
7oN4TE6OxCyZoGgUH5PkmkgMrIaT6mZ+ul0aLJwemoYB4nO/jLcAHPGWe53CpmhrwhmLQHMgfwfT
VMaQrSIkYU0UrbnWeryaGDOy3DlKJTCdiwW90pD81gAsy3kd9YDshRbyyu4Q0UkigPyjDAWfFBzL
K/fnLGUY4Xb3rzKIpOBWFTuTj1mYfeyaKOt9VOaJs/YTQMZGK85JqedK8VVI8O7ChVd9QaYe81GM
G+lxH++HrvNtLkP8eBQ5wW8UAQ7H9hoDJnsfvuWFPYRwhabGESqPmqCVCxrmJXk2lxE3PmilnyB5
W42xMbsVa/I7SYtmbKq+/RK+ps2/7ap32WzBr1zGJZovJWyc7nihVo/VXohPmJWNBWCI6H/8Y6aj
hxyLrZdW4mXxyDeBJRba3yY1G0gDFrheZ95xUkXb2Q0UEaKVGIEkp2M0Bt1MKDkFdUgOfqwViOx9
94x+1TapEAqBGSQ+qHMJZ+H96Jf7YqDnnX7R6KYEnokgs8zDYv0AtBjs5BR4kfkRh0i+ibQgcD57
oDyhAwdeOJk+uPimdYHhCTnMfi2iI6de4lnc7I54Ae64Nia7Kc17D8nr+gsWyPNSffOviXRITdZw
sz8yy0nTZk34N8NqmvMzI/WHG8aUwctdGPoiXHBcGPKMQ8llEmbi193sVq5IJgIgBVKoxr6luTgN
u9hnQVNhCYYPPdLImaaxfPcgjDYbyaECiYxiQYamg8WqqvJPPR1AoZB7+rXoPMRZ6O8uuYyKvsJk
Ei3TXXxdrRMvr8SJ7gbbOH5AUXhM4byLmwUl/7vVe5l4Q/z9oowEE79q2Ox9APz6z3XscLbhcQAu
VLiG6s8XNAHfUxFrVoE66Rzb+wdTwmQYOFJCS1ALTTXZmi19zWFU3gu+7bgoGsO/uzWzGa2ryUHG
hMMC/xl3AHqdpULxAtUKnKURAoqsW+WMvrcGnGhElSHY/4FxQbHdjSkSJWUNvjJdZo8dH3d3IuyN
QateS2U4q3s/WWxYhi/0KG4wFQ/yoJKV7Qp/Gb5qj8DCHrPOd+N4i7ozKtYIzHK2vcZxnkajIU6t
gObFux2tarXxAamq0OYZrXu94BxKIlbPscWcWwR7fuP04bKTzEZmWVMx9mHHXXAPJtX2o+3uc/3T
CWBAKi4vmsFIfMwPqmXRq7eLw1geFUZN0qV4j286gLJS+IytuR8sMIV2J3cGOA+kN2AcoeVJpZOI
R+N8fF1ql0Ow63+QFOj55qg3wFVGVBFTy/6p+/kKzZYB1RtBGoFQzy34NeE0rqzCG/FZ1fMGP4Yw
IdMy8jpeq/QkY24QesggpwoX+TYWudYguGZ+VhVuZcQ7rrqahid/6XncPoN6YXflcSqQftI9PQQE
zdhtVu+zNYnIwmKRSgGLVJwDy7y8F6k7AsIR6zYRvXdqanInh6goSkIte+9fmMXu8pde3vjoxQl8
6MiOD0SOIQXdz9EsUNYT+W8Ga3t5dZrZ2uI5T6O6wvuzjiy+Nh7wG6vPqbeaLWBCO0vJ8vVP7UoD
SMOzoe3PWCwdiowrlB+JRif6ZJWhQF3E3OGcpwcZ8cdVyGYESHvqWXOVEK9p0t0gvBE66mki2RMW
fXUF5u8zTFmYK/t2ihIOjhxW2rj46tl0I5BNAdx/I4aTN1PiTBPOVGL7+nZbK2S01cwei+x4ZREd
KqBnbkmPUh2h8f9iGscyA/9LW68Z4wJC+ILpp+N5+c8XqVu03NxPbIrWtWT/0syBVt3ke6gqRaRs
1RL44mnfYuLFen/KadgVz4gs/93jVHS7RHH9DOXSZsRBmkJJEqt405v6rWirrA0sqEC9A7xnF9dV
Fme7MCRk7nQdqqP6b/q3MRGVnBNC2b3ji03n1MjshYNG2XwYM5TULOmfOYy2G6mKXGe0p65UxKwI
NxNCYDL4tM56MD/K/7e2jDi47rNCrjENE7fzXnWb0/6aEDg0HhGPsEfoRSTBkfC0sgpqrNbL9sVG
VyEXhBnpX8842pps4TgWB8lUFdNMIq3kxvAfIFwVIsAF8Yq4QODdyGjnpzA5X9+RvZEtk7a12XtW
DWHb6SutJe6vnTnmHGghw9kK5ywNE3QetDjtYGG6lX+5RjH8tZToagzBRXuywJZjip9DK5hOmxPm
/+fjOVWfdgU6EOf9tGn2mwCJo839Hh9qF8WUCwIrcIRbS3l9VtACVlndPXYGlk7gNoXjeZ1D8/35
4+ZPRShfpngj9BMAlNVKDBLIUsM3PiCFOFClo0+SfZB2c2y2IF/7GUBJDA3zgrUqFwCUO3hGdaXV
JmlyvEMdbucROtdDufpVDrw1vJleGrR4QP3HtDrsskGPnhGaH7ismHdx8nid9PCQ8lotSIf8SxTg
K8cfDYQ45cFvoIDECTlsfj0h/8wxLkXP1kvO8a4DS5/xBVQzPmvEnulgnjK8PHXhTVr3YbXjCujw
HN+DZwf4VKBuerAmga0E5p1hm8oJYdv3E5lXTtNDnGV1GsuHLUHxcLGRLz/+c7zp6fIwAv59s/qS
Ef4B4L9WnVr45ibPOY9M0OVYXiXcQFmDdi/q6sCVjtk9kfL6ki9KqhB+Zd+Spr366NjWKhQTy5Dj
btecqW/m+shpgZV8uAQFZLA9x3eGSJM9AeKGaJi9otmioGELwpSXRFBWjSf+7xJOqV3QF95cbdVN
lKslwS0liVhifpCjpn3JB/S9hN22elsEDJRcY9x8fcntn/y6SzXlj9Gw9c+JNo+7jwryjQE6X7MQ
k5bkWV9kQVY6D9Erkkk4Fff/2bEPLScxvyoMV+3KUB+2S8jlInCzv5bliBb+lSOPKFF+MnlBRTnE
wff/EYD8Jy39IPmcOxJ8z3pGS5cHaSQvhD1W96kdolzgRRozY8dVWeVsEPSnJ4mncLpJ+amv9XSh
k4nBUeCItKGW37XOMhYmL9iDuRENs5/itHrfMRs1oEIYdf0fO4I/vd2ZuWB1c0VZ2xyYySmwTzrp
4dMUOPGerS9ERPQfVX6KgcavbYYXlABVHJaABBQSxOa9XIiMLq0F2Ro8DXwldD7V3Ztg00185QJX
LrNzCALs+SDDwH/yc1vpGo2QOOMNYGggYbLbj7A6dJvO3V5WgvIaJtTWfFhZObc9pHxgztG5MN/F
r8d5ybEJHx3YoSNPZeljCUzYPZnEgKsvAvAsIDDsQUkM5UkhfgmNs3y0X5J6+DCFxBbvJqtDpaqE
tx+2DfmUE9qrI/wz73erivXA06vZcvejPidE4lnxGKQheio5ftFMjiJbfEhEwEl7GUnjDjQoA7Kz
TLg9Kr/qukKkv/rwFeJbHYOInke6RjS9B45AzaXLnovAKF/zZq/u12hGeEyxLw96nLzyNThDQJeJ
071rj2bT8SKslDQrFU5oqSvvpmobSh+I+6LioXypBC8QCde2wCMsASSOmtCLZn19d+bjzuz83xvc
EgnrzpS7wNzEJ1kr8pN+ZqAYt2c6xbaqxoj/viEK8/xUJm11xhk9erlK3HrcgGKZf2PcAX15wKiB
sih+osls8reZYYSle7h11BILldebFgYoi+8z4lKKP80RblnGVe7v0QG6Sh9w66jbybRlditf8K4L
oCVnHDkEa2ccNTxen7bHBp/12nR3LBwOU9Tqnmuc81UHu+UBd5yVuWr7fTc6n/FAUj5IR2Eo+pUc
OnuyTVm2x3VfKhtRRTBEdrZhgD2GZ7KRKCGCm52Bwa/C+QZUsrB1Hm7Qqj4/UBKLDblHQ4PAOzQy
JVjfZl1xqwzYhALgQc5dy7dV9pBe/njyyNXxr4V9UC6e/LGFXm2n7DsVtiSbLDKmhLKYb4oT3blW
9jjjwhI7pwBle57gF5aMvC4hz0zZ2V4t/oq+1moeDdCFb+cqCqXVGF5Y2FBYZ5mM7aFFQj+oOjJA
rW6nQva1kxk17aJWizrRZTxONstB1zVhemi5SwYpVEqw8F2Nb9Gfk3cDTBMMXNiNUBNXbXh7wUTq
xKekmYQoS54GVWbbwktki642TkQaLDkpK8SGkJRDgKXVjcy38FozQQ31J47w2AILFc4KJrkSFmqu
r4MSXZI8knlR0v3Rf0otnIjCcePfC4lR40W1PMHSuFQQrAvnNqZHW9sEZVnWhGHAAtfCp12bWFSQ
PvckWBhmOMjJHIeKpPtVBV9Z7iKthlcYBRH+bx0GcJXcg3UWOmfuq+05KaF5AtGQucrtUSq8MP2e
vcVjK3hikKT7d8vHQh1c72s2LfDZGQ7Yv7S8NdOB46/FbBp6OPWRFhi3C6V+6Yt/IEEMf237mwLi
26q/9ABCwboGOHxU1c/Du3+nOZn/gALrZzAdhU9hX5Gypg7b/GcB2jTE03cDEhdIs1XONDkNf6m8
XzO/lULAO7O0jDiXu0NAoluKoXb7OIjjwlB+EoOsxYnKDsTUH0xFmYTccMQ9KZmvTE3k0uMgvJjJ
IAy7jlwz/0SpWXKo2Pkr7dnHB41wBBPQUOyoM9B251w4YrE4GNwrq1oZjZVaBMQFcyEa3j6XVIhL
kJJBRunIu7QuJHQ39zZRUqwMHKgI8weIKNLjnMiJJZjZYOK+D17veD/riFzvdzL2PjhzgeChnmCk
HkGoPo6thL4VA/rFemkPJdm+fX2opa5r6WhpxHMMcoL0tN8XvY11ZnXpg0WeFrHhPQ84GfXvhVWS
D1w+sS7eA/JVKl+2cIA2zRe3zGkn8T6sO6mhWfm2GfR1t0HqLyKohww/WpgyPBV2Qj5RJcb1rIx4
8/TGs83SUbtYfZAltL6njJ+VnWSwOEPDlHLp0ZOn9IX0K7Q9BnGzeJtT6ulImPfDZVUm+iNhVEgT
plKCuUWIz2piVt6gIwjF6J/eJUjH1cfvpH0r5c7KU4wW06QaLIfa/Rbr2qa0jXaYK3Bs3HOYh673
XJI00ZEohY0AxW4txEHUo0gMXhi8GhfUKdxkOQIVzR33CiN5PJ5Ac+sFJl3DWSLkZP9cObWEwr7a
JvQmIoKk5jCWbRb9Q6SaAhLdC3my5GB2oMkKF/pvHgWX33WiZXrr974pi+FgnJsf1toG3bH1lVje
VKTpTFw4gln49q6Mk0gTQAlQZtldqaTL1oyn0qL61lloMgabWYwLRLohb8wmbDoP3uA7vjJuQUXD
9jy9hQPaVkSdABO2FSIo3vESSyy01ykddN8Xv4p5Y3VEfT6O8P2JZ7Fk5qMLZAPDIOsK/74N5L5E
Kpr3zHkSmKSGYXI4/NFQWyHlVA8jnDu356biVXE8WsKRG/Jvr96Qdm9zXedjiM7f//ZaEH8rSrlL
C36i7upV1SIlikdx+nYRWhPs19G0RldfKHrAGXEocGxEu31XyMeO5/Mg6lFsBkuUZNEgW/RoyGA2
d0Xk0DtSI7/AEyvEChl91TDIQUOHYBM/vAzIo2x6WDp/0kuxPwTNMkZDfFe0u0LzeYcqy3MrerFW
J/GT+UrBlXyceXvATTHtpYJVfZSCXH/2GVS9osL2B27i5Uypwk9g5rI2PyXe4P80jXk8N+O8fe29
I7UtnrkwI+YrNgnibWO3tGp6bkhPQIJKypC3KpppklUiKUKSoOAO16PzOBbj4J05P0J+8EHoUtrN
5g2pYQDKCUQDGWOK9AQSeJYsXsDc1jmfUYnSeiGcR5e26Jfxf2fotQckipasYfwBYndE+qy20/G+
wMdFkxHBXph/1NY3CG69HiNWDhv30Q4Xvt/TKkGD7Y8k4fD5QNJz4lUUrDVCd9/e1jpxzHXcatfF
gXO83/XIvytDOSSpsmxrys/sjaSsxgb2w+skVPJf7kMEX2rP3bBp1a85LAOvmr7FTcko8jtJ80Gs
aU3NFOHv9bq9UuVezhj0lG0daMluH/PtVTEms/CXJmQCwomaEtNZ8GKXqJNxANmUmP1TXjo24B00
P+usapLuSckbaKVwo6N8304ozRY13gCOvFCOKwW88VGrYniTpjBbECVzEZdCjxI16W/59tEOibM/
nrRTSdzoNcqBTV+Wkp8hYx9Aborn2HX3yeqvIopi/7i5KW2gMYH6Jf28wAJd2A9CEKbalh+s+tWY
hnUxhUEaZlNlqS6Yh7AXcaI9LMIeUQyCXgMbm39OjGDmwoyQlg3hFCjBGPoUZL84Dtzn9jIm5Qsw
ALdm9yyxZv1MOk8u10QmpmwQcpywOo6Jhqzlb73wG5bEYjEP6Do13XxHsPbQ62w6Bvczj+pKkeOg
fr7zd4kIy4u0AOgU8+D/6RrsuJ1OfVWenkG/aa7JVil++mfqmNHzye9b6Yw8F039yCpbkhAmIcVm
GNtPpIjjjjwGMqQ/k4PH1Fd/KuN82DXNGPARlImlsPYMkXcfCuDBQGIbsuPYCxFhJea4bgTNzXcK
3xrckQ6MtAwPtwUNjJkhpz/xntpT6fSjh8gLHnqewnWglx38Somfhb878J/xZLh5bL2sPsjohcTI
lRXD4aVOyLvNQI0SPnA/bFE3u+c41zkZqKQYP2piXMK0jlIehVqIQtfvhzDgHjwOJbqWVc9Mv2lG
Ga0gc4TjQaxVWViexzwsEiXIsm6zWhfe20wDyFav98k7Rk2fNctc2XBwhHkn6f8VVHZbD/B4Xq64
r6FNXK0u2khmghU2JR/nh/fCQGCHXvODdstkIYgRU7/HJDy5GZV1fNrP6pvyB88HqvHibyAfYxhG
VWbT4c+toZ854CQ2tS2vv23BAmtu9KK00X4qx82w1Uf8YgSm1VmFapaZh9MHWevQVdcl4M73f/CM
cU/1Pdhpyw5ikHwDIJ5NoTP3YLsOZ3OuVdbh2ywDH7k8z1624Vr+f4Y71OBkkRkEA7jjoG9gTd4B
p1BwJ93OSVH78h39Tt/ggFgJKqPuwwj5hlM2b3uLVCtcd1zRfe2Y4tNUU7Xoq14gNS2E8fhm4SAq
6j4iSYLq2tkLB7kbaxdvmTtAr31Kw1c8g/nV9uXG475Kblpm4DpBnJaxAyZO7ze+79WIfs9vm09G
s4mBZYT+YpBdn17qeyZbLVmVr2p2dKL9T40iyh7ibN/ORjhq6Q+jGgB1g3O/4QZGKwprPbx/YSNu
pl53lsWAUwo2FQm9WxCVI5LZ82nTnjaK6Sh/GgyoyuimCsP/FIogywaaApmdEv5x7KI36x4+ySj7
92n51LBQVzobO9u1/7FqUNVssQm4Lo/QjwqenINcoWkjpq+MpNrhkebN5WF9fAj0Cy+BgLAs7YC4
BmIfr7AtieT8gMJ0DUcii6UdMLlRYrKrSe0VlBpsVCyMFeUCm0aCBdrI0wuGcHWRnEjwV9DkpWQw
+RNBKYar0KAiT+HuaaOcWL/jO8tI8oHsOhDgAn/N5abY/lA05i7TJ+VOYCGMEPVmDSdMp3FBRY9D
+qQQBpfYEMEzWz4iqp7Itw1Oa4UDS6ozPu32LtEMfAG0kKFhLbQ24NXTqKOABxZtQNq76zkRmE0w
QDHXphfQaXw1a8rnBzrg++hCzsVh5v8X8CglBx7FqH7CxNyz4tl0WFStI/Vym9Ufir6Sx4rZkD7y
wr2PRwYxMBcLQEfM/K3GLgQ/Z0Tqpi79iuMFW0z+TvH3fBeLDavwInwBFvnmz7CFukXZjMu225aC
jlqYSjkLwKAygnJSlhN6pPk/6kICuZ6ZgE+8f1PJxkKoUavEVHfyKgvvKjBzqKJaP9JRYs7eH36Y
us5ZoIGOcJ/BpWaRdqiGXCCIMXRnZ56SB/iFhBsvrJUVTKHg0F9UczxXrpcn2WNtlYNtCDVeBgu+
jkj+m2DaVjetkcCNRQY6kItVzOGOjLcJRhfwIlVy9EHARePOzINdEOVqZxLyopXPOJ3tI5L8KX/V
e2jTrcdUty8YS0lmFwqB8vVzZWI7fQ4TfZVtvKMeswAqAz3+D5b1S5ChilWWypDT0CM8paPslDFk
4dE7zRrj2gxRhuOOJujQaI6nGh6QHmo0aBiv6ogUz3hOI/IcxidNzkR4BTxsm65Y8JIifAcaMBCo
uVfG3L9mX95H1B9kV8Ko2qcvqCNH1HVg4pVJK3Aq2KU0kI8xUOhOzSvnls+CqIxQdPZ2ZK4t05yE
yCxezcsLodRdG/Yf/UTePTkstvnYPXpOYidSje1pYKHv0GHq44aC0zcMcnA3q5K6GRQLOxiHiGr/
BgmGo/8USZLTNorP2Opu6Y+u/Mw+6bwncMizuvCzMLG8QSsCI1jQkB0g2svyrsw1AQJO1xINj6BS
AzuYIqnDRKRF9Wc3wWq60OvJmSY5Y/YsxfuOx4oYZRJWi3a2x9axXeZABhmDqlTeUvKybCZORrG3
LB61JC2A5UmkdOrTxPr25UQf+TxBEDigJGNsrHA+I3S692lzDgmRfEq+KBLuVuAgFXaqxnqcyZXj
DF0iuQiH+Ol8S9tccgdE+g0ZoGyIODWiJRPdUbSQzmOKPmIbMI15twuNcVFZlNZY4xgb5kZdeOcO
40Z2JL69L4IrixE+zearKOq3KI03G3JvddNMKq8fCzhbChGP5sAs4zjQZglUtFTttvpZZ5BpI+uf
FVOz73QbF79zaLo1tLhS0j7+EKP3LTQtA/rdJJQs0MCplhr+bHEHEKdjy9gTduBF9SVN0z6MQwQ3
9MjIk+rEOdDMHNpZ/++iwTVShtMqOhQJT+N0KDaUnAjLiipwB0SRvEF2/AC6lrjVSsbDU0eFZYoO
eN63ZPU+tC5hPxqvi9DSRhMJhPVVQhJ2vcEo7rm8F+VRguTkDYfg6U4vlpVqHAB4naRMVl07WMQQ
7DRGjR62Cp6ctuFGIivZ1CESOAC2aTMca85kE9+l10ThoEacQTRcDVoLT6Yxi75JKyxQMhQhMJDG
QHV+vBIVral+2iqdPvQUqmbWmO/c2CARPtQMS4/xcC3ECWF5KMHBZBR/bl5LJrUdtf7qr2wMkPhh
hvZ4sPldw6sHsksPK/V5SEoefTqYcEOtGIdSmAzTLjJXzpZMk2xfSz4vyT0sm6kfyIDH0mpuC8vv
JWzNidxlOloRocPvNm+O1lT3r1CIe5vtitn5xFU4otJQAfCFkCDSPSX6bwBGVzsobHsk+wD8rQVX
yBIpzV3cxoomGmWV091lVNa/FxT0q1/3il2TrjHS/nyxQitlqerAhzcraLmPPaKLVOwykr5ZIZrG
sceSwjwpWNWIO0FK3BjGipZJ2HT9Fp+YXr7B2NIIwYbCTHxXvVdc7YHyYOvyXLrMp6FbPaIq91Up
MOpdAFMBL6x+luCRakgT4oebmIaMC/7v2e/OXgqN09J7QiYsogV0+RDvEyWRPOyCptZrCEzl3yk0
YCbpRKNwaFrqQfyKZW0hP/nDCH9yld6+BWcZFyO3+122OHYkXi4AicrlH62vURqZkzoJgILQvVzP
8TuMhTip6th49HtNNU2WmGVZOEKXvYcUAa3kFPOUJ+zywsHx0Z9L+X/6MLYpIEDOpnXLmxrcc4Vu
bQ4EGuYYwmLUt+/giT8vTkm9o8Kr1bi1Yihb1GL76SCavmsZzGbElxd5BEO23YCDzUpgLMMX2HB5
qoYkJH2+UsoNsSNRYgNgbPDYN7xxNQT9SoOzNSlZf1+wDTej1pYmVEHSqeRfKcWBCi+AN5QSpg2/
R1xGQvt6Iwvgx1aDnMkt4kU1peb1cAnr8nAZ1rFAN56kU095XjLIqqel+0GEG3DBRs1uJmeiy+MX
C1K7QN7LE3zRaZZWksnVVP95ykLwCI9vflXSAP0+r10Au3p5ReH6FEU3drfPI02puBZK1c3cLZp6
OP9EnsledwMOI65ZLyYI9VAtOyjv+3jfyiUWySnCOh0JUdIwMAIbIvRhjaAeRltE1BfgTJKsnnqG
k09WZ+LM79X7N0vXlICv0nQcixCCu0MdISdq50ZCIazEbxzy7OLOeMPDqgR8NFSnpqo7wrNvxkYy
gfnTmn/eJCXOmFpsQ6I/S1tLiYPAQNAAwcHCAGeJsb5oZUIx6w7yUsZKCK7cezKB7IEfTUMenwc8
zOsvJCLrx8KftSJciJTX3he61T0QC3x3jdcJy7abeYnBtV9SVtLeR/o2ubQKaTzgvd+UPoEZYs3o
bWlI1gTGZQ4S9w7/p7HJXSrotx5eO2cYTMlKdG+lDnA3ohZhBym3erWny+08067n8e3Oq6vTCcfZ
abhOo2HYnl3GPRpSZL/NGEpLzPc8/KIuK+cdBxBOOC9dR6OUOB6n2s4uPg9U9FcJ9OAyu8x24sZu
2GtMyeRS3LazX932zf4dD1oApeITFCyl2NiqZ2ZBOXLXmhNCu8V+XybVT67zORd2uMu45cv33PlL
6zan83929sBlVAJVDAsKgk+af4nY83+ojIT6iRhZK5383k/4aQC35SkAo5BYAFeCbPKS0vC0VqRr
FmgofSTaoOH0DotpcepmW4yz6RFZfsSq9PAOU7aAHBPLFnOcbRq039Eh+Ye+mcONak5dLPMoOFX5
Gj5SqkW2O/iJbefbluT9iI5xtzxssf86kMFtV/O8LrrS3yejDldofeza7wPpLNmE7sYZ1nZFbzyf
zCZboYLwJxE3DlIO01B9HpyzM8iog2yaeM8jyDJvt/4OcWbKZS+BooGM6cYM0+zG6OWN85626QDX
a92gkpOYTfm+aOv/ebgXVX8orIdUx9jaak/Bz/AOA3jwgFcEZPvAXV0y7u4Oh8mlKSXyz5l27zX+
3/3DSw/RqGM6gYn88/HjPyZ+9OV7gp881eDRlK2yvhSgeJNbzxcSGSklG5nIS9X3OL7R7ONgCcFE
YoHdusfMQ8SZ2AYkXnom4HtrqaEjXdle9KONqair+WYGiuLifIqMNZ3Qesjlb3jSbgPGln7ADFBe
BYvQ/R8Q1cDN7oLm2wq2VU+nVjrziMokRbS7zWQ+9Au/Ks72O0U71Oc6jtNqh6NfT9nlDDkJLOpq
xJakxcuJ7G43bbstmjFH+FPod3IyR/5fvVLkjIvh2Y2/VDysywNf4GVlxXj1JpM8kKMhxTDUZoP8
5xl7oBKB49yak4HwDQYbo836+ynJUirIfnYxs9bB4emlvnTIiCOnGE3eJZ8ZgH66rSd1nJaeSnav
Q20bjWAO3VPKcWd4kl3ciZCkqzDgvLahgr2WraubX/iox/IHYtRzZvKdmOAyRyDOrAS9VWX7wTxt
MknVzykvLUVrOC3HWFcW1obpsdUs7CL5FfSeneDCo/a0grpHD3YwIwjyhrcrhWChSORbZYQVstrL
MjptZEfCacJMWScnTmLh0KdMhd+BrUK4HtXHaqwoA7YHRodpgWOjevCVHP83sVnyoCDOWh/yu5ee
Ub2Ta3qhkwXVP2+CJKah2qTt/FvkXwpBGDH21QNj8eGjVF0g/54e0OrB1US6cbeifTHCjkpU2JcR
MPdggVHGg307v8HXumVcndvYi/7P8avmVn6uQZLqZEc3tPTn+p6Bp6T0bVDMO+Topy56eDMTgW5t
jKWmgQDWIanKFdRwtiKv25z3+Rb3J6QOhowY4A/k8JRVtrVL15Q0xECwKSOaLNJm6vh+0j09U0B6
OqqnPdOl15RuI898/zY0qxaM8mhEGaLDplxID4FhoJmN1EZfv4uirlhXqoVtaJx6s5S/+ItBdN+9
mUG7bNiiExSeIv0S/MsVYxoNUk5XFb95Fls6dl0M+Gf0ISxAfAbD77L4f7aAJ2KE9J0TWGsQr0xg
Wi568THXapST/EZGw0WtWgIiiDDSVawENNHdXYfL/7i1QfBuIhOVKIDHY0ZiM3OxHSLBMm1bpsb+
sKcwxYDTE8GPRGjwtD+lY3tZWpdyOE9z5p1pbeAQcwmeERK7R9maoCdDkS83J8g1ZPvvR1M3RNOC
+oxjXumh2LkXjw5Mu4lCKd5Cv4PLvUzJYSNb9K+t4lHwGvQXaf4Jd+XcBOyg5kKiRKXglKvsxTWx
9VWge24kX9Fw0ln9RQRc8NlimTVaGlMKVxe+6qywZlorTU+UTZPBuQ0GEiq3MzvKZB9uc9YPVu/9
z/IMA9hnK0KiDfae0gaAn2a39NcvhCoxfqNzy8jzgRrl2fZzPRfX+6rGG/RxmD0QzQ5bTBvrP2vg
0cFgm/WISoJzXpAfEdoIwnrPv/hZZgMKPbN9VStjElpLkvZPd9KP671ng0lyqyIKTUPsEa5dF5Q/
tftY8xjNAoybXzQEaprvwF38VV7o1w+mIjXLn52k9aaJ0bVWDvq8Nhe8PkkvzQlCWHl64e1HvFIi
I/Ero8I3taXjj5NUf9rp0SfU1aLmqd0T80aIN2RCcxsuU8NEpNfPCR7JsQ7g8nDGkFs7uyZYO2cu
LnDGhAjQ2cTG1xFujnfJh0dByBLQ9lgWEWIvj+VsTrfUftNK39KN1ad3RmOZxdwd/s5kzaIzOsTq
GmBj+uDRap1KGIyTMW9M8FnU9SniLXDP3i+iqt7wYksNxC3h+r1CVgOcreb6Xl4A0E7I+F26dhiK
jp0hP6VbHZGYVaizN4ieF1KfuxDWnW7ns4jDWV0oKNU1JhB7Jdgt6U3ahU6Ob6P1DmDG5xgNAFaE
P4SewQfiNySXGw+oxdidwHgnq4N+btkr5DnuHcj8WUSYsc7teXZ8mW27p8JvESvngY7aim/8Q+Ll
wYkdwutHrUC6og8xaVBsSbNug/h0lYJk212iCQwB13pb07AcGyusGfExRFnoiAN0J61EqIcYHbVM
hUuHP9cNV0/Skt7v3EsHZgICkte+RR4Ax7WD3oq0OdaoxUwhNnlSZ03KN8ptjEgtUu4rtu90pUlz
xmYcaxx8KjZ8PnU5r7g0ot+a0yTg+XuQ+Y96dPNAHfUpob6QEBEWHfKfc9+KgSviQJtw9kplDTl9
v6JAXrc772tJFhHK7uItBr+t6DuepANi9JtA5V3UBrWCy+Yl7ARLGtUl1CuiTtE5azxLS0jEuQqY
Y4PqlSUmsWhEyLfnl9JNVhRyn4vJgOEakCXJhmxnZkn3q7UYr4arij0krptBepmZ//QdR1+0Xyj5
kXeHrW6+WETWOHC0iQ7d7Bf35G+45KhwYZOyzAngyGjMGM5q2dhDUK849VH9Et8E9noXDAI5P9tB
d1y33TQLvgv5bhU2MQDGO6Q5RH7yIxx1fpFcASmHa7HdWXYkQOvni1TIC60/LULZJuZ/aXfm5EIY
Xh6CoBXpgvuh8oYI3jpxYbdq+LusW2yQBMTS+XnD08mWy10QN4HmUWCoX/6uoNwJQPPvEj8KtYiN
UcXk4itXk2AOxh5NjRat2odk2U7SYMlw3gJ712YYPRtQJ75+YWhXk1ltPRBXhUJ2WYGuuoBif18z
nysKWDG4mkzwz1Ndz/ypOGaR68XnnLlpU4P13hFfIK2sjolQCmD4bCFc4sjfJnevwA2uX+om7QYq
5fZSkoshRgpB9QypbD/74WQWxAS/I3gOSOZGiry+DtX660Cl4dGQ5+hjjBD6h8PBNMargrEVIf5N
AgH9TJrxyWmpgPfCHRthaw7//jrws2kimXO5KX38v74HWy+labRLxBtgTdHAnbDcswh4IgKVesHV
p9ZJuWd/RCnf0dfzwDito0P2dA+Yej4KiD20odyZT19b9PmyO00VA9iIv0WrGD4xtdq+uRVF7uKi
+MznTUuH5nG7v2i2kQxtuNBQ4TqEeykx0AVJq4/8M9g3RRssgPTVDpqkTDeIFBDx7LUpfFJFSe5w
Vxgn1ewQUHoMVRcalDXeF0jXV2yhgbATfNqpGvROR9zwCvuQkIqRoBUXpgbdLv98/vaoIQ+FCz7J
aVpQqUscj9ffQ9ntAmD3zBYPgvVTxmmsY3XMMFrvGSIdk1U0WF8c81AMxabGTor2LMxorDDgOOIq
cbQvYOX05MPxlO+28ofy43zukCVpJkIRT1iwm3Gt5QP/wIFAZY7qXiavLrneKxgpXH8e0IbckTHQ
hywh3zExzmLms+rdr5OOxog79PaiVfJov6RiM8xD9RRSTb97WBh+XriXZHX4zRMXRqmyRmtc2O5m
dUUuTC6ZKmCNamlEpnJYGjOdZSMaDdRU8LRvT9Wyuwj1hb+/N8dDJdHPRrxItOEENPc26pkQBDvb
pOlifUTHVmgdhF/3/m2Xbv5hbo4tb8xdmPkEp+dTyc0iF6tFVwk7YFEP8XeYwfbXhvGue8lOB6eo
nsrCPf4EMpWytI+DFJoqtRSxFdVvFVC0/6g7cVw5RkGPO74w+nHZ4xLIl2jK3g0Ftj+oBWSm4wA4
Myi969FdKvFAgw7+Ls+AXUm+Enl6X8aKMe7sN7yvCRRwbgltcd1oO7pDQv34rk1CcF+KAa5PNaaa
pmnZJCqEMwuVscB9vcNocnwo1v6W7tH8UIqXxk6Sbod9Z0W+7HmzljKpOz75f54+yBuzKOZS78W4
7aLv+NFNWJHZah7ssKMHHz6ioWPKGfH/49FUUQgIQAt+w3uBcTu0YNxXzyKwyHghqu6JFcLp+7Ga
eLO+Q0TNvvUQpDi/V/QO9r0626sOZsz45cJQBmHij9dSHPvmIDBfp2u36n64S22/WSgF2fsE3eoY
TsR7g3hTOE8FqBNylXk2dFIxvwi6PDL1dhybS/kuP7zNI2JVwHqworMXiu/A4VH047bBaN98Z1XJ
9/LWyqOfyGdPyqRfzYxCE82NU2WkZ0rMhjCnsWm6oe5upVShuwVyr82A+tr+KgaVe2aF8jWARHq3
8AAUZW03uTHBh2BGfZjxN+5Ae/xwelAvI8W21Zgr3TJLbEPzq3jGFT+0aXqobvfkBSGwMWxf5Q3J
zm51kzM7cpQaPtIla9/koZdikFnvGI3GCalzJ2mcjDv80OQD2ZmgAzSDYFk1+QEj1+1MKm1L2j5E
EHbjMMWI4lodCUFI0ZUFMt0vy8qVKy3ppEGbTzQJ4a+Jz9byKmD0MLwbpTJI2xwE3IcUe7q7PjJF
0qFJyNb1Dp59bEMJ/HHFKqgV1uPcB72nsdJCcfVE2qaTpGYWFnMGrIEe8IyjCXowXHRq7i7MljJl
l0V26IFhj031g5ZVJQ8MFc9LAs6AdPo6Z96H6kgvBxamkmmKhcxkg/lXdLIGF+Xd/8ga01esJEXt
yg/NXJFvaJPCXr5sOI0FQjGS1jsVgG42kFUDBKZBSUPrWTAOh5I1GmE/TS+nQTR4zhVPb04k6g4h
Ql9Rgcs+zLJtbMrg3bkHGZGEAodA6VTGTFKjUpn/ijrZ0p7vW9NlqP0TVm/u5YgpOL/QcETl9k/O
mBg01vf85ETDy1/XtqUEZwp7c3hqo/c4Wcw7XZZo6DJ9aBWwVtgj/Q5Z6veREDniYxiEusr2meTf
eSbr/yuy+fIpSx0T7oKNQYWZqVeyt/ScNN+iChGArOBb5j4rrDGaLAGbNbdKkrvQQ5Vm8jZlKUbe
YTtiYLoXjKA+pmVrS+DXxYZ1jbWTi8Xg+JE53N5WQozWix3JZMdBsw9D5s7wg3KUE3zFekcMdyTW
uBxqM2O2uwiFH1xci+VzcGGiuyKTl4OtDN+wk4YhoSV8feinxAHF0EH9IH4YyzjSw2x3/xZu71qh
ciq3VXbRkUlgbzwB1eS+HNiz7YS23gPaSZ3kb8fy7F/Eu8UWdTOqOwXFdnG4MaMSNAlV3tHJbtzk
WmO21i2d1DmAra62lzdErZG2FJBVi0cZqZ57R6erzVYHb5YpjLWVUVSC/tTuXJAArEBtCXQR3KG2
go4lAULsQmvzoOb7WHe0ppDT1Ntfp3c05BnBJWry/7qO+FJ+G5dEOsHMR10dVSLpsaST+LY6kKQs
de7KSwP1k/Lz2cudHQDM58J+KpqMYQLrEKlwbnHCZYSTjEjInAPkFDfWCP3OC7kQshyY4SvfFbEe
p7ELqOTOWJp5KeP4IE1E8UqDVleyC3qEY4QNvvlsJ2bbC1NL5MNNkxPSsrMfSXw/UIRQu3SLI646
yAtpnXcMUcfa/r9/+COJXVR3NcuSjgvuMbG7FaqnAo3TdVhQEkn7rduqrqis5Adc7PSdsF1xVsor
bN9DcLXkoNUO6iJIQ32z7tx/Jezk22xOGRmxyrnPdzYR1HtQy94MteMe2mEO5Rm5itS+TScc7oQ1
0mzNB7ExUHLlec6ImqcT2TkRFZeZQLs/K96sN4wJH61YHADRcspTkWDXmDLSGLhRpM5AAaLbeOWR
PEKrbG7DvRjaVVL7GCpjvxZtNUmPCkL4qwBSVykyg/8MsS55KTP/dMAGzH6+KtEJTzlX9MczPD1e
MzMMmIuDsLyZPL+sLyMYaUIeUFEuwhw8JhS57lDZRjQH1SR7HKTCTi4sEQerIH1bUxLnW19/8png
9Cx20iWz7cWkAOWTePTCg5E6tQFTPIVxNYjIZ1fQ6DqDHQz2VCMIiCx5dINfESgNSFG3l8oJKF4z
libyRr96u75teRHHEJi1fybXaAC13TFcTotExROEaEvTt+Zhspe9+cft4yfHYzmE75Jn0T45iUKD
ZJi70TI1h99cKMrNGni8NOmm/0u8jDj90ZzEDccTjm9R7IFxiH7MbnefLE+3vh9C1MJqnaXbFULe
sBVYo46IyuOaWJ05DzUIDo8lxZf1a3nVoq0/Gqik0sKWOvPZerqLdHm1UhrgdCSIJwPwPudFQHX+
60iz+gDQ7uP0pzIDYvJhLOK07+wU0mZGBDKNbJznvs504rtBIzlebdyc3MHm7v2dnlPAIVf4PBHW
hBH733lRcKrVO+6w7/cx1Ol8gTwrIfREDroweCZijF74N4ysdr00EGw6PND2y4vBlDQQ5HQbRpBx
c64ISC0vw3A7CclZBvPfuSjqBjUz0qt10tdXibzXnY0QB9aShEgV77CAhOhadsz9EWN77yawCH/j
c2RjrHLOG8Ieseyx48GhALLqoSOCVnUP+pzJYhDH9JqnSe2xdAgygfjRoozrrn2rpaSyvPdpuOTN
WWASM/mVo0bpRWzKVA1271gIb0H0zHrI81T5gLycDggEz8xJ/ES1bcz2PVfnAcOpcLsjlxvf9TEN
eO+Fd29XCfEdkFK4hJUPeDnSNQkCe2RO4C+jLFC9QBdMSDOhTeOPARcBPMahec233l+xRRgZekAg
qXuZkwOGy320xbf187LOwgMtaSyjrgVvEcCUvqIw+0+w9n+neK9f/5QXtLE6Rvqn4z9Ii7CgTBwU
VX63Vi204Yt6UjdMf9eY47BMWEcete7cueg/2Zb1O1qydMQdANGAG15ty87cXcvViC8q12G106Ox
tfB80MKkoV9UZv8J/n2o4l424U4Hda6UwqrOIBuJ7lgJW6ll/znGxsJ0+gCkyVnjVhYYAuYOtQMD
TnWs+ucqREoZGYXZXfdqot4ZYmzYHMWb8Ql0K5Yku02Xr5rHGfL3zB+4jQ9NEyOdywSUG+btZgc5
FS6ml2TjP0HrhQmpTCW/c6DKPI+R9sQVFuEO6vZaHICFae4OGnubyVFW1/nqQQBuUWhXVU7HsQUV
lKm73vyyHi3jnc0WP9dYINeL5Tyo6qwgex9zHhitoKOtDOy7OuMUBRwMjO0ExcJHl6QN4ZrkbUNc
tTRbFOJ/JmEIRDpq+TAwiB0HNZ85UizqP/vDcdQ2X3bCNo6D8e4vRrZ3xO0d6FH4Ozgzxs7ljx9V
rn5qJdACQbgu09AU4n2x3Q2Ncs2wV4ql9rdZUYKWrxYnGCwlgbNOK7xqflGisf9n++gUefJuk0Oh
ZnTHdRkr6CVp3//U6jVfIAPmmrIXVh/lHu36eypXfpi2jkj8ZPdCAvsM69Qpu9qQZWXDAjbDHss5
KJeeUJOfD+Z+INXLhPWY9LQo2bJC/XZju7oqLPHqjUjUbRCcmmnChDb0d3zgg3Dkg0Jk3aBB5Zhi
vq+W3O2YOtWvUGO/kR54Mv2JziHt9Jfr86/PvQHSSzz+i5UyB5yYh7Y0JvfzRiyh8Nk7nqTApM4K
NQSciChYm8b+2XnkotfUI9KmaVEJ87+y0diemNlkJiQi0umDmRI4RuYpIXKWlFRqDCDel8RDclSb
rwscxIo34OfVw9R4TvqH/qBJ85EOB8LfGP+z3sHx4BEhdWnwfLC8Ot0x4J5ZO0PdiLWRcVgrwurg
MuJGVIEajzXpkwSZvzrG8mItdbhXbWyXX9wh46g9K8UnwLVq7cpyvWpanosVN4HOzzCYnatU7r2v
w5kS2YbNR4c1AeNo8Rm3niAFEKu8q0GqTt5e7a+OzFqQH1hX4yqRLPrB4Ue4gpzJqY7XW+DC/omI
ClfwuyFPR3dZ58bZ5IZF3bH6ppM5JK1JPuRZuH5VuW+1NWklN8gEyGF+43kGXQQdJsEezlREPw2Y
WO8LcZ5VEkq8+LU2JJDmPe+ggtGRUgW7KEnyl5kCdv3FehdqG6Wh92zzR02hHele8iDvi9b5TG71
AJ8WDAz6xVJpMUnGiiWo7jHPaCmSwxec8C7MGlL7b4N16+4zVVgwDQSIquCUvdnrqaJ9Uah3BWE+
ESa/ll9yAHn3K04dHXZIP3tH/NS2/mL4KOSzkwn16LXb253CRUgJnFW1XoQgTbagw2jm1RoZmsUD
TAvCJIb6yKdMBBn8++uTfGigNbIeIpX7NbojpYHNGnvBhp/YexoHv0GNiGDAylEpu/VG4WUBBVGc
xeLEsca6r05Asj4eG5P9JIvN/D5nicBrOQmB0xiG6D/Vm/JFagcl0+L+RiRXaBI8UeiXosb6znNo
JF0iOaSA3Bl8OBKOft6JF+Mn38mhQLIXIZ2I71/OvyHiYrzAUzLncDU8D+nQfluXCAeFHmFSXIzE
3yzwSnUJM73WlXrpE4r8JWQ4ShlslUtsfPpNXaf7YLzOXvdHKHTftAHKuM2a0BoQn5/5IiH5R534
OvjnZIYC10r6GCKgZmvLRxyzPtUutcOhD7us3A1LjppT6jmdUWjk5JqPQio2r+yGwZyLdTO8avTv
6x29M3hAXZrm0RgWGwYyQOGg4rwoh+tYcTm1XcMW3z2FqWSdohDKC3QpGjFWKKsjCLUZdUGDXxiK
rvlbWZig7jML7TrzuQEMvvG9GLZ7cvLgkKpMuolbPl98VpftMY7hxadu/jOXHPZ+ZE8Y370phBLw
+H28Ukeql4QT517gkTdNlUE8rdmzVSlSWwqdWzg9rvuTQBZp6o5OCM+ND7up9WN/8ilypzCcRKph
XQsIGaoBkJj3sBjsO91keSKNdg9MxV1V8DejunaNA8iNKiu16Bd0/UA2s3nn/Wiexz90SerKABUh
PfYVveEjBUDXpuG23fro/MIcZIdFeZECtDbQnv22+wd5vKFPEGJovN5jUWbTVbPctwRABXnaA8Uz
L5HeGOYMvXTAfqNY9MS1PruVYPfVFrWrARj5uwlSRkveJq+88OZFyDa17pxf4niGWYEX2rhRXRVn
IQiPTMHziJvX9uCGSuJoCdX41NhKilVtkz61GDNKaE5lFgvQnB2HtukvmRK7lOJQR9ld7rGZiTL2
TqgMrR3CJBP8ky+T2nW8+3wj63fz4LjujZel0kH9fZEmaaZ7+gId45vo8HmZDtWEhkYOXmRAhivD
B9yiyM13ZVGDoPpl0Ebbu1/POvBaCutPyiJBxBluZWAQSWA1qZV5IaWyBUD9OeWdbejYHFUyHTfQ
wzgiDiO32HgUSgVIea+SErjDkopqK3GOIEm8xfxBm2xeK2cKRUE20mCfdGTqbVK9EgI2x5W7uIt3
WIoBQIxsgx5F74EWjY9InoUxy17aU/CsJuowCpijubHKfMFWSVpK9OmPmBCegr4Hr5IjuxIa4UER
/DuvwBwrNuUaf8OsMnjQ6RqLMZZh9Rg3i1yUqfKa3332/YgfAkW1dKDfrR62YMHvXJTrpPR/h5Ut
O7EthAp52algBo52JL88xZaYy5/ULE0WCt0UO1HHQ6ZmleFHDca4y6YLdCWVTq9kMBfuMJHa/1vn
iKWSXzLaUwj4XcOLP1xE/w63Bzg2BWMmxPNfSH++xtFFeCrAVmzP1cn0UOTNvrAOY5PwcqV3aAq/
OlL/DvyBzZvYm7KKdL11colqln1ROWCnbGg7H2IU+TuKG9Jpq6l7HIzEh4UDBS2MYNoZ/OLwfJ7k
FXefPlQmSv7YrV0VHT+qEPJK/gNoOEWsGbVEdIboTl+dOOY6eBRlaQW3kuJrYoJKHYrUxJyzfjHG
c6sJS+2sUUEfh73/h8dsej2P+b21S6V7ayXxXR/H/KG2Qw9OC3Eq4Q0f3EYseSFjnkg+JKCgi1IK
ptsgpLRiQrnVWWuEfahD3J36oZrxoKMftzVdIOyhmHabCakPHFMFJuhkgCf7rAxrvfXD/53MtRNL
xO9yTntDv43VwlGDnbLeBOfhulJFl93rpmAkCeuUhNW94OKAXvX5X0Su4tavCNv1uvQesv1iXMb1
OvlF7Zronfq5lvAnWr5OekTY9KGTL1tsztvOrEwKtD0ZfhaTyRcstep1jJ5TpFpAzydKYa1GS/Jz
KAnxYLg4mCx4pQuCNAJlrJi5EJiKWAEBOaMgRCapiNQQGM2sz1qOZBoaJi/UNi6Le+dmcbNBdRgi
lyuqSJxK6yz9CWnPpEDhLEdh8L4jdvpji7oPfd2GD10gFXko92UUFw3eHm0hrfcNaYggtzkI2K6X
CY3lg7TBWpIHQUxvU7IU/knapAKQBfb/2wgw2a4k6zxMtq9J8q6bugPamDyS8gPQhG5zgp1nMVkV
IOhFe5u7MoToouuWsJ6soX+tmC2G+aSUPfvoL2e5YHYzhPU5OVRkPYl7pQJYkFVLDJBn69SYDiso
cLZBPFuzWV8H7+/BaaSa9y4g1iHfLsbZruQdqyphha2/ey2G8veVAOqswYOlmelqQ4etyWGBQKmk
jNwE+g1ETpFtREbUZxNUZ6oQNow/LmxhObLPN/N3gViH+snsAAMcQ2vQSJwCZ+Hhpt6w4Rcrn39s
xSMMJkFvxcJGVwGlJh5KFS+z4cuYTPPHe52YkCe4FnbQR8IHBqgy9aT64pQkdczyfxuwWWWn9ZQH
NVqt419N2QXeBEBhYMBTFVwtEEj1+5ccDy0q9cSGdwKDVgrs++IPS/KJ/cttHJZVrP5o1puKpwz0
rwJUK7unD+m0PuBauum2JHlhjWI10cj8lljamTe+HEtiOjN2Hojx8PD/ZWyGh2ehso1m4C3ew3Ok
4dxDP9ePKenJXjDTIQOELk83e80Kgb/V/XOc9APObbELoblTTaANhVsG38b6nQWTaa/+ubQeZvpU
jriX+luLytfblbQnMqjx38BiToh70sz7WT/kTVREaypBraPpWm3nOtF7bpaSW3WjLLx8gh/v45J8
sdK87fhj+9rz2y6zJ0n73kSU1reu6EVpFVBT6+KAMB5SNV6Z4gU7pFI0St6HLE6xGYEYLKVpv1q8
voawkBri7fxEMa2uap3z6cQIlIyLK2z5BPT5hA/AieXVbHkcw988AXpOCQhw4ZEAzHVqxkowICcr
e/ZVcurmrJEE/occjGzN9xY1HnUYRCu699fs9DjEhKFVChW3q1D0o4byb7pKoPvh5y6MNjny66zy
eqlUAChg2HMSF3djftKfSQKxTi10IbQmRs44Us1Z0xTh/G/rduJLW/76qxo6I3vgc4BuYs40M7Bg
DpVmA6GFr8Rb9D09tKhnmY1H/NTLlA1aK+dXhZ1TuFzg9XdRNqNAUJo/9np0w0VdOtEsI65UM5Er
kxzgPu4kMZ2YzrrToMTzq0S2fan35jRMakPXzpMd0caFisEXKxszk4D7DyXEtJc5j3v9BpkL6Y3P
5crR+0s+mPNXROgGzZW+N9+bVLrS4C/uSxWWE4QN0I+/laAYgdnwmk3a5Gbgs+3Pve/xRMmvfJeV
CStAZe8ss/DF+ONOe3DpT/hN8A3ZsE6S+DIIbtGgPRAE9yeylbxlpCNralPz9q+nTsa6/mKCOAGf
KRfl1Ut4MvUvxOVRFneSfAng2aepJ6Wx7y4ZbQtn0gERorTlm1X8poJfImNtA8VxuBH4X24TzJIq
JTrM82fPGl061k3oscoGu28T4uMp2Em1kHllqq2xT2Pv9ep/u8Kyxu/DhBN5cNbU0QtQDIzDmk+O
9Lb6zw5CK769ZmYi56GSu0L3AghqZseOk/zr2MeVjg+Z85iZ6165KDzVj7pJccvvjM/KuVJenkpg
tSDGt1zOF63l69QHN2IdQ46A3atC9KuuYuPM+inQpU+P540HViFF94CWP9p3yA6Xr56N535YcPn3
Ndo6leuefxty9USxY0MBAi95IMY1BuPoCBWKjIX3k9oM6jXV97NgFpOzzQ20fzQni4iC96SrKtte
gmbYDRyIZjvu4R64huR3lTpfCTfE3UlQ+t5Y9ijSC0OsNygjxCt3AzsPeYkqUaUyDzVP6k7PnzVi
VTXHrkXuLDCBDkfz1J/EcxQ9uJTVhVBLw3SzfRF+l2IVce+O/BbzP56dNarCx4HbM+WyowfeC3/D
yLYcIMclZyBbdPFxkNmwOTAi3hYVQt1un/nl50n97QNCtH7hOAVBJc3XwdhYswIYkuMhCBYR1y9p
yHhiaFADBgBc5QBQ4npGdJEOmZoz35glouuHB4z1LBYGbxch2EA1woftsGXBikGMw8i78hyKC3Iu
mMjJ30ZdW6YEOao3TLvDUtd4dEV3b+Pn1Lu2P8Ix3EzO9GEUwaGuw8adBwLmFaQK+Vx1sU1vtGB7
a1mlTpnrLTXEuAOPg9BxNzbxoK1I1glfOIT9YgvrbZGZPV+0pwDLioFh572LxluF2VJqTh0HqGON
lYNzFOOpwlzjoVoxFf3sHX8AKt9LF4k3GdwsUZ43/EOBXJI+AcyXt3MTtYkGVNfqFFxouZea6VGF
QeCHn32uSh9D6z/ZwjGlVVl2ZuZzefyKR4FiHFtCrIwuprcYB9HMGcKE4NqMhQD3gquTVCN22W6f
oIwWqCsdtxWs47LhSFWvj04Y78H+D1wfwZEYT8AJTVZ79KpaKbXlY7NCbHtRoZjbf4nQbe9LJGGw
FqldTA8TNLRUA419ypChz9WUs3kbvNruWc3QVgnsTE+3lq5y3QMsTZybdHpHklXmjPViNxcZpUXp
YHZlCg+fyUXdjANTYI+FO3plN8dkUGQEcsokF5fULy5Ozh/m5IzpCOwk3OWmZh8LWwE29+Hiovin
IIvr+0Uzsxf1btPW8lfMsx1ml7VnOm4gqVyxysmSzLEfXZSe3ZaAbg1KxsrZos6jVRUnVOzyJ2pD
aYFFczTvpM5N4yQ2MY9tIiAOJmajmBROyTLurwtLupV3erS6WkIK+N7I48vKanIB5Gd2jgqLjoIC
Pfm79ChNDci2KDF9ABWo7O74eYxvPBYMmE5uG2JiIicZqLnH/CfLxIToLChBfVoXppTfgOhLn8bo
pmqhNNpWyrnh9VgCJCwuf3EBXy2Hv9oLcJMveE4WZB7hPQimlfj3qoXAZBHzk3s4P3bbm6gnr98Q
ZbOg/dm+N/o/9g7t28WdY7r7KOrbqrspVgRPHgw8vHmD1+muKsd6e8K2o4yd8SFH33WHkjaDuyo3
mDjlV4jwDwjqvLyv2ijEhKGF/muPHHhCF0na1vMeXCsQZdVOMeipk6gmP9d9p94wNyNA6m7PfDWI
Wz9VR42chEAmaJx7WuyzGGoRiWkc2r+vMmO9j61oInMpZpgwM1erkdEyr87d/ezAgNAp8cpLYbhL
6GQ4Pgp17Puv7ZWC5Ea2LsHhMW6RPD2NW1WLyor+W4Jlhj6H/BTqHNTkODfQMwUyV7EwZzjMm8G1
6tJI9Y0vUvP0XVlO5quueDyHSuT9ugktvSfuftT8nsArcPgEQ/uRaNy9gVNKM+B3swdQOEU2fnRD
sHgxBxqIGMdb2jIQPGGm9ZrexavG/wIezYNSIztEirETXoNl+qx6HEZZ/K3ELdGMfar1nl4xJIo0
sa/p6gNVQuzaiyKu8TMhSrKpnmJN0vkoIvWxMGkt9PuZjJNGwaaKc3cJkA5PbW44QJ5QIaH0KajB
fbwAZJVuhqOLzcN1qhfHRaq5ZU7+qLHI01FmOq4Fhd/0uiaPfNbkm9Eizodhqu3rfkaOOhic68nT
Xr1nJm7HAUoR0mcGsVobnYc9YW3BKD7PkGBAChUOIi3nu/N7AGoGoggNG+8IDT4cgvwzoQYYr0TT
WTifraNY3gKoKxQBYv+NIKr5NhfK2m/t2wW69ant1ajHXLRrDYeVEcWGqwxdWKm+VAnhSPTCiNdY
rVFxzCjgO4/lm2J/IOxwONSgP7giJulli6amyM2DFQ1Q6qFi62yn1a7pOPJKVlFHqNxItDTvN7tz
gRxhsTazsO2kuSMSDB/sAzkYzJ7/hTrYf0ZhnP9Vo/uKqioF0zvntvWXdlPB2rFQvnzw6FYfGTU9
RV8R+Lc1soCDmsR4M+Xkbpgj6VE1boJJKx0RXYK+IZEHRwRPQ5aRsi65fsC3vMQ8RVwVsP7YvHGj
yfWBAUKn+4bZPqW28zbN+RpiHmj7oIy35ZfT3Y9j6rVR6FoUh4Ak6WJ0kkSml+wadw/8kt2HXzKL
Agwhr6ZNTlkBl7jle/89DNSm340S/7QAIz+GHKo9CMvN8e93U87VBudDsKLDLsGHX+fPVyvU2rsx
IjY2nWYv8cLc+534fQ2bLcDQvDUxSZi4QpR8oAGfNuaBtdr9bUf9zg/ixIcwCSCizStQ0i8HW1vk
NX8pA36T6+xiTirHxYz0FwvTYZphJh+qtpx6al+jsNN/d1vNwlVZWPZzKUzXuVTmTypFjvOOj1iR
pBcH5IxUCOGtTHRWns/V9mpc97kAIw/NJN1ZqwOgE+DbqLsSQNFvKUQDfeJ3/F8roKNcJI1r75FI
Mk5OppNY5kt+AXs1/pboVGhzTd7OrHU5N5CaBGyhIDyl0rOnsRcmeqjjx3xV5ho3J1mfzIYaBl5k
iyePzdtwidWnPrA+ivdzfhSPyY1f0NNw35fSDa8luTjGIlBGNCJxUJ8i2X+0w27tT9O87NK6KK/U
ObPv4mDBLKerfxIQzPv6Su/WEaUX5CRKIO1oo4I+v4nX77E6r2Fsk54MztCvqKmO1fmW9y2AUUwd
bOm1mo5VCnrOlWyIp+WpzTgMb3QysIiJcRK6BkDDhPnXyAQ2iH0cHm3Lpwsae0ueyQ2S06Rxg8XS
w7HEbqrEPFzGhT+dS3EyMQG3P+VN+h7plu6Sh7iQdq9X2tNuZCf+y854dweiFl9NzRb74hUy8zeq
vtRq19lzBnYECnyS8egEiKUF5hOXIGuXtXnmsCiacUMgMRTvyYj+sbbNOz5bp6m+090J4J6H6Uo1
InulRjeI8nAEgUz3qOT6hE6fj6vqrVyHlLG4dgGMu5BTrcj3y3XrKzkRroyrKE1aHVTH6Vl/s9eK
qJNsjyTcRCUBnEZJG8ReBnfnMX8G/Vosi3PBhVtgMS52/gRgjidaewUygJEPumfrvofbHyWEomHE
t6Dn/BWD+ly1sd7Jwq6dCfVGOTT7NkuulsRny3Ol94OCEGrYet52p/fUKtmvlCk5z7twGDGzFbPG
SQHCbnolSW28LjSuYUQCgCOr2Z95KCpezxhUsl364BwJcwUP4D5JysLew/Tk0vfTd4+CLZGWr475
dpWMBATKt5tGFK0aXTmqIsaoxavsPzc9Y/vdB0z+ndjgqrf3F2+HDY+R5l/9g3fLoirrktp/nb45
rZ+Z8iGB+XjJ8wHTwOjyEbdIoLOzfD+Ezc4FNTrLZoZxRPAKFq1wc31+0jmPQmIrqKP1axWF6fmO
Zi8mHukcjQz8sqOVa8fx+OlplWMrwqv342Hsu0AAnxWF5X4bMJTWLCk0q2+bQldR7sIsp5y2ue2H
7A/7SYWmGAkpUDGXKPdovQCmBseuPiqHlyn4xN6palRcZ5QHhuLhRc8b9uryrMS+wN733QiYc5GO
kpllP0XeHoZ5JNDjeni5+m619bBsKKT774M56yxKJ/SyuN5TDUYjvEQIKFM2M9AZo5rcgapLfVOD
57mdRu9JqDini2fIwI8JDEHHlEYP3IJUI4SbomML2SKp+SSO48DPlksOV1cU+OgBqJz50LdS4xit
CGMe0PWny/VnvqbJSIqA2fvVKwPoH29RPRuKxi283DrvlX0xyBelCOroutOaN26bEs+LdUtvyfzQ
bOlbGfFDNFqfhZPLqENgIW2rDprzJK06+8vaNZgE2uvjzsQAzx8KelHcb8s6b6o/PF5akg/qv0k3
v2mpRYKmcKZdDFdPPrNUWXW3YpSWqD+FU+QSHfaW3lgnUpmPSWwzQcsCD6pamMoUheVwjNNYwnJR
8qKHyFSwrB7mOCEnqJSHOEbNivFxCPzn/VCwajAqXOR0+32NCBavslqp0TFAz7rS2qQ2Wci/BcjW
89/Gxd3xzaGSLv49Pb43CxRzmLHfgsAxfysPcR7JuNiOqAhgg4aqX5XCh2xqxDe1VdlP5/T4WyQe
l6YxNeb9VNIArIoptxZW3hQ73WWao4vZN9h9A2rjLAJf7dUC6t0A6OUgaKxc2ANR1HKc4HN2FvFq
4ZFf5h91s83GeIy7XHZd7Xl+xlFWu0DrHGN82iNm+LhUDVoKWyK6/eeuHSPz3rWgw5HnhQ7Agjtc
3yeI2UCMcCmaYtSjlK266NrdqFcU7dpp0tFyKCP7TJMcZg+kcuLyrWfQSG+e1VoXoud8wKqNE9fr
MiDEI67XGpu6wjvev9UDN84o2ceI3bcc58JsXIR7bKqVH5DFpLgnU1EHnMD762ugN6M83di8Cyyq
sF2g8h8WI1MBxq8MPscGoqg9RafMGZk9UAAACktFXRxl9PLf+13iv39acQ4LlHwebvMMeuGOZ4TJ
/W5TFOAJVYccDE+WYMhnojqVRaoB/d9D1ie3MIfdf56lrMP33GJgorTBjs+CTqnBM38ApKi28U/2
Q25VmOmrmI9jV3q7kmP7v0Vc9dimueNYkYopsJzRJ54KRPyOmmtVo+9tILKPsRLnpzUFWTvKiyeS
E48Cx8827zC/HPyp5jRCIuhBgmFc2wZ2xWPmVPu89RXRE6WuppGkDecu+Oec73PhP1ssDOaHN7P4
JXlhWJMRnSeKu+KXvOTdhPVw8Np4QmIthytyg2eniJxOGU28lL27ch+U0Ho7DesNLY7aR921iAIN
wpaRPj4gT0wY3SK2scNfbvOJ/Z3jGHMsci7hy3s3Sa6uatVDFDgnQiJwYjdDnecQMRk9XWQ1cxOP
niPssoHoeSVA+2ww/1M0Dw6Z+0Y+l2lp5AobTV37+fv2lWkd+183lMtXW+SunRPExMl5D3Sjgd7M
hIbsEyIpZnnTiTtOYtrDHNtdvO+TDYat/ozenhG9x0nVt7LGMimiN5LCHH0YH9yf8G9JbGJ0wRcL
EkOBrrV8yU/alSr9quZLw40K1lskA8Idp4WFT6P/K+w+b3Ta/WpIHHgP3NXzeHpBnUdwMOknj6z9
V8XcgOenJ7b8OTzlcjOQYjVilDr1FwXkMreXonEynwuJQwberUxFwk/Od8SMdQpJT+bcSTPZ4esK
0rDFk8BUKBW6tEIXewT84FZJEcIq7TXiFoA0NagUPiug4u43mVeVqmIs+yR2ZRc4qfeZUHcAjczC
sSgqWyg/fV8O4eu8wKa15gezsXsJVk7bw6em8dbuE1oSYifahde5lCEOH0rBRCvTvoIp4c1tfEsN
Viyq98BuIBxKUEBnJ4aqSGcpo8SHiAZ8eB1kUhC4DhA5kmE0kl1+ehIbjUBs2iuBej1DMQwroHhc
VfabDep4FjYWviLCTktXiJExqiftp0r+LnuLd4E0qryCGABnMJCOTnq4NGxikNwqSXJInSyjj+sd
Jsicu0CiRmNknmEBYrt7yju13yumfxdhqxXrEEz200atUZDw+iKAD3F1ruVdbKccqnuaPFOPNm7R
GM4t8C5lRp7GgIV570sP6nbVSk1E6JpUIxrqp1Ui2eW1BTMyo7YegYbzPDnYDH33RABUy3LRd2Ql
/ZCmYt5Crhs3YPOCsG4mkWar9nqHXX4hfHtn4dil0br+iFa+e0z28t7f4PjzerI1k2WI/7V8n+rt
ajz1P3QpK5fJcWA/JHMKE0ycSiRFY27BqxcXUQPVxabfoR2aJVjmzCI4bYceu9OyTh27bXvSEEzB
+t5JXEXhXbuhP6Vj+RpOdnfFBG4QSMvbVOP/XFLlQow32IsUjsGgpO0EFlmne4Ht51h40Y3lpwwZ
8a/ax4lHkL91ANobKqXS1bT+E9CPJQXf3ZXb6pjLo5HQgfbdTCNwx5cBFlCT0KxXt4N/ysZBWVkA
kq1dNQwGazrD6hAaYTbwEUbqcMM2gw96zFNip4afZxSatN+StLvLhGyJKuiqeYN3UAjR+9Y5XTNk
85NI6AfxvToxl1ljd6l+rGOhMuTWrpuno2dJMxp6h7hu4AuW0H16zJDF8mpfB5N73Anqx8KeeEV0
Q0mbEdCtvXyKAen8EQdQHQuWHxSF2sEZCsqsmjb6ua7+g2cLdOYFgF6MLTzNXN1CU79sCIppcb3S
XtuuBvq1SVVW0q3An0Ck8k55M++uOUscbKB8C7YGMpgo3klRHJ4PstLlxCwMwj64NMlMhmN74Jr1
pAftwC9umNTltH6f+RCuCRufzU97zFK9DbqfGTisckLiSHIzsK5Efr94qf4lH69GqpNueEshZb08
6qSXk6nD8yG7RcvhYJSKZCf/5wdSDavDP6LT+/Lhm+7678BZORv0a3QgCzKC4hXMbGVVj1anXzwk
c5ddgjBttCLnpdM7GriPRc8ZoUBS1LrF7eZbA315akTxfxexbZ++j3H4X/rNBnK4wCO3kuDfSq4K
44iUPyQbMA55TqsV462LNzU6gKoDsxXgG1mDWTkrmTpUvRlKkI4O6lFOirftONgyp68xsTf0v0BI
4pksflEBevGJjoW5o7jKv8Cadi5OrwVBj7+d+Yk42o6Cm5f66w636x6pxiMOpeg6uZtPtZ70Ak7h
OVXTRjD7zdn9LDxgJ9UWwuWocILC1Qr+uNXCtIhXbpx1riYAdsxHv4TLBnC9bSYODqdEJBhItOL1
ZO7CO8l+od+2y3kEDr3uTkoreuvDgG1vounRyuaf3PiX4+r8GSBKgLX+a1RXIKNnzD4+qrWFwou5
iKoybw/n6ecLkSqTALDJDuP052BDHRqNmyedS5LY8Cmbjuioaiu+TcnbqTrzsbjL4K4PFJMPz0jm
hs2CEum2l/WpPYcK3ATQZu8D5ViDEDX/VYyV0Agi27u7DKxjM+isEp0Oj3M0Wbv4OlmEE9bEYDsM
7KYJKgMW0YUFpYxNbzv9rIDupZIASHtqnL6h86K347Wo3maXyvCizlirJnV2OllAQ/lFWa97Py2y
f8ne3cuKvAguboPdfDIJ9GknAE+T4K2ikOyEi8nwwhYF1mQw7WhMw5qM2vCfs1K0yDf3g7/4sCYI
5EUMJ9pANP1W9RYrFYbiI84uzg65jg6+a9lX/yipGLAptJ9zZI2qmRrT3r4H/r+8m5dlZaeUMFwW
zBAoGjMk/reaQdHjhNL3dxqZchh56TGQ2VO67a5VEM5CA0g5YMWvcej8AjhrmjLW/c0QmApwUKSv
ypJ12LYUAJtTrNcpjU1lCKAXPBpuiidm7+KGjMAdWLJmy06xaqZk4NS9SBd/rpEp6gbSAtxtWsEb
8g9eSIoc2t9Ei60FmkwDGOyYNZAKPlUdWeFEMhs/dlDRKOrJOHW0dOIYA8pAJnrkyw7oEu2C53dT
97cWQAqyXSw5n8v2u7K+tNjhwECsUtnHcPNBgSyZh/Zh9TLqU8iBt89LpuZPifSxBZgn8Z9DVGv0
qGHBRGdsWHDl4tSZUtsUsrEnzQBWwtRtdgcb2p219H6nUf0mmXAzmbpPSJcb/ljyou4sXtERvqiT
5n/EsCOI2XUi8MDAHrcSeShhfSpcil40uac1QR0CsSLHYKN6VNyD2+np8hiok1MLGceHEOw8caTt
dRE6eB5aA0JBUsxp2LMMkKGpO5pNk37oaw665HUlcc0sd47lJsfAmBQqmm+xN08Bgvu2/RcyI5Cd
c7ICMPJlQgSfLyncuxPKdCL9XPxIsduvbeWi7Z4+0CjoKiRVGANf7FE+3FqZxvPXeiKLEiM66bar
phDHcmguVx8fC0y7lBh5dTEgMNYOWJy/bw21r6P1QDMIdmtDDU4ugS5DAW1TgnpBxolUSQVZ97U/
SBYXEtGSfZrDRHinbKmz+iOZMLZzF5qlVXI363AqIjFbsCUMdeqjOPlYlVSHmHRkiLn2GoN9dESG
8tu2K4zZPZehTPldl1khxQTdp0A02HXemhlIqR7xO4NepYNZ0gaG+GyquzfwTlhvuwq+YArueES8
MGt659UVNRGnRkDwWM9vsOap1Zag+vwBkx4Z/MLSdgP4PEttFl6HPEupMSBpx1yGacYiQUiM5WbM
xrpMIebdATOoDm22IKvVr+ZQB9zKl7Q+FgwCxYyt4eiSoUdGwglimD61aqa8II8TmyFfV8AeMogV
uf42x3uUY/BRHaJM6CE8fkjFKAN0dG5sssWPrejeuqdDua9UBlemYT2WM4Q5+1OT1u6n+uDaXi+y
ekiXptDagjJIsEgzLnnp287jNKNshbhPBLfmiFXkg8/atJALHqEXc0cxCZXLnPEUDHMaxO17LteL
bIwCukX3bWgUU1MAslT2TwnJyG0mIcequfeH/SbdTcoW4IOCNt7da+92Hsh3wySoT2G9VUhunlot
qOCcqB2Pq0fn9q3t8DmnwvKCEI5FeheUre5TRNM6MUutP8dhOPYDwJZlz4Sx1NvAmjBs9k/bUh3a
fiwtVCdARFd1HzAIJ5uWafzhIsGW4DkPgON2XUrFe4bpOs4l16wqnFQ11sQV3TfTArXVREm0+ND7
6iIrt5xyR33+rW3DXlJqEPD9LNyicG68WKaAZUc22rIdY/lmRls0jXnpIP3KVRYux/EUkD3m35Dy
mSUuoLQW4h48YV2fF8x3OQ/GZYPvB2Bqd7xGpF3N6wsj8GOIsmgmD9Wb/c2fqTapD3Y9f9oXzvDw
DAhjqtlNsvCA9Y1Z/iMOBT24EFnOPWjjsDf0Tpnq5VIU644WaVF9wzch+Nsx3EGCkwouGzjqCSCw
uXpTbsL82vyXztpdr4csISrnFAwmieQfUEf14/VUOwYx0xgSEy4ZC7Il+1B5Qd1RE44OJ8IqOkFB
8Hm5CYuk5CGEQZh643Q0WaIQJpWlLnS+sRlfR7FgNuxN3168Nh6MptW4kK3O+08jduFJ0bRwkBEl
GGnqdr4NKj/yYIM14rJ/FFta2QngrnkWpalIijvUTVJsZ9eQXsTEebLpt3IZPIDhiHwO/FLZHS/r
W2cKKS0RXuXG4z+iemD3+wm5Fl4gBEdN/tXWTypdy/dj/OuEfTTxiRfUBaSA+VUGC3JgJT2XA7R7
3bKJrFMpT221hTnUpvQ5GBATX7iEQExqUKUQkHMKUHovE143doybwoUasGpNuBTFPCT09vC5xljz
ZSywtxCWeHIUNwf4US9SXn9Rm5XNBp9tjO6Th0TUhJL7QHmXHRjnJuC3LadLwuEDsGOyS1IwsJCM
/rbNNErk9NQHw8vy9ntiyXxhnCsrDHJGW1oM9XVMp3EY2bgwzintDXdMNozmqilzI88Hmv6uIL5x
YWvJsv+zMUx07qIn65qarWe2id+37Ol6OKMXeVfmRgRHijWzybcIVCvU7fLnTyQhr/1whU4tZJhC
UOExc09E4JwXmzGIaUDryhzkAxQRux2yQoY10WEwbzRpJR3Z2PLUyLTe97Na3tdfXDU/mBfAtedg
d7+8bPfWKtj3fxPtvi58xULAn9dhN7dFiJEYLtjCKIdVXiZ3rrnDRJCoHvGvOf7VYQ4fV27YoaWd
sGRT7r9JCVgK0cOC+Uszya85pXeiLFsE6RzJ7aH9MvRJYCCyeeGfn1hIL0vnt8zCV5OIbRDVgTNT
qetI6YP7K41ciXGOvgs2B+jfeP1A6NaeNclxxcOHfPtaTthnMafFrWrtNwXoZhWOfFp9zB01TOU/
WMXA3hTPzN0Uvfz/06ApCunAJMhw3bekYpFm06aoqv/MfoSZtFggCw5eV2aEUFqN3BcvUbyt6Lk6
XE36nTm1KGNm5XWYDoO4spkTHYSW6sslt5Dnj/IhqiNtH1H0F/qKiruBzVI7K20i0TG/1DO/JznL
RL6vBRrJrhNbByJ1ahVl0EwPrnXoqjcstinmvRuVoLRcneQC+m/uCWtFrUjjFucWEeIyZL5W4oRd
MQVEw6KKdb/gKK5jwz3AwvIj0nqjQlb1eNMN9f6L2OsBgNLeohbWI7tS9gKY7gUUHNtbP4FyrUcG
QJFCT4HT2y52893PT7PMWMoGPfKWsq42+1o+9SNrb3zQEx0VnR9KJje7Pdp0ThK0QLoCVTbEC6oj
vX1Ur6zNDCH/u5EDciAqDPfJmByg4NFJMHKnvV2SWcj5ycivAuYmLWbxWLar868Mvn5z2u79OqVl
yUJFY7AlHTN69Ar6zOhvOz0NZp7D3L9a4HMByWk3RAruyCqGPMCWEEN7oc2G3XjkqmA//hRtcHej
snaEBGxsgPL38zf1azI6A4OVW1JFfMQ5Fs6OPTHYENSWlGcRE1rmxugypWZU347i77oPrwsIItM1
7T/FyGkLrvOkqUkN7TpJ1fAGze/jP/rWdUUDbH/eee605/hjQbvkqfVYfN2F931o56gouM4EaXRf
SfTNKiki09Vuy1SFF79FnZ24cmObJsQBqGsTYGLawYC8IsmYiO3ZbEA/yXTvxpopNSXyYrDXHU2y
Lykj849b8VPjoNOOacRKCiCUACWXILgrrYq/2ieLO/vCmgk7y19WeiEVbl2UWQZ2WypJ2SlVEmYZ
bKmjjLFhITSgxWt1i7Pn6+g64+Z/vwi6MDabKRSIcZmYVOrokmDdOa2Xu/5PL82VTrSlqM4cDFBv
gn3yBvg0er8+/+VZMqCXxioaWNQx6+9pCF6o+fv4lJi0FDrBCbY/kc2zpWChvLJNzMXFOQVV8NNT
7+vnVSHqvA2dHO5SOV5Z2VZ2RA/W5T5FgsPSvaSbvy/QMSGTEhuQuwdHXKMBjWSUrAJg4YnlGhYj
oElnmuX90zpEjjf6k8lE1uzUg5JynGmrTHyn2YBwGF+veY5yVZ9yMlOI39R3VqR/6+2OBxc04yv9
MDN0WjYHhrhIXGm5QwRMfVRDrEmtibiGBvSEeg+JXjpT8gNyNmgrHg986b6qPQj+LykKLnjrkgl4
/u8PdzR3rdhBGU75R+2CYzo2DMxQNvFCp5Mjx3YbmEuygi32v0j3GSWAB7l0yTkxlo7uzzKvt2/Q
/B3XBLSlMGkUEP6+biVh8FzMMZ+NPzBD9LH+rZZ7f+EagEqqPgfg6U2B3u71yqFtJN9shHyf+8en
c3Utq+wmZZr0c4PEz0NvAJiOaV67pHmoqeP8fNZOYLdWX8P7PsOVaZvPgSA6nB5bidJJUd2r1fpS
KlXztKoZbeSBYAXm1o7SpITqgSE2ub1q2gZ8wIyQQQbQ6k6OD+XqV8iLwDU4HhYy4mk/V7bzYltP
pv7IxBQ7pMiRGiMCvjAaoFJCAc2ucuYd3jdVuzsmEA7xwZ/7BqHnEirMC2lKLChJjHUZr5SKocb0
SDmVVAn7g46bxoOrnEfoi6H56nXP1EDgM1YZIaD0LAUHv/6B0s5tGULMJgK56wSgTUxBtZpVOEh+
ktGvgZVbk+fs8KLapbV2r4EBATeed/UvW4MyoY866Nz7f7WXbHpjVD39SsUrHwL4yF9tV6CJVorF
JNLMbAn8zAPQEN902lH+plHN8RaQwXu/iKxRVE92TxOcplXfuNkNa8opM/et/dAxxJWDxxFV6rIi
acFuH9r/ukZKarGLSAmXDTVaeBLvwXHeUEfUbYqTOX9yrNCXuatSuyDVbkFP69868GD2ItH+orIK
ZXL532qeNDHEhM2aWBMZf4g+yFbHTpbydfL0efUoPjWAjQQi/0NrXfiP2DZWseChw0HvIQ7UuBEd
AxJckGdi/jm/KnLA9Fj6O4JSk7kn0aNz+J8SYHEN9HGev0L+BTWajpu5InI5K0FmbAWJq5V1aWIc
8/z+SJ7gpGw3Q3EfAcnqh02oYHevJIO8GMr+NDSiZYAuMlPF3QdZjCwCRQb9aYa8haVEGByMCayL
IWECNa7n9N2nUgmN949WTFHI1JQ0PeMRqte6WcYjPVAWkxQCtJpx7LcZUzp5ZteY+C2bFkBN/FlF
EBAdSGeIhPzDppiXTFmgLamztIChtWDLxOOFvRywBPYk9Pc6PkwpH1Fmepsokwr71Iz0ZOSP8TXt
A28r31Bn/au0yTas9Lg66Q3UKHvb8uLmhBVY2LROxqUFFLCUKNp/ws3NVlAC1Q7dSg5Pbmw9qUk6
lD7sMtM2u35Ma2LPDc9JD50w8InzTHqLYCzKy9lHUbosYHe1kIr3rS/93okaYfSZK5TAAuHQGSkB
vi/mW9Zi+u+3wtoCpiiGsNIfuExuDB+oCkZauXje+VhT9OoucTpzOkBkQO0WlLVf7/axGP6nfBWM
bIPXz4uuSf8okJ1H61o6Fr2fcTtHSmCaPDErkciZESXlmQ+Gia/r5jJcJF3t6FyQHh9wzeOTxfbh
ymEB0PJW0/EyEc8VADRB4761p9QcpwQCpZgo2BbWmp2okXuThLocj447TEC0t+jbsQT1wiYaPVGF
eeb03IDdHyR2Ggem8TM2IDTxgv8NM/h7hSQsMqctMAx6yJiiZBXlBigFpot02baS44q2fU9YisY+
zrtYUHA3WPE+HMwd9MWoHzZDZHU5HD15Jo++lDioZ2RNjuaARUFpouWWwz1Fe9G/pUuQbnCBofWh
1e3T50ZDUn0gUCKRTY1VEpBpjZpEGfSbAqrR347z1h6Vgf0x4P6k3mHS1FW4Z3X+X7pf/XQIcoZM
mpCtN74xE6MgljY87enXVCiusq3uf5YuZ2HixHYieqhZNSKbEtbPbeSNGwEn32qaZGUghrhGihaR
zkstNpiQVyia809gVI5xQl7Llmv6iw0U3Jx1C0bWZNo+NZoiUIQa4qOKqiX3YLEwcepNOxlid+eT
gwfos24r4ju4Y21pTtYo16tj1XLZwwR1wTeb46hnUIGbfaYJuQGQbd2wCjwZYmMuGk3HYK8A704X
cReiYaP44zuXfes+DRttchYKPEnWyYnymkkjwD8LyEOeWCf3nYQRcbIDsNuJZfdSISII26JhrsIi
Pzg1smfrmyWrTNo++5fqGLFxked6nb1/92dofJrh1V464pshxnTQ95sgnJG3sY6I0bxFMRm+34Gs
XhTt2pKLDTgCYGglfyRQny2XS5o6AFurW4ngn3vfxd1qBTz5WhojAEfPZaCwQiZ4BUP+ZfQ/bc8I
dfc0iJ6k22zf3yRcnPYasBJc4idFkD65dT8Xu3Qu/36HtKl55o4QQHzfK2JtbLW/5SYmYw94QGmL
ZoYG70yVWgD64AUkmFvgVuVvbww3Ao34wmGN9kA7CmFocOWfoBtPYTGz8/ZfsGYhpJQB0iI9ZvZE
9liAVm82U0z1ufS+N7RKO7Y4Yibv8k0yixRLCN2FjRCzjcbQ/ZhTwUzOb9OKJ+zrTOOdvNz8WE2+
FmwQ+L3/me+WEaCCdOblNWfCuAtzzXrAeMvaGAB2Rwi33DTkPDwbSDW5GCzR0/0d6C+Tc2DHfqKG
BDnTXg9QwyUj2Vkqt30zmhO0KRzRxg17NwNeVr/OMYxL9VD3HDapq7HuLi4cVtfnoTAbd8o/VpK7
HybJWxp+vJS1But9E2tZwc+kl6peDQwWjLQpd9PXlv2+CnsXVUKePxhloz3gVETdFNa0gUQL0a3y
dCVow8xUBth7LIia/n7JPJDW2ctFqCZ7FXdj9EBhurwbMNyF636p+mH16f0zSOuNn1B2a1I/QAM/
hTm0OFuWoYQKrJ08Quq4npR6wPXSO6a5lMEGncSl3n6naZZbwA3Y2e9kB9oDVzmKvmiTqA47Vjix
ZpjmVz95uuk2t9sbTa8s7pIuUk3KGh9LRptS7ybBntNNtaJ9paxsq6RztLrv1HSXZ2BnzDtVdd5j
3UlLarolLJOsAmV1t2YDlsF0RPmM7gN8ajWD4UwrSAVTqTPt0wY/WrH5EzZKwo2iF9G1JFQ2sFHr
eibErt58LuS5u6zZYKTPoQnzNQUl7A6IP6e3/+UIVYHbv2Up4aBWzanqKfZfHNbIxxAbEtCF2EAk
V18iWPSjZdLCcYn7mrNkURZZmZ+GpBtcYDQqwUV8ElmdjKEidbAolbrKzIECEg8C5iKC4TB+X1SU
Qkhy3Vusa1p3GqrzOCx5ofAB7WxfpDDtbAeNO1u6x72XLzzuVyFqn/MnLD55mWg/dGO6ty+HNLvJ
kNv4pyF2tfkMgb4V8e6lj+53634d1tVDW3ZPE/qwfljEdGlw/l0y2zpDbdhSyVI/Z30hwgpFHj2N
ZXEpjlKj2UzbIInX1B1RWGiS2auaEKzewDihakhGqev9ODoOYzKAyU/onz88qs5XdhwZ3Ex+7NqX
C3CivJIkrTGucW5IPKLaHAocvh7cNlrsA1j0uaPN7oGsvL+3TlbxMLJ+eRxDkRsYN2Asu4EzpljW
fQjIfvk0bQj+ykhxjh4NzTkaKN5eYtbzLgajgcoLJLI8FpO6j5K4zRalsldHzQeiWoAwaV44PQCI
WPuIqn8Uo3NJQ8miNE7d/nP+jSUywPcuBY+U+P5BjWGGEUy6b7OTN5VI39kW7QG/6DqXOAZ6NDYW
rTnGuA4y1Mw6xhGFGZKivkR+qbDNThFPDkl4n8mtlMgu6HWT9ZAv5A+l+HK8czTgm7snGTBJ+cLp
wfVvcA8cWHCoqhE97/sJr4JmFIT1e94vxJh47e/ijdVepc3+oRUw0LmyWVVMmeug1OP+VYIry7lO
GzVu/RPj5hKox5rhXOk5G6wsesfW855d53lffhY1Fi9D34RlhcbhZq72v+oRf9KbhdYTLoDuhdN4
+fEMX+aYcG8fGW49cuDCl774GHVegYn/trBcpXiEMj0FhzIWTMY6b9iilMVIlukVe/UlDTcfEAa6
PmK9pNRZM1l/mi6gEfYhSG2BcET4RQmvUEMiF7YYFFghD5lKJvVP1yuJRTvxmi1l5hcUxUyQYyS2
5ppAgTE+wAUsMMr8JqUVoJ/XBCyo2dJGY7Y8bcMqrzctEs2Q5cMuJJImef5p2eCk6WSb78lKc8eO
kNFRc2cP4mjk4jRINj19jV1YlsECJnHKlxqki3TO4SVmhSKxUz1BimxpLga5RX/ulqptaQfswBZK
0+JMiFuKWC3acD1mTUCckdLTcigNsoYoD5eJuo8sZefItBc+PIsVazMQxm/pFwSHw5tKH9mDMdvK
a7HtSEdj9kP+WVbrmvEr7NCwOOfEBndz5DVmLsaz9o1y/anbTJd27aJiKlTTNbR1E8xd5p48BiLm
KqgjOjvuTBvSILE2R2H/tYe6KdbY4arJbZWhaf4Tzn+5s1okxCGOAiQgz+pN3zn5aQJEa36GBc1b
HRnRlovxL6twnxZ9dGF52bz22EcSWlYZ068hEcjOSHTvngoZKyI5kFsgkKAz9s1poDijhcOmpWtq
zwGprRHsyGWIyC90GV3WxZROhOlh32LjvqxYhJ6FMIovHMlxbscXKbEcPfxKC050uCDiYEpCZydx
cGxG6Hc/owaqqjZ8vnJX2wqkvsgjRqa/uPJgpig9oT7zCK7EnYf3tXzyhK1nHb6zpVGSG6XmFseW
5dlAwCSJptHyC1mBPuqPdNscqZzB+MDZoLeQ3EXja9NRNXp1mxCaELFAqbrfIAor1BV063iR3u8I
wJlAeldB55uuvodc/rVfuLLbIuxfkKAjPpHSJFejXe+gA5wzlcWcySSy0qOE60rRveogp4mQtTIN
MpoBSQHTIioSBF3swaIyrO8kyIJBXGvIPlNEiRu2DIhCcktRgtAC7NQClpeJj4Jf6LzohXEPUNEL
f5PzBTEnDiapX7I+CdF9HNbhclblm8O9afna5Sp5QyQMpLP1G70ph0VREWDuaAArF23Vh5RLk3sV
WzTAk/ekS0uMkrHp4A+p2ZqMPh96StIWBLkWvsrXrslKPOeg4iNhEyZsrBD1puQ7sPh2i3uA0kWu
piF9hS9eK79GZjRXbXjTxn7zedsmKdDzc2LiLXO/hZtYVHULVBr2fFMphVugcKMmLpA48l2GI0fi
JFRfrEi+CgIDUTxBXeTZHYLswA6Nk3BXjx53t+UHUZT5nFqeA6Lz02VrwuiJyscDmiz/WJl4qT9j
D+lKsXD8tuwQwfvzEO026F+hgTkEok8bg2ZwlS3tWuLmTsldGHwTe3HAK+/NjlotrmCAWb0up8ps
d0t/YJ0ZsJBxH7pDNWQj25v7Aq/1SPnN/4woP1MfqZ02RxBlsZuSV19NncLHBIEfVf8ewPiWlrUc
jCWB4CqMtHESU0Y49NTe3UCTTgSGBQ6cJikZIHWvwf65rWkmFLs1OQrGXlgI3Eea2ZJP0cU5YtGt
YZ6ejmw9bze6ahZ99l5U87xINXDBUP8fvQtTFMcSK3n1HyhuGYMbcT5G1Qtx48s9I1dKGsqlqU/+
Ttmcb0db75YECdNjcmx8jMOTLzRkvR4Fj/O+Z2CwXfTsLgMQ+2Im+FCQQHgmO4KgLWN7Qjj8gXF2
F76TUXFC7gWDZgW47tKmigtZZlGk3qS8/c7qc6wn89VIiE9Ix/nzOASuGICxAIzyCAHSJsHr3XnW
x2sznUscRmuASs5r974/Pgnnx6m1VMEJknsZeSgQ2vD7YvVzwtdWQIXLJmhSc5B3RLDwt0/3F1pX
QEfQRXPqWHhYjTN+vJw88bvcd4nItSS/UHcoNWNmjokqF1laXvUOAC8iBYEJP/LLcWFCvZDviFL2
jMhPG9EQN48s8SPWPL5tCXO7pCGS5l0Lx1iEC9cdItRmed/5+Cx1rkwl2Nfk1M+dzT27QHf2Epjk
DlxEcwNl4A/GiweoHpJwaLVVVj1lSYGzHtihvWWSvYh/X1sNsHwj/JB+WQfs+91TaWiEPre4/0C4
twe5+7qTO/yNGPduEuOmdf/jtmE0ubIz/W/B4DP+fPcVovr4zFgwu50LM0X13cFpldRIp8jUZ3iM
1MIFLrGnztZAgk0yvK/+ePXuFalnavYbyYkxWuWLC2g6LR8NQWSBnPw5xnAlkKEXYuHprPdwxnwD
Q/8I5uNIp21s3Dwu/w41k0pagqbNjCcoMFfwhuSYnRk4ti9EoixCO/NAUiMsJA89pViHPeCE9EfN
mZ2C0NK57LqCwiWKUuZh6WVtONr4f5eD6oFLLNpVcAbfysjr/MC69Xg//oJy03e8/OGG8qNlut/z
soZOSaEBj+GqHvdRNELL/GM2uDusO6suV/vuAX0ANo/kw1ukPlCdAqzIOEnO1VEUA9w5mKEyMIWY
BZY/rAygGhp9S9m6Xg/cWhAM+5d7xngWeUKYQsR/XepYQHXdl+iefskK7475KG+iLtwC8PAeMrho
Iuon78/dIfJg5vSdcS/RWPX75XdFgPub3hEyHyWBgJhiDcdR8jOWkQN19i8hNKwlDAMUpGEedjSn
ubz9V0+ppPpl4pQ24aVr2V5HjHONPOv5Vy3Ys3IVAH/Qban2Dv5q1EeQ8vLxABRCcjrMu5LcVIKD
wYtMQfPI9DivBYlmFz6AjXh1dNP7JVF1EQp5/jP4gnQQMaG4bQ59QyaXfBE5ye2sOcnbKD/esMy2
aUhBUBvo0Y7BfYiqtuxP7zajDNUVjhyZrK5wE3Z/gkMw5lrDfQbkidUEMRZWNIdD01ROo5VWEN8c
8yNA/dKqaKW+gNuGq4bcT4kqdEKvikC0E6mwJ4U6nEMmFkPGK5WvVq1mBcbKUM32xPEXXJLJ0eZw
cRabVIeGopcQDZ55Ub4TZ/rppZFiIJ1T9gcJEWUcnaYewF3CQzPGucLDVbjqwXmN2SgdfEYY8FTY
DpuGyuG1qIiXTfIbS1kVkTQkHRYjXfPKYYck1/EIeYFWp0bwE2ZSqfBCdN6CRGiPBdDG/faz0P4U
SfgVtKnxpAndfP3z3SMM0aP8Kswjzl7WlPeGdGnar/RtE1BewtRs2NDoRFybMwtI1JsZ5Fb2mpry
4HFMwwgP2gTv626ZQoSv/0sr9YprRAu0nwD7FV99wHWqiCj4zKTxHlPB9mSjYWHtdbZASFTXtELD
QEuQPbWNKkGTVpw/ucBlClkHnaUcQV36t3xqtjWYPu9lpIATH19RNMS7WMc3HdlzG40EwB23Zwho
FuLxiDMuT9flWl2mSQydF0Yy0Ls+jD1EuzoLrbY63qBpxtUCEGGivRZ0ODShTIR5xGP3FQ/NPa+i
Hy0jzyJEyEKbca8XsmPwWMpB6YQF1MQU74mwtnFWm2vilo00PB6vRB6pLeW1x/4s0LUkiSoNIWk4
MrW3kOTSLBORaOOeSY3+AeU/ugDUbFsE0DsHDu71G+8ZXQPHzMu/xo/WaGgKnnP/pacBocOX0ZNK
O2x55WZcF184ZxnRuy/dNN3DyaSt6KvuyYvXOFiml2umgsdwYpmPsN+lu0VflunPrdAC2JiD8ZxO
FMN8I1lERrYJ/0VHT0sAf4FRMc3nrLKUu66f+ZR+OG9YqC6lK+Cnhr+BMCC6USHDHWioYe0Dr99G
a6ZGbqj1ejy7ICAcISTKTo/1JOP9faX/p5QGLhpM8ehsZcmwF1nMHkuC7WOefPljNkbGKz5MeZh9
T9MlZBceHtBWSb2taAMde1PsReMkkGVw+RqT3kYK7GB+XEmiRU2RVoZYxJdj2Ee6PdiA64RXZqE3
czcDYmEnvd5k1mplMOTeoubAROZfbyIwSRzhlFZeDXfwXwZ4QjsXCTES64wFudq7tQFGjkQ2F92G
GterRYrdwT+wIvo2DH6D0S/a1YXGDCHEEFxrDOapeaEfgHakSKxUSFOMkxeb/NEEvZOew4s+vHH4
lNbD1BKxV97/nFJrbn+qfB4AAZzOWd+2su3UE3OjGsfDy95FoFTF0ktpNxacgAyNx/MPgyDfRD4l
zPQ59ZGOzd9smFLMPYkXvEJr0Qd9uSSSIjTsdBFAaK3hOQxOG9LOeULvZY6BnrnV6idWHuUYbWE9
uWerwcvwkTJBDxT5eUlX4PL7aDsxNSRkcl3FaKyKg2A8UEV6QnVS3rO+pgPXb56FTSCxPJgQgJr3
uM3FN7qbkoLictUnXIR3XYXw/Ea4JrCyLF7YtsulQ8kYjA1/JD/BRv1Mv1Bxk9ymgsJVHFxs7vDs
NtxDWS5hl7uZtJpa6/9OZC/uyiDkp7/+PKN8pt0f8Y7nxE43BVb593vithKWGyKLptvaMvSJ8x5D
bn1W+TRKKfKLKGUP+O/xs14D37awYKQ4FYiTDtLrJJCBRzKM4+81+WbKTSzWcgGE/O4gcT36wcPA
Yj2n/CgIxwVfqjcIGTPWHtQ4mofLERRLXpDuv27JRNBJSljt8VOIWh5cs3eDpbJ1NZy/96g4m10h
KVWsSGX+t9tsNQy+uw2etYO7e+8Aja/JCPca7TAJm3K/rVsaHEkrYPzp1vYNPpul4lJiPx+KcvYp
ric2JTFyiThuFMt67bsM4GM0+OBMsM+xlG7sygAOcpc1P149USmtNyp9WJHqtDNNNfBcgkp611Q1
VoYPwD2YpfbsKBLW7iOBHUZGvnbeUKpkn0ipCrRXL9OlUI0OGlktInZHWzj1uSwp/3kZWtgDtl0M
Eg99+VXf15I03rTQVMXgABzVfJ5gLa8+HJ+cvdVTaFf9ZgslYSgnt4/tPia0wHJBoZ/3xVcIx4eR
/leR1ubKvcsKNkiTqBVWJ3PZdnDPbyoNeiaSPs6MtcuWv60ic2UJxXeS9HtlfDPJf9U8X6iOeVW+
VUQXY2gKe7YcGV9Cwea7wkz9ulJqtNJk6vZh579kAPafj7R6sTuBiU+VyTLTjTmhaSD2Pg7q2mX/
WSHSo4OMz/sRXIxLMGCMJ6DvbkgQIdWmlAGiXt0lA1ZjEnLyxQyLUHi6na9IBvICaQxNjML5hn8b
EpsEBk+qgq7Ky20DRHv4prkyYIK7xfELGNGvAQghJGOi58CK9A4/LsC2ZRnpPsT/XwlycmVCUjQi
Nd6PWvxM+3qTQLmGdBQ9mx23VUUK1ysJHXjLT8chr7rDxuSI4o61hq/T3KAEsQBsbaLxZtDsPDf+
kyOUYalkIKMkWaYYB0jdAnt4CZMAMEHpZEVTWjWee3pzX6CW4fNGm9KXvOnV49nEVKnJRn46NmeO
utaoEj2yopet3yPHg6TE2xhxwCEVyus3bCFwhhDOGuRjw2HNnTewC80CUzncNfVALwkOKgSWqM+Y
0B7rUKMAXqNl9ZmjqEYOzcENOP1RqD9eXbHfP0RVZAyJc3sleGFZi2oh2RyeZRiqCFXnzPXRtF5y
34hFW0qo2D6Z2CB3TMeXYDJhQ5vcjqQ+HSrsxQCFeGh7YAlbzoUy+NJFjGw+MkAOop3fgtXaDSYg
v/y6gcGWb+q/KOgxFo8TN/xYzC3whUEutIvcKdIih3WiJpJb6EJW/wj86eWQeYy9W+ReASoBOY6w
AZcrp4YmHeWEnCHsTxWwVkhx+AousHg21K8qY5eS5cZhl5wGErjqnwGb0DcBi5SII7iuc6FM6mOP
mCTrbEeBvNR52t7kBJBJHzi429E4QsoweKIhXbnedrj/y7FJTIJQ8CjNnZe033yx0bmoBVdX7q3j
s8ueXNarguR3HCrzLobPR3hzgbYnje+I5FTTz0MiZ4iXyMlpdO1uT2UoAEP1VuEhnw4kVOoLMu8d
vggwyY+rR0ptzG9WEigyKNXc7NlhoiGgW//ob6WRxJu+b9Rv8KQe9vzKsy823iLgLChvLIw616vt
Ts3xtYg/naZVSNX4H6j/DVVGDXf9TSqOtAVGeAEth/EjEC59cpNGtaIaxe4IzGoWSk0lD+9tU4Ng
BI2zmNLIrz5I78goFYSGdHCvWDTqJJZvkGTNkambA6ag2W6+w3P9qALR0OmIe+QEGD0n0whgiI7N
Nrd4EuaGX4fWggcE/74ByqQRrxjt25adOiAfwUV0saAhdSztG3nHzNd9TTPHKC75O/rwFT6osJ1+
FNV4LM3NBVZak0to1Ax2vHQ6tivy/wb/nAgyBblSa5uKODK617DMPrbTeMDHWo2JMDcp9ndRFJEc
eWQEXIJR9HnPzSx2eFgUiaUvhmTVRdaHrzFbmilXJqKPL8elsK85TdzF6mxj6Es0eYedqlZoJjqW
jPElrMBH/b7BlbbNPVG24ba5jqNAdvVde/PkzDsVTNpyKgokztVyn3ts+zNC7eqY3xAineUbIYaC
rIsrpeKEnrlfxb5YtduP19KGCtrVyjbhXnjeMvPh8U68xu+kcESujfnglgoP9NJaYaDOxk6iFOGE
NNU2EbJtL0C2Q52LxFTu2XHcsSb05a9qNUzlk8gNYUHUsCiHXTWOhb2KaNYdE/yGyLdu6Nb6jfy1
cR5wnciVYhhSwBNiA4arbDKkrNyvOxWscH/ws4pu498A6SJrjVAICd3jeJ6c5xf1eC/m+OkLcYEb
cJekokwn82o7x+aeUPDy17QNaWEHDfAGygdnp4LRfRU5p8DSsejXH9UCU5UPlqoY9oFzmlIAVc8I
NNyiHDDbiHUSEwgRO9ySR6xzkzb9IOpQopif0gQ9DuSmPuoH4BNyYu3tpuRi5x5TDWk4NmnlPbKB
7q3ByDr7vlMlZtKgZzJh+QTP8VANk7hDcdPzKxhWR7WGrUViy0AOo/sYDJBimrP4Dzjy0A9qkSXS
6rtxa4MfHy0XL1/v2HLBROFth7ExQjpOl0EM0wICw+ML65WVkCBqXUwmOIIuh5OnZ4MoDpqz0TmM
EmA3IYEe8YF7D0QMHlcZnIOr0cEoAp2uR78ab8puiYS5Gi6rIe3Qk7N51tMRnLPnUY3gx0pav9GX
lwkpl7ciN0lO9k6Mlog9iIWXleCQXIv9jIKaPRzrg3Q+LO8fVpJFK/9FqyEugqUZRAifIsxRaweM
FHyjwfIc5mBdFQFvjbNOlLKzvmgvvdvutFTQe0g6NVtHK7DonPuKWUtEvSdcBt76d4gYCRo3yfqL
D4fIgehFMUI6c0aS90xL+MQ0Qs2HNzr4Se6FECo18nzQrxZY/CMf79f0z7W2KGj9tkC4z0+20rPD
5lLUBr7XdBZHVS0k1ZS+0VZ/acA0DlBwIb96nfnSurxg6EOU4MN7UGYc0BstpQvV0KFcHCc0MJ3r
u8+p/LJ0okguUxzYaPtBWEuRslM1FcIPDRF3E3UFr5N1juMCjlrf/ApKTSyLabLlkEMVMl6RomcP
tJG0InUXhZQcCVoqkG50dywLK68+j3GXplbA41hR+ABTyWyi4ZB+yfXhzy8YjYYT/AjIZn14BGgS
fV8NV02QudTNB/ouG7PJQOeW3j7F5E3YemprFR1ufdz3kBIgIiDwilzp7tgBsEV68qEbwpkhSASw
2EL5tp4iqcu8Ia8m9ZzrEyCldFLwbeYqdylxVutaIP0g1Q9wGO5oAuz93wxvun4tty2Mo+q+EMlU
WqJjOGnFwsZKNSt6wI07UdluEX6KxG7RSXO4q9ATCPhdVmSF3niCN3hUXkeg/7xWJ/LM9eby8wWa
mxKQUgkUkmkVNBLPHWOGNxA7y25MpvuucAjdiAeaZKSefhBl3B7vncj3t2PMd6m6HG7a0emVbgr4
r6xHwwvuX7CLLLNRQxmyFdM7ghf7MG2aQi5jcl/kLnnXK/ByT0N5ELLLtwkWzBtajOeclGmUk1D+
P/I6Cs/v19kQgGV8qc76fQjY/jsKTkXttuM9O/BE+kX4nQFTryV8RpqSMVloQNDAaGEqBL/SoC+D
Vcgtf4C4Mc83hU5mMo9q9KpeOaKR6IQ1uk5gCQ0kb44tcGgd4QZypOPilvYvTcUYWOfMm4Ve8aPK
JcETrQibPgUUXRSrOc9sY1Q6LgHb1v/El67DDifY60f5Qn4nKl4mxtpVBweCto9Js341ix8P+s55
14ZKVIhXniWwHeh/QNiZ1RmyryhYrb3m25Tfm22vFiwtB9PKNMXC28J4mEXb/lJ7dKy8WN8oGVV4
0CWsPgiTBGwCcw1LJPAe/3uGf8EILo0iuazrbsGcDdajyyrmenncr/fvA4JwO+Zxfy//K3+3Fxwv
d/Q0G9djgDioCSt4OY1HcZ0jlwhIS1KVK1sGKuLoBiLbypRSniClFb/o1+gqnJeN+deivhneIrt4
nWixsXqhB1p5n+0Jiik1Zzp9js22hzCV8bVW7NE92488IDRbMVF7vqkO2qmtjhgv4udeoIfX3ohU
5JvhbFiaXMlcY3mzUBuKv6vk5sn/o3ZQVxXi6azgoiuteUgdK2dLDcwk7nynDPrUjU072i9ceiC1
EnjiQhTf1ZuL+aB1XrVttOjhH0YA+RycqQ4r5XjZTKR7cDgRGzL2rOdz5UiL/TwDqL5p1oa5fdcq
Pp/Tfkh5EGhq95HFa8BFWYyP4Tf2d4zy21p2Pn9KWseHVE3otbM4ir5ME2lwvRPAzwCo19i7Jj8K
FsW1f9Y8TPJczedwZ0r+4newaaRkJECcFVK0yl9VerpiNcWC5Dq6uEhDGVzB+0ekJ16BY2mR3xyB
zKJC4jpOLX8AMZ7s/7er60s3SLspL/X4e3qDHSoHIvX53noLxW5YzUY0DYb6sklSjwnL8C7Z+FUo
a56vtmehXwRSQL3et2tr2vUWCVkfws9ybApPLq4QszxLalNxZWeJoN0QJKPNORd02UeoJxkcugz+
K1UVINAMCbjQ14L6KEzdn2caA9sFcvsVBfL9vnzSwVMWkWA+YdHeKzxmXDz+yREH9NY+JVR/XPfC
Y28aG0bDf5dza7e/0r8tRDZpL2+3+A9qUscv6QNkfj3dx3RD3V5xcN+geL8Za1Pzsost10zIobQ3
+RBWYlZZV+P5PP5y5Gkryigcg5D2GOrrkzFeLfw5LV1lKlpTgqgeJb8AVNn0W/5pyIuxgOPLuZtz
NFOEFCFX31S33Bthhm158NeH3rtdOn5PEIJfCB5YpYI/KZ5YHizuVoHNSoxipgPiT4Fi7zwpP88u
ZcNGkJvz1aclBuqsYl1rsU1Er4APIiICEBhp/7iLwvajsGm+YYW6CJFcqkC2kB97kZJAnY9hUErk
aeZLLtFE1vEoRQv+bwnYc4EmHvcABuBvpsmttn6fhzHo6jINDPsnUYM5HUQPWZp1S3VitZQWQsIn
dHyDqoDt0Zv4De36IN6fDbrsrrPmtBvLy33/lt7H67LJUIddRkna0UmwwSwL/JpbMC5vhGWy/NZ2
NrYjjGvcz/fETGRXu9gPi32soupRZprtTNGeyAV1bsXK12KgIuqxZ62/gOx0MFOO3gcZaySDORTP
IY4e626ptEquxalGsdeP+oPYfHrO5Tt12Fd5HKoeQoUEi5vL4WY5fx2N95zpSuFWCMLQ7m82rSVg
10/1CZccghb7pyYqGH7Gc8XPuvZHV5UgkfuxYmuwAmvqJmcKvNlQolpeBBJbzgcnGXJEiFliEHMI
+jOAgP+T7T/h4LjzOtCZwLLinfW0Y2Wm+SsO9W9aD/QBHgfNRy8Z11Fw0n2aaHjp1z89Qh0M/0Bb
M57FDej+2Ax9/doKQzVyb5nz428aQosTRqSGy/LcaUmxALGfTfab8VrYAr4lbs2T4WHk755fKkA3
qbwLekrAT5RxiXlx99ozIdlEKOmKCp9D7bskCfscuURvbur/yXwtYAlBwGEJZtLjiA7B+eJj6AtX
XMV7Q3LNkBjh7esyDNHK4BQ9IFeCj9ND5NV3gWCGuFdPHA41Otja5W7v172CFguiOnGqoWUolKsB
V6CV3ZLK6rkQruBSeJlLJDodDufA6+LoBVjd/EzQktzrebk8oH4f/Oy9emBlo/mdB8WMtLfziIy7
SJGHRlUbvSqMo4ZPHTeLW8LX6RsXNO4hdfkxBlQ4kG+2ULHyG7h5RYGVM66o8RTbDJ/ltzlaTh92
6hGRVdNRJb2L2hJ/nLB5aAoztYyGRqGJUWsfKABF7OHnvdA6nQPuJSquqILTSBcCCsohb1Du6ewQ
FpW+1jL9zpOdLwi10UDs35acpcY3gHiEClyOv/sejhMNexNwdB3Wp0O8GfRG/4+AYVRNZZASjFj9
N7WxBgiOt08fVz7dPFst2rncoUtHDyMVK3Urt2k4zDuU5TluM9tTpQzK4lL0saUeYReQD6qZ4Zpw
Q7WBXsOZ+MrLCsS9Ji+3YaAlYN1ojkzpoblXcE/Gf2lki92gb/2eKorMGrYOKG7qXJ1Pr8DUAr9s
7TeFxE5E7pxIXiej0N4iBEmgCiqHWiaVDJEAuvLZVrDkbrNisiJEa70w9YlOWdZfYMwWplHxkXtj
Z6ZkJiDoKPpU87IaggaQ3VTUm/woZP3A7AseWIQKFvoEQNetJ5s4GPZotVmHKlEg1jx+1+Le+H3T
LDUNVMq9eomRUZq45hhTXQaVT6zxLhvbTZ7QeBT5xZuV2uZwNHgnk45eXavMeVgxXJYaViRmKB1T
0kwriz2/25sdouQsQ7LvO3jM2UHlzkV/el/RlmfugrX19WZZxCsGEnTAjxifXV65n6gn7o7w1z0U
E+tAgnfBP/Mmom/xM2AEZIgz+JnyKWFtkyGkRrGIm6ndED9iMrBjQnfgDT7D1lDRWZ8wDXd4xIDQ
js1Ekw4oFrewmaZJy9OS+Hwt2G318C8RbpbvTzKD8llcajGkTCGAG9pLv0P3QbrM0qikdIldouRt
GkCkvGnSChfRE6NRyVhapdEfgopq0xtuEmYmAK06RLkBWT43RnRWC34mQxXuLBi6Gu6vMwQfSC/d
oBK27NlhmfJ7yFwEGpaxoiRqge/+3xgqifF3K9PTzcXfOFwopMZFPJRD5OamFGnS7BedmY8rYKe0
YJ/1uUplIwaddRiALQVAFUlLFXaGJ/uH8S4jygWbmnfzHBzoHmUk3XsNoQaw777/hx43uzGRXgUN
0DG84avf62NMtsyhsVPt0Jf+ldHymDILz/UlMT/G561EK67DF81ACkd7RtOREYdG8HcVHgSL2GZV
p9EgJg0m/E4v2mQc2wvjbVubjr1o0eCjzv9Pqm6HeglVgcwbOLeuxbEUXmdhS84uOYZQwA94k4de
g8cGYVKy+DOtee1fhfoDFVnmrHajK1/MSD8phzy5ka0C4zMi9NWQ7u3srd846FjVkgDnsaMES3iF
1Ix+H/CSlRp/M5wGNsrlliZpBVBqNW15j8GtTglGYs39XlHmeumjHeXbX40jO9ocpOAMKq6nPStS
JoxanNYJwVc41sbfbJjLwWqLYGnnL8gkps28WTqFNiW+sCqQZ9kVQowFXJ9I2tzCwyrPWfdDE+e4
vk2hN57816uO7aDJZdllpmGrtSvLdb8kjTNz5/pKxnAlQqeWelmhJBTUfK6l3eNUQGPXr0BDIqnP
CtXaKPF9nbUnl9a9kwRpswavGxJtsMwTRgE3IgCz5mMNGGM1cQVhaXR80vvSzsJA8MomBVKWaqCa
RRhH8krs5oHFe61n1TEn1zP93EsnIK9gxh/gPrsggjDLr4dWSkrsheq+IwyrGwUrw2exVK5jnd1Y
c54huPtoKbBvsBjnZoD3dbErw+JSZ98H7rZ+1xQG85zasbSDYfOdz4tURM9WN3rFb5Rr8fX8aK89
iJN0leuJD69wNqfumL3aISi+pZVxtETONHfu8PyhPI+b12epkY63be+iZV4KaBe5NDP/GDFJbglv
M1yv80tO22Vkq5iq0qcFPpZ3xc0Ak/IiKwhM3rV4ohCNHIYswg2rpIO9X2bIiZ1raSWEa20j9xez
qsyIUcVAtoXybL4RCDEwPBBkSbmOSB7qjL10r0vu7QO8PM76Y8PLtd7evl+JlFgEXOz1VlOtal0B
cuqWZpFEsBSXKIkCUrjzQAV6wianUsn+BiwUE44LE9zp3FfiP7Bs3MZLtiPccR9FGmwMD3N6zENi
3mc5kyEZ+rPRH8P4gjxVRk4mTkoMQLlK9t4ni7CGBdwnGqSyIIq/nZ7xngrOOpdpmO/8VbClY/s8
RZ2CDkcjaxet2Wjf9voR4CFS1lHgPKs/r95rX5jXdkZunKIqYwJxfoRH+hGj2HJRDjGLvFwDZIMA
K4CjeZpvcNl7HMpopgtNFasGL4LwyBbNGN5Z0kKP7togm628KgsaGEdUrFXkfBQGd8hCJuzjGDhU
jjosMW7B0dqqc5SsUfqanfWdR6Z9JPGe7rDqTfGWp7WU22rEAJlmnGZGSls3brkE0AbUAW/DRsk0
xXUaQC9clepGk3AuhSrmErx0TXP9T4Wz34fExsU00O8tMw+r3FA4oJDovZ/MAa4NAu53szCTyk7c
EYmUOLPZHmEnmtGMqD2yclLp2kbU6YaIA/jLsjc6GyTMH9gyoaTN2SD+aEkP0F8lX5SHZnxEKv3v
vNd5peSQNosg60e2IlHxWfATS9KqxgOc9DQXoaqqrO1KfERhILQFDXnDh1vEe4EQ6b8jR0Y+CfYp
BkLDVPOEMKpNRgh81uxY0AX7neoY+iFm4d5oQDFVLJc9j0TnVPVkEw7wp3YDLan1fFSoRiiySWsk
oz6+zVZXi7Y5uHnX6KBqtARwpHhJf+mhuTSFwSrnquh1uOXLWsHQSbeVaZCJUW3/0gxgvvCzDE3h
jVnyF1xN8L+f43K7KkhNGmsxE2tw0jzhTFgUKNulrsHRggUzW47XzicTrL3r4i2B/fxO8Rd7Jk0h
99C1Ti4jLGfgY6WLBGD/K8LAcyJLhPjPHGjQxjTepdbcNxOJxq+5qeBi8b1BjQzHzwbwvP7dLD6b
niixrt7upUafSGUYT3Tz7IGhx0A6VTkEs3us2hMRuNSGLaX+oDgasjm8yBgocfEFHZ64vXxedmei
reK585sCVgKEP/jj/EP4Tsek/FQBtV6qwYwnk8fDXoSakoV4TJJGyB8RK23XwgP/SASpn/m6zRHW
VYDwUZpe8nt5wFFCP/qy2MmCnr5qnU2oeFyVK0h44ruaAN3JO2zC4SlozV3GrkeIXPim1L94jfcY
MatFR06dWW5Ja2MaArFXTupAeLvAG8JSacJxBakTLvXl+GgHIIxCy6fBB1VuboqAIwm8FMaTT9cp
fXVUX0Ggr7zWEHwBeTZ/WPzXSw4HaIVCiTg6Q3QGK5merr9Inj2s5AI1ksdWfcEBfj9I89c7J1Mv
SlBUwG665EeJCOxg/veU1iv99/nETQUi7MLPFp5Pvj4X3T4WBLDXAwls+HIFkP8Z7E3VkY+Pd6By
/Df2ed9ihXx9Ig7FNtUiSt8r8olnjYIW7EEzAfXbpiHCAWuMveXpLAkorgL8dHzXAohmD7YpHqx9
kFopJTn7EhRHIwpBta8EBq38x5b5+6GySCAXlyf6swhIzm1SBJ6qlRPvt3wdOI1JD+wHkep32JAP
YnBmm20IOR6Dh3Njnral7Uttn6eH213p/SoNuqIiVbVIR5/dDuHrGcmH5wVauFKKphGu8h/CYLm1
83lrA6ES+XiftVlEUEb8qyd5cMKC82U93JPOcXQQW57dmOpYPZ3NJ2eXu9Qa0fIMDPQBlYpGaO9b
B3OTpQwEb4LfW9u6AJaKbi6Rg+8c+KvIKF33n2QI06XZCkA2IbNgA3xzF5VAApnnd7WY2WfSMmJa
24pAmSaE4LA2p9febKgBke6kZm6ujlPml85i9uXf5zRxe1FJ3nKKYtCWyCtxMnZaKi1WFOJ9btHm
caMgjPgBZRXmEKc3qX2uapdzGVDKKTHdPmv7tLnekrl2LUOiUgCPPlK78KjTJI7/Vvi4eXwePTiI
mFqo/c1mq9+Xh4KworMclUACApQHlQg8sloBhzsdQBmkIYfEjkWqZqe3t52bvUvWgnZ7JU3xSarJ
61Em+hnMkLRj2RBPt749Y2A+q/gxZzu1GlaKY6atx189Ee865VejjOuTr3U9zssonFBcZn+c0uIg
AFoTudwY3QVDc3d2mMd0T080FuRPjkPFPyQLyCo5U6/Hy2M+Iou8fJdkN7cdx5Di89UBrzdM2LL7
GEOzYIXJ1S5zwirwDLBvZPr0rNwW3d00OpRFzuq32sxBQMP/GvBUIW198r0xYjPS8l+OF+kYNxbJ
e2sfZcdhStY8LYZgwbhwmPiHtOAcEapvJ9eKAvVjXj90sQAUj1SuCT3kN4igcllJCrFlQ25MafG9
/bfnz/m3hBwaO8ds8wXj+6EdIesHpg2dqTy5LWD6wHGmsn4daJPr4m40BPJNDLYRTfRnqfEd4Llf
Rk8S5ALrCnoVEOkrulGKQ+DPLHk8FmUD1EFzgmiM6Gx8cio9XFGAajAEwKGU8rMQoZejEoPnMBT+
isX9unAR3TyLQqVdN4ezgASVyEGRN2cRn1YrP9fdJ3l5bcO+24Wdm3ixP1rQkJQo6O1WtTIlpDAC
qlBfkjVP6mN0NSUoqNfBaQwmVg/j1otCBHZE/WZr0vOyabwCdmXRLjF9yhZldfDxU7xRFXad2R2V
SkE9UHiFB2YmWdETL4wJSZH/90w8K5vfkzNDcDa612cgYK6nfWZ7R6IlSGEmSMKeIDo2K92xuerC
lOh62HvvLKJka8zuIbh6+nbJDa+GK2W5BY7WUXBof9Y96ZlcxAjgtVyHVublX0p9pRWUeS8Cgsu+
Be9WwEEVJuMRrowMxW/qruLarP38SgHEVGt29dz9NS4vI/xdUIsPnTSKA6nm5pq7tZh7sI2Ub5ya
KTb6FzQdQG9PCCU51JiXdxQ3dHCx8NOAK0KDFJ1JKnLWOF4GPXRFcuVDAupnFGW3RCGoHXOTcJjJ
S6a1jgHuS+bbgtxs0++s8utFWkIhXPDCEOwHP+ABvLHJrG6DgZkH1mfNt938fIuTeK4iIu9qzxm0
5WVxVUcgQqHeqVcQwdPBsah1xXslqZ6sKBxuQpV8jgbnO7To516XwanXC7iS3vIIa49/HADrlaYN
eEsxY5xe5w1qUZnV47r7mQsiKZkteNuyzWsg0yS1gNUNL7UNlBC7hVx4o0RR1pjbN8gyU18H5oka
iYKOHyT/oiMd7apmblJSeYL0rQLHJhU1GkLHVIIygCOVZJ2NOuXxc9je6wdOoZ/XjlUvA//3xQvi
Q0FFZZd0YINO9oQXSxPGjFW43ZKB76G744Pu6h+xqle3RryGaD3hjdjuFHGHSu52xErAS0H9jO8f
HUDHjECVfgOjw9UWdqj0UIwJb/ztAmOq6siqqabHwTyj/oSXeaNQqYl37PgiVjP3yEqNqIab26tw
mcOWICg1pvCHJVQpnf19j8a0dFMrJLqVlwLp7TQ6Rgq4hE7k5+vTqIdALDDIXkvI6YKl2FrLEpwP
VGed6sWVfccQJoxzd+pR+DmmmT8hA21rkP/1HradsAbdyefvd/aRH149ToNE/nZeyoOqFHqlK4pD
JWKzfrnUfqNhoA5s/eLXzCWhTiegnYisIyJbMOvJii2qaGJpVQs/x4GvZJBqPbkUE0gMHNEhB6gz
IuhvMAlHIJooo/Xvq/VSHnlw9v5O6d0P/9C4soiwcEY8AsUOrhVaQ/QQBKGe5YLzPIJOKkKlDW6G
hSm7T/2khSxXH267zMfnnHX8TBgKtTWj2mUeuHxjx3pXHZ3EElbZfRLR0BzSAyf0ZqiGJSWJlOCR
3TJCWOkclVG0jtzYiqTqmzA9RHgL/zjdZBmP091ny784wwBnZi7AcSNMaqNcfz63FQTXUDXuF7gC
06b2bJ540jDkxXtmO1qIOppE7e04ZGsms0FD7oLks02PHoyzUMETMquneJOsDR8lts7bbuD56NW4
XmNrtxR3ps5bWT5FMG6grdWRjqWIY49c/BC5Bg8g+RpzNci0iR/chLyml5i/HjTfyXWRnX6pDeI+
u/lm4rs6kTtcOHqqWKvHYwdVL4cADKrW09imPhrJ3n9qY7AU6pXjYhilLNDMPOOKASgpXdKEdR4N
Wbf4hRzQWMrIjwd6Y86vfLTk2BiGkO1km/wu0YSX+tESGzehi2Jeg+Gl53lv40WISeGXDzb+wbhQ
eufoe+xbmJA8R3J5nwmU0XBFY+29U7UwbSsG6QKjLhS7DpHDXM0AamHhpPHS4LZ3030rD42p3FOt
3b4Nv6hQBPciSRhhp4UMU0TrRsuIHqgWIpBexB9UcctX/R1MlhnLJnDuk7Y+XQe4Ff9vmBu8e+LB
hcF5i5UcakHU2vM7stP3c4VT5q0oUJgZPpxiM36fKWlEAX4RXuLPr9KRuClsboi1+wprP9yIgibF
lUwOLjEfubb/KX7FsXP3GIRqvHcSRY1aE0HraPaT7UKkgVKlOEhNCXiQr7g26xhvG8PHLe4aC03W
is6xMPX5kFiKzaJoHaLZNvw+KFLIHJmJri302zl7fTP8YOaJWKs5i6MYELTduT70aVsqyhTtc3AO
VEGVINqL34luFiOhBja2c16NEic5pJWU+C5U4JfHTOmQo1XWohySENWtx0uA/Hq7m+DaebS5wNo6
Hicd6NJlSV27aS7g0BVJUI+8DtOvCBXBfNXPeogXwO14cSNXfia8d03eUAn+rb7QhiAWVnFq4xfE
q/VofTs0NwlJk4FayqvgrXksjKxHU0yR4v+0J06FuDcU0t7SrInlOe3xOhHoGTsUoLNus592enUD
ePhX4aBDkCXTbUHYCQSiLYGzBxgHubWP/gyRn33zH2HqXP4seW61XZMBQf+RA/z/q243cSDoWjZ0
PoZ6BhfMXL5HBglczEcGqrwILtJdz3OZCIa6J4t3pN73S4LsYQO9FIdGOnz4d3f1FGHf9jT8RYa3
732jOatdI0F2nB5812/8s78tejxgYTwGi8YAzn6QD80AoE+xlFYxpb9bbmprpGwryO0Q+MCk9iJP
I7KPKMmydib5iCaZeKaep5quBME0bngb2H7tHumitUOCu7vAr/iOsv3/unZA8zu1wy74eNho9Ji3
hfiR9wuIxkLN91GnkpbmeMG5z8jEBtFr7/LfXES8G0UIAeS0amE/dqpBYHn5hiChJsoTf8A38lg5
fx+GukoXNDjkZ893Fghz5WpGeNAKTnSV3i2RyG3elyk/uLb0WGxCn3XfFyQzqGfDPuMwlBbxy7h3
yLBJifhr7+GiFb9RUgHoRShHt/Tckn79BhpL5n0Cpgy5J9tLtxuf1HPs6C7QAuJsWYdqJbLTpGGj
WwuTlrrJrAAe3nLUNoZT+gESsBXoZVIcxvGA3joRohsWZ8iqKe8tIOQpcI1dLdCkxEqtypPIU/5e
WHCqqzx9kq+RCjZG3VyUbruI+5XWmUYi+i/McFpPTe5bJRBTSfjytGplREATVKTbUAeAeVOWhPZu
nBOYSRwhJP7ZJzPZ/IIPmR7Lze9YDEb7gxybOhT1le+NeZ9Xko10/pY9jYlQVdIPL0Hkoe5ROfZY
ZePuLkdF5JIqqA2SGcucWyJUCHxbBTh/fKYewll7FbqBK2rSGBB6TbsYTgZ8z+eyk1epD4mnlW0f
zaFgsNkFjlei86HI17DhduN8dp6bAjWMc7k8RuDYHpvChETWYkBborcrG9N427UQtNXJsnAFmqml
vq1ueyy8MaT3pYhKnPVTITqsIM/Pu3nDuq0skQBZAXW4Lb8Hji9COktISdzAIUDsu0eVd/gBrLAm
LnoaeFd8tbGCFMNjF+7cHnjYr/T/RbnwW+DtXDfInEQtZIuIQVSHShdDzF/OdYRX3KHbYj9nLxVD
LxyJDRndis6US5XjV2mLVNDfZPK+bdFeO7hZ8CP+M0SsNepOQeyHQRf4zabud8H8mCyEqN4UniVH
bfxhwvEPGCT+8oFxhfAYkVjwJ3puTMTSevjNabWE9Exv71J+A2sYPBlYAwRdju7fEeFzRuZsBFac
PSfiouhXHuyIQ3gSrIBFFwfNK7vSTIlBQW+BerkpYzzMuaqlg6pxr5MAgOXfeKlt293Gipb6fikx
eCDr90XHYMKsBB46X99z5sclJmJVr4RoZ42b7iKHSR+eleBHDwCHfQrMaHkVcWEenXlzcOOqHyFA
On+2k3MWspn4qRhmkPOIofJhY4idruwXwy6MUHiqZOrCr9Ox8K4gUJqIEbfHbuqJeE/MqxXseU3h
fwVJXj+sCYNxl/tuVbrXFGHvba5GqevDaNslg0JRnIwwL4QCc8+9WWW8eAUqxYqqdYfkxHY2iMBm
J42VE6mPbHj/ofc/bsIQ5yYEdo9LPNtBCFgTaCyyrMe+V0ttBBNetRApMkZPBd/H7e+XKhHvcpdF
V8sIYD5g7jo/UdKQAHmzzX+lrsi45ScTniTVOH6+ZHn1+kkXmocRGoYEdPO23TFEjQgjnEovpZ47
iKvPgkCyrbIVHcVFwMxHspyKzVrBwfXDJ8X+75l/8c8ex+1XzrIUdyfnZNGTRLABj62xlfeepecs
acJ0m6mU93j897Y/DVMNaUNTqhkUnCSlv5RyoMG/lYlTT9JLPxOxug+MWRSqGviXGpsp6/PrUVg1
OPv7Az20IJ/8DY5MgS99RN6pCLN0k4CwUK2Z7NoSMAypvLEOC6jD9Oisb5Dho/OtBonWvjfIr6a0
ahUrQb/G11H8OBcWNgbmDY5aQXWGFHeFiCe+TyndtAP8ODp73Ebqstv/xkWPn/d9sOBJOQskxzT0
vPv3ThpiHLReitcpI1txShtR1+o/c2vJsNM9e05YkaRyppltuqiFKJCQsJL1zuk9dup8uphSRerl
eH0ejEw1Hs5Mt6DLSB7EmBbByzVVP4qxXubVB7SWDvkbckv9h9jOZwLHXejZ/PAzbYxYomJHdsez
8eK2ptzrykzwdEhw4OzLf5e3KcuVUkj9l0B4D4kllcQe/DbZQyW7spiBtydBPgJCKzdkXcUgXzxb
CuMQBYzIgDyyauL6Vp5KHTj0H/N+a7kYhP69yfe38FZ26RuxksLjuCLzPXVmlWwJHuI5u6UJ24Xz
lAkAt/IIv7CStXKA4Kdqv1kwgH2zzNKSrl/A0aJMyY0IH05LbOqqmFvIJ+//c5K+bkudmSDQDY47
ejxgF9Ups/YXEHO3a58gujz8m5EEydDMXudVpZO3eWinxqM5N+PVwpG2dnkk6OvZjO/wAO3/6K0p
IwZBuD56IBQlr1iUaiHmQY01pTJKSkU0KeuVXfAIHM8sX2SD//wEKfyvoHksGau8IpgnLYXssx36
MfU9SeilS8a5F6h/sOdsgcTr9LzS9WKdHcoveO8rGkA4OO7vz5la/H7IarjdL6ZLCTBZ2mGkhC7F
i85yZgGBjwq9cF2FRqIgcPS+0lCz8NzEXkb02f1W3k9DLuaGBVfiA/O5pixaE9rCQZEPe9pvG/Rc
UWZ66bWH59b2gqXx9P1hJGt1uJNx6kv2FWMu6cjk4pMD8/7vXoWHFVQiq2tEcysUNwzlKnoB/gOf
h2N/UAQgFF5y+j7hYsFEZwVub+8+bvG0lvTQTnmr2BNfZqdxG/MK8+nVRDdPlR83tFKUsedpdr+E
Qov1sXvcbY2ObnlY7UlumBKmCcCsCigfwAMfYpvG4GWDK6wXit5EizdiWasKldHbczo3qH5pciED
APY+Iwoz4/u3mmE+E4kgG1SGHq2KhHsnTf4Y1U2RPiJ0mhM7XiCOqd6v10gHAYaAEitYLcpZW56r
D1T9jrsYkL3AFXWHTVniT8ZCa1o6GghHH4ZcqrYfiILkLW4moycCnuQnm92Gk7xOcwJoLXS/N0L8
5krz3BhBSZmC7LvSfGA0UgPksFQEkBXoONKF8r/CpOdia7A0OoqUuTKlI0ckTcMv2q4dh9ElEvHc
cToGhGoOulYyCXjLivoKSMlsj6Zs3bpUy0RvAApFYcfQLyIm3vAeS44TCHK1EskVAO4T/wRd1Rf1
Expoh4nfHORnNhhtZvGxKrUtfUWaU9oXwIZlpdc0QL4lzBZxx/rvy8e/AiwbU58YORp9h8kNHMQK
ypRQxNrciG5SwoHKMPEDj+Wr6pXdEFLKGErg4NNRBZqe64ms0b3d5FA1P+yN0xR+93MgGJbeAnut
xMzcis5ZuDTE+ZsOStyCt1lndqu4BqQsw+qgUB0J78DQz8xucsG6Yecyx67WrUpY0uiC1ChtI3W8
470N/gcG+I0sMHn1p8SaIcTdZhJyhUk4orMgLxKKm7IKhjUjPxCQXnPY855YVZgVQJ8FLyjZ7idN
Feu3iZY8SPRZn/71U+lTkZyWAxoe0Yu/CTp1aZzF1bASloi2jjt5h7s2Z6TdN65xgCja5SUfu7q1
xzXtr/KD0fhJtL7o9wJhlkkE07JwMkwThc24i10Ory3VoBzzilYhSnxa+GyU1r20BR6wnEA4tkIb
q7C7SpG8saossa9kc6BPn2l7eoOGqfXBwu0ymUrDfGP/lfjjDz/+MoTnfTgT6FCbHaEg33oljk3n
5HNVT52IiArAhqcXBVrNNLI9MXlru8/LATUI2cTZbf5GTOGAjnDEy2SQS8jHtGu9fJuN7NGzsKcu
s4uVsyYK6DytTkxpNOhPF31nQlxpR9qsQrhwQfWb7xM6h/pEBUmPnY9jSlBZ3meNVYU3rqzTGIcd
Hohd7dlxwF/ZSgvHKgYaz5m1IgBMMHpsvD79Y5pXJsMxMrapWG0D8g9bZpUzs9MiEGvTETpGR4IV
YMdNl1AsRt/zFrsaKaRt5qP83qIASTT7fWCTURC9tqqgdRIkmmHaMHyiLK8WoNCG38D1g/JxQRNR
1OA3rPe6txmS1Y/0ClXjwApa8IAulOYtmvumFXyHGCIDB/utUnSOCuRzfgbwv1J7syNcFb1+a9ZE
NU05B96QEJGH7xjLT/rbNW89506RUfjdyl47nf6259GWPezZ5zwCPVtrxuiG05ngvj0HKOIN4tIa
ruraYYUmuMF7NL1R/DsYe3Qf1ZHffajD+rKjP9O2LD9NRGhztyvbqQzQK6dl6lrVpzQ4QtLoEPQn
5r1zzy0DDoTBy6jU8yAadqJ3RcB2KGAJjftLqoQODk4vCsabqptsqk/ILUgpkqJPZHcesxyvDiql
BiD1OLDmRw6voS4gM0PEnq3bal5xi0FS6OZSMN3dLdRH8PSeFvI4KwfNZSGQ75KoOTIYp+mClsd2
nUwLAS21cr0y7oMF6rkvbpjrFStrnF7B5lOoQO22r2nKLn86y01jPcaTnqQ8v/h84iq77hoFfhaY
zdnm4WLBRIxmpv/22/rnh2biZHyeKPFP74SZRB1VAcmc4Er2j+7PTiUtaMT0cSo/1eX74NFac8FX
cS9YVnX3XwopACFaXq/awcxpUvBy/O8hABPi2KvN4PDLi0VWUQt3Jh7kKP5Rxxx5fT3uxfI6llYK
l6YTPQvbnyOHwsQ0pV2yNx7yH8IIGjQr/RmUY/MrVzfW6cpxfugBGwNYZLyjh73lOKSXze3nrjkn
B+tF4xcWNs1QNm4SP3PCvz/tk7IX0kdxMWeitsrH/OP0IZFGGbr+gh5baWFWJXAiCuaJnOdW3Otf
MxmpRd8DdQNeX89ODv/EOWYvDk9IcJkTqHLHlAyfcaBVA6OknwbSC5QxA2GkBA3wtCMOgCMOJOi1
tLGBkD39ZQ7T4c/RovGXq/9N8BdXEGfPVO/QGyQT/5tCGRoaHi1uBlb5FiFWBK9UBaQZNKCmm+ws
HbFFCmCvPPwgg/13VG6DPT2IyZGNYt4Eg/Zb2apEJ8kEALpj4/pvLunsjM0BP8cltCWofkQhKMO9
PfG3sTsGIAupgkRsuTENeKlZQi2JFNnUvCubZs9rCWj4dpVUrJNPNwOvtb/hLRjplAJc+Lr3LrWA
uhJTcPXwM4GM7lCWaSxh/u2Tg60dUY+rtwr0zGD1X1HqYMTgwa0JY91D+6et0O8Gv+58XguRcPmF
ok3DwQV6qeVRc80QdKfSGUabamIFCo/cPar9cfEBNjNC8/zLn4ydsPbR6pkyf6TECIYCoYgh1B10
fMuWskvR0RrgvrjFd4H3yk2h0fYV5EPo6ZPtwYlklTfHNRFP1EWo77t/GortoWVOfsl/M1YB5EOB
GSB4QIif+CzYp97qzc4G50sLU9C0iZ09IxDWT7KSw5dNdTW0+iV4wZ5atjVWbyadb8eUR+xypB81
KCPm3c2moVgGeEzbbpSHPkPVoeJDZkv6tJHcR1hj6Tgo1+T57CoiPz19sDgPEdkHaglzxRaUNVq/
3Nihhal4wWnmq416hkzYMB0SEtaZRXUDklfmSC3cVTCOfxHC8qcl9bzag0WC9083uhvCR/U3hGDM
enPsGFxew7nw16DE2Wm8DVzn2dBQOcLaCtsMiheQMroxtr9y1gFy/x/y2BVzn0RAS1Ru4MYcKqhu
40snoBUq4CiH/ogZCE7CrqVm/KtCtBFEv6E74febYWqsNMDW6M5ig3dLPnrSqdm1/COuFQeiXRBU
+5iC8ReE+Pj96UUhRrpAJWF4J7XJOH20ZMOvw4DeB1dkPT4ecgAx5NXapuBCKwnpZLJXt6q+IkB7
T8PV7gkJzDf9USwiWftpxckkiBJmMgdxj3hnJgq2he0LArf1OlNJP2gncOgPls1WYlhgG8uRow56
sc2CEQ/N/ybbw0bzzPn8/+RSJKdZI4sngUf4aM+RcICuIjASZa4BKJQsfHmS9gjmBc7Rh8tojPjd
Xiu2uYOulj4ckZe28oUfQSAVpqqTno4lqhj7vWsfrCxkmU7PSm7a2u364UrvTON1YO1TNKfB8JY3
6BK7Pc8Ei677dhLFOZjXdvPjWevuBZxq3Y6+hBv2ZSIU3RsZatXwbYdsy63eEg9KFpdWP4ddUMto
3ky42yTo9gcHAgG8dvQfFWP/l579DByXJG8QDVq88D8f+CPlk7/TcV0ZHR3OjH+DCAdRl50mbH9n
wHA85IQrtk4cMyqmaX9w6gQTP1/j1IAoC3lrcMVYKEeciFMFKG756POHehlPFlLb02NqakwkTRZd
BIlMd9SCS6OkoxDe848r0o/axTxBGZ9TVITSnuTnTcq/f7GwGMldTAXUN3Fcf/xZekx8IDkk39eg
7QE0xnG3aP/ALGbLP7rR5i7Rjv+q0n2BD7BDSOQcGnFuvEzfiaKgABTDLtrexCeTLqQXSLoYn4q+
U6UP4+3dZdRU8kH5cKLoLbC+vAyVONd+iOsF48wIbTjtjwVQ2YRWxxlyRywZkd+d043KGy9NQ5sl
inbrD9sYNB1U5rI/FFhqamYCtJvcrw92dZA5RcqvqzSS0B6T4mTr5iiKvosvFyOtf2LjfU+B9jtJ
S90rMALtFvGwPMEVMVaO1glaDCltVHjEj6ajIOsSoHu3WzKSE5LEv0rpwJxDWEaBctKa3g9WoTx9
wwGmA3tq7v3gk0LqETlaMqTLeOFsCh7jL7rv5rfshBChzHgGlt3bA8zx596k961WwQhUGbPq4nG/
sD1tzZa7akVRtV67oz0UkPO/SXyofXJLAIPyY2z6BbeT5lZ2MhGX5KKexk7dchehlXzU04qGHMZS
1oggWrg7Ld+q6KHb1VS5t5S53hjlgmpZf5aHF1n4Yf0T0T3m943+UbVBjCXkI+Bo5SI7fx4jCK37
3G7rUiQvA0RWLXZSKkoI8jUcZOfj02UDRbMShnJ6ZvOPSBcX/TyMhy87ymRniaVpYMqajRUKLzKy
KjVePy1tPFq0uXRAoowELvMLf0Ye2mXjeRGAaDE8e7S1AsgkOb8hneaI9FWygXDB1WUSmBbEbjWK
nT5AP5v31Kev7a5etSIu5d23Lbp6WRDujm39DeqzIP8nRLwZzC+2bCdtbE/FOiGZ9tJw2mTAsI06
Si1xkMVT/TxA38cNiPATPwNDPI/h6/9OVIYQsBfbFtyfTLBPtYwHgvzS+ZJ08/gOCjqAdzxVUdGz
ioJkpbwwnPJ/6BzDxnxPlNfRGPbvTeMntxwAfvlpD2bmm86kdAAoqEXUEd9OUW8XRs/Ea6GFfNvU
iLBnrMTUpAdsLvm3ofNP7rsxu3cg9ZqsqYByT6cF/NoObv9t0AzUgI/UKYtvfdBAHdIC3iN1kmJV
mWaKeTsiBj096mrhZvI8uQ/aCl73bGSnyZZhbNkWyODi5b0hixKuIIzopxx9a0Cny6yhYohqnByK
x7hYwyUKaloRP7yxNMhmphgFwr+rVeGozPmEuQFroFqtsVd7p8OgXryBb4vlSGACYstbhcwDgU5I
E23aXDiwS6MUQEq0mQil+qYyWXpEyVdeDG1DQUjJbWKUBubMixSKkG0ZB8QuR3FBPbnAwXfl8EZq
BIgXCInGZ3pMQZ77hJlbronSj8hhgSqFGTEZZQLctFU5lOdziqUeD9IsbweHsg6rWFu3rvfSUnvw
YIaoxU6xwbVTsY5QJI2mSDWxXciH6HXOgtfr/fmjnCPs/+reA425lAR3BAgsflye9neDyxbrMX9Q
VCUWTWIKtPLpCJwphLnaU7ZyJ9QE3g4/3SqTZbYg+5FNqHG2hsT/1xg3CW5alo+dTf2jO4LQpxtP
5OKY5iG4yWH24I9Pn4lbMDdIYvPAFMsRYjL+rj/z5ME/16IxCr5E3u5iRQQKME9JwNSxC1nilcH5
5eZ8GQ8Be4FWOs9Yplj2PLKIwbPoEwD7uTk8KMzJT4PktcWp4ptDZrZF1WGVZRLI5brqGlnFgPpq
IlbdAbCrF2rxqUuOXmuiHcG0TYA1fxM1kOH4zwBQykGWhPrvX9LOPXOFPzxmBTKUWZltIa/1J9TI
DuiEZVoYK6z+B5gIlCua5tPAqZC8VBGvUeX3NhRkgIT7j9Wmxrbz9ODId885oY/Y41UtY9mqhqTc
z3SNlNt1ILVDQeFOEN5R1azpq+FcHXXqyB5dZa2hSo2twOqQg7YgXHrUI2blxmYNsAaCo/PWczfK
uLRXfjTsSQKk1G2fzqKMEArq4wQSJu5muYjmPISnfGcuEv24DoS0DH3w/GHtJ0UbCbAXffnSh80z
aIJiIrdQPOpaw7f6z7Dc6YOvEgDu49AGNdd6wmOZPYxAaTP/jFu2Bh3q9SQq8jG4ZHTtk3A75LOp
4JMMkvZh9o9ND1pMpsRlKfYfcUffWy+cyC+lNANsWvfwA6urVmgdgwapTWecv+WyKRKH17RIQIpn
c296AlHkdBfrCkzR95AcrWIjZ4hRQQj8sLQRHU0gR6AQWaKkdIu3fA7v7OyPSn2pfKviUzqe9Ejy
mg9uj92aLUvvKNYd0MfzNsug4wRTt2oFU3d4WcKzWFBusxYknabRM9WcaOGg7r5fJgLG6DJvd3k4
YtUb2m+vUNdG/K3r6XesXkNp1sTX2tzcgdDX00+wFT5t/CoHrN04a3/JN1/sfQF0o25/N3ob6k7H
ItaRCPLa3R7Lr4au7npgOpAmVYpODYTVdKoGCi10U0Djl2AaZtb5w+0JsSb/rdTI1r7fYejPvYhC
c5JuuZQltwIDT3s4lblDP6vO0EB5hgwPoMDEzhK1dsEMgfWQz/YC45xegrEtU9vm7Qht+YvNZ3G/
QcChkGT82EIGQeNyJB4vu9xQzK2weVV6Wnpg+R1POrsFKABlr6FaIo21l9GvmjK9ldQiz4fqgmsz
TiPVeH0dLKTGl71k0h9u1WeOo0vbdeRSsd5UnCT1+tHjwbwe1PJp6qJd9XszqaCuzqGptMdEFroJ
2fxkdW0tNbZGYN68Lx/QPRgxL4rN7FPXxeUn7Ob7ien3tHEJpAAg91B1cGJhImCHHcLWnSj0VtWq
CGo58BBvbGwZpNsVzsnXLmJ7WR/c9DrrPwfu+dQ1nbrn1/QMPPBEkiHg3mtepN8IvsCBTSuIm+uw
1x3Mn4cWq7igE3mNv31vnTsrKUD6Caq9PAQ1iafcW/+d/F/OtwSVP5B9feDFkDtSdsubjcNo7rff
2JEL4WNx9uU6Ad/oSTTLCWwLfacs1Eh0ty4JYOVoModdWHTVThgBSgbeLUekngZJkSYju5CN0/Dj
JpDh0gE8S1BsBaequk0CrMiPzukqsLeqAcmRWNqLDG/AqSPub05YhSp0BgTg+ZdAjvv3zcgWCDb1
gMV1NH5LHp+Wj5CcgY9y+VK6+YRALHLN/x0QG5yHKzw+5haqSkUBf2YJEWUwn1vCfEXYkx3AAlR0
ZMkYFhG3e4NKhccJyJF1u95A/gNCG2eWVPMV5A8KCDSKc3dwhfCFEnjZ7k7OnFyShv6h5Jo9ztqP
HQS3SDAltwe7+++2mLD/VXyLwhz9i1L6iepzUaseV2d9h/fP+JXqg8ZU/CPXri4SNWD3lYdr88Th
O1FhjTwxmZSit8+jQ8zxFgAefLhoeRqqJT3L2TPo1GybzOf1RfhfVOOwCzWB+JUP/lmzV73a0a/Q
vzTY6sAa93dJ7euMURUpgKfovES+f4h3is9EC5K0bax/a5Pig0N4Jp+Xp26WK8FGPWtxeb5ylXl+
C79J2f413w0mJN9nQWvhoOyprTMXEq8YKdWNbY3uSe+rXFLqZzmPoYj18O8PZZREAL6R655Jekn7
0QieI8d7HP7WDDqoSUn4NoAStygHFxGepFezimA7Cw+dZmstcqto5GunBWZTCA5HE/Lock4K9U8W
lSuAY5jtNLm91+X4n4TrSz4Z8jbycDXD2HVgHHl1A2LJy5p3N14xbEs/4kRRbzxa7w0jjHwftljh
7luSYHM4mWiNIKKRQ6VwYlaPASuc4cVPIXFCoZt/g+J5NS9/irg9Z1F1eXzOY7DP/b+y+491xrDo
BWYw6stwLa/vLocHJI8ZFof/k0aVj7nY9z3nzDTIb8uYVZmuMAMObxk16tIUChiL9vIv7I6BJbFJ
WlfsVt0ZQY0g4Od8Wt+PukhLv18/2G2a8lsMkFfTGdFv/jI8e+p5/uTwQwdfAdQCLR3a1ipL/GzL
wEiXVC4E5ff2Aj5JzVpPZlwu69VTP+RSBYvtMG0jeb2CGM/5FLMZ6exsJ3iSl3wZQQqjSJqaHGtl
i7qjP9nrGPd8YCLQt8AsdEiJTtJAFYqqrgYeIqi/GF3Izc1gCCZqYLPCo9lx8Ht7OMKhG59tdLWU
9lCDlYp4byHygU0mynLlLNunENujJKbIZHHrQEQolBRMzosn8J2nB++bTWLBgIr5ZBYp3k7rtAg0
O27XKpiMKmw9eiCBf2Cgo+PiHYEsvXbzcr7n5lfJOqQWP+r2cNn4FIJoSJFr98LGQ2myPbqKowkq
LFB6OfmFwyLtQMC2wC8PCOVrzw76si+JZAZ7xvLgcHRMR93HpRiMhH9O18AAD8nBrChanayABN3d
Lbos2W3qKRN+9A7r5V9MXoXFItx6tZKuWXnTjwO8ZsswGTE/iBrmZMEHyZDf6Hgm8ZhDNxAHWg5x
rxATU+yj/y2shGYk7679XhlxoqjJZOT02WPA+nMH2hOilb0xTwWaeO+r4keDGCB9CEd0v6AGHYr8
zvNcV15YLi84Tf8+XueXlBIL6QqNTpEez2wq0rWQ7RWVymvSkjHsIzE9o5OKLQwtKUfGUNFVEQTA
y5hAwg8BBmVdSOjUhS4kD5XZ5uryE9Go+ww/OpDdI31TV7ANYg5hKG8BSdbTOXxtSkSDlxgQAnOS
/BfQ9+EIn3Cz7aty5e6yOfssqpzt0NNeKnC1ff8yqNH84V3n6OlUzqu5064MmbCylURpjETBA7yW
Ex+fnTcVzpoJqcZpYv6w9X1AoSpR2OMvKPo8OsDiAcBS6KuyOw0GhbCFc0yJl6P5+VeujriGJ/Nr
tCQKpgWeLetZabrgEBKaOXRYKxMhSytAM7RvtcwkC/CMH3Wx1szs0mrRJ4OmILfuvGQOGOSTkHNL
lGz4QOdmzQ40XjY/geKbX5NZaGDjHxbRZNXZPtlLt9ihSdFtoQWa8EErktnL+SwHxoJfsg80mMPL
c8765qMzOpL8yqiJFu8FmGVgVoQQ7mTCXtF8azde2wFMQXhmkpGaKFRUvtTyenuMko6HKy5joxBY
qOJpLkDJ6CZxskglP5tD+PJIh78oLxrJFDJN5A8atqp45TCgks7gX60GhFf6Bm3Pw4MnMR5Bn7N0
ad89JdcLCqenLiBKyILM6iKYvWicCc81V2N1l9uOru0NtDQKcaiNhRu4qmFrR1lJPRi6mfDkfCYF
KDnAMSV0w897jzmrSvoEPzev+OUdxrWDn4zMekjexfk7SP3aYeLaScGSA0P8PNXZUGAcFy0loJir
KvrD3NzyQG7l5CS2fH48Q0H0qOUu1893Mhq6kJ0+rcWEn1T9QgAAMADXxHFpWV8xIXV/joBZK5p1
QdZHM0q75r8jpYJ4JNzB+qfvqwySZcQvCkLHVC9yIapMnh3McW7FFMqr5o7/AQu5Nz1cQow3+OKO
bf80eHsjPPsAz2DxUQWIvOGw5EcGkFpbX+iCPKsTHjZMsPhfQns0tFW0y/vsspFlRJo5Cedz7TfR
8lxN5LrAbU31/0nbGGMfUK3TE2vn9H+QaOtSRSWR62Ws5NNVzMKfoFMebbTHm6DJOWSSmOzOJtsH
kJbaU5eOvrLUkXHRy2Kf1P8wx4RrRZIlXrrZyB/jdo53/kDgZm1yYIkxzwt7q97eBfQtoAFGaFaj
PkS65IBH+E6ZRh9bDczW5I0MpCYrBXDQP61iN9yjTqBwnhbQ9NhycGBFXafMXqA4wAvkpIlQa6qN
C8fw5ri8u3N+LUjpo1PH9E218N2foEgqZ0iLwL8wjLdNRsDv8vTUqaNSu8vLgDBhri9OtE2opXLX
W18YwXf5nz0i6Ut2fmgoy/s9rCIx9HP8gc3FocJQRHefaPem1IfT+aoPX4kazX+vb3fpkyxeLDsd
pNpHzw+1XMELrkwXrV8rIDxv4jB2jWU8LVm1/vdrFA2vwnuhttEHnfS0cD7X0Zr8+s0FQEcGOj9Y
gI6/tylsJ9FGPKHYWl29vm0Ng4gFgCx4Mu4S1NbWoLxp2Z8ND5g9j6/wKisZoM0a9mOTriX4lynr
eXLNGLPFG9i1dh3/HR7eQCLfGOGMyn2Kw3YvjrLkeY1zSsYKdNWoouYuh2DBVixTTyjmXKZPWw/y
uNxsOOobanaPDJ62sMhhd4jZST4s26ZorJW12QD6ReySFLPq47rTpiW6UjUEoXC8W9DKQ3QoM3Zs
g7AQD8DX5oClJDjlkZLMr/1fSM5kb75F0zlroG8maZWJqM/DD/GVzD69ZfCsaNEqXF91TJJHhIX4
CrnlDXxi60tfeBJiWs+nHCbXsHO/dgdELnBclnw9z9hAKh6MwtaZvoi2w9JiB3ZwMagRIveDf2gT
aMC2eHuEdaKENUtyeaBTfqAtCba1IgbnsjCaQV/eG1j70DA45Bk8NB2a/+rfwbzLnCmKwmzmQsBN
Nr+8AiZgljFQFhpqZ1R1qCIuVYB6dxGSlPkRxIHeLrxWjySv3MN1mOADjb/EMDn/JUBECxdOuPMe
5A5bbdsmSDMTJw48zbGVep33jIUwc9tgy/LVEHjT6PjA733f5kaYMIdwdCwNc65v68efduytWXqq
8le+HyZXly6Dwv9BdB5EjCEAD0kP+OfMvGuqddhBLn/GiGi9ATqIcTpALe5CfpjKzdMy1zt+sa2C
D5QF1gO3MSn6yGe3GvnpC8ydDdTHSq3+cs23QAbYc7C332iXvYyumwDcEFq0ik/vY4+tN5O9ReJj
M57dr42jC72axFTbrMVrEc4Bj+dHEFAHhVjp8dopb6x41AO+eAFNTrW5H9JcrWlQFi66AI3P8koh
/IxwpGCpv3R++YIP5qzUWlXQlSm/Btv3gcHvCaYP5sSMihIky1z5rgfyrWna1CdiCe/6hyq2E+fk
OOWpzUNBYQmoyGBEkoBfhGtUpGKoAvzvz+5oKd5n7Es8mpB3ZSUANp+9LpdSEH2lDFc1mcEzuPv3
TxO45kgXUmYIzuF0Mv7OhMQZrnNDLCT7Dl01eKEZIyx+dz6pqyo0GpuEVE1T2af6L2bhfcOGTjYY
nAfooQCbqwVMJ5OW6kCwyuiDWTACbumWOWQM1r9dYahSTlAWCZ0WhtOxIOwUFKUIw69h05BiT85G
wx1jbTDRTNMRarVmp2EfFF8m7w2CgxmrwpGx5hSuidSRcAOuQfOKnNtD3STl8y9L0xBRxd3geqvZ
b2BEHGXP7PCIrKU44zMNTsFVSv+EZ25rX25+1F7OKBs3amhrJt8xbDr97E1guHBiDcMdZLbGpUK8
kvzXI6fivXJLI2P76BpgCW8Ys4AZGk5X4t/NujRgoM9upsQYIa4T1ayYXYBx2zGwzenwtrb+AIOu
Drez+DSiS3vDDH0pHi5dvjxYEX2PStwTgGo2DuQWppoAyNvTA2d6mW6HFn8kMN460zgw0V2R9z30
DN+qKKSu2RhGTFu7HXAnXfdK8ml0XBkABUL5xE7W5SRrU/54Xl5rvEvzhHmnJ48iTaeLaPY4Mm1H
iXksX5D6KTMfmpRA/RUDq3LGRlrQbcUKVrj4AEmShweH8UT6Bhu0QANbeUMbSezc+5O0/zaJhz5/
U9ybIVk/ODMOXm/25FTpuZ77c9roZJLkJbuou1LDz1RfLMn9w5Vlaou8KulUEQSm82K84lHsJ5+p
QiKotLeemz2pv+N1OSnOQsN6QiSnnFx89jdkbHiY7sjhyx6JKeJKFB7lOaNB8VeHqCmnzgSB+ueZ
22GoCvx7KMKYdgNsrNEBG52wiHZl+keJSoLGSDeS7zMnZ6GmJlfAaButRk1GXMfGf11ceP1GbjhP
XxHUiaggeWUkapEa6unfCisB63OmKtcSa2HH5f84og4iBOiyq6rj5PbFrJH3MOAyAe+zeM+HdrFF
EbDGd/YRiwwKWl0sOKG/rjJLAYUYDat5DX6HuJvc0HkhUZU4xyMa+p2pPZmJaEe9sWCj96xMze7A
5rd5nNQohr/aHuaDbXRZ21Nl6HN+pGoTl06A8gRK1HYfO80OhPmwSg3IPRKkBv+dldZchzP187dV
Z772wjkELWwQl+BPDXGXdlPmHhPbUqfObM3u6dYx6I9p50cdmUK/G+yesG0ZOydXr/OqJ7snMCb+
8D2EmkuRd9vZzxQ36JpMKavsrBUVz7klfeL5jhm2+G4quUX+aup7kNFKXvSAM5CwGpV/csVge1Jp
7FMJPgq0spDOAR5V2+75IgxHIRdGF1RCxIGbgmd4MLVtr7x/6LPkNmmEXgc27dDxxJAd/Q9a+80m
zDu1+lyWxztKBv5ENhxIizvUw/GICxqjMsz3zDoZ6pwgJT14GIbQmZnoV0I6+wJgfg2kyUyO0VcS
sxnGlGCB9Q5hDXIVDp+JDru8eihc3USAxkd3af0IVr7NFb40ZeZJCsG76wzAzfmE9sshFUj3whQP
tFS4EDLtuv8KKQ9hxOyhxVa9WSqOnB+P7YU2SnnRZZYLaoTWcvYxHiEaoml4FIXJCBc2AjswFk05
opG1zIJTKp5XNUlo9+EvRGi37uRZyJNaimJ9Q774fuDECO1YHAIvhXTxJFj4qs7UyCEaZtpQX7o3
WOqE2UvqpoKCI233xp//XDVzOwJ9iSPkZ48rnG83mmVZV78Xvr42NG6HjAGu/dwoWxF6UpMlwRsH
35MbLuAvwVD2RARzmChhXqWBNWIVcyanWWWdqi/SJbvdjzyK9k+PE+WWI31BQ7D84xYk1BXeTU88
3z07Qlnx5f88F3wcXiMZDaOhZe92rk+1JBKEXZvL8Ph1ao5DC04iCq+/9hSRvKSNlUqyzRhmebBl
G5wtJsu+mh07PtKKtMkeXOz73C1CigJ9AXaLXikiXrqbAOousJisz5F5bUy/rT5hB2MlE3+S+Cv6
qOnSJj9+XerAJqEOWNbT/4PCMkyEk6o/QgC7N62qhWNOvt9IuUK+9YSSXPJh4FayEXJ87uc+fwO0
5GgHVL6PAjsqtNWnTwi+XBc2QA43CFCqXDPPs5Z6jMwf7LF1nJJNb0WrSE/ot7h4h/9+wQY+cVra
Qqqo7F0h1shnXy1a/dKmfgF3mhip2wjmWU3X+W0DY6n483yAG5R28NCq8I3Anug+kdRzpWNzK5qc
r9HhgJeS9lWmFbms/M81AUpNq/CDulflFbaqr6kpTIAuwmk3Swze6AR9Zve8hEP+LViymhQ/LJWR
Oy72yr2sLBzlFUrHn8sCeXQI2RZoo5VdNoiku8MqcmzBqui6n2AZXZU0iZxOC3fOxSGqk7YAodQu
677Y7JexnVZJzkwxLJKaqi+T3m/+g6lWktK+o7dSBGgUAvEzVZyelRLtFz0NGffFawtxhjRIH/tf
j80jdXoDJQh38Sp1x2w7AfCyYu8/HnQzXZIqAPcIumIoklaAL6E8ciIjeUBlSjlOGij2LJrtLtd6
ktnmilcE+HvE/xaNwMReAU2rIf+RgSl7aQASg+rYn7ScYZnnSDNvkgYbIAjhRNsR+dyvuoiKZWVf
llK2xN0K2HhtW86RMo9tt3oPr7CNtmD/vuV7i5+8Fb7mc7rpUnL7QNsbcclSUwIdN7miOKVn7Goi
WEkaDolk84kY+Q4aLz4nJuK0op1NZvCbrIjvXu2dcSgmy4k5DT0KLRvnZATzTH+HRFzM9mO5pGy+
q4Z3xGxCU04K7LaokSmsx1sjx3GkX0dU/ldxqTYMUe+one2Nbc1sS1dMw2AdsQwDLwnkrhzHWA2N
z4tDLGjBRzO1sNBqXmj/M4XN8C3Odzepc6KMsLwFqeWEsUxJ17eh8+J9AfYRqZaG3S/+7M8C5Gwn
XeIkvZUxinTcSLy1ulkvdLsk3N3xXPIXtKAjzWoD5tMsLtHFPx1EhO7VoTsJ86cTprhRJyVB+zHO
Jn29DfnZFINWWKebEBXtHRf8L+Vc3OxF7mU4qvY7H0T6MDaZSwxbrM95hBmaC2NBk7NL9vfEhbNx
rSzKs1B4dv7JznJSE2D1r5OxT73mdsSo1mig6K3WXeqr18kT3ozvAAsG3lvtq2FZSsGzEiKIDlny
wDSdJWgnD4SpNjAjnVaW+cRApT/lz+Q7LBE8NVhSjApVw2M2/siVS/F3YOYHsA2wID3WD+VKtHCe
JNGreF5X9ARvy5yDdI/dLDtVQNbm7Rf+Hep2EeNkL98IEiYetXRIewG87tT6Sat1gNIbyDWr1p8y
0zbC5cOBAEC/F62fYvg0y2CsixulYLwXNs4mO7ZvaRKEadKnLiY7aCaFis6Kfgf7yR+miOQgTuZ1
kjTjFO33i2rG/ABioZF+MCeJWYpce5nAGVWYr0fDIheqE5lzFB88+HDqdJw1ueq+1MFNrXnJN9js
dOvFPv0J2S7q1G8LU7O1F1DslNyAtKhj9t7K0eCyaA1zGyLK7tEMEuL0JUvCMAszEtnXjGQqfdsR
IQEqoTr9G+WvOX+D0W8i0ao5lQ9Et5AQGzGQ4gj98YMiTBsJOIABc2lxIXSvYz9HGeL7vA9uPwpi
ah2gfaT2IGGYEBzt+DiUfGHnOOYnaqgZdak6V0twiUoXg9W//EQ+GGIKu9dc/FvbcV8Js+ldr+aO
MMAx5HW+bb+NMPxdQ4vr+uJJXF7N/LsRqlcdOGNOz+ATCmUYUmFrRBnuogkAI9jLw1Mb9N0rhIHf
kwJAlNVSZ2/KEbIkTJcxaG94vSSykoSBxas/p7XNHpVwuFBG3WeZrRGZ8dHBMJNXzKTP1+Xr6CD2
lO6hjwd5wtPDIvub+wDEMoeYk8rkvsfLGHSW2aOjChWN4TduWx/WRXR9U9FDqQtsZOjTLsi6wc8F
VYh7WS2GbHVGkjKbfmQovpY5b1Ij7vvf4243ORygEWMdZ6znnl5RLeBJc91ZcOcopaFAlys0gTJf
McsW4TpkRG6lS4w3GMU5Y3prv6y02VVHbZHO2QZ8mK2IfDc+bhaIDuitUPJqbpfFlLmYrI1numWi
lOABCzKFR6E3pbonjgoIR7c+YX6x1EPTudXIDyRMI8vqm9jBisz4wmEdOo5idwMjyRheXOd7kRJU
uoB0EbTYN0nBSmnkM/pl4z13kcJctBIoTtwqlx7GK7Iuhot0HoxN4XHCaSOCBtOaSTvjaOzoW7jb
uiFj7LqK0EgMu59Npt2UlxP5wQYcQ8Cero6Py4nkyELbqpDlSMFFe3CgLXHSnowGMFgONaksYTAQ
RIzca9sFjL61kejddhMV08GYgnEwPioiHVyRB65wwJopLS1ysccgNLzvl3NbZpn1q614K9/VBI7q
4rB3ilYj1WHAkU9Q9MlZYFBAGD5QmLFb4zclWfiy2elzl8KaOR9jucB+CvLc10s1JiJe/D8Vj8x/
7eLUuWpHYLGSmnMbJRzbdBITmaGEjn8oIYDs3VEtqsHrfQjNuRrWn1YRzC9ieGldj2c3Aiu2oZ+9
GiJqDjc/zxtWUkFrfZakvrmqLs1HldmB9dmfftos/tK+8LVwGV9JQ6TAQZO+5oqiEbe2KGEYtZ9U
kSd+TtdEE2x9X/SJqAR6qWujVTFJeC4YqKB7C8b2I65FhUqxWyWfm6fXb6w2fVjpXT7M9SjMNeHG
SJ/dxrY2qrDdSzDqkUH5LyFTsXXLWz0k2LPCP6anN8pAho9wEKP25GPEsFyoBcelBirkpgJFSx32
6738izugMuFIVTRjyxmwVoJRWkoGAXBsK/cmy1OgYKf2r1GomrHpyFFs6vlGrtfButg2DoGS932s
ufJfIurcKPUq5m0Isx0RUuhX12sIO+CNvZA+06y2JxVYKJXmgIgpHIzQqLHSVQ2AV/9+/u7w9z/m
vFtCSgwNowpNwbLV0bNz2WbcKD0ltUEhQsCaTfY+pPiDatbtQ8wAuFJZT/RIKQCEp9pbcjQeBS+f
VuqrHUrx0Xa8z6fYPp4Pvi8Nuzpbp0c/B8G8ASZlZBlTBSIvaV4JczjuVGk/SgG/Vy14GB+Twgwj
V22tbbsnU1lpfXNuWpWko+8WY8+g6QzPMaCZOAxMCocggh9YhfHcT/g1bNui2aLGnXOd9VtvPQmi
smXbxwnHcExGXw/8yAYsk9/OIVRfKuNIXVtmw0SNDSZc7+J6BmwRvsPQEHAXlmO3c322mL7SGZla
Z3TOYg1cusqlKutkjr546qWChD1OybLkR7+T34B65QrmSOIS3TTEVapfhKcGyMZh1Y59whhl2URy
0lxydIRRS8gFrz5TbXw1ASi5RyvwNCYjcFkjqmXHqdTVVMLOQhLxxhehNA4yPyuxPVnFjUWuWRU9
dgyAJbbM37TjoEIQ45wRdKhm2y9GOSzFhMl7jg6JRlEzreE4xRD2nEaYK/Mch/YFiVu10YuMFYPD
Q5lw01dRNJOhnTlgTPC/4pHVTJorgIBNZDgQ/nE3bDQZ6KDIXJBUdI0MtfJcf4Vh5cSMNZwXd/Zt
wachbWnFziBhYzSoCxzthLYqOm5zqKS/EWzHHfi5ys0kgnBO1V/rvAdifxWue/XFqXZpx8Edp9f7
Fi9A8tW8lGbbQU7ls+IkOZ03RpHwaIeTZbF1MWM1JDyqH0eUXNmGIJq1n6SJWKrp5KwFPEv8ebs1
/tsNTNoWRcDnfB6/j/ANHodDCYGoHjSdK/qfS9afgUiUi77H5fYYqZCyH4iW8cchpcGTGVyW5Win
usAmmHjkI6Up5FlwdA4Ap0xcPqdTK3gWBc7vIngvIYOQqUI8n5TWxIszVx1vnn6MKTnUJsv+CTl5
BKT6+W1hN6lbbhKxWe4vAKp0O7/ErrdNsl5RcZgKc5OqwYwnpor7UIAtfpGzI9dXO6y1UHVTsHSy
iE5epbw+YvY1HdsS9iZZFUKjhUPJFCQdp00k1Ls0lM5BOyqACkguf/FJBWek6vIvoiD5Byf31A6M
UCcOix8RVqKx2IQnWdrB6XQ7ZKiJiYzHyk9+//KkBSfe+q5qrykS4kEWdar/0tGziRDcFEzGyfzF
z9g+zm5WtYVn3830wdGiG9Z4uN3bXxELlvbzBLImWmC+Yx+EVZxLlz23eUM462SS0pgLM6opQRBI
JOgEsmZF340AK5IWel2+oENLZZLbApfRE0pyu88/WlecYWkeoBAgrOC3T1sjsE/TmspRUetvLt+k
9tRQPu45y0Geetni7Bg/5Zhj/l7LwjH2OYn2nIn00PZ4TpAEoSIyF9kQX2ol4apH4pOXwQ/3APxn
jidOFMAeC3mNFk/vrpMC165BW5NdwsXKHQSOgWn5RBd1JffPVdpKx4EBDLmjMUvjPEPgBNLnQMRv
FcgUv2FpDSdff4iC3zVXiLcgY0gq+o4fwkA0HkQdBM6kl5PoYfIjc7wqw/WR3eeEk5KF72q4T1Ex
ONB+YFn0cyD/sBfcccz9RDmVJn+HXfMHncOhCPAXAL2SqMkbUZMrINhy373o0j/9qqgUL5A35A9k
2N/KgiqPphkujPDSzSCwz4V0pUm9wv/qepZd58YwieUH9JhbDrv7sgLt/+a/OTVcBdrKi26rp4Gx
RBGdPme1/7qD/hTzGCV1N+nsf76vixpIYhsBIbRDFDFmwSBDEOWAkQj3x4z3ytLnaOWCEl8du8tx
Zh5pLsutm1PkLh+ZeJfHv7kTyhSnfIkG6KIOE8h0ELZzDZwSuqRe6Qa2j4fu7vRZLEExllNtQFnI
JZvsB5aYIluE/1m7QXGl/CZEooy1db/d21OClP19JoAlnDHZhqa17r+ePkGwwq8EmSr2rNCb+xbL
UtlsZqc9+6wJGsHPz93B62Mi1KOUuYwMb/AzLE4ozYIpgXn7eAvm75q/nKXwfAhGtPajMLN7v+6f
jVY5UbNmLQXMxIaBYOJM7JZ7OefO/7W5+CyXARogyvj6H1TRaGHPTmr83roozCSZfT4fchqdj00l
x2ssw1K6qRMW9be3D4cZH3njc6+Aw1s1WFoAac67iLy+HC5bZia4y+gQIa0FahSVRGZGAkQ9dfIo
phbfOEz16D3yKBhHvNlrpzS9qXkGtxhwnkJL23lQvNz2p7Wzglr1fN0hM45SRMh2LHLoomI0lMuP
MR6+GaridhGYT+YQgf+FX/R6uwsmxkGpJAoHxS2Yf0Ea2sh75BREDSdv2HwfhYt4ulaEf9LLCUj0
l/up7U8/YR5D8c1EGjMWG5d8ILiqWo1fySslePKmNkyfTZTabhzHJr1mumzPd6ydt/9hc8Y1yFu0
Fh9V8FCUIkcwFQDYiDze1Ra85ZM9+ZEZgLo36vhe4nhrisIDGUTR3K071QMWbhULfpc+VDqRxACS
nWUui9MsXRWR2ALqqHZdHlObZPk8adEJgBdsDjWfthVgJEN8O7momNtVsyaY8Z6jbGBeXGBar14I
bcpNNmOPze7TySVqM4tXEX2U8xpLi6sPYcBguKLd9APGKP0Bv5IQOqem1muTNGccaqcZkmRfJ+Lj
Tj5RGmYi1P+HChtMstQUBB2Xd/nBw2WAMFDoCqZ+azlWfoQz10XBoTKRILMlaiqFh2KpvXKaGf05
kv7aepaDnk0n7Wyb3h/EqlKAQX1tZX8AbWX4AfQHxrar+1pJ8/Im9yR6S9SbvfhIS6b/6UDApeML
IEwnqD+SOMa/YIose8MXulwIY3f1sapIuvb/b0jw/r07UXfddeQkDZehW/9wMWdnm85IpnFWoq+H
DhkcRRGHjq34ymzFZ9Q4imClJuUrv7Vwrpn8iupHpg8SxVKuEkooDkhUUzP+Z1siP4HtW66BtD0Q
FDYhHmHuwdyzSRRzNWXdEl3uNivrSkIoSyUhTqSTzEd8d0V9lkFvP6ojuymQzU7NVYV3G4WLUTCc
CK7+iyDm+G4xNwuTzz9/t5Wuqyrk6ftqd/jjo8WBaQ41q8caTEU9uNsrP8hFoFj7d/Hbh6/w050A
iB5ozeGDIJ0icfvqysUXmGk9tcNLjwiqA5BLx3slo7qZBmuFxUwkw+HejyZ4cl1eYCbAdY851h0/
cxYcqPY/+5zh0Tq6q0yA8oNtO/jwYjE0jqD0nwXr0RdfyeEwI92DTNb2zBVwonruTk0+Wb5B2VAZ
lDy/yNQg+4qlhGG/47AvM0NN3FQRBDkWOaGyqrqeOkAATJCw84qwHSRPUtvTwGiMfhMjVVc0KwN0
mpzefxoQTWZvGzjIa6p36Xhk2QDh6sH4wgjhL4QGmSRjLEuia40n7qO9k6qmjeqd/fhH4iesxqZe
jo5AW0FgSoyrjZ7Zs78AhHMk5kND6Pj96ewMUnLZp2NxW5iYa+6jUdO/BBbh0TUTuJFjeD8RnU16
MuYyd8MaU/wlNCzd8Gnh1xdVRhcs5PhpKZS+PalcYKFspNp8LDgnbd5WEUvZP7XXF7RemO2gZMby
XvF+vc8Ax9qqSo6DRvU9jvn+Gbw/qry+gzXAKSeZvJrRdz1AudhdlpMFATkY9Y7fMurXvmYUytv2
zTroYJymY2+M6tW1oy2jSS+Ap6pa/zeocqqeGNNB42eMB1NIcXHh4f4DAm9PqQS0dnCx0qBqt0yg
G6D+6X8hthEvqFoByIDGWTGyVmQnH1u9FytMSBcIBbvgFrXvmVmuGlC/U6ocqBr1CHsYUJe9Bd2j
uLMNnwqUk5fRcaiWIFLAH2H7aaMcziQl9eMp4oHoKCKnXXB4wjhCbVe7VZSDaZqya8ZYg+g6GEAu
A4LdM7lE+1HVQGMyJzq1qBVS05BxFlZQHqrPlH8AG0p77Qd2Mirl1uM/B9w9cKGD6+C64cDBkcZL
fCHmO1dRZ8NyGpDffwMHAgCOOj0yQp1mF1OLyKW1OIvUJARC97MWcv/RbIYqJPu9FV7g4i0Aqp1S
amunm+v2BLlEcxWeoOkyeOeHwmQ75VHkQ4nsrJqS5pnJkxfFDcwHLaeL081OygawsoxHUmY7yKMT
cZAMFJ5DmHazdLBEUDKysxMEWCKaDVAtxFYZWnjBa2cY6h9xh9v/sujnusCNlTgSLYWsEJVI2ou+
gGS7uHBE0Fk4nyhekt8o/PFSqcWJ9wT3c+s0ft0a82FjNYYXi3CKCHUJxiSGvHM7b+3OzV7QWeso
FqF3C4l7C+nfEUlkIeRqGqHhqSkCeZ67CprR19AocOOkB9sy2ZX9j3Baaton/WjUsgP1EJJXC+UR
TxUgt5PyeJ49clAorfWd4VuhpCZU35Gc5/s9JZDuqdxTLhQr1j7YByMNdY8efVNCaK5bfVAKG7En
f9do1682bszufWPNBUsl2AX+CJv+g7xdkavMwtYfYYRiScN9nGJvI5fuDtu92TC6BoSFGBuepVUb
fjh/wUWMNUHoeZ37tpUDLopAF0gac4RUNuhVNW9lt+uiCiwGXSSrPNe9Ot2s7mzjNx/r2l1AuP9e
D6lftLZixP2GVrSdBUOFnlEkAk5qvbbrJG9QD+5n9haTowA7N2rPYMBM3vOYHRIKsEmSLZ5C74Ap
v/i6Wlstsqd50CWIHniFrbTMuigOmtNaaR6rop3Ipg3GckcVfmOxVgUe1yPvRsIed4g6BhsHt3EK
V0U9ZZjZggPNaMM6Haaq5JVRAJ1fRX1SueTAaTxEvtfQcyD2ye9J+b8OcW1UZKO9kr2MyEscYa94
QncQiNkSsSfKJVjuFSQeaoVqqo514Uec02VUDV7BaDcq9pKPXHO1GqDV8mcM0FV3hvBolWULjunu
T9r2NfNLeR0/xve6RtMS/soVp1Nl8FCD/1ZmJ85qmNUYDq7I+/l2tOun2P10VNLCU0cP8/JI2HED
b7W66xQqwMksA4vk7bU9brnjTlje2Nvoj14WejGR5M4cDgDFtbuXDhFtCWBTq1iZvdMkMgTo/ktG
tmQp/1EtD7l+jx+I8psAIkQvF6brGxMwB8ZzQkHCXflzrTGyShKJe9VEMPP1Tp4GE3/Kb0bvDRb2
sVMMXEzb/C4cT4JxWFruI/Q/+9SLJL4Eyzuy4sduxHY7wVN8Qvd2AVH1hflk0jZMhKXwo4fzmTVG
iJFWYxTMLRwVHGpVlSLntQo8G50ZE5Uq/lqQnGbH/KH+xJFCsoPgzxExoHNB1gIDU7GVtMB2CKOy
9yHroY2yPG23dDH+Fcq2djfuMH4tITL+tOJuatD4mj6zridV7Ch5+/yG2QJ3MJBpkyhJRBGE9mL9
/4nBUlpC3/SBYTJp7VZaHTIN2ycT5zJMv7p9OCg7EzVdyZakbjowVGCr/e6UH8IKj9Hr4XAn7olx
zXP03BvfLPVhV8iPSMuTR1+O/707JT5ENpND2Ya4uGGRlQO5wJmljBWI6hHMHDrtIrS5kInGewKY
sh8KoYI5xv0OYGpQziSYB8ZtXamll3g7+JtvmnAJiIKFNk3xC66LFANnYDMyw+YHDTy8OvuZtIUF
Krpq9TosZPYHoGJUvQ/7g47+Pvp5PHe0bPmgLlav8d/OZ3zE3McstzRND/dQCe0I4J/Eox2i/zco
HGp3dr6G9XfTvzdFdOYeixxtUFx8lLxjh4fd7pZuMkIGe9/BZLRbdZDRd7qgjN0HgiC377SyqmkK
xbclRn+Abhg3FmKt+K7Tmp+eEWq35m1O8/rromKo73EHF3ZU35anOR8Rli5TMYgadQgKgg2w0xgP
5OEL92Wskv1gV52lmG50X/6WGQU9z98a55vlWA9A7sXH3akLRWwBLUfzCGVfEHDTjocpQmNGsiFc
W4ECmEk9zsGplMJA534iGjU2k6g2EBvEdVFqLaLjSRsjpSbogozMklYBB42r39f89PFw+G/Tjhis
cRRbYYX9cOh/Itc4DqOv2vx3AedwUYn69I5PBiy7eux/jBtPq6HIKHzdAMTk2OU0Au6WtVIkdsng
FjEbtYE04OWlNsn2fpScYmzheZcYKBxBK1t/JqRbAXLx1EZ5tMSwJ5+XUrCw5cSg7CM6qLHz1ja6
mVYtOCWjlv1eNwObrYvj/nN4rYwFhqT9a03kzU6QKuKk0JcJ0qujGqn5SgQLfIFZaG89vvxpzybV
QZ2JzlX03UWxoQuGfjPFBq7A/BSdiOuRb6weu+4kAFkIp43gKwHaDVJm4ODtenJV9U1gUcNcNXR9
1GCBgxxaJZyAFfIOdvXLOPxzlfCDMf5PuguA3Qy69yMrG4JHcEjqe+cf7WOKMEbWrAFPsO9qy8x0
6foi75Zqx0nvqRx8bNFRPi+/9SFfjsuqxaV71RfvLwhlwvMwi+n9JLl1ABjOJors4UWs7FiCviQw
U4UMuUCq5Vz4L+fpPN8sSOWFNPzJnYLyioBliaZS8cUlqmpsbS2VgzSZLTkpUsI7leZRuuEnVZIF
REKYd9KmjLpYXfbXQm5CQP/+0zilfOC7whOF10Nl1NJJB5QOtefaZBL0Z/XxCF3x1MFkcfB0mi5N
5G2t5eW8CpL44JjvWSmzlbu9lj6GKJd4WT65+ANS76ANYM2J2xrQBTRrIssBHUzFMtGsUojKeHR4
4nSQGKie+kicBH2qpM3ir/1iWif3G/zGG7lH8saH0Pfq1jFutLgi5V/BExkTaQz9SQrX7hZhMiaU
Aw2CjJijZHixS6j6d69n6rMquqlpq9lLbwMc+C/VTrj21ucfCUpwxKCaMMH0DNBXU2jSbS54goGZ
BJ52M1yuPhZ5RF9mZlszfWrgfvnnqs8TMCNRUo9uB1JtYFjxat14w74M7MIcTXUBPXuzDpvv0B1E
lhVJJRIBzYUISZHa/yd/xdj9DvxjYqvVwY6zaB3UbYqyD3s/THhluRiTuOGrBhmByoa0iEaY5xPO
VnQuspnRl2E20pn7wB4aC6qzucg+FRGEiQ3IcsUabiufRaS/EsxVzK0jLQTWApKsA4g01WmTWzvN
Lp80M4zW93mJHYdGfW3F38ESk44YzNLWh2S+5oMr93mcr09QjILnrNrPgFrHLXRjlgKGHYPXE5GD
+iaoxDu+Yl0e923+/PgCNmsGrhi2htkXYP3uuzW5PdCV/CgBzjdGqZIoXfafnd6k03mYaIuSg/MH
s1FA7o7PP1nmwHgHdnnPa8SyDV1pO2iHOtUJWzoEUWa4VK577/JIw3GkksDPqCiM2KtN/cK6Bdt7
YF9tF2eViShpUdXMWwK5Pkm9KnVpOWSkZBOkDrUHIzyC7ddlRXMFK1nrzOPb2p+LNWc9rcVobGob
OuZxaCTUduCnLW/r6rS7AXnSoa9hSYr3wA2LuDxa+zq/AqutNV9WXuhrcvwQ6IkzwEF5j+NCMV3L
+FMZP0JJj6PTrdmfoSqGlceabEHa9s6dX3X406ZfcElhPhY3TNOoKNy9EEspwATfaMkCKFlkCLZ1
DYfKmbqH5wAtNxFpezSa4obLy1hmGB2A1zPRdR23cwggQBl2hfS7bCgKXjhrLkSeirYVoAMc/fs/
Pe+LjpAmUG8OOKHFLcv2nf6GOEJcPevZrvdcFbh/U9DNERuRwIJQmdHjNFO01KApLENfTF1gZ55I
mLbMl+5vc9shQk7z5X5BAhILK6NPfZnIPnb6siQ2P5FSE3nB+z82vvquUOdwqHmUPKYOvtHFbUos
h4va55cfvAikdQLB0HEE74i+syBmp+a1rMiNfKy43T2oMe19Iz41UUZ1w/8nESsVQOtHDlNyZ93n
8RMrKiidjfNtRPvdRjX77wC0T9BPc3BH4W+y8aHMOlPaJEa+7ZCTG5L98MHjIeEZvdNEJmXNjuCp
ucKNTYFij0jpDmgxLLK6hz6W6LLRlxRje2MdMAK9VyI+wBVN1UdRfmJF3BK5ZYo4nNOiq/aCD65K
s4W2sDCRv6ZNhXtuWUC8hNxeoZ7CD+CeHsAL4bLjGp2p00rVZrrV2jKB1Y0gRzaiMcaLAScl/3Qr
h8bOJvocGCDqpKWbRUMyXw+heU3NqMlW3glYIDQt3bIOBCC5/cDyxQ125qWLRXgpBj8CDUtusC5S
xumHqCqX+aTU7wXyUEk8IDKLRh3f5o6DfH/8b+c6qkJFwkMGu1G93xh1bUUCiWIQs4tMDgnckl8/
6WLGe3f7po0mxNJ3AxKi7+C9ALS57XEr4unarg3D51+G/y7qYqT7RSu6QCCnvfQMNB9Ue5ZIcC2a
egwOkafjkxqNPk0DSXinP08etTd/g5J62jkz82LYWO871iFjTLRO7kFbCGtUSGxvfTUBgNZsbXwU
7mWM8zTOyZL7HGBvljmVd3GXTPmlxPVTeD1Yf0+b03BrmFoLpyq4XCR77jInLNI+tM/zrHdgX8ha
gLNr8FQhfHF9Z7WNDUVBUZUgTWVROyZyBH1buM0WmqQ5RH93LpCxX7WvGG5XotsrLdKogmc0HSHY
u4636B8E0z1q6Bq2u5p7IQFT9rKzJdE8AUT0g2zALonzo2NIg7KH2/e82OReWCacG81r28J3mL53
Tfoqid+D9B02DTzkzVUZHJlNdUcbo/oX7p6bmhzNKkj5dkZ27tSvEuUhaWoSXjjrxEFFiOFY0Gf5
4g2szQI7NI8mhMp8rD1gi9OUY/BGzav188mpyYiDLYfIq4aBd5tSPDswlydAc5W3SVgrAYMX78tF
KgjM2WuDAyR3mVBOLY2s+LwACgLtoWLzW9Pu6EGDusqJzoCU9f0wBsaBzGb3Pnx20hmTVoPArnX0
xjH7g665mKlgspurDrfcwUbqTbzsLgyq4vcDfDtVlcbIcR09T6vBhQXURASG2rfj1PFyvABM1GL8
A2bMBDILi2a5xAk8iNdZoT3Qm6Irs/vJRU9kR5xd35IhvC5gk9TNrQzfPJCla6pitXRZMyAyogF7
sWMJ9w8z7rSqhd5p18FogBpeYJiYj7JUfbfqpLAjMs1+wjexKF4H9lM9hccE97zoc7qbG3spX0Lt
x8qOGvvM+QnzTE1US7gjo4ghOdZQ8m8KcKy14zb4rQGfXm5S0Mf9eGWi5GRId0/Brk8JXM3b8HL3
8E7b7ImVYgJ/Lh+ZRuUPoVZ1+qZ76soxFw5pWzJq3rE/NvdNzYX+5P5LfpoJReGeEx091a/Ec1vD
uqxy7/RiQkwzoJDF83eJtn2L2hOAzme0ZVWo9nrgNPO1FiIOv123srgjyq1U68dYgS9L56AxNNFR
y6Mg3Ot86qLlV0Z1Kf64MfejHG2TnJ8D7WO7TGFEKqt+Tu1eNYk4RJ47Hlf2gnrxsJfwoMwFbXqC
B8p2vuB86s6cNG5ITPMNEMkGtompLMz0g9LXhvOsbRNwe7+bco54q6wSIIdfNIVVFGYVvsaDi/AU
6Hg5RbdM3waVofOoXbL09Bos7THH08sZ4r6xF+Q3ubtbmW56OyHRgCmLs96gfMJTsvjYRooIewnY
k9zyryDEr38uFmGUbjMplUsx8aL1osW5YC0yRyYhUZ6Ds2OO8/ORc7RwynCIMhpaDSb/nodLr73a
xUnapu9juLmOpsV+dz5hPqOj6DXmvDNqglV4M5Rb/Ks0LmlM9cfHiXdUgdx7QZW1gN7HC1S45acc
yzW4xTYbYrT+42CgHdLmr+ybmzSgfjvMBM8mDdGDDXaeO3bgt137NGXEma3QifyR3w5CmYKMqOoD
ewwSg78wGa+aBIfVca3pardDZMSoWmfn9Jcp+rL5ENzfpGfpH9EaTA0UPUqijRk940XurhMNYADQ
HaP4EVKmRZFPX5xJWNPEmWAh4n/c2TKs+Cwc0MJ+n5pNGe6EMhcQIF2D4S1v1TPFGBua85gVf9zN
SZvg1fDq5CyB4ol0lRGNRsBqMh8R4uZKNpdPNUtFXurjM4071dO5e8qJyT4Wb+ImLme8CL+j4u3o
+UCEGXt0OSI/z9Kt74dEjS0u3pnJuKx3ZNmVxwantreajobbTtAdrlV2NoP4f4/cNMd9iLRkoLSy
T2eXAIyw9rqks0YXbsZET90Z39DhshP+vpEZIoGWg5wflFG40oqm/54gnpghXs7XMI5hF+CwVlVN
zijSyuLIyaxMmdJ43/ryeJyBWF0IqMh0iU0vzSZczDYvRszYChISR3cbFilvZflvQEuelNAnKa2G
zsldWI3gTOOoX/nIzL+Pclh58Ml6LTyRc3frNJDYo8t1vuGbxkJwE7kVWF3uQoE5SO+TLwbix+pj
bPkafx49NKM6NnLPODVpRHYgTZ9n3ArHbvQJ5jjndm227w6NtqCfh8UgZOx82MQRvxmc4E9djOG7
wCMONxcFRwpXevsVKb7suppRCiJGgbXPGzoq1S6k5KZgAT5S0UM74nvLVvGonvMwpta3hSZzAdmN
7PYZC4cE6BxI5ZWO9km5RwJ//68Jq0MUQJuK4wRm8w609lrPTdNzbBPzs7pitn38UaldoOb6nXpW
yhI3DiCNVFKeGioNh6XO8kVBoEvQSQMfoeUWLv/OkaYyqgh238/XCbeifSErxmX+CAKDMDtzX9y4
JTRrPKXuh/AQhtAHURoWwcL7UMGdzLGztSxuNs9FT456dsJC4jKmrRZFLLzIhzM/PiEEfstww7jq
VO9pTQ5OUNWqcyrXuy2D+Ec4N5taox+G0g/1cx4gfIDD3GpY34Wu+jlfvG1yUU5VgY7KKXNR5NL+
vStQiAVt8iocNVqvr7qtd3rhxBS02Y9LzkO++EYMsDqY6UeO/tKrEpMt5fA7XA5Bz7RgEGuIxoDZ
Fo74Ibf2IAUXZcZM3OP29A4BYeNsIWBN+uR2YDwgsi9Wmfc2pU5/1Chg4MEpTbgSsONLK/w88Csb
wrbwgZNlQLhxMoDxLayhbAzh9HYSoOr6/+w9S96+QLoWF4Kqry0grFs1/p9krGJjummdp8Xpos2x
3btuUFyDtcReGJwUmScxUx6m/+3JB4xFxaL0W40uk77e5cgACjwjLe4uEO8ssNUGOqgK4BKhAxKE
rGna2ftfnBDWLyIbQDRvNlpQTFuZPGJPPZlk/1PdJR7HhYxTMMXYZq6LPt5eAbbmkYIkltK42ccZ
TWgkIJ+9RqfOfGx15Qs+GVeTXXVjVVfsBL4c1pt9EbWIDmHfGwD2BGi78Ir/8bFMxoRZ9LS1u++B
UV1h2PDOJJkO5IGC9MlsmRnW96nS6D4pAM/o1wrTF5ECxG8xc+XnoS66Txameklz+v5qgaBULRNO
03hGxaSjvh4TMHm9G4wGpPyT/5LluT4v77QaB72p0fs2YnVviolSMOIOJqpFe0iT2LIHv04I77WW
dse8Po/0dUmS8bQlKFQN+s5YxnAh2QmrztGb9aHUsPhe67vHW6TKN0zgAm+4SvMd6MtDwIsv+OQi
OQBdN0MBzZeUJfSprDPBqWXpYvWSqyjhmElGMVCp7pTaYPiJvsKQHF6mU7Io9/usit8FqnJmzMPu
HYAkThgnJFYMxB5ZjY7+JkQdNKt6LgoJxzyK7hZWqyOp0bypdUGGjusJEmh/O2X2mwb1UDNbKl7t
F1uOF47/tLgguzl8+5q7+JkdlMD4Jd9/BRUIHhrI4FbT0Ntbtl9zLO4i7fTCoMjYIUlr8EJieCyd
r59dy91M7qmoBV5n37eMKA8YqPhRy/YJjrEP8xOPqaTP4ymKNAUTSelldIo2YHsovz7Y5+bbsUHk
yV8nGfegp2iWpG6yi1iJnHq41zxduggKZ5VCWcbf88XTlP1XK0rhvayyGunsVVsZJ7p4Vg9Js1Wt
Kmk1GSsEL0PtVFJxzl6i9m/QyVduKwU6ZE5aRtjWAZFm4LCUFdhMJz07sTd7LAIpuHNwOvdUwowI
1iD1SvUdTcE/5c4bZ9Ggd1QTRxWePb/GA19CERYm81oQjFxm2W0uXJDf6enH35QF8nqyZ9/iCOCT
TSyDz8lcm+2eZutGV+pNdoj3lyWOtPNGpkwjGoxf6eTpgPkt+HHOF35qy0XeSb/QGZkRXBuXgIsh
x7e5Zm+WCUGvlk6dFY1bYoBb13yIebml63AizMabRPDfukCzIYScgjoKjPDMbFFSTbLRuYVlPzR+
YnC2bowro+YKBGsMB/KEOmCJlbfXUYH6i9lulTGrGThnhJnlCEUxULmT+d/tXTK9MG7CYd27A9lk
Aby/5vTIeIBKSAqMEqxWfSn65eT3wazmMSqxAqk/R1yyPM3JM6tmaxiKlqYUuAakfMRRJpmmbPfU
1mYFMAv7yCnwGxVI2TUXW+82O/XmtO+gQnzYmkqy8JoRrlYJe0XMkk+Wt64DCIeglN3sdY+bpz4h
zLBH9rYcbEG7Skwny42Ihe53LhBVSEbjGTJ9lkTRemc3FVKjHmbRnPEWceMYrmwfiGT5Rp4Wh3iY
x5M2dLV3hM9lc3gF+8YFhaVMWvtQoZGAIKK1Z8mSA3SJc0spYc4dYkOWUgJ1/O5avG/9LUuzoxOj
s1VtSInhouhukYr/1V9wEI4h/H/LQ4ejic+HBGyajKRjNi/dA+QoiHZ+qOIHB/dPEJEZps0dIuJM
mQukVRqGiVcI4sa8uXLTzOv0B9kiGIv2SCcl/NcncyTYM59b6SdyjCRl4ijFfOVNw0kjqkwUnRHw
vjQqB7l1RUiJywUqfZsmEK6Mn0wx6NIxjDqTu12NV4B4EgkjeC6yQZgI7HcvVio4k86C5JbxK3Ga
JHNTpcnO8EAa8Wb3BGI0C4YyigUnuFmq4RgLFhf9r5TkXGuicuOCR062/GVrvPsl5yb1yZ52LYhk
QjRQ5z+5l7yH0UbHkafCrrZOAI8CYedjGMSXf23vziZxaml5tLCtKFuXFUtTDBQS9wP5USqmNr4t
wf60ENf3FzHhM7nBsb+HhcD33Kudb+u2gRMgUtAtE+ZGX4Zh5au6Sz4kG1p5UALrRN16tFaiB/Cu
g1J1+FcjhDkEYMi5VGqXKp0YwqghsDSozElf9k2zcV8NrLcD/+2ed0Dnp/6h3oiyr3nUdmP1aogy
+jLgc/d3gupMzHYWchK6enQnmwDNQsa1WtGdH25yqetQ5oeWg6SWVYBOCYnSmor8WIds1L+Uy8N/
gA1pTilG3WTRj3dJkbpE/fZmezQY8liAmKGgkjDLZtNBN2O7M62ZBQANYgY89E039PE2F93A57V3
vz+yI+1kMJghZwLVR7hULtHdGREvS12GwNAJLT8ki0jKxC5dgcNxSrc1fTvlmbHFzmdmi3bBaFc5
bGyXeWbf8M1znPedrbfL//9r5SKnITZ35k+IqtKxVlLfB7nN6BgkHjs5imlCLJlj4k+QObTe2irX
nywHGdoJhce+FVINlh0JNOpTT4NY1h8viSsVEhLxxKfLmsWB6D+RkHEwDNNH+gn/33ZS81KpO9Ka
KJo8Qljmqzyb9+V4bNUUxlH7WHqsyH6usBI68lHbXc8e2tClixKlOvUA02RSGOoQ3/NDeuDkl95g
xgLj5mDDOXgWYtgvyRNNVXKe2o5LLNO8/v+bidtNJdaYclyR/2cwgcs9VJSVh18cw7rEumga1Zs6
eAaTMuXrLyzMQef9T4jg3AG41yDwmXwbc8G0tIHX76cydnSy/zJvLVue1GXg/v1HNC/xNrxFx/+m
qN0FhJQ5mJJco2Uy0ugvLNjROoL2JYqdMH4a0Bk5n28NQH2+n3rFBAVh9tjp8MtLsD3JiCYPweaG
6esNEX/2BX/xcF+/h8woxXLTG7CSMLc9GpZ9WdEb6wFjMfNPrfwfi/yuYrU8rb2y0+RibzC8CGd2
pWIcjHjt55+uS42SY7dweQtbNr4Uecybu/Mtza1pvTwcISY4DI5Y+tW7M5+7mCcpsna9jjmzyZuZ
H1G8csb5nCGm8E0uGBOqGnF3894AaPeKkRHD9iRQ3ewBuW4hJIRM9fEiviggnUkZlowdrH1oNwgH
kInuoV7KHugg5/u/UiggdnkfgvN7euAFnpYkgpkXf+nS/1LMi9sHVbXDlU1zo+K8n/FzvShWvX5f
C1Nzb23ngSkcuGMH0hEhFdWkmuQZfFoeqBGZa+EZcRvF/giMw5+cFQkfOe8RXrTRIuGxosELjwLW
vchKC7nSe6cMyS5XW4TEmUYnmnf82Tr7XIF8WkoQPMu+D1IuHp/dD0+sN4JDPF83VGlqzF+jcwZz
CiNxCKB3dRkqgWhRMv/Bs8an5fK4yuQEGKLcw6emI/BDLxtt+s4NRavbs4UsSl/sGww7TnvTQV24
fMXd4KHZzdxBZen+I8Ay9fQkv4OBJlKU2MOYYvFLDSRqO8usp+ynpLdTKO1e9FRcOgToVEmmrMH+
YtqjYxr1NShHGh7pHXz73yzpP51Ip7iEoJIEG1RHzY27pUpTxgI40UyewMe7Z7zsA8XL+jyTK2lC
gFLaqjyn5ZB5EU5t2iAg33gNiWn/csGBFLhckTVR8SfbVnU3sm2AtuaaBtixYD1TVoX1+Qa1x2Sc
pi16WUpP52zHq3WMs/xmM6TXP8omuwBjl5ZK7yUbU9zV6rjTW9FzoYfaBxkODsAh2Xqv+WfOv6/x
QbGA4jpM8HjCUaT2POdAQMIuYLUgzYMXpue/Fq35FfIHtQVzGPODAgYRhq3V2Jm1qHzhN1rPBEM4
7ZnGQpv04AR/3w1bqKg1apV9DN217p+l4fB39Z+ME8jtgo7iKA+5P4OqITIdt+pa/vU8GRA+FUBi
/N0OfY32mn0oA86f7ogBhnU37eVwlBZPTLIrl2VhIQx9GseGO/V/UEITRnEO2ZYXBrcxuqibyhny
PkuEsnvxQf5DLAXXzp2LwqlHHawuUfxrGME3wt+hUEYwP6bCSqZ4ggt0vM9Ym5GFWLweTk2LTxCn
RWEk2x4VoM3yMs5X2SPsOOKCiA+73QGxVSly8GVRYCNQ8CO9PZFVXV4+1/L8SyNFZlEGRXFxwyMp
mbC1c1k1v8hqjlbxbC2TuwaES7EfR8KG75dI/GDhPF8mXtsh/Lhat1B1+jd8u7k9o1goRK1AEuX9
oivr5rCrhfPpxqJab88FEfeAaM4DU3G0szGT89FqxSeI0G3PRN4lGnG/PWLa+xFpb7C9DDiWXOi4
g5SxV0OzJCMeeUvGJYKbD7EO0FLgXKa4eeJUdK6cWBsMm9FK0MyScGdWcuUPhysBIl1ZJLXkFJzn
zyDIK2TwHYWvBI8Mzext1XlYW9XykDyPQ+59wtn8kCcAHimYREgZgMQVcMmAWdIoEGtzj1CId9hy
vqssmiUfaG2BgNHD5QANexoHtNDEqTPV7Cv01pRidTanrVCzz0yaEZzOxmZtKDz5SZTu0mKs21Qu
9h78HmHaftu8cvfd8929yDTYkqIEsBJAl6LJ3hEVXdh6cZ6HOJX4wniv3C/w80d6s/hXTSBHzwmH
ifCJCEzmY3/S5ewv7z23gmnvtuj4aVT6dKX+3mwKgjn4J9OP+xl8hcteEFUbgW1SYHealFOBo00M
d8Sx4lVznkvTjpRNy+EFnBhlXSLZFqkuVjAr9xKVm+Ap7ZRqdkuuexudu28BDVzEDgNZzG30uEVI
Xmp7d2g6luvlnZJuG67JXWl3D2c0tJ6X3gwQh7NjNlZfxWcs+3XHRMVwyH6Y2uhQtjxRHob99ayS
gNa7Yed04Go399REcCh5T8X3TC7iM6PLNd2AlxIVLlq16Vq9nApfoaQ2gdiYnkjT3wegJT30xrms
zlDmh9EbKBhRn4aEAy28NkYsST2K7WiNkpP6fCXlIv9+BZQ7XgJk1l8UOS/ydVJ6xu62rWOuLG4I
XlGAjfKwSAG2h1uIt01nYbairHreDZds5zqlovchcez7oPpV+jHUFQraW4Xbn/jfB8/xhyFtHKVB
mMXw6D9YbghP/niTQPgo+W4OICAQKJBZhMgsXUtMrQN72TKprZSssekCQYOr/dq24N6s4QEqTr2x
L/JCuyOfH8DQmHs6D8+Gh5ZNfxkfbacKE0ac9EDqAkS4rIv8lUgaHyMVVZcUfIl5CYMKu+nrSvA4
qJL9+6VloNuZA8P+g0B9PZij4P2zd0Jm1yvkrWxoqqRmuCv4T078vRopctbYU635F3ZBuTC5aqMU
QZZ/fJClfvrkfGlzqknriNS30RevVgJ4RR/OAFtvuwUOb68qm6bYLc4639qVWsdFLZavw9CmuX6r
+BKyNoh86h+UkIxrCccc1wwpoz/41x+BBw6V1wMgVRqmXBADrVQkFOJd47ebajyVLfD0v7CFal/G
85bCHll3ZYTkmjE35xiOYucLZsoYk0ER9Y1Owy+aWbBc0VL13Q76q6TZdwQIMSZzq9OUD2yIj90u
CsqoB/b1vhTFWTIBF8bmcmO5dNa21IXIDPhv8JFEKg7Gy6hg+1tMqC1Uo5wZWQyhXSWRZFJZZkJc
jZk2tnVZmoBtvaI12wlE09XUgbSPE7ssQC0zi1cpYPYsATI+bKWOnGa8t0fYPQzfWbRPhjkey77g
n6lOTnVAh3qs2ejU0HR7vQiYccihOVCbpB3ZM1ZhDwPfeFymLCO/Bp7X9zFKQIauRzRZPBQE7Xje
FQMjmREcaQVJaX/73axVtcL9xNDTywRbugaS7HLsL3obfFrNRWeiTKmKSsNTu4e/vEPgs0naSIMo
3gtPRRbvT40R/anhSCPKnGpes4MOQ/IwFMgSSTDEym4ur3/9cQzE/86mDF1X6VqsoMqQsQxxGcvA
l9pdQFD8AnN6ONEcS+BHLRPz5RVxuXqL19pkEO/5jzDc1orWqFtEv88CVFcf0XHx1u3xElGPVn8A
LWsxRU+oDDn+VgiJ8qJt1E07vqFTrSMs7rdfeo4nDbXe/2YFfItRHrUs0/bJQ42Ufe7FnQoqA1wa
aTz74ilglZdiOw3vxxT97sUGE7efBLT34p+z6zZBm1k4p98Y7dm3qmhzyoKQfq9EdeYTkDjzz9J7
erieHEt8NuefXVqc0Ni745KrmmCDgMe8oTNExqflxNaEg8wfSjZPWOZ4IgyAnwzk69nSHcLccMjg
rArBLAZGdmo72/dMX8OWhY4FclyLm5qlu7K71vmXS1zRKE9bE99fGmuEPS2Q3NsCW9MJ4cSg1voK
pvIX/3gG/O5EPwhGrT7qCYO+htJiiscmdqotJR/WBB3LUzPwNXY9+JAyOCl1APpmlgJkXREC4eDH
PLAaTXP3ZTIASE0rCzK17rER7+U4yDWlPxxkez6KFuQ3esHrUtQJJwyXp06GqVtBnaTUf4S5gutv
G5RsaWtGVB8Rx8jK9+XybtfL6wj3CH0ad0HVM0t6EgEvcOkpUbxmR+CP9ddi8OZWY63yzGm5r2I3
NS9T4XjECx6fWqBvXPUPBseRfMT30tZM7DWJO0J9CzALhVxFfH1RS17feajvEBp4UGjehEHl+81B
7XXl8z03jFgzgUjDKjYahJxeFtidxS6rUDzMygR64BnPMWuK510zv0iZH5bMv9XRduWwrgEjRLdJ
sSCcYMgXN85DfpGBokJRgPWmA6usn6R2xjVvvlZn+DnSSJh/Z5I/+g88w9NBUThRjylID5PEDovP
Vt626s9vBJkYDKw=
%%% protect end_protected
