%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
xjdbY9/v49pGN8ywwV6vwZmzbcdLRFH19GJqpQkXvoJjz/FsWmlGBTenLA0WuBQ2GTI/CA4v5m+T
yGBLZv4ZUUsbgH0URmZ07Hj1xPFn76mZZq/i0Wieje3uZiR+QMRATf+Nq2lJsysJmfuOHxUIdj+p
Z39ENnRbm8m3EzxM50ktm3BCdXgD4O6MhPuuC57ikc7W5iatRrD5Kk/fRU56tfH0xcroxDiB/YhP
0LvkcdfWLein6z6uMBm+1ULSsSxlnYCkCXnuXRxx+qj92mxoAUExWn6AeS2MXxzdQtI7E3KUrx15
rR+SqT4x9MT4+C3xsRpxmIEKSIVbMOXVtUUeWg==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
nWUj+zGku5OLxPsU0eSgPJMWO5yB/AixuayjJFLjSC9v1j7EIJdKm+pJ1rKNTOJuEUxipzQLWaBN
x2mGO735N4qxtR5jRRr7e7PNeNUFU3j62HFVxPNrc+okp4P71p/ldBuz0Mth/7FF+gEpz65gHLPR
xHr909hs6vKr9CU7KRWaeTYtAvsoTA6yrKfBX1fuKba71+13h0dLbwSzUWOsjPEiGCwtetkiEwJC
XpufsfYhzz50hQoDun2EO8/VuyzzBMZTaacTKApyV4T0DicW35o7OqJ5CiBu18Y3SBfVYU+1wvcC
kNU1LqqWZnvWtsMQD6zhXhgH5SpsnUm7LP953bxJlgiC82CNID/G1pQKb0LVbLQDSZsblX6dpBdM
ToE442Ov/umDbvJsHM+meg4rW1X0tmqNCj/ZqMcZZX54uh7AsC0T6gI747cFgAAitinFoFzY9HWr
1berF7ZRMCCuaan/UtkDkTfH1YMCqcyRCosjJmlFh3ehwLHJtxd0jCn1CjeHKlCwcr/1wms/u28Q
jbL0cDfLjQ0Wi5k63Kq06eIvck72Pc2Ye9IKIGLe+eDZ6PfHK0LKXQGMHceNPRum4JI4BAL5SbQd
ZgeBu7AugNnxRRyln6R4fXFSQ0w2AmsWpPcexkqvnvvPOAxoqZZ4FKDxBU8D8hDlbNBCAoZFMFJ9
c6YP3sfTbQBr6ZFvDN5MAkJRXyDlj+oagvfO+0xQf2GBUEbDiDAiNJk081mkA+JXFVxbUhO+VAak
jNPwlIjk+rqFq3OfonHFOVYq06gPXuR2px+l+8IONPJobH0xAObnL/d62AhGEM6ilObaG/1Hxq/d
/XOwEiV7tfmUCM7fxOAuTaJixB/0Ayk22cAlDWxxDpzrZrRcu4P9GfBNC0AuDmoy0sFYKe0kDvLY
QXAOBe9ILnW96XVBW32OgvYqOtb47rt9IOfqQDIzq9ZDe5v2rJ+bGbj/CU7/w4oITZhhXCwKo6xB
4bUnh02ySeIgHnI6CbznsQyx9ktoFlfDjCYksAzWAgQR5ta03aYXGMZ05YWcSRAjSDSaaF1e5jHY
wVeRPlzQH4TCPK/+LevzcTHspddawl8cQEZfFlJ/KUmUBM7ISEIKdwuR6PgvYYxi9ApWvbMnC7Yy
+2LbFQZpVY90X7CBjEEWQa8LI04i3hl6ZJ+ymqVpHwCSozO2+Q/wRHgvom8vYl8C4cGtrLrHYNzO
OODB+E1fOgVdNffFqi3xvOS+/tbFTkjcAXjyPPdUnFjWfU8rX48YIO/7h38L1dwDUhFkveq/H2L8
wtYQS17nVJRMVBEBEPMjEPsdOyzY96x6dAfHVz6in97z+tbXNO26fhupRHgaklfuyrjL+CUIfnsE
cf22cdetnscpRkvVBW3WhKZN1fGfZxCJbywplMTPvEIQIRBoOpWiXhahQ1goLYBbOeXBTb/aex4f
MRFpJ9UEDN2cj8kLfKElorHvi6wOujf1pBv5/LPdaJqkoFf3uvC7IG1x+X705yMEUYKE82o7ygrl
mvFjJxHiHyIMW7TygbKIFdosfrojY4YZ7wDYdr7viChXHbuLeq1hlF28gl6PHkiJBK4cSARm+Lpe
jDp4WSCIJb3rUTVfNOXUXcpuR/ykJBxwK5ZTQHxpTo3ji79nZwfrrgcD74lCw85V/rJ9JQl1DMjl
+DLJTE4KphtuFp8fzrt3VjP+zPVN3bI5gnUliatvcGw7a70h4HB2NZrXO3pb01kuyqwz6pKRrKhY
kLqYFwOE3N8uBoRX/t0qHH6aC3+EQ7BIneLuBh2h8PYhlgt5tZXGUaM/7tVdRgPPf+XgKhMNtBdR
JezKc9HC6XpwYtxMthnDWZjgJRl/0IUlvztxXmlSDNuL38RRgznbo+ga12S4tl6ZWq2UyVQWz/tI
S2Vf2uyF6Jhf9BejoPErXFCqqs+FnbzUWQT1e/8M8qW9DqBwEmtoiXAod7qMg7mkcZmhMQ+KHsKv
GJ6sJltqinBqhPrEo8AOErk86SWh8GX2xXecUqp6q3JGwfH7m7dAv9whO3Z2M2MlP6j1B4NnpzJj
CsXb5lVLuvECh+mIaXxQbfghtiJz7lkHYDfOZw+Dgs5bYYezts0l/VlAy83xaOAQ1FHLaK0yAM2M
9L83D9ixHwI2BZp5yxzEe3+cL7CU7n+XIn1p7mnZKcPB2P1JWnHD3KiWA+b5N+hvdfyd9pN4uI9u
oN/U9xBrKIsfMYyazrG6g0YTIO4cHgHuLSwS6lR//ngLRWlDJd+nZJfw7pw/nhYXspKoRm6eX/YT
RgEpYGkpqLwO1eA+UTAv67v9C97f76nWkriH1F1RbANIvAS6yJ0igep//iiBuHbe531lU7fg4dXS
bwDiDMHI/9R6j8MUk5mn//vZczE/hpQdktZAYKkGIj5RuJWhYRw7JMwXQdIGEisLa6Rmd3Q9f8Uf
l5EomtnAFw5Ys/9ooppTcLdYbiLeiX9mF7YRDJLdCK4fr72yHaGYltCZoE+oqP/2B5njvft/FxsZ
QcpYPkEeFFrtxzYCymxidleGm8IAdVQfljNHZsjYUshkHeLinf16GA7TZmoJVyT+QHEY9Dyn5FJV
rIRgTJbkw6l7jfr1F/i3Yo64agMVj8xxkcP2lsEsgaOle8qWRvu3auMGDGPA745xVdNOPhqH58aR
MIroLWN/tHBm+YCVCV4fkuL7fnR9yiUulOn91si0fXSfBc6lKhv/W53bWSgHL89d4fsKSNP7/YsL
VtDmauig5hxU3s/Icf/46hVz3aY68ZDnhAt/B7IB7yOu4dNiKNXwpOjRweoWllwSnRe8oXOtpgzz
2M/q5q2erqJSMjYS+47nm9nVKtBl39U4HBjbTGtFU6vrvpp7PeLM/2M1d9bx0431ctHF7KXCjDTM
YzBlvoJKUecQcfy5Z0fGBYm8H6SFpb4OkYDi/jJPamGABbsdEbx7UQQZnEBFHR9mUHTWn0nWpdi+
7qDuo3qHh1vhWmaVYql8LCRIAjKsaurFtKfHYjGNj5idepGl/YwnXyDXrpZUTtKzV1NZQK13TNRN
cvp6Asss8QNCTZHa6aJkQTqw3kGb2L6iDNsbYlyRe/717CUH2ni+AYa+dIY+qF1FSSPuntgbhNp2
dp6YVq59KGoACv6+yzHDufTzNYDfsPUjMwuto+mDLX8gLsH4xYsgnrBRxaz1+e4mcNyc5uYTf+BX
z3XqvWiSUfg5YfVYPc/QlCogIe2ABxRuwRIQH1rGMFN+TSrJ9MuQbHyzxNfBkMqURWgvXoGnp7At
ZuNM9PDe2+UyXqmsGeR+VpEKcilPB52pCK3l/9kxeovryZRs0MeEcnVeMzN3JpTKd2ZxCKOdt4/u
WRnRfcJv3lFvu2fSnLtNFWFuzauU+QIoQKO+yFgEIcLYcFgofEfWo9A5AT46Kfk74pdST/Ztod1P
AykILuOq2w/og8sYC79b9hxIM7FO+teY0BPe43m5N0AdobopO0UF2/f6X/+JdOnZ3l9w+qdjLJ6A
kWlGLVUsks0IOenmMisBrqthNGPw+rYK+ySoq3A93ZL+roII/+5kUSHE3avwb2xClM9aYtKxKlVK
G15oLdDF7jhnWaQmolIPrlChZGMIXEFFrETPg2gd3HW3ChPAmeVNc6Gx5mmZhiz4GU0VStcmyBL0
HoDe3sTyQsxnkDVpdj3vgyFdUf95d8j+SLyj8LxH6i1rze7VudMjiqtMe1/6uWio48RaJDy+nhKU
95MIaIOFl0E9gFgF5RPWFw6wSOWYdn/9tRf6+bOlpxZCzFx5KiTR+GU7RU772LzcX9kvkDCi5TAf
QQMgApGEAcG9ppkQBhXXzFNk7TrBQxXtWEMvUzg19t0GsM5H5dGrX3OdLH56gg/KAsw+hJsfaS9D
D910ndO9s994pgJxOnSPeoEL+cHkWCoecgzgpB2FcWe+1Q4iwfSBQG5MeK+5fUv+GVzahFGvzU2p
v2qjTHu8/e3O7tC1UqDR8HpX+ya2k9i7Fwxo3i1K8VuYMDwTdjbtN+BXCLbJMO2Nd3N90wPEFWTJ
yVvIzToprabftHc86RbfhYPZ8CDyVLkCxyUAQn2jB8Pf3uh+mmad2/gzmVhzd7nD4nftakqNVKRL
ZIq9J6iBEe6xHMKLCnJBmDIr2DrwHkuelQowPQIYXSmS3WJnq+9lqycPoZLU1EmxUVtfKrBG4zB7
04RlmflbNtKSo0Cn4oy7K/PJof8SQTE4qE7BBOy1sK2oIjfdI6c4J29MQCjJFvJJ8noyRUjOUPkx
KecX2LxKnXRTCkSdY7YpTgfgKPC0ynCjZYP/syUNR8HcKC7sQfURMt3TW8VPBYwZGDL8OODHHr9s
Up8ttxsXysfx5CnmEvEo73yZu5RX6fLoZ19tnWTJdF0le7Wz/VI4G2UWZTqqpCD+eHuMjCTzFhfb
eHLgEDx7tP/mPCCgUOyDxL6zlVgXWdYuUOaQwgIBUp2n6SA0+UsJpXGoo+ZOL1WFPS6FCuCWOZCu
Y3v543+iuMl9sREQHIRsTXFldvbVuRNsNOUXTTsritMZVqjpXi9xNOGamCkGqQ+e38aAnylqVrPm
Dkp0jazHvrTcyZgNEtlX043LYjGN8q1D1TSBQS2qEWYJNHGG6IxCF+P4zZ8ktQGGnCRADYLvIpAN
sGWXnLRkvutmbWzTsSwaHYi8xmwjkEru8/UvUALo7uL+nV0LPN+jXnUNMgcilHVIgM1nEymVm+IC
+HkXbsrsfzgUU8EkMlL0A9o8bTlwXjitLOUrWSY1m9Slu8zwCZ2pmbxN/jUld7ozx3KRYLPvsaBb
SEmmi5b6ULsGLM3q3CpOcNomGpKzObG7/ek4OvX2AOdooPJyHliWSKNtCQUAkdjDspWMWroXsbYV
v6c4KvuG0GoYpLj8ieUJP0PJaXmEJAqMnz+cgKEh2SUqKi4EpzOvuubyhHRONrLnMa5qhIYuYbhI
QZv3TsDjfzKEyBG/Ews7YHuOXggl0n2g66oFuvygRqKvUZbJ37gaOzT0mUyVJzu8ixPqAcPxzW3A
8nON5gRQu45CW0cFqmRqWWwdLLTik99sfVRS/zlTSriOPsqod3ie+xZFTSnnFS8p5jTQcycVQQ9s
i6VdilP8ehVj/epFK3vdOt+fYGNRfzvC/O/ugiyVoDLAGZEwZUm+ozPQnWOSsM7fKR/pO2bQLaZg
NSaeJHB5pxIdVOqygLaiYmtol7F232NJymnC32+sYbgOxm65JWvzrXWbpFPQx/4X61LutsNt7zWk
63zGPv7akiTvZ2mlzI1a8lRUq02vHcyUyp55fCbuII69DGmFzwPDDWrx6ZXl7rLSRof3b8iZRLoA
vYpOheXmwxUz+1ShKmoetQkdhTY1fJNXDQQ/Yek51/8yaTbPEjWIvmB//oyomhZazD6QvtAz5X3r
TuB1Ehef6+pbr1mQBu1XbcNobZwy8Q4eSaihs/D/IjOK0H4GXGxCrYBdy0uXBf0DfEkKpv0gJlGV
OW8UP8sRmNotR8eHRlksyG1pNNPuhVIqsEAD6uRT1B5sKo1gtB7dGqcn05QAGzHdIg5h2jYmZS88
cCR2osV2ikaJ53/1MWShDAzuIZMck3cwuRKEv5sEE/pHS5051i99K5mS7M5Te7fIN21B0jvASubY
OJWFNYH7vVRFpH8NmK2TZ5AhB5yPs4SU3Y08XZwVE2QMACWHaJO5NtSjskjnsYBOGRhK+3gxFjx7
GPCth1gPwCcLN1fOUqMfFPeqB3SEE9U3HVAfKk1xBrF9y3RZo99+g06zc9qADu63FiNjASVb4Oej
R+IRfk9weoPFAxuxcJZRVmLAr+KsBNaVw5aQl9o7JUG49vD37eXfDEaLQ/30YA9BMuXKUbtWcKv3
zHgdd4eTpkIUD5/VrXryhLNfVnG8Z25iO3hrkIiQBaiw74OsLMxc2C644lkSgNcT6RT+RK7j8KBr
/n5+Z1Z9lf1TTrmYd1gQiyUCAvaq88ZOr3fGkJD9HAP8J8XYOW2RSzvlhw4lHfHStJ+G0+vZ5Thq
C5H9uWMMvsIhXO1IMWRdSXrVPQyb/wWynwmtUbq4Hx710GSstI3/ButiVnXTAKmIrO9ef23wsGyr
7VwRAjgQQL2iYGzdeIbC4n+4GkAsdAcD5LB00MQBTe7ftpb7lVKrlVRuc0kmyup/WURYEyl4BdU/
60m9sT1+IwZ3oMWqVOFxJi8/HWovNAbf9RNfCDl1e6MA/1u6Rh6AW3wM3xirv0kjgo4602VYkaU9
VNeNtgBdTN8+Pffoa62YSYs+2yifolYgb1GDim5X66UaafLbqKXXcXuJGN2DqIEzNJDYEPbgvnva
Y3UoSbnrn63MEKvNvr6F7HlRczR+GL6qOsTyeUuIsx6RnxgOy91wpeLopadpfuXygjmKWgfGotqk
vDORShec0YShlsBJ5DrhmVQ76uvmm8fUf+gMb85o/acoStAHqschoRh4R2kg3yg4kac01irocplk
ftcZgMLL+IlRZcvnz3EH9HZZq6eUJ9HA9HL84fOwM3u71Ia0Bo1iTrgMl355ImvCpRUZaUepWPK0
u/GVAnUjuxuCnidlgP1siB2FYKjfPwk1BcGdLXxRgV3DycwMAhC1yp243Uth0mYFYmgprEeIkq2i
iPeMDl5dLr/oM850p0VWv8QiiwPsxOC6580m74z/njjozOmsipMoxD/k51V2e+fZ73REAqchLkab
+TNZ8468kIXbzhjQpqOBwMIG6de4iH/d6I34J+rgAWz94pXxy458AEO+ENaeG9nRv/hH2UmZVtPm
ItCbeltf2FeB8XeV7iUT7zQsIQ0MPecFIjNFSb4YvU6rQxPVIebl1rvQlD5yBainh2NMiigX2D4+
Mmx125zwT6Pago6whjX2yBd6UFJY0BSkpFZY81CYw2ILkAfGDD3P5a5yAgBFb2iGg8iLp1vWxv99
HyZdIU1UM9mse2/Rv7K5pwU7iO+B/0+NVFQ3pnaQEeNIPjYQI7f0x2rv6QOOyjGHbbOhy4fO35HE
TmGg4/hTr89gBE/lEPB/ZjNKAhD0wvHFaRdSiFcGdIu9lCCu/CxS48l6qbv6D6p7LMO5qspiEfY9
mzG7124cNH1FRIpVPpXmZvu+TzOIY5jYoevccTc0Qm6aAbu2nCS9Ataoqi7RmYh2+VE1hVdKGcRH
5y2/LSQeFLBHD9c3SGW6N9XjNh9EKXdDh/4RlSopXRtcb11Wjkie4NSz4rUwF0mKiFKAu4AolLXg
AHoLKZMyU6saKMXbBAyVgiDR4jUIJDC4VAlF8KJr9eLnRx0GW6o3eMEya89fZMBbY5xW5SHSg1+6
BM3MQMr2GBcrt6aEu2s8+bjIbxmci0NMWE6vAK5TYq2ku6DNvgz87/VCLmT9oYipdKPtsIoRF8x/
pAmtc0sh3rRQ81d5+bXfhOO/nkpvx7lFRqIP8rPerNehs+FkEcwiDYUvsCIYo0N09BnB0nEdLx10
rKbygc5CjKET1ltk2HPFH3kwjVgST1lvqaNFTgtq5tR+7bDZM4vv6W9UNXQum73yknZjkZySrB15
/nSjHfTUqv5jczZrxLkxomiL0p9Pw0JjnpLtFNc6a1w/zGjMbXjQex5Ly+NJdCxHtznVe9HxXvVN
70RHXzn7yLWnz6+p4dON5XVKhbgQJIui05G9iqnBq9XHINtCniWR+blQLrKug+jAiB2ynvi0/uRl
rXP+qWeZKQ0fMpaqbWDkCRtCw0MbHRSma1kOf7+6k3QyHFoQFYbzB6u2BMNaIQm2fq0ZeUxeQgb+
szVf+Qvr/jqeVNKESV5cirwtgTY/PYEM1RTeAHUq+6k4GfA37m1Up9u2ZT0XPcRrxqcS74+HnEkr
XJRyMpOEYmwGIE1nWuu0NwwAjTuGfRUFoDYHUNHQpdPIWBtiP+yHdbW+UFxqc8N4M6tbPx7hhgsL
Kla6abgdBDu3ch6t9KSJLZy+H9Srxpi/dvPOVmfRtGHl7UmknGIKE0X0yPerQPtLTFa3GJFqV2QL
vg10LpuFZaqyEkWW1b6bkUHVysuc3jfog7GnNpfEM/yXs92Pown2EgVXJSBU10y8ZWCjiW0zDZfM
8quTRuXqcyBn7moRnJYjksrN/wfwAGlYnNsF+6gIR8uX9Hy8Hx6DOKvPRVmQnuRu4OcOdUGuxt2f
QbioC81z8mQVdPtUuSceYYGt5OfFDaaZap7GPJGRmDbudH7KIpvr/NyHeK2H1v6yCnPbC70txWDS
O8i4Yn4FWDNMzuDNUY84O+J6HYj2DkDih2wPiOHsZK3T+0RUV+EHqWQDf9553tuJsLsIYxGeAvXj
ep1hLGqSDO+CYwnrkwNRbA6nqoJIwgld8qMywk7XxVZeII/OqzRacfwDzm9NIAGnuE8kj+/CRzIl
46rqvOYgkFIHN7Wf6PS2xPfp45KJ+YJbn3JLRYvM/7zUhGJJupAG7MTUXzcRJ0qQjaWJZTLJKoVm
NK/sbUJFPNZmedOKtnIO/ygXuDl3ITLBFH7QLtftDSP7jn+gxOjif9O1aGV7Ncj7O1y2tYVUr9Tj
SeeildKadoI6wAOdR7Ctu8wVkCo0WZlRu7671Rvm39Z7qbd0Zfxl/shGyhdNFdsW+Ei6qYCp8gKJ
SdlVdOTnJy13Z8loKqtx/wkH4DS/ty4iZn/HAWDZr4jp6/I76lRU2XSaY8ZFwRqe/NTLXLlbVGg9
5QDbHWZhHExqUAmR0OrntA3K1O7AfQeSDJKYWGELtRJT2lP0Oea8kR4U+81xalSM1rdxbwjMPhTg
odWBdaINc0gMGvDTeRefxcqc337Woe8rNMU6MCqz1B+KKDxpCRmz1A8rIMvUjfEpwR6F9UA5424I
QaX5ruKKEmkpWqAcE8v6ytGKmQuFvdGMoTeP/ghs+DoCE/IteVGitbl3MRle2y64HcN0EhXlwn/D
8FdBsVGNj6S12ChLC3UjB3aAoeEOXgmmXD0hCLB0cHVr1O1yoL6RuHlAMhoFs/zEKlOV2HV/5DON
pOogFS1zUiPuXNI9V/3dSeEQ9T7Jw49FQPKZ5/HV2CUBonrdOS2yq8g85ZgPTeBxE9MrTdbyl/AR
v9j9liu2FJSdKkPizx2gQHy4K3mKr5sGPCp8hZTueHew+/HbGhwR95wZigGy10k8UvqGhNqXIkqn
pEl3EO0oMHiCnWE8hA7PeQy3S4zHcthAp7K//rPcnXEplZWIAoc1SW+E5SirIA/kzAHxO17JgkCG
0pLlToPLf+UQ1Cw7yZmqQRB8UDPQ2cksxmD7bUxz4yAh3olu8qfu0czcXy4gj/uW190uLUJXKG5l
VoZ8zpEwnOYeav8Wf1ytZuISRgafYAPaH0nNuc4n0dDJT+hsXQutJxwdGu4wvVDcaSRHOOr98i3X
zKIxyKea0jktdK6QkIMvFh8C3JYSFYyJudmJTGABMe/XYLcLrCOc7fP+W56Ob75Q9lnrAGQTncDu
OaY9658ef2g1yuQF2cXypaxK5syTBcsbDdlo3xG5Eon/30VgX2wsmlUDa6/4PWKbmYyhw36H+Yce
m8TQLyD8m6m6Klr0GoMIHYD80vrjEXhRMJ6Bik+vLOZomgNOC25x9MG1Q2ZjbAyZrPBVP8Ax+CKy
c83/vmMQYFUoakzDAdqyIp35NyoqYjRhbaDjSb40DkVvM760hhMbf29Qx5lckih4IOj0V/JRuHVy
d1X8I5Qa5sknzVcL7reKgXOQN3yf1xvovt60vmYMW7EXu+TirzJ9ntwGGwoBFCw7aIAJgNrMhJ75
B27o9GCc/QRUlEEqSM3DDpooPd5GdJW0cjiJiWPdp6icZBSfdUtS4d/vUslDJqz9GYA9V5gSylhB
hhRCrWNzLGguCwlu5oTcC8W/erXv2Mso3Q73iKDcvnVWMAWz6hW1wawyXQ+HwRERZCNhfYkmmbdD
KgVSQIKB+yODMBbm9aJbC86pr1TSsC49QCjdxi5EXk74KRTw6fpPM0scepTrFSfKcCeozJrDlwfu
QETmQvkhHhf9VF+75J5WV+9PQ4C/D9Ij9LDygu5vYR7ibrNsS7E6uHQ2ZW5Ggkr0z9KDfGizWm2T
RERzhqiOC9ftXlbRUa1qrwcRS9VhxlG0R2ecrMiYJ8K7hV8iwJetHczcPi6Llu09g7SkJydejv1U
1ISYP/QB7xG/ksFWK2EBNyZXgyoM8eBFo1/dU85E3Wh0iqR1ojPUwv7lWjcCoaeAtSmRkJPVY646
V58JtOC+2EmTTXpMLrSfpji9P3pGg18RNNBxTs22HwusEEO6qE2eizZM9HVtsztwgwvTnjmb/7+U
Ow7Cl+Vrw2jXlckdUmnkEbMfPB8nLtglyjHKccNngyMCeaIMLv3+B+VLNTfxUepArWijiZEcA4sH
dIBxQqLxMVbKxrK74xAHxCz872wLwwyV3/n0kltDJU/16TxHDHxaRp4hQMDKjVyMRqjPHN7tQnae
KfWtfcpcQ5MsGGKIqKg+49b+07M8K3GeQSP7O6UN9KpwND6yLKRTJXT8+nxN3GCr0AEO+Y7RHpSg
qasGdi2432lO7dz36g+76UPevMT0iYg6KhwdMQZuZNl4Ws72UZv9Ml7EBOGqU43XqdjOYf1Gr7sg
m+YiM6xgdkMosoJOixD0zBqyfJw/VDxktI9Ypv021iifdQjzg6UH3vpcsYIGck++GKemB9z1mO1x
ufvgJytBxy/cyR1PnGl3qP4noTg+TbynHhEeA8jV0mRy6VNWukqAjSV99/RJzDof5ioO6vQyf4Wg
Zg03zu0JEq7atOXPDzLdFdfPct7tZVSNT0YP0jP2/DQuizao3QRY7ZjAxH9QSNSL73TNRbvDn/lG
C5fhV3J7mxkIU3cyuxkZ91R4tsssgrUDDgh9qJVIT/vtKfN+a/CnWyK5IBsx9ZPQhftc0PwzuoF3
CpqGBj78vbHyU0pR3Pbn1WYtSUYDUXSOLWc53WEMzqlfiBaA6ZY+hr8ralwcW4hv3aciYs9rT1IZ
q4QNTgMXDwbXCd0ZyCBWFKdNjZJIosrsrHIaUqJzme3diC0HzQbrhSqJBagOoUdjInEkVHCtpj4g
+N8KBKmQNZkhcG3vL9K3dVV6ce7WiJkNF1MI1Ej8lueTj9fz5R3D3KhGxLCZRVt68gghE0Iu1wLH
ec5nUAXO9C+4qOhNDXYkzX/dzYsCqYxZIqxNqozKrHPmITjBK+qRAnlB0ZtxjA+DPVCFf9eADWax
uWknzhcKo/mNUxeiYFW2MwU5jag0yQm16PCfUjF/TckS+wpp4r3Pvb0klDeUSqbM2gtix5nJTVgB
DMhobFH0lJ7dUgudOWyztzBnA76affDZELoupEshsnPA1y9rcl4cgxV8qX4xxbN4/Wdu5yGEBAOd
Bl0eZf1i1T8YkrONW4ptGYQQVhYwVkbEfbpvaZKGSHy0SbOzcNNyAgE5Mx5xvhah+vL6vFRVqLrk
pue2W2PnHG3UQJY5S7bfKb9Vd8RRKGafZV4OmLiCfT+m4zBG+Oi0UPplI9HNnrIlvN2WK5OCYmkn
5ZIXaVr/EPUSZarwAoVV4Zd8fYaCMFT6KjehVz59I1UMOhIB9k7rz/avtlOnkuzREadYA9X+PfMn
QVZiw1tI2Y4YSD6n8ncrEgYM0ec6eCb6FZ4IWzX5bh/c1Bu19foJf5DqCYpMYqtvYg36Te508xrX
Cr8FeXW1oMK7SDNi0X/uziU9JfUofugzrFYTpAXWCxucvIRlAeA4ozZJ5FhBDsIt4mfhZQE5cvmJ
fSVFNsnSeGu7QFdZQCJaLqa+/DIABk/qrL39W1F/BhIWNGAKLpaYJg0C3NR+o44x9+AljI8Lg/EN
HdPxDd3gKO0eNI7T5ii7vWlnX9Q50jBUkZGThu1HpHNw3ksKFzHLFjHLEs7oiB5CGuhNWf6Iu+ve
IP2y3cdo68+iGZQHvebaBDFfoy/6txhWlvdr6KG5N78AV2zbgYIjpWrAb1XF0PHzgZIRI7Eh+Sgm
2TVZXHpCO9Do/t+IzIDs67kZ7Dck2CoGntavMblpR1tNvx3ey5agctHpkgEFdp2jKiOkaBHFVUbd
NMLhWQlhHyekLia4+69nWZs7XM4AaJh03sBNzWH62TZNApKSkPdUxe1g+NqQA+Cs0IXJBjJ0x/Ld
8JHPOxGGWtOGXsSBECRXSQTLfYY+sx/pVmLdZV6ULtU2uwAqrjnxwsYhIWV+EjgZJxIO+Ds6hgil
E0Nh9s7NvSpUL92o2RhIQkW9+3kejZ81+iKTIFNa5Anb4EQm7dcIN7JKNwcBhhY8big061ZlycKj
3CbBlE7C4gWCFEK1bC/rWB11rbvqMcfNoJ94iQ1zLUlBSMKZBC/xNTK8Yc6IZ+ypCUqfeZv98qpW
RVO63LhwCbwtcLKQTvLnhHiVF1yl7LvX7g8wAG07a3rMAoewPeM/Ji3obuJ/Q7ySPlvN5pIsgTPK
0fBzxi76o4UIvtUQaCmTi1evybl2wJfKjSyfsUJ6N5q0O6dSBPxkFrY5jsjnZ4EZJMfrb6kgfe3p
9lHUoGIasG+GQF0sxZ8m6xnGQcjXUcWuN+czGkro3/Q1Uqju5PJ2qraIMlbSMzuISe6o6hBmTvtz
jHS9BTk4vMPpykvcjmQQqqVXBPFylC7SWq4lM2TlwzAHwRzjWhJEn9S4+Yb2EdzIbch+Z0/BqzZB
eosjov9dese+RuwSNnj7J0t8Bj9QdRiFZbo/o9/ADAFW5mn4Kx/ljQ2ofoZaVfgjdQNSubiaV4DU
EHT3SrWgSt3GaLExWCkjZa6Dx4BGn0EbM2rJFAHEGwqZ8ti7HOeNEXAnSBzvP5QfWhaMu8gtMFsx
EdTGryM+odeJbZqqyf0JlzcDqJIF7T2YIUyZ6h6WhVeU3SWRCvXT/6KVHHxoXUDslQmiv79jJNJH
OLCzJ70tgwQ3u9/vlFPGkC3N2eLGOBlERWCpC8gxbSpOD7f50YLrPTr7YGO+WJVB23oZHCXwadjY
LzoKk4mMjspk8uw4cK1ZbQktMeQM0AFm5Lz5YHioeM3ZrxK4gmEAO5T1D8OynWjHWVRFdbP14S8G
ycP/A06TTYBq/tLaBa4pAOknlfSYJhf0WlwygngX/2rrpKdY3OlN9CuXHxL6/Pi6/HQwswJu6PyE
q4fgcPjyD50ly3mM7aW+k30GnE5TExMRiDkNTpFVta10zXS0v0pLGeKNYLT8mwxDydZTcqr4o8kh
At1aX0CJeaiADVBDa2n6ECJbRt/6dwGB01AknwiVOHwEtN2Xq2h0f30qhCvFWuJIXPTQJUnYHt0i
OGD4Dc4qNVTMnyBxitfD1Kr1L+Zy1dyZwDy8GaZcBCsuSTs4ws5/l2bWofsra7zvPeIyExIoNwVd
NKq1zw9PY9n/MTWQpDHEfGLmf9gdSwBNQG1OcZjLMT6nhQQgowTI+ak620JmVScDEKJ5+A2tw2xb
IOBwny/+jvhRzqC9JNwdTgxgewATBGYi6IBGf7EwY8Tk4+g+Nrd9F+RJKezVzXzaTpYXoUVS0u0+
KNzExUtbH2lTHfBi67d+izb6xW9Orguj8aeN2kthQkUdt/t2wT/aoi4hH9yrSxWaLq+BevcxWtVT
YbmI5H9HLlh8YyuMSg3J7HkuUad8SgWczvN1rEzed3TQ4gdIGVlKROO+Dp2NK7jxDFbJasuaMr0s
NwtNedhDVlWMt7zYCaAUheLY4CeMwSdHdxrX31nlYnvFvUhP2brOTQti5am57P1QJFN4PrOm2C9q
mYGS5ivx1gFwmuFoJUxwF/W4h7lYIJccQPxRgbguF4QzZgYGbX2InB+9d1CKw3pHzeMRg/xzhoDL
l9NONlk1YYsq2YfXd+08QCGIEdDNzE6454aSmGHLkwzHXBc9pKDK36+4lFn/YjroTLXIiJLR7i8j
fUONdiIgoPOc0jVnU6A1iwF3yy09IRIuoPMRyV+eDHzJuuil+PF/NL8Xsvr6viBg9dIJXC2f3I4z
QbSnjcBcyCeb24TE/AC0QKxxXdOjFT9qb1xvDWRVmyjzwJOProhNrFxffJcq7XopKAMjKg9cGZIR
hdSkO928wWcHBMcZ/omdyJXdfMULnEx7PBqAaeuc9rVAy8CLwUQLs/672wNeSMm6PFwweFXFf5Wx
tVRw7Ksjd44mIzzqLWXEEIkiDnTrW5G1iPd7qGPZPKnXSY2ImOJnF53p0z4xQ1IEdzyweZJoq/hW
Jwfyz5Wq2700FwDpcsEUT82nllQv6Htk3F80yMceFAunpBPnvSNRI9FbyrDWHxTZX0ZzI/9fEV4r
3IzuQz0Us0nPb/uWoZ/TlBXobEl/oI206srBLPUcjzSadPUsvzW9EZufHe2PNiGxeZ06TW3SMUfg
j/XERnTm9T9YUGh1OPQRHd9uCiwHFoSgO+E1NxqMK5w7jb9g0rnKKQoPjupnUgiFFVwROwZPGVV3
kum6ms4LR4R1lIAyo3hy8blKq3NZZP13eXwTxmHiHZOVCLBjsqPyEVvjIkCJtLcBxwcnVIpWi1uY
yh7Qx6HpFrGu5eXDbd5WoYicPpaxgfZm5QkYTP3mp6SRnM3eOJ7jhkDpvi8fiTNWsu22MP/QVqJO
VbufKJlCT7uYs/uhIYZFqz6PsmYdfItjXqCWV2oWUGjJBhQ9abdgpIu6QMazm8TRvWuZcVM5fsXn
g+LLdf4S+X6Dxg8LWM0keHFHTZr7HJoi0uhuVMH3iZOZyGAUCgij66fq3s6kNYoxm+KQmsmHsyqg
aESUIW1yaXKb/kwaiKMrQWStrXtDhGqK7UZMKSqbzP0gJzo07etXl7/TDAuUasjJPbi04uuc4OjX
ivlvGshM69LOkVVohLlLuHJ38avTqOWT+hBXvceoCxDo83IGItz0pLbdOzkHqSJbD+h59ropVVVI
IjvnYGY1+f7QciB+8kQCzGl9uHE/lmNnxqNFjyHHE7wh9MyLCTSI/t9nyk2AZlYM8oR0XEC7mY03
vhXpP4trFQKGADjl8NR6xIFw5URpL/t0cbE5ufkj+UGAftw3gwXe+BtIpqI+Os4qZN8BtNEmVnrz
q/jTeZqpwhkYaXstOAXUOrMmWUdJrRMR4DmFmXnFkaDwDOEfHFBv+NmwfvcySWAEupB58bsnbhWw
KorgxKV23TZNP+YtDsAZrMWz6gIquX7QBnV/F36xsUbJXwStSeRSWgig1PFRJMJx3aD/MSOdFULL
sjROh9diz9sAnKytGZqQrjzpg6ApXa8D5oDxGz07hbEZs+EHO5WOC+oNyUPRLqG9MQEHfti5mVlO
ItZTU/04aGRWnxSODhCBZT09sGdE0uzJnWHDcG5846lRB5kAt83lUz+1YPKcWAXyXY7GYkYkfhSG
cA/bS7IdFvP3CShPQJT3+cYF3jIZpCCUIsckH6SG3zpQ/FvB5nOwvAhKhNvoGxeYSSd8pQNpZyEh
RzQSG1dYbBbaDkXFfIX7UvzKh6QgpNbdTfJ7cAf6dAvHVFrBgz9ojnLKV70hVE5SYNS4l71QGAd7
4jBBsqbMAhKeHEaq+E8xkMKesYAJrqnnx5NQwpy4Dy9EmmRiM7+Jf0rVypZpunhII6K2v0PLx1oY
fi5MQ4yYtYSEpChj0UzjyNShSCgCm3ftsn+E3dox+s0zKqeGQ3GY56AW7oGPKNEaxOsQ7Uk6YitD
1/zMhZC9q6cmsXCrgZZDqpvXD1P6+DZLYHHHl9VxaiXSek4sJwoFzmnKcueEr3qXi2pezmJZMLpa
XDG/nOFIoNwAnWlgbtQqJxvg4WgtrsW4B5bZ2V7uvn0CDvyrm66M9gexy++4x5CorHASAMMzrBqn
WVN5b6QMC4BnPNhK+EyLlhToaFx0gZFyfRB4nGgQv8fjJijku6RrOd/ksWmm0uonpOHTD3EnI/Xh
U2bYnHMX2isQDrs2M5Q8WyOi3KvzuFD5V+fck8PlcIEqxWot9/i4tNV4Jx56Srw7iK5jkD0ugJ9+
nmcNyPI9GY1WYmH4vWl8kyJ77N2j8MenLyfEC/xKDeCilH2OB1Y2XDlTmxPyiIEzRDi7BGrnRcYI
/iZQ9G0S9SVEpTHXKms7oNVaAFjvHXa/uRj8h9aQ//+Z/VGYSoJDOAo2lwz+jjxcE2YQcwJ47LYM
peugSLJTE0+rO4a3GSkcOUL+KNy8nCpxCwH/9slEOltwQQLzPe/iZcmR2/GWK3hwLAQsiwulQwVw
yANXqmXnHpZQv+1SoBEZPLIlgn914bhDhIAAHerD7XjcK3thd/cCIqOyweiWN47cneYO8Lpy001Z
BC09PHzUAwmR4Yh6IyaHBHTEPNGJoZsZbmXh+ba7i1HY8ZEOX1WSr4iT8ZeIdSsD6c0MmIaQTmXp
/YuN/j0CRa+r0dHvNX/4B9+cRN7FvZo3miFZ791j7Lfy0PZ3pfXAYp/ktoJ80nOU8Hmpr42epy2Q
f4MgElIfH1JriLhW/uiWDYv0UtE3yZhUGfiVocDhcwe1AA655DrEBd2qhOC7ReCPDRUE4VDKNS+N
AiRh7Cy1zoZkmqQOxPNGCLTWg/FlHM/OYtMKLJgLzHEHeJjTgN7tZCUWObRlLOlQn5qyc9jKC2GC
jEnpPBYGKCI8Oo6K3tvTKyslThCYbbyUQb2d0VeyQ/mcuVorRK6b7RSW2tjZpxGkyZkW5heB7mTV
d6RbWrVNWmzs/Q+zUOcSBVw6ZKnz3qD0jlBKTB3DPltQIfchIlmnVAw/CBIhAAwuV4/n1Wd82gy7
4R29jIte2tLeJEA6Oq52u56NkC/0A9wmpbq4gs0y3Oy3++kkUxjNuxvM5gC3yFZ88Zx3JOPwmUOp
iWCRCaVmApAlcZLVbtPli7icrqrmbXUsGIAZ6trET7KKQr4FosKXWl+lpmJZOyPCtEUsWRAd6Hkd
mw5eUygfGy5rnFEiUcjM3NTatipv9USplV8OsIOpOu6ALAmVYfHntkYitPw1uTXFfZKwTTMbtikh
oC237NzObjE0/r5+yt/oeSSlvEO5wOyUq31WSgKZ0z1aofB+q+mq9IaS3fQv1xRHvqiysJEIUMFb
p//CZSdPRAal20d7+TQLuuMB5KkiFXg/fJryKvmCI/8o+oFhCgOW157N1MNOiA8ujqZHhCLz88bZ
3KtFtPYi9SalyFALsGGYOlmbBDTYEOBl0qm4KL4iCBBQTn/8f2giBt6i61e6FwSz0ktb1jBk1pdN
9itloUBBXQBXRruUXllfRbAD7cvlqqmQ9o2UVQTqFhHmyTXemaIcE1HPe658wjyMjX45Sg6T9Vzk
jj1nWoOmhaMhlFO+yreGyfH+66/bdej9VOwZGgnyXOeUrsq9+xMB7Y1nblp+K2EIGd7fDh7eveH8
u8CMGAj3OYEeaVF3Md/51bmfogJPaaTqqNTRslAX3Ol7wzwiB/dl0i8Z0okKtowchHOqHXZtmFzh
yecQMn2JzLiEEAGS3mVyiXqkvBniAcl0It620tuGinjskr23simDbQ63vrnQXn6ga5BHw6VyNNQ0
3cd75PKaUOgOU1R2n2+FSeiSQTGFkFm4fdkXBprYCmzv40IzfxorKAeEh2xF7m5iG7J3dhuY9Aa8
iMkKLvgHtGk2+QyfXlF0JZ3+Xnx+e/sbKhZPGn19fcheypHQxvaTCpNY9RV9AXKQilP851r0uXWE
bzQMBqoD2qlY3zfgrbqHVAhLt1/EUlxxZKwYZETlKSlss0wd/dFCcJ/QFt09CQljeYB/TTj9fJ6Q
IYz16XqIcBsF6zapDnOCqDcz/1LUKVAIgf7w2jeklAaO2pHXqDoXEvAxOGkNRR11qgiz4u5snSG+
3GfjVOEVzQPvHmC2ZmUfoZ9DLnF2vFOT5sqzMp9UfumDcguc/RXAn1o5nnsj3DEMkcmq7OoiQ3EX
JEMiubNeWsxSYoh6tPDgFdG5+RpXZtKvgpQTT23DDjLqlLx2timn6yKFcIbudFNDafDZWexpHI3L
qdJ6cqe00jwOwzT0GYqy5IaHkyw9fHpQM/m3iuwkbofRi0IwFgbcDQT65/H2953+kMbFyiYpCAyS
ToyhLv2tph1ZRVCHLrq9H9z+S8Q5ialGzZJieObaJh/bcAlGmOTCjqTIkahf6tFDWm6toVdaPxAK
LJ4IaXU1PGLatiCvSas43vzDxUA93pWv6yDCeXIXrE6aa7i9wo7IxryVNDdKG55sKRxsU4TgjKHn
5zKIM4e6PR586Opv0tEU8m7NRWVBZjtVf64E30Z0/jxTU2EiBily18yl14q/Pw7OrgBky8wtPFMj
vkN+vArB+wPGeYVWFX281Z7Q3X/ywR56kr6OhnOKVUiwnE2HrGCiXGs3oqvFEaF51n1q4dch5O7T
eOinpQG+vZnvnz61hWStZ6VW2KjnJ48BvtJz+c4cvpI1JqtD5q+9FdHi2s36og/dFJDqjzTO7IRc
t7o8xja++VSA9a5Q/GKOEcZ1+xiFE3CUcgQoAwjYxkBB72SiVOjW77lUe11fYNbt0h7uXPcsGCao
KZ8mqHEeOc2sb7JUzjEl240v0y/tKKJ5Nj72YDi04bjc6+j0cYkI//9gt31L2DeTw7o8VULJIvtC
LGeaPvgnrtBWRzKTxxE9u4zKmlWFcL2zfvK+RP2fkMGyz1V8d73uAcGVsGVvYbfYQ3Uu6Xum3WYL
52DNc7m+3N1Ss2i6U2UzQH2Z0keObWWsEikKEM7oVHBMuyp1pWlLszVb4BztgVwCwi+PC1cuNKg9
EvEDyIh0+Afta+07AcGQo3rdcxwb34QxOrRMpwmOXdG7AgBBLvz7sYbmBEbbVZlDQ9RZZjY+2PZ4
6giOcGVSiYci5+v1fwhS18mG8eOLUtEW57UsS1c79RyvJQKn0j8qZS/HgjlGHEVLlz9obKGouUKN
pKOSaeHXrO/Y7cmuvN7i7UZ0okFxQt6e6S0PP8DtgWxnFrxWy43H7Xs3tXRGgs/AOKOueoAaqRtf
irXDmGY2j2e8GLGB12xTJGin20+pzK3Y2z8YO839+2R9VQGuKhcG1EyOoKt+Wts0RCkFXPya2RGJ
++Ge+/NQGgziry3/SZtJ5ORkWceA5Kxhte9bC/7KitKjWuHlizPO3wmGWhFGmK8eErN64gf6YLtp
1j/XLbwYOZ8b0WyOInl2dkGJ6kJu/Q3TgoRGLIp9JqZ6YqIdbyTLftnxVO7jTEYo7jmgrmgGScPn
F+ruhpBU1sayAH1H1jiN+bJt9ZSrWcS7+URlLIMuvQBuoGwqNVlVpdzVCb9VIXQe7cXr5SY7UZSE
QW0lBBuNUJVHbB31v0Zh3xGymhphHVQOOmNxTBUjpAmNcxOMTSIOuZsI0eSQiOJQ7KQCe/EOo6CH
L0gLhar2dOztdowhI3Oo4qGI1Lq3fNeCXrlUJIyUl+xoy7K7fyrbKa9NDhK06zA45DYeVWElgpxN
DLcakO6J6bB/PBzf49CK9QzeYoQPzT+WUatwgm5HbKTCIYoqgQZWZmTN+SX9eU4KsmiQC1rluZmE
aF9+tGHz0HvCdaLYOKaSEtmTirPCVcpV+Ly+vZNvPEcdlp9c5Mfrg1YIIlZqWR183o8N6a6JoYWE
+joqZvvpqz9TniGRlLehQuwxKGe5lY6qFl0D/lcV2I43/LTlMLHCw0kydOrsVp+0OBWmyr2wXp5V
+EZub7EhE0KWrZNrE+IYcn0Mt+FbqBcwu+TUd6yW2hSuHfjyWoVEzTaqz8DTvdJu4wp+rBKRBn9V
gaZGSOJd8INxn20d4c2JcgdB2+JFTVwljYPZWs1bNhsUY4nytSs8sDkCIiEC6hG9uWZ2A05q++Bj
xeyz4Boeb7C1mULKnufYMQH750DSKhIanBocpKoA5mYXGfepiMhxdMVApInkgje5i8R+84yJ8hAT
QQIclRGoIzTdoO6pFAGytPVVLWkNtOSoZ4acZ8Wewue/yck7wi0NZdn9q5aiTo+u613z+MI9raQB
bNmIkCtOgMXe/WuHScR+eVZVhHwOX3veapgXmHwRmHyR0TeXdM6vJ0CyH1cxJuIaWr35xPgAG1We
AL8q/c/FYnYbUEYjdAyFPFO7yYAefZFt7EJzmY2MK2c3ZJru/s5FoKshtdgehFXKsAOounC4ySXZ
njB0UORvuWuayYLTuIWHCd0kUbohxyDKb4RjnuW5kWLIH++xgUI36baYKjsTjvfAh2lcfs1V82ty
K2BgSDGX0wbce0ldpRVOfcYmuGTKZylr60WHZQ8vdLapbgbU+x+tGNrol0jv7VkP6YR4SUZ8um5P
3B5kfXAlGqXw1Rl12dwnRYVhMRfyzp5h+7Fd2hQeGHxnru6H2cKlsTeAftHMJQNPFAMxDYQvZGbx
sYqOSQ4+BD8U8CVjrgHXnD5EPf7u7mQC8NSeiPhhlaAOfYjBgYEExa9irFktUsaCeUr1i8Bc0Bv5
vhmauLbzx0ndMOXwzizdlwlNv++TkYuKktJ/AETLP6bsiV11rtrivYZVMqVudOfm3Vrim8ITF4kT
cAjnCL7s/D9hZo4bwgqLHqL1b5vBnQPLLCHFyT5Vl6dWkT6UpCisd2CC5UMROX7ETyibBCPPKtm4
isiZxU3zDhKAR9XEViiDsxnXR9sUyiOJ/YTiCkJBHofmrAUVBIVE79qGgtLooGyfESoaxBzBOngK
gJawaLC6oQ4u1wEOm8plkj60A9Lj9/5oPHMsImuLuVXD+Ejrue1eEVVUL2hwLDYajWg8PChQMde0
8dqDJDqlhWA6dI8SOSKxfBuOWipPX51TLK+eySknl/I3VN3FmFf2BUGQIXSouSkDE8qEt4Yefwyr
HLZ0pNJgmVDgvd7d04xPM/HKPMY+jRwPRr1c3hl2RpRK6nIWJM/kNQMIzzsvrPKeXdgvTU4DZxFw
75jJSxTcWb9/jSUqRcjg1FNatCjSPT0Ag66SIQqhLrV9TxgLgaqr/HeQkgV4B8gkBBnvh6x8WLcM
6am7VryojOkdUVsdKIM59Er3CzUvwXbeIOXGU9+lGDqmWtKOUM99CaFJ9K2SVembjmAJnXcmACJR
ePLSYMN4rU5Ubn3KVTns08o4IxxMxCNRhHnvZs9lpIPD6IY38s0rS9xfvz+gCnMRSknLfkay7gAC
92Cad013GWKOmO/MtpnF3kJc7hA6NUeL9i7ajms/POY1H0n/KsDfMvP+ahkbWnu8S8k8m6oG01Qz
MzMI6Omu/SVX8sp7kVrEuWiEGiZPoIThd2vyHy9+3szZe9C3R+zGXoQy4o36FOuCph1fylhhuGVn
pAo/FcZBVeKoL7NrbgAmnsBfqjYjIWjINmWEbBB9JvaArbXVzTaYDhPmFMpKR2nYPQOGO+zXUgHG
62aDFAvi+OKs6oFRyP+hPCOqhX0+2Q1BZ1hYLAObiILe4g9YE/2ZZ8KIHGhD4uYuTpJ/KOp9obK3
0DrKJysRTU9wSMF/kKAt1CMqnD6JnelZFYjr5GDj9pPNHLAGbR9dy5oZedDxcf5KkURydzItXE/G
+vXtMKMaXfeLGsLjIi/YmnSSH1jcDcIAT+USTLFL7ihFLgZhSrvsX3SNWOrOhA2BL0wTgkopxoV/
cOmG/Hxg7bYpozHaGYA0EdQDlhOzDdvKI68Y7fHtRry2Lvc8OLNWuXO+O/YMhtnEoazPDoCIWsbS
W7K+0GVn9UjHupqF9bLQ9cP10Lo39XYU3hVdLMdmnj44ZcYTMKQXPbNoCvzAWarA+CIjZ8wAgg6d
N8+wI+BD+WOfnm+lzOkZ7IwKX34KkOuqw7xu0zmv+q5LnIHDAwNXcM5E3fihNysCBvx/Z5BcBL7B
URkBn24/8j3KRQYGnlvqMMZ5SYhycoQwo0+B8S3YGMMXwPm22CPLAHJ5Fku8gVJUUS2toy+fdj6w
/HUWwwlY3sEBIVkXXSNXbOyK9hmaN7KPbQe6z9vhRx/9s0XIR2jBPFe77RL3mtDbd5xgBLzIFbgX
UWPO/jntqRnpYSU9+IaLlX7vi0oLF+qzhHn8wzn09c/hpO+NUbCYSF+kDLNcbH9t7JFb/87IqdKG
iqw6ROg3/lLtaf3Niux+SN+NdXmVBLfmM/s35fnJlkUXf5EqqvYA2XMjJC9Sj7kaWlH2fn05Q26x
zdNN0kaKKKtvRJdRth+6obEQNB+bzx7VweuYJ/FNBizk2oakUv10rQ71TACKBdWchhVAiBeJ1tKF
T8B/sHbE+bx/9I9x+3DUaEk5Dfg0laHoJewLA4UEwZA332Ca/l+kLIw9N1gdU8arrpyy9Z7I0KqD
31E02DYP91C+iH0x+zZ/6uau/Iq7mLs/ku8xZHc24dSz2Z/BwzjuAzRtqqiPNWqoVI/Edg3g32bU
H1qzRUp+4tyZs7EETwW6hoVesfvUC8RWmRr/k8ukbr+p4xLJJ2euS1oujvOYUDtPE3HxBsGzkIuS
//S5GKfXvj6OYQFsJz0Q1YgtN+7ggB2ASFm1cRW53NnzXAkjBQPIKujzBldpaQVpLrOgHylqDwzc
CUIm5J0Ca6IxIjvxQMCe+ipI7inZdMBEcsO40Hl3eV1d0WKOCIQoKv/wFsuKGAQBawOn93qI2bc8
0jqg4tZZBt+hO0s/8kKgkQaefKQe7RaoDp6RVrwQyueOg930U7ylNvwMm8XskIKhT+8vVxQ2DLAR
h/+Q6mHc204B509hatRghcwyW+A673B77PWS3vZ3glKh//njtuiHW2yRHBrKoPMGlrsKvjp7XQSx
4tf/HoiMUZGMFkSIjWSUJIpZ5mAxPGOkPL1KjaTgD5oFi0oWtq6HNWsYi8QxwpEL4BdBAkFW58O8
Si8PatRclKUPbXSMdVHcvjjsKI8KqTS7O+/1fpOgkGdEjYB67BeUi/PIYxFgpA26wxziOvfppbC3
Csn1rBbeTyEFvHs80sf4T2EQ+aJfl9h6CdtQ3qoJs15UuMij/Y5fC7PvW70ATzt8/VlQ8M9tzKs8
xrPhVgl8akwDov4XIbl2Nq76fGvS54P5dnAab7xxRHuojqLLhGhVQn+8wNxXa3tV6P8jILOYBPw6
RH8njv/vQUg1fwIdglBACZQGWewabK+mTjlmB+dxHQh7mgnIzQPvBMQ7LSIGcqHRiYpOxO7VbvMl
Dt6SZYUdNXjVRO5+Ol2tmHDw2MNeU/OKZa9lJAJPSmkEUM29jhf6DJqK3x1kylcbbdk2Ozo07agC
t59p0aD1qOgh0lPb9tD0AHfJUdY43lQdbZQqmu4JI9ZzU9y01ewiRhbzRMrhIGQJfgMA2aYoShQe
QPUt1nijiYbzDNFK98La0gra+SJlzPupxpgVPAc9AqZMJgpqokNBkiW359ZxFDpnCU9E1wz0RPLj
Q93q38QgQGNsXClyhqTpXQR7PxiwsJFidcSM1hewFqIiQTYsz7Dxz1LawIxfeAQNSCbi3qii4ic+
yQrvc5Kslu7r9GFN894X+kDDfYiHnceVCk3B6AlHViTgZSPSElPR2mFa+tleTVk91NEHUWUj/lAE
H9UceJUFLr3rUxGO/LeyzObo6vs8R4vjWsPrTzDK4b5sSOld5T8GK9PHwxjWWXAGQcJH9rMRVlfr
5YZ41c2gf4dzsqrS47esrHsat951Kdg/bCe1uSSuOQXVwUN8qe8s5KaXnzQcsiP4hPiTvYZ9hU/4
mpV16262t5O5n7x80oAy42JfvvM0NHZ0mr+woOsmZLaDQaiC8AHFsaMViG6D8lBiVKJMhuZkA4Kr
8EDydLO9zGWMZvnQ0tFDb7Af5Ghci+Wo8VJCylLBQpwK6NcjUfLEGbRVwL9aU2apS33qeiVuCGn2
TES3rZngSAmnkqwR6NpYGkcPlyxfYSIgQOssgdWpt+2VfAeJn7523gpDOFK9U/lwDFVdQ+aqFYUN
ZWt5YPXuG1kxpQvRac2ZpAs/2GDqsSCSnzAuJ9g4TiZM9rQV0sojFzkhw3ki5hcAKMtC3ZvNLxi9
Um5Vhci7KgkGgYhS32OFN12rPEaYLz1kBg/5791J7GCAkwu0IySr8KPTpmiyxfMAQqiZBsfz9WMg
WZ0XQSjPkXGJaZbaH8OB8Q1qTlnK9Mit1Q5mGog1su8Js6DgXgaRw1IGnSWgJBTIxQ2FgtYpMwWC
m0a4bV4MOG6OxGj/mrGi9MWc9hnyBHA3l/s80SBWuR8t8/40EglxKeD4hOIkRspuOs1CE3Q/HK9f
ydxuBXOmX5a0wKagvI/Yikbm3WZDyup5JKFJwmAnwWG7QgYhnuwDvLQxmQOnoZkZnrx0pIkSOuvy
VVuSylTUvLN90Vn+nekf1qSMmF70lAc0EURCB0BsxDAdnpiiagPzb8OQGG8DFrc1eEVl2syoz114
PqaItCQDVc3CTXHPRX1e6gYM0UG75yP0hD5NR9MSKmg/gHBh41GiWNbNCg0W1N+EmMwZoDTrPdy9
5vD8Kc3Tbi+q11G5gPhkmSo00T+kRUb2kkbe+FZ0KLxdjjT71ImKzM7GokYtwoYfyP0ZY2O1O/N/
RQhdkYBpD57lTatNUucV/tu+F3Z1qSoJO557WnX/OySa5TSKxaykkRlgXXholAgzSsMdiMbntabD
CqZfMIQHmnU2WObFZSLXgAapuvW7QQ2O2phjsQE6VcUd35aBScaSf47lgYXIs7S41bK2+YE3s10x
TqWID7EqbYkukoXHIGE7G4ivGodxIoXwdsNHRawqXejzL5pkH7wNtXQiOTh30TUZBPFtCRBjn6YJ
Ky6/2rQlg9uqSnypYLwG0ZBCOW8ROV5aSHaXGMGbIvYZTgwe0/zZlOMYSKfS23bnHFkSVC/7Cgny
AIK0S90+9z2uRsmxXAYG2+guauWIpf5p/MGIw1ZLDhIdF4Iw9rNxNxH2pLPVT7T8wYZ3GreIAaO7
fHPSCeJ42Nnwjt1hZOPeeGaC2Z7bWmXFklAz/p9B1B2xTdzzs4E1V14Un6SIMXB1AuqseOR+IXy0
n93+XM3e2uM5eWayx1ILKl2GIWZucxsGy971qYjBKSHi4xT26PrIK7H1t+ZqMyqOfCX8soCcUvBn
jyRuLNQd10y3vkCDN/gtD0quOBMD4+PlSWfg8dzo6BKUx5L1Ap8uxih/1mIsOwpPKeoMd20BY2UY
swSUgAaaIky5qYizZ92Hsc8JIuCNuSkf2++/3ECXa/qNFvXGAIRDEM0SYPrJPacuy8x94t7t+Fqd
ynVWQi+6YVvN81TFDQHeZH2SAXRXDEnTg98YXy0DTKMlZCm4UpzwUySts4xYZE2dMO4g8PZ1LZli
hX75s893ugYUpfmgq3KKLagAlEYNcm2JwOX3iCsk6pBUoAnx5dYomZJVRQirKI53onaQfavQAbWw
b5U0RLNqbR3Fc7vp+HrS66sDtbfMOeo9zdeaoeWOGrjMyT21qKklwzJzwKFK50dZSN00q6V8cfZM
RHVa4Ae0sNP33whw8JX47OtpSVDjF2Hx/G3AGUjrNt8owaI1UbcqpLxDt2rKV5l5xm1e9p5hfTki
YCjnC+Zae194/u/ui8+mH94TXGtITQIb85NbyNTtiDwCJjz5R+6U7tFbupsmWQ4TVrY0N+eI44oM
ubLK99J/BZhYbkrqhpsJPPIUvt44gwXqLbrYkSKyR+xGPKjZq6HadmEqeQ1lkrJhNOtsmjQ7dkJ+
sU2IYLYgevWHzegGzVo2dcEPkfeLI3IQ4wVjAqESijkwaOLtE0IoaVHuliXWk649xP/vP99Xr4+v
ASgrZX7CLeEPh2pDTW5UD4GwaR5j1Cu6wIZcf+4xNOKTQ3GxA2Xv5OkL1+QeWgbOkHZnGer4pIkl
npj9u74sRU4+7Xpo+wW3NlLiBH2twfWu30hH7u8zKC7bc4YpsK3KQNzQ3IopRp+pbEC86osbzp7n
0Fis3xG53J9ZF+rKi58KddzdjfWOzYUEIyEn3bW7kpe2Dslj4e4exqu240FrbOROL9GrIOJJug3n
JdcFwidYeNQpMKVUb8mp1Fpy9zKnN6YCpB3GyaldGtrcmGTmric43ebtdI93VLxvDf4vdMM1JPYQ
x0svaOKOP2IhNxtnB4HcNC5tpb10nN6WRqCCrjVgKuP7+xtCqj51O4FUcuJVA2GYmVrhE00Ok09L
U6i8ldjFe3OFL6hu+NLkZQGDFKzeDn2+gRCQsNK8xxnZ0pc95h4j37eox3n7xneIyRxpo3O/tqHr
C9UO2yHFvV5AlKXPS4JI6sqQkHpEWrS5kCzYkZpLQSnixWRvs7nN0V14FDhhpTHr2FW9bUdgaNnu
ndnCMrggymJ5kNwlxG0hyZ9gb1cg717nP+GkYYzGuHaUuNK0JaLH3wlXbgBzFwEp4h+m+MalnPqO
/MmHQs+e8XzRem52JakFHZogFX7RKxqkZo2+zF4FO4W/XhHuqjAxFAxn6ZdO4aZUgO9fpSvCmbII
PsWWA5thdlzfO0zulT0UBaa479IFMuSUMtbbk9zRZ4ZkMfyOZ2FcoNzpA701cq27PEG53i3x2gPu
XiEeuJr9bscdr87r70GjdvglFfLcYuTw4W7OXPVWBRqXt6rUXenB8dMa1bLcKqZ3DH/nQAJyVOVc
kfcHWW6Ao/wbs4WWYlYj+X8deBwiTAxDdvS+mldruxWcNgZ0iuzYtXBiCPyiKwnmNg1Jz2a1K1Wq
VIHnHha2DrRPxTe9KiVTRPmfVBX7BqlSRFg6U9CSfSVB6vbTQXpjZ708dfDgJidvLxi7FLLVAxze
tYZbWQUrf/PuUzWDHUDDGGTtRuqTCQAsgLr3VxETt1n27JYbViE2cWHGzcGQijfuXcro4b0eaYvU
KYQiviSHhzNQh1LHayVKX2QMFg4LTM8245hMWFlELqdI243dpAn696vWmck05gm3P+hCTuoYge2K
0PGHhqBLbtlEZPGvkR1SoRoe+elFdHBSyPXglzSYuLWAszwE0y9oN+U6Qtj1T0iYKCkosxm0hhEI
8JL2Asws0J6/0aqAnreC0dBAOSB8pqH1WGuKWS0MRMoqWPFYvKySyBbgEx0bK9p5+srrVdJKnrsT
C1lVg9L07yQ1IOE2T/umYbpFOAbXzVtVCEljJK31623tqahpBgebN0AfyYvd+Yk+ykKSg1WojpTf
nVMXihv9lT0C4IdCfEl7nYZOp0V+Cl/Lk5m+vTezncv/+60NVs6gCi7xnuKds15rjii4G/r1VfxU
J+FovY3B/t9b+1DXqD91mukTSC33Zmrgdh5Y9GYRBs4+T8Cirq3O8LXRP2Sjlzk1kcbNXFo0i0NO
0k1tcgqMRJPopufx/V3MOBasXHJP4BBlDjW+2YJcBYwpq8DV1BmEhLU5pgAzj7/2Dy+xaO9dSnoU
Zd1lLNgoWH85muFPRxQomvYb5/M5IT4GEHU3k5QeEFKnBYxEV+XtWMv/DMDQn4k+wIdmCFE2WBEV
k0hd5wkNcbJWas1i4y+8P2KmJNx28f4tObGjhSSLHxiFETb9Zoa4tCatSwuEpsRLivGNpxmTDrWD
Gr2cTmPE2FiK2Q24v/G8LWoZnIUcgGdtStF62ge81UqoPLcbPUjqbDFBxQnxph1CYgHpSQF/jcjb
kHKrCHxzRIJE2YJ86lwxJssvpDJowUgynlrTs8fomPnpgQjjfZTOTjclzKj4XV+g5Kcis2oAvkyR
1Txj9H3VCM6cuaOc9v4q2tKHth72M2fk98oaJSmZni5lI+njqfLbaUonD2N0JPfMprL63iSN26MI
sxxjRtZRMNYKWb3gJ2cf+WHOVc3xfchNhCpsBuq3aVbLXDMmvAk0aveIA3kH+HPv9Aqrbr5UpO7V
y9TfpzZtVrPR9TJfmmHGaXNEJqJO6/h4iqfT4dOuoLlLA+SV+GY3TDwlD2NwycKPoYjAMlvyP6Up
zc+gMvi/DeOnGRL3UbogF/zB89tItArCPmWs/R3sWVLif/gRTuel96YGsQNLgZZPIp+BpgVodZDN
phFxJ1VxVUw4A5O+bjTm6XtcTlQoPto3XnOGV2gAFZMkUCrMJp0pmPg3ZJdlgVM2VNPiyKz7E9zS
vsoTuzMTa1qxk5kHROpSKyZVK5x42XIZ5OZOb0fEECkIu4e5kkGd770Jq7d7j7+9NKhNBHFnQud2
bBcLvQpFok2anrMdEtUYnnc4+ZsEA/7+enV6npvMm1CVaSE+5kcyheC8geeI+4aNQbCZ5e3jVzuv
j+/UY9DqSE3/NzIme9+GWU0xuFtQd9ClFw4qJvnIOSxPu/Ncmtb7SkoRNhPcnKq25Zl/YR2a4ZLa
Rw+wHW8IS0gOWfUtCZM5f9pe1f9dGpi5bAAIVJyIImS/FWUY6X9jMookXACv8q/usHzH/wxFUgOH
JA3oemtAy6i61ApD/3fYY1ass/0AW6a5zeHSM+QWdUPcTzT0FERNMjpZw00BROhvP932kA6kUZqb
Ag3sUTNyrjxitkWxpzgZy0cI1VhXMKSNGLzuGJjeOH/3U3aZF2eDPRK+PqDQ6WKE7gwosau0LRub
or7Cv0isFfNiEhNLh204Ui1sFp6wCMtNiV4QhMPvY2hkIMEw3omSTv90K3JJqTeTTw+YRAfR/uVd
zmkp2cbfiOI8HK6Xnmdp3vmoyRKTTYIYFcxf+WLOLeVOrLkd5dwWQe5471UdrbGlHp14VtCERBQC
fjGgPBzI8CtNOSO2/2z+bVgFUBv+iJB53Seu/VIWW9+7ex5/YiYpXlWjEFPJFnB5HiFdsakS08ou
CFvLdQ1Nt4WR7xSMKjnepZTtZmPczE6viGML/qYmzVbnrZ3UDWcBseVGUXwZ6CkRa6MyTkbDA+qU
hyJZ4g13iysrGlf31NrDUBv6aP7alEV1z18FnFEj7MKaHVKY5pCktUQNlcOVNy/GV/oRLL92PDVM
xvoOB1pSZhZOC5sOb5yJj1OCJI6shq066RWCaRlkknLfkuMrPQRkGpuQB7jgXxh/OI3IlNo+Sz2o
9bDj46Mvct3kMzmGsZDRa7pEizYj5CK0f9j+GcTQDfa9IuYx4/mUkNOdGL2V3CXoIN9W4kmBCGj8
OsTumAXM57BG1DZyte8ZgogmmRmm/3M2wtOF0ZPRkDAT2IBF/vNn7loPWAI6GyTa07bcxGWLf9x3
62oOEaGYFoP4icJBfucdVpQxMJxEddAeN5VaXpDBFeJBng5g2zWl8Lr/TsDpDw/ioWGdgihXyjcz
b71+0w0qJzhDyLj8iRHXaNOU1z3KR5l2rBOV/aqUWNgv43PtLZ6HpwdyEg2i7Zhe16dBUueBQMpP
anBXQIHvp1nfsfLn51adZOK68ftxjnvkvIm8YNJY0WmBEw5WKXvcyUvMiV1IPDEw3XwcxtlRSCM5
XLSs0i8brz2dmD4hF9lAUM6c0tY1pAPuQ2fbAYoPbiv0KFL1/TF6V19tbVKCsoWpJ85V2ZGCL4gp
1yq8R7JggEzzH4466sp6N0cAks/VK1VVTik7davX/fcaABU4pFTHm4KSah9SgWDWm3MhFQXhTgKS
S1JZGDzdOu5NGAMmMyYt4/1AcLU/ZJ/Yigr7kTHBtPqkfnleaP74BzLTQdxD08W8hvxFzs90PRjd
tLAjdFkjcrApKSDkbVA5IU+USMHMwq4SMDchNP063kVQEPxUVBF7APgUip89E7WubUqGfnmIHaSu
cX5Gr5XYr9rgRao42y9Vqw8eAByBUqmNfKVsJbgCRlQqDC8EpmBiGZ4x/AkO5mT1kzTyPEKKfbzU
sMRuEMO/Gb6zvKK+yRw+eqyP8Qo/s/99n9LHUOktKgIXkm8PD5MYowFW/sYL5RWUeMRBzbxVT855
oyHbu44T3Nhv3P3s2U1+LJULlhoE6Zo+/tM4iB246KZnJzbf9SZi2w4AcdgshD5rXpJVk+p+8SVs
f3/xy5JlpkLSwnaIyAggSkZPTQo/gR4FBpNGBwX75AXUDgONT/GQhm/8ZJ/cNCoJaWbctiITCovS
X02ijuW0xfI7HAK5HecZdtdC5lnhKv6UZaB/LcuER/+Icw9MWxDg17mP5hbCqiaunqSBO2FeTGwM
1nHCmn8mwErJOuimm2dupMk38VF3KyTXGR476OBYmpFr6QCvSFXh8Sw0dcyF02tvcLc0LoSumfXs
YRZnmQzSgsIZ+/RUBuNpvWPCPm/+cjo2XbmPCwBQUDDPlkPxXrAtzMNIjZVZtMoi37sAp6UFJho6
1hTxzlGxxh44Z+uYPAZoH8ZpYWAPgNncPy+D7pjOWlEtpkn8i4yz1e4r9nR5pjxflM7ZwCgDBND0
L8aDfWE9MOFOtpRO9Xhgw47RRMmdj76HIjpzbRDuvjMJrnXtWcoSFmgrcxzvneChxo079YHz5Hq8
P3oBlSeGrlCrDRSbkRftdrz34T8+z7kfTh22iX8Wr6WoO/72qxiOQCR+Q54SkuI3bFeqXPHuFwUD
ewkdJF3KOqhAvQ4oShr0NnWfGqSBaIexOPC9rXvPCXAe2yQfiZMBOkq6PgWxHTUA9VYHSmoika8f
AzjzOxoxh9Yt2w2tqSHBAPSK3APH3W/N7fMyvsNXQrmuUkfXG5VIQDMUW7ESrIBDMEsEfloK1By/
K2/WRvlIJcORahwYBXniWEyP6TIkdl7fkkB7e/RsWLjuGci1x86FSAsTxAeNhkUtPFJ7EWyOMXhm
yL/bJ8jNz2RjXgkrn3+xap/CpPV9qrpdoX18j/Dw2sOewvXHp9o99bJpRL0q5qlyaiGUIizOdEJ9
VWeNmw5jMvgpb5wpIsCl+2ijTRrz60GhctEdQKmmA4x6QkVwhs93ljX+1RD7dnA+xKvPLPOV2gu0
IuKCkCIwjVbtrcFhFdsnFFP0k01Fbu8c07i0P5/YFnxG21rgOizs9jjtNuyqgmTivUATQg7Rk5eu
9Uqlv9uqxevPGxCWI3fMrZPONi0sO1XN4qZ1tXm5ciOimJYN3EYlibvzkwmfiKRzfNd8JoeDIhxV
ikCw8l/DBGvySxPES82hlpTnoQV4IKiytrE7sYM+JP8quqTFL//4NT+Q/H5HTWBtLgNOJNuhoV9e
cw65BYQ8ji7g/jaHOmFk2gOddWvYTb8+7i+sWLztiYumEVZiEFLykKy4Og4PkCsukhbR4zzJmhr9
6k7yKTz0AbYgnvGRddOJtwCcp316ZHS4Ea0dTCiqc/fc24WID2TsYF3ZNGp/0Z8R1ChhvcfR/fKq
NrphkmKflP++4QRY26H3QQ4+T0d9Gr4jjPOlZY1QZbQFYbJjQQd6I/C/medNDkaMYhuvb0amRXpA
AElL6bvFAZgu7y/B4zKpxexg7wNmJvTcNQjlyFoGnxel6iQmZb3i+c7FFDw0cUw2nWlnh0HBf+TQ
oXwLGSp991OVPtESm3si2AVzIqiI9jSH+NqrIpj92KuDfq/TlGI7JLRjTTouvgxXWYcQalFqRJ+H
BeIgRGS/bhNNPIt97BWrn4xKrEljXywgSh+JFTR3G6e/6TfI7K09LTlblI3MbKGwgYl5sd0+9f19
qznKz+xlusonpWXXrv+sb6n0EKKOQkaNsZ+fSbH3IMlKloCcSuEFXB0qqDiQQffxHnFr9rpcdznl
u5U7LCPPGHGGmGrIRDqxMDGMTng2Ax6UIFS6gzfAeEKeFqVeV1VL7JZyKrNiZWlvhAhWjQ0l705C
9HEBzq91ARA4o1Xazf3RGNYc8gOTb3zYoj9ZF3K9xiON3ad8pQSjkwCYC04mz0rKq25f+JBH5tMq
QTX9sPpcjD1lHw2//Ln935jcjdMIOyNt6xZ/KyFExudVn5eNziUOPb4Vf6NdY7I8iV7HDJqXB4L6
DeN1bIoTXWfmTeNpWNP6K+laeW3x57ar+7QLg2xOCFK6+9FbdLsDuKfVD33PhR7FndFdmHpb/tdF
VxuJY+ciFc4TrMKMS8AAHmrlFE7sa6wTGpo7qWl/oivXIor4eC5T01dfnRNhl1oz+8GUxSx+wiY9
yoy55wE19axqmoxD48MGtqzuRNh8CTA/KLMxAh3OpN7qvVJdOnajna904HGD28e915K07RI3xW13
k+ZJHyyXaGrwZmNG0nZFgE3FxDzR3QeoEitO4G4dcooNUHR5oiQDRPLzUZBQLuX+biCLBQgXerkj
ICnb7ZivgML0N1VT99WF+gPWvt8Ri0y+K38tE5y/a32KnP+tcMKu/1or87Dq8rzg9DO+o2PprX+x
Zh1YvTILU24XyNMjVQfFpLlz+reBZTz1fyT1DnqWwgRdmPOdXbualdugDFiI4pStpXy9zzdlo6Na
0EZgjnTNAI7AoNc9RmrlLlT0bU6G829cZTIU/jSy/RS7d2W6ZuOepd56lOAwXl1av+HBOZKvIjqo
vAmCLC+9S2XHUDGjPLSXZFkdHTYC0P+8MzwVoOu8EYhv0MldpmFIWMe0xj11UEPZjvdxReTDCoVW
mKyuSsJQeV2+C8vqjTK9ZVXc7WTi6MAq79UMcTvsHHDLQEZxN3T/QTM+Vx1bJEfhJGD3OM/YmXsI
JZpHYSk2PpDN0a77YMjK2iO4RZk+ef0dVVSzQmMScIaRRupm7oJooy9FKDl2yT9SlB3vGqoXoeiF
DlAR60d9tjkGuNK429QzxzPN4SeS14eqjp9UP0NV8ugVJkZAfuy+21InxIomv9/i8k0CBnRRBMOf
z4YBvLiSMB548UT6n+kPtO7tljtCX3bY7uLSzBFIrq4eDsIC4Ju5TsDxpiq/oWwRxwW2weGqWkJg
6q7EvpYD1lK33+mAUJoDYxrTbG+x1iM2I7dcQw0axgzDcPJU8GUuikxOVcdWwej2XQYRSnn3p2vV
bI4mOvoQG57LscrklygtlRCTqCpSQNzMnpFQn6DE9ecaDJKcqZw/g4+uNxuzNooNpvNMtplTgoqY
m9z/7IEb+xVHZcLvkyAI/wOF0FttNaaeEb9nPFowrOGv2LBo8s7qtEJLitaZvl84GkLQF49bPnuu
eeLzIHoBTEMzDEIx27OmRRe2BI6oUzqKWQrBdxFYsI/pMeOFJOv1qKgEhWNsZWnTdvuR0Dg0cZ4o
Z/DJJ52Jt3NiK4UUgNxpnkyLvbb8Ox0Jj/0IcVEseA1rRJa/4TEj8JkB+j8Zlbvl7aLP4pbL0pD+
7rH4aD4AHoWASJxwzyNI/Qw2E93/kXuZlqc13Z+uCn7jZXCXm5zo5T3fdtOO3dYhAJbXqd339zDy
BEnooQ0rmwSGRUyHxmoQHZoMj/3BspOXg4fhqx7J7MLwD/8bntdgfXOHEBqqrPV3r9E7riI6HES9
Ud5RTrv1HTMqvJiXwLT453EqQPYp0OYK/LrM6hVg2FyVmrZzQ4ruJDmcadBq5QnWgcqPiRvyLSB4
hzBmWLqtsfCekgGHvI8TQ+muqtVaDTB9fPzHWGLXN5C10/W9M7//o4nkQBEqNS75VHVtCfhtdaLg
LIDeyk8VEMpw+yyQ8tNVFuhZ9mKnWwfSxRFTsqrPhqi1UN2AzNE0gY9M5Lx4WUCqmzWmcHUwzCR2
/JKRL7vy4f46CSkzq7QD/Z/8dydoJzVcDdGPhuMtVmbMggE3VVGuumajw+C4F6gJzgCXUVkH/AbS
TSlMM+cfXszhQZ4r/L1xNMryCqy+8lM21/EzjrUAAjeAdAB7h1bPBqIIbg4Zx07LdmosL2Zp6cJF
KIHOKhHlVtkYEsAgaBSBVHJmhZVPz2F/UAHdSgCr+DVxFWkXMHuHXHtA78g9opQkXFxChasidRIY
p9ApJ3p8TsVx0w1cB2tROF19aoaiw28KJzgNbPV2xL+6lgGefIE2eoHDjmIM2uSrguMgOjsECi/Z
57+jFflqwmZe8qUekdPk7E/F1FwA7ZDEv17eflTsWr7+Cvm1IfKh7tQGBoJKf4rUdJmhVgd4z8qH
wiN5J2T6JkYAeIxXtTwbfoAgVScUStjrzpLCgbmfHBIaOc2XpvhlrE2Xgt1kBdnubh9Ohf1dT+6Z
VM6V9cj/N38VRyPfv6u2cdE3C4p7kLRsx3VUuZKhVT9QpI/MpeK/hJTg/3lvMgcMxSSAE6NuRf2P
k99Y6ofy3MRztJqt1j1/YUOxbJ94JUCsJMTqunt4mOMQ1e92aARKN/Sc12WpdNs76ep5aQ3LcEmL
We+O0JzzwXuzTwWl6K6geUN4YKlwagJ4r2qzZO7fhnT+S46rK9bmHiZo3LaPtAkS4X6sslnhb5Zu
owlHf41BtcuLgEvRGrpYdyTFH3Zht+Kr+NaFAXfxw817m7b7I6VmsdZNPyezqj1zMslOkAF1MVNA
vIjbWu3AP1+zEvyOzM2iBnKNcDZxb5oJgksVJISZeaDO5nx/rw/nQohVn3ehPTXNMag1ADBCvXZD
nx/ZTQJ4pDC82zvbW+lMmqz23QRqxi9fg8kvUQ9l2mfd3zUClXFUzNfw/x7kCNUUXtQL6HMtohQN
Jy8kdyrYFjGBx+T9yU3SQSFIQagampm9YdCH2mw15f/E6v38sLID+PkeTnPWKKD1zo/CDg7DqBhw
I129gfK53CBRJM/LclNwf5HpOQtz4ydIQh2yA7nwg61x02n7uuZ7vacdEjeIIAkmaMVEzpb80oC2
vXLJi+vHKPdkxLGMvsy7doV/q9x9O4StH6vWuJDGNLhMf35bzVkUDVClkamwURxrryg5jnNpHTHH
ClutxjSFqTkHH+53MSsDkDEtfUEKwTYUyT7h8EBIPz1oZ4eMFmCZ1/pWmfjt3rJsZYxFtNCOoiTs
taM+bCefime6b94PpoH5N6681FpYBGlsxee2jImensXfQho3FHbGVP3QiNAuR5ywYaGZHHihSTyI
+84SqQ1E8JEddPbDcbyCmMzF4hTfg6jIKnMwrG0N/F/D6pxCWaKQpS7t6+ct5luvLvh4lgW93hdi
4Or/CZ4RKdWHis921sz8vzOw/GOQ9vRFt5u1sykfpwTrsiSRg44OhvpiZPdrSyuQw6RmzHzrX6pQ
kb/FYDe1alhwaIemqwnL9naE4uhUg4qRVYL+ZLQDD0NXyLZ9wSRdAthSVvE8WhEuWy96HKDy5cmH
apViYPUfYZV9c/Lrq+URrV1d52L1ZS93TdQE5hlsEk+cbHiUWD4r+TQK/izvbLZ26tETug61FPXI
sWp3s8byL2C3KZ2YWMnHzAs0y0lZ+N20cCwatMR3S6aTotgKwjKifyGVDqvDueDsUUapONf1X6v4
BoSxVO9GnMN48//mF4ujYexvSZCcTbu2IhJJ/bPfskPiMO4pfO9Z3GhmJA46l7oLHX9wd8qeI8mB
/AepRb92R6PiJuXgRcDWHK4HmP/6vEML6X29Mbf4AmGDUttc+wXAqG6/eWEL+MzNYcd4zcLtZkA4
M8P8xkyZ2peG1jvMEAb/SwRPk3r6Iyc0RKrUq0A4yGdf2DIa63SAlWcrxWKFWwcA6Lnzwd81p1EG
X/o2yHCOLBkWpmeuBxCtq555V4zUwYeIQMFKtSAgafIuMkbJBrXATOywq6shXy0qkUaWHjZtIpDv
XpGRpfZO/2ROG5pDXMrophHj0RxyoJkQkNKcTl/YoQ8U3biCEEaNQ2FwZDRvdyydpXsgPsENoyXL
9ixg/rdHCmI9aVA0me9iH1CryU2uaHa/DSTJ7DPMvnhs0KDYWQ82HbDW8TzaolvESuYOPzBYTvHa
VGHscEkAyHSDQRCrTCl4O//U+sKD7qFrWBH6AQuWW3TjoGOaTzA+M6kcG7W/qIolgA7W4fYOLz9h
0PwWhlxWAPR9OoIRN6bP83Sx7ErAQDRmSQgQKBbP+CE2mw5Tk61Syk7sR7f9fPRhzWRo4n7Vl9W/
BJKkOesIXtVtnkGqdqoCkwh8MBhNTDm+hoDEVcNdhk7Zsmh2pA/1Y6WKgyXSXoxhQZ/iT/Tbr/22
N1szIfLHNFTW6QcgowCkSkfYhpGfLo9OB2sJv4jAs3qwjafV1paMRq18T9tVJuv6mP7hVWLj3uyV
m3YCweAR7UZ4tRKLXb8oHT/MSUH6I4dAqElHEAMn8QSu3rs2WdYUKqLjEztnkgmtw7P4is9UsPvn
Ngvqhz/CN3vuuxaQHeO5rKt1WlNfusN3NC+4sFMQQhWe7za+nEaUfFTQxgxNRuw3UnzIN/0CTAV0
axZEbfbEp10rkTpJF1UrNZxK3W4pP/QenA3ZDnEogmcT1NVhrlKK1F6aB7e8pFo0L5bJKtdiNRsG
9N65N62ZVHmLrbmKFfN0WoA4RVuo3259iJC9RMYWa/ihNLZ4t8oIobSdh6n6sXjnwMcYmkt1LahS
zgZF1Gr5a4JkdeYJkZF4OfH31qR/HfU24sv0kRRxcNu5x/tVDc2R26SHlrb5XqOe2ALDwivoL/L2
+QfXtERF1EV7XddMhebJwuQDeb6QJQzHT2aNz6q1J9lp/3MPGbjLWcpeVa7bocSvdBKKK+Gvh2IK
WxhE3gBBMJcsu2op9sDsCG9NiRzk0MJCy8MlYzSD1N7DtOuu95zpVwq/hbMIrUhYAI5q2Px3AHDd
w3NfL0H/F9QBrOR00LcYPFbgDONfSnMKb0knd1BwBFC6+R9Yb0izgvZWHFjhiuHevuzUedK5GTT0
q8E6RwTMK7LMtWU/Kk8Ft1n16kyXzo2aIt3edcmfd2FsDKh1LuPpQqtmtatEtOO7ZiSGdEsONzpo
tkCR8H9r5zW8y1HBZG2iw36W62lF1l7WdZlAx6d1bemXyjGZLYo55NMUwySdIONbIVxckXcP2az8
xMg33eHuFiVpXiuUWbRJBiM2GHd0kh558PCrVGHADRp4LKPzVActjYmWe/6AwilIPTC88FxRfYku
d4RgGWAoFFoT8iGuOsdFGcsd+BfLTRzfx8Q4G7wTWa99HMtBpXxtNYiw7e9YRSn1nemy3TANhN4E
liAO8KbLO3FO+5IuWy52fJ6gTn10iuEWUDCVa7ijO+zPZhSkr2jHqfmSNgl6aX72vUn3KQoazsOx
Dd3a63ZeYV6fSBNjrbjPFEjCqqXLG8RFJj41ZPUmdVzs9hQ8y/v3nlpA9bt5eVicSFZdjNz9dPt2
xDBcQt+KrqdZEQ2nUNsHaFmG4LDGcE5c1oGaNB5ITwsMPiuVGZ8qr5sCI5hW6oqM3mqQmW/jDqSi
hKcO/J+Q83j/r4OdsvLhFS35UU+Bb0ZiTrIIuNKXjb90NCH1P8Urzr6O+eUJPv4c/QIx9Y5yI0dN
ueqX4oRxczn6+1+tm6UrHrGWVUEBve1bNXyZFORyCVE8WA0aDELrXhMmCkKIT/9AS27YaPI7aq6k
1ktZnheIjtm6lZOk2v+WIbnCrV6gn90ANpnwiERvrzvYt/VfvWIVmMMH0kEcmeB1efJhK9zHyOJI
z9ya9PJs24SBS42fJ2ht7pptiUbZAXDRoG8hbeKqwwA2C1ZpQwapxPCHFDTIzRnkREJVs9fuhOMk
scUYx9gMM09xlSXpiRzkH1nnuYPMvTvCqUKD3Ze1RjeLRuqgcIMOkmrWw6lrnRWIppMuHC5DZ8GI
3/f9/gWiIp8wTz9g12wpJo/z5G0JavhuUQvXuGuZLXQi3iFjkR67IbuUs4Lu/viaoCMCbs6yYmrn
2+jSTH96mTCETrvENVNJuB7TtOW6R959Ve5M57xNlWcgertDVv8mQMc+z7hVVDyus8bpVFGSe6Yh
ryrocMOjd6PPqQs61tJs6iXg1Yfe5VmxNjHrqWw0q800GjuN1rm3Chkx4VBi8mlljSnIK6dmAYGu
UB0Sr7SZhmLZJFQL5xo6Dj/jYzeTtFAMcrgXzmwSc5gorAwqWDEsE0zSJ9IsjC7xCfPL/zGvxITZ
IZlso7ZeHkPgN3voJvEFm76CYZWunmw96jnTmT2KfbentvlcrS2QjFCwSYuBEutxSmYGqwMmi+XA
OOqELtoKZBl930A7lfnyBeI6JGz/sFD0aKsNIH5cj4X0KtU8K54UTtcrqUWFufVX4xPyYaeV84Py
25pgA2u6OgtDc2REvNDw1gblwpR+n7aJDCRVJ5IuxvxDgi9Z1EHjg3VKbn1zEloNLbcNt9aWZ0Rq
C5LM1cC0hD5mq8VCya2o8nzYEmjLh5/LatXjRnEaP6jS1wRsIwvMv0d6U0DGfJLImp77GhHiP4iI
+xuQTl3bWpBDjQ4uxbCTn8M0mS3GpHT4NqZSAiXyiGLGBBf+2PKPQLAOK5RWaG646qRqxHdMsIx6
CEzkCwPzMXU6lR8GQakyu63cPf+5Hpyq7RNyjPqnwhra2/Jxbd1HLaDfVg262rn83ZOneUmj0DeX
d+qv7NYsHi1emDI+jlDZlLUR0ixHqbv+LjDbrkZvNZUSZrpptQnasIaZ6eKokan79PSpYnSzdPfQ
ExiRztnZvRcaYbhp8aILLz6RjXBxYsFqUqqLw5lZDYgytI09Iq10QYD69B2Ug0dnutlwUeqbJHdJ
issSbLPrLWFgdGykOZR4kI85qHjJNbPas1JYSWFZcJeqAdTmA8PrdIDW3GmkOhV/HVMrK3Wieoqv
OwBL/v9rk3UlnJqBuW8u+KVW5qMCShLs4FnuyieCw44oREnygYUZlyLzVxZ/VplhpYKS4yrkkrTk
WUa9yopLbQtgte/NWt0XhRKa1ukvE5dqOryVse8vHiXbhelc7LtylUEx1egz4fTL+LlRzaExwRTn
p1EVHqw9o0wK9T2XBsT8CSZBCx0ozRJ3QCdPM3sKB7oF8siaOsmXKT6bNnzsUuREL0K2KYsuBYW0
Op7e3Unp0XfA4j9ldzjSW4YekU6lcOs308dD6lrd/M0CTf3zPwo8OarG9sigUD5SdiWk7+YToXU9
dnxeJ5YBMupBlaCvyXrWWJ+iYNfVjsZ2GwLx/a+lZt6sU0Oqc7dJB/9F1Q/WAK946mTvJ1XHpvTi
7Kt6JTWTEcAXntzoMEu3CyJmCM/9VC4FkRNtJ+GJVlivs58JjIPF297iaS5EaBsZBEZMSVngGptG
4eLAF8e76sJnOz1LqzyUJMQhfbh+yGKZmA3aeCcwsqafNyUjVEzLMzCPt4Wc7YHu7bntZ4ue8LGc
hl5x1jLhlBc2HZ4KsJIYFBlKu3HNmebSThylPE2c+cX9GR+zma95VJrQWmivQBBVjxc1aM2nxcul
prhhpWTi+wEg3ARTTkH9KdxfVUmOqIPDbjykBUd/GD9tQ/pifvcOJxoJzaYeHj+U6jfsgpsL2OGS
/dmFKphvJK2gXtYFGD609ekn4Y98e9x+Tq2IM1uiXEZMeqREDC1qNLWtmiNLS0Yyv6Vsc134PY0l
0lhwXookJSb9e6ObAN1rZBNFOECaqR3oWO6tUxbYkNJhxyj6auApLm7ND8pmgFg02mnIqU3DNbSW
cZQsefNvBA4aBxV6PGXZX40cB38Qdb5aWU1ybJgsfXIpv0aUtAGfwxwxnxZU38Elkg0o5aMUOaAm
k5XB1d5DRq+q8N0n+aVXCLRHhxPKKuAmaAgKs6D/5r8KsiVCvIYUPEcvBCUlkO24PY4p6VXwb6jt
QIFic1uyIH+6ybcYfZHotA7k9Q+Q3R1l5HeC+aXkD0EtDiSTGcuPGPFbUDSMaf5WBr9aUD0MFoBi
W09jVlWlfB4M2aNi50TnA+aIKdFSTg0BLnnfCuncm/LqQr8DQU57ajYxDko4AXty25jkfwKPrDrR
b4JMJ2uE+Y3p10KmVG2EPhy+oR5Wn1tfUpAWLwy/heS+bZmGG4PPeDsSgbvQT9YeHdPl1nRZdATJ
F27HJ6UgFn+tDm61lXbiIuN2PC4sFHod0mh+FCbnQsq5xnprZKu9uE+J/4oB+IEcdpA0mTnIam6y
U1fzdvF+NMQz9exh6rzXo+9AHG57Hj+GonwXlrj4e6/wrVohmTE2H5s3VvWyscrt7ypGV61sUxAP
m78QXI7cL5QuTUU2c5HNX/1p9VwY2+KuU9WE4BhW5Ytk/fGwdKj87ix25sRYME4pFy1SZwkBftcH
jmil6zCSrWoWOKypJTIxcoZlG+8RfpFSE4GVgy/Lke/ZeX8a5hYoy0DWuOWJfqpIz2bqz+1B2vYh
hQ12dpE0iHO6+1aer6BSw4PhgWJToNzZ2nvTvBcraf1ToDiqhU/AdOl7N72Ft9I94a9KZ8kNJJCn
c7uGPmKbck5Mp5nM42uUYeXMiMaREQ3SlBSC5GeKaKMd5GBpe9pz6fov50mPlOJ/LeVr64HFT3Av
+I1KPTZFu+e/6tziiu/s9TGBD/2BCRPQE97qgz0ebfp5NtY5butSM3PWZ9qGqGfJL6pdET+MAv7e
Hm5cJGdckE66u7ULz5tu8/n4ZNAyggZRqCS9f1K/vT68A0L9l14h9QK2XmKuwxh3k2GbjEz1OTnm
39Oh8cJNZ5aKkJV44yrJI59FkNQjY0NsksD+1QsHLyX9/zV/5OSNJixaplF8/EHeGybo7WQM8FwW
8mQ7jpJQmu5IVF+EzI5yfPSn9v27B9WvLgiDLi5IqmGhOiA4fQ2RZWYmKNZwrYT0CMxkwHLrGqwb
H0qMUOt4Ha1rG48r6xXyaBpfd8w/QgDmYXmIJLoZVv5xzwLE92dEOZJgJFnKqupNVl5UNI0Ka/lo
EIw7gZqHqbR/lD1UzNWrtC6AY/Vk2/oIYLzRZu7DFwNbS0uRZzSS7jQcznogeHhUa4ucgTLGgbJU
2xzAzaJtNHmEUoLWYehrIeRdN6uD5Q34D/mnSpav2lZPUfVAjBzmE8ot6j6Dob3ICNEJtzMkOYuk
LEvgJKufH/xbAKlwApNFTg/4LmLB35PiCrNtzTBEraOmi4WJDfvlwlHxS5XHO8ImO3+e9yK5trRD
CiyCreLTF3/87BQL732EIm0Nvdch01uo2oIwzKfy1VF7fI8dW7Sa7wuWRZ3WptRzAEnTKdKGc7n/
Q9cCGrpatCr6bmWFaPcNkWvFMu1IyWz7mkhc4VQHV5quZRnKOOjtKQMfjtDg2PjTZKTOwTyZffzv
QxnxH1CmctWy86VX0f8KNseXJC1GiTbkjEM+OtU79NXNrifD1Qj84Y3Fye5O5p3y8XjOcZzawO/0
i8ZSBo2sWpJCy2MP+CQr1D8zeZIy7kHSKgBcW2a+peUcIVtkXeTLyICjrgpPs9XAfyMN9sAcXGbi
8SfHuWZdCiIbSUNwb0AY/rKpxVmx+q+6FPxhjsIPO1vluAEZUU9uZUcB0wRMHf2K/A5cgkzqAo7d
d33U5LPeJ0LUSrEgFPIO0NK2kJQvEEPXDzfXH5p411wwyPUwlsKUpwNnwlRb33VqxNLh+QzHLPrh
I8ZjugIzMssvfRzgQdEOfr7T2Kx71tDuof5QqqoZte24AjT8KSf92yrbzKLCPiLpq3vOn9RBmadu
nobt0Lph7JJMtQQc4nDg+sni3t5pz0AwUEsdn2NIUpQyYQtEFQ2ENin5he8zHhTMxE23uPRUdPvJ
snd0yt0PyWVPjJsxuYJxowyysfUYjUgexMRFBFp8ljEWrIl/tVz5EjrMMDDzEfkIasNbgjXwC3WI
Bgx30a3FVmgtArNbAmOu9u4aGIHmOV4Wj3hkv46zIvJWfzDp2UI7+paSt8TXgZOHiErqbhttvupU
C43iypRB6njVxlykcpWS5gfNCXr2XUjfzVqDedNpBQxqHv+g3sS3qvhQUiFIdjCvLMhCHcvX2ywc
mUbAH5Vlg1vPaEnpZ+idza1PC0qDfWbhb3b0rTrvgivq++b3lzdPinUr1169S7Mg75N1V82KVtly
BMd/UNdPM/eA+ibdeUOcaOTEawgpgjpFQVkwXzGOGQ/53PVUfRS5g+qsj594/TRVgKOo0XSVINgI
A0qOnQc7NIOas2JPQwAIfSclgzV/9lEEdWRs8zU1iZavj3NbDXh1f3IfpghFJPhPZCWlsnFSrb+q
ZDJ7mOg1u8DVhQOv/bLoZpbqAmzKdV41mMZylxp3VjJH43bjZGrCck3UoJOzkeHp0W+soP35a+wV
vk19rs9ylxvTKaJ4l70pMt7RVfr2Y1W30ZwxIoD+TPKhScTisn0XxgIxQiX69MDp4R1wAWo31fl8
wFKXuFC8guifzOH1+K+TGkLgHcPp3g8S62LC7wmDBsBk2JVeP3IUeKtT/0EC140QYswHjskkjIy8
RGdkmxdvhmbXTe3TE8/VpUloqqEzrvh6JiNNZZ7vCNDkzQYuG50caxceQTpir+TE930rLDwUVsWA
nE3wz1HK4AyfLD00tqzGPKP0SIte5+ZR//77kd9+kYM+yq6xwZiOdnsuxDyVPlQMf0SYACQ51h49
aXUp/j8BTjUHNKih4MkyFHZUh0/vVM5gTsCcOTu8WDifvqGS5hB0lUAKGKGH9bAAIcPSQk8kwjTB
Jp5N4Mupjxy93eknQ8ODFFLaCBRdbr8aam8uGI0WzAPLnxzvJaB2h2551+LZ6DQyMIw+pcwJfpBP
102/mk/L+sGDYGzptsWQIJiuayohySHy/4w2Otb8qCdfcJfvBC9kiUBw61Sua7gHBg9p9bL10ieD
ZamlAhqaoU0ufaoKuWLbHLU2M3qpavvyAjPjJgWfYJCut3m8rqfuT+NTV6fH7u6vz7d0wetkJrqA
6f7+wHdZpTQXsdxmRQpHrvEV7K6JwE87jRWrO3pmRqwACgRB0aK9dvk/OXDTrLtVJGiYj7r5rN0X
Cv7u572Rb+lSsB+HjgDXKVdeHHnW9qhwvkiDXCQyIgjGxJS4OXV5GYZYfsFPcFzmRxAjTnUyB6yo
C+A1wouSegnXRbc33RSdi8Na3BCkvLxHyR5j8d5qxBGXUPvwRTqhVo7jp3YnW3aEoYpefgw1v4F6
Ni1oeC83gqvTIkstJE1+ZW++mpfx/dZtm3os5/8FyZMCnnWRa4xUBzghLqzFnOSnHfPaTI6BtJxm
m5lZzdJKgtp7gfk87P8k3b5VMRUXNxVnssjHQmMw1DlvtMfwa13b+mEp7CCdnNvLro8JDDJrngz8
ntcoQ5RuEDczTjlLeGBoywyDgkq/N+6FUuYlNQh2fbDccE5CtHZR+vliRqDJok4SW/eBDC9b+Kk8
olYDkzG/F7fh6X1gwHZNTuV50BLqI6NC18gI75rUlKnCEWqmPUPH/cxUffQ0GJKh1Oj1jhJvv7xA
ryZP+VaJekFo1JI33bnref4RcudZuZ/+pZmVskYnKuUHnjf+67bbBaX1cKYUMxojrvEX1ETlA6E5
MpX9aMXnClaVcJwbraPBeH/nrwBIGE3yi5xr1NOTUqrfNcQP8I1lPBA4ZqVIWViiKDXFPLivwR9O
pzDJ5wRAzHvzQckrY8aYgbRaaDWeZ7/MM980SRnd0djZTFuDtCU8R2+t/tdvLE5O8dk1bX+Cagx5
pYkzXfFkLx67LpLGFBeh5TXGtj9k9T5t9DG7cF+t9uuLeaM8SNBxvcIHkYAmI4WYkOSK5yTXisYW
RHUPmVYWt5XedA95QZBYaOjThezi5dIPC1P72Q1Hs1SAvpWMGQXaYzHSHn19IGqGM8/2RzpmqWFo
oYx0IBqsCBS3w9gyjjKpg2EUAxKaMWcj8J0c6f7FwncnJ+6O0NqiF+2+NPM/AXYnlo6ZGFSyhAa1
AVSIQzuEBbHSkLwwrKDDttKqkGIHlIR949jJafBvIWNPEYmvOUmu+fr4yVSoUI/qiwJPu/AYlEBg
LYgxu0LASXbsl+tRM/3ZUmciFSNY2BllZflP0xcI6CeAHdXehCf+TK8fNfHy5GWX/Kh2RMF1OiFi
qRvNJL3/Z1vXp2yvp5vmGzpPoq/6PIcmGNqKP84g7pdKj7/5Dpj/xVgnDP+6nj/kZOtTEooR2d3m
gml3s8U5/04CQQxAn8oDI9brrrv7SUAhv8MLqIWpGDpgHftE2KuebSwAcCDGkwgHNEA1Muq6XBJu
KZ+bys78rbl+FjZF0WFObFsgcwnboTmNemMqlzh2SSKVTL9d+AsTW0GdXdxHJ2uYcRAIgE9eVtaD
nQqoLvN6ETN33HQfXKlcp9tqauD5pkvcw4H8TsMS17MPijXn7Ckr1Z8XMut8NEAeaps5u3TjUPEW
nA+qFwfoQWi0ZOz6ujKgNjKC2OYyM7jsIGpU2BDLe0SW1nuq9o5/EXoQ7ZC1mRySea0O/Lh61eYP
BZiTc0ToxNdNAMk+k7sAbB0TiAmO14Qb6rT0+/0yXsF/hlrxohBz9v2zwbsJuIN1Uv/nSRVT2CP2
cAGltRDho7fBtXQW/QwR0MIKzgn/hmbNsTfLAtgqAAAn5EGpMSKauJJ8CliNoa8E/Jb9Op/pnmIM
ydYMa0vEMePlqLhxW6Z+9f1KA2SXzGNZ6iJSgUVKynx2UcVKWvOzomzXnKTXY2zQw6CJh/OXoAPb
Z8rXvOOrviOSuPBj3TXdfv1EqyTLg+8nJ0SX1r9du93wcyh5dEoLhkTrjFL+xzqkHznaxV8Bd1fU
o/UQsEMx1CfkDdReglnWf+V/2rh/UWlLP40Dctp8Khk4J60ax0YdMaYaO7/42a2CjbgbX1P4S6p9
EHIJAV9pNAYzN10RWKt2gblfQ7/GmZ5Ul1wYFXwMNzQfZ4cZNSDITBsnggW81Z4ippmSH9P1fjag
sNGBWpftOC2LDU3uZnOVQZG6mnmSOFA8cQ8FE+7ATeYsA0zf5QQLFJ8UDeIzjHPbxehAwJ09be+N
0TCToHpptIC8s9jWcZmky+CwXacbOdnWicUzls46IfFHt76tUt7tvpx2qwrBHREN5ggGusFYqff5
cCxFG8zT1yvxqnPr3vIqSIKgQwmNSn+t5xChnaeWU5mHpPHpX/V4738Ae6AK004obpi8ZixQK9bM
5vksVVrz3YXL23XMEuEUwmjGgc92ZYaBN4KOvg7lP1Y6Ar0DQ19AEkT8X86uDGXgm0WxPmYlHQY0
xu+ic7Y8u8vmVFa82lUqhV6zUS0rjv39ycEI6e8+Fk8QxWgr7OjnIDMxURiVbEs40CLRkNVN9n6/
82SOrO46KXfxcKVgC/M7vPQlyTvXZ1lWORLTm74FAuXIhXQfFqZMa9sdSKM6wvNfs6nAsnAdL1r/
l89KpA0b9AxmQx10fgml5NfKTie3ZrLmu+uzSVZQYerCL4/EJLpgZEBTTq93y3BbXDPc9/OIM69b
zqzoKnrOI4WDS038gHlS+nB7hquauIG2OUspMu1Oe8fkl+frsEbPnNxVtsfOU61+a60qAVTPB/W2
zBo120OXQEFgR0zEGi7f3QnfBNwd4WVVCcNzTE4MJ+9jDP8Oh+seB2V5lB9VKkthRxeb3QKaAVvZ
9yADmozzWUXgxz9xqyjX1Qr4vRHm5JImlVDEC3SOZ/D7RZIwiwRv0Xb5cMcDKPEOrWSQO0ZrksBR
J/IUWMxG3arkrN+4CdSzr1ppOSQ5NWoNaehTvtUMCqO2CUAd3Lcd47ndSQZNLxNicN8tC7JUtTbx
kHern6/hfkr29inPUlQOsHaL7oc61hSEPhtnHvDeWkHv3kACGmPFa9AQjiSCl3AKLRjw2lhLx4Ac
cRhL3f26ReMShLMaL2UWLkSxIF1thzF25TM2gCZUjlFQV0TSCEfDFLcSQci3OKHV7iQ0H33axCF7
48YI+nv79vvOYLGiBVhlgJ/XQ+HWn7uc37kFOLiqpzCWm513k2S829Es+f0in4l1VgchTvFY3r3c
6Io7T635uQnvkZ66Ez0pFgVhy/6KPE0sWV8fD+qXaZEEz9NrL+CfhTlVv+Jvo05lzqrh/JyzXf6N
d0ORoM8cH6e6zJqhU6iVSYgjJlCfGV1MuDXEJEWCl7p+tG/Im/pLSZVBkClPcPtBipcOpcmYrKq8
CVNFGLPNPYrvv47Aq+DjCp9lqaSzUFCWnsfnOd4C5E5yMbp6sHcGTTCuHVDha3d/FvDB7ZvrOiXZ
5xn/S2cnaV6G3r3kCDOUwLkp31v1qlJBtqiCpbTmV/XHy3mRF9h/i5QojWB8tphBBA7j4y15kpoD
1btEy1E1uuIiqWQPgdmW3VX00G9UynIhKzifXbe4zKsB+9AN0XvlHfRXVIKzKmq0nY1VD7jsJMRj
0ExICjSa96wkrOI92tYz7jair9BiYlP4FMNaJSiNSbZVmWScsUPGbjZ8o5UkZuFdAh2vNaWyR1+y
eaYwlT0UWFsHmuIQ9KfnCozjm4SZhqBnqrwAnedpdUV2xjBhfnqQpllJ9T6PqE/N59K6ukU3AAFq
iU+Vl8mytb8LvDeULoIBW8YSXKzCLy6RmsDRnVLKEascjCIL1/PA2+7nO72bko/dfXJkL/ylvZIB
FAzP48ms0ZHXX3rWnj6jEOk00LbhnGyTu2FOb97gKq/XmnGJ9i0G+p4brOGgSQEC8vzErKN7XR12
MC4SUKKcAmTF3e2aNSPhc5xxlXM0GXXTM5DwYtNXvfr4EFEwftMdFKoYxQSj0Rww9ulhfmW6R/1f
AO5a9gwKLyjoNTcLXgUWJiJg8BvT0frqbiD4m/OauBOlo1gpWck4y/hftYwSUMIcHy7lasOY48Zx
cZg9WvmsVxC+n8783+1UUG0kIfpd4U0EPOCFLhNZqQRQJhMJ5OQ/yQV7qqM9Yz+xwhUZY8xsWNDh
2x6v4prHIii1bh48MfrG+j0trtQWqf5lxkiHFdg9oQ6vLM+VZQ5LTvItX32wj0adLGY2fCNMqnF8
PV0DdsDVEtLtbJjoX1WCZYAxyXB+eBpuuxUF9OTyU/d0xqkM1woW2LnXBikzmzRJcImWxeET+JZF
eiK5DcG41QjXJz6UeQdyc3zNGbHPjXR+tcRaSCjcnJd+wI44d3S6c0CVaKTsAg9ljWXWAy3k2SpU
TyMayY9N1fJP6h/QbNswoymy9+3IQSZ6m3kSrLmkX0Mnd0dBdWKu83z7e26culEKRkImTwZiyo2F
2ofvCvw5FbCv+1N3k+Z+aTFlIK4HhHtLs8FgQASG73UUQKH5Syj1HTEZEBZxsf1AFLXivoKJjxOl
YkRP2c904sdQfU6k0eRybJME5eHUuS3ollzzIJxi1eA11n7MfvDLrT/YnT8ExGRJnS3iNdaxsins
xcYihfWOT9cO4A9EQnyPKtXzVDKtfdvyIIwOtghY4FWf95EH607vjouZ9T8/gnknQyQQAP87f++c
bb4F5u6P3ilXZo+pEnxW7NcKPcxmQ1ZS+f10/KO5tZtwzwVYjG0nqLm0OFMqdnK7V7emJJiNiamc
ZY/u+C5mbaypj9YQvvs1RyTSbxrzFWNCP9aveXpbUFFeBxixcRVpnL/5qqwmIlapD3+PvYWOHFxl
Ys/cp1UaJu/LuV6RcFbCzZ2MCP16pLraSfmtUZjN3I55doPFzM6h0sDa7fk+4h5prueLwM3cl1ty
3nH82q9OR3LNdxwYBpCrMtRasdI9UMHjnih//Rvya7UibZ5yDi+sy+AVM+CBGQN34iMHfmadoU63
wl54HfOBCVtFbI3TKhLaoc+6pq5w521vooC9hvDxlOMO2uedETRIyOTYq3CemV8zE7aroJgMnMsp
gcz5IzNE0DhNu0QxWhzia43KGjUeeUnTaaqsEbKEr8+ZyscR0i5+KqY5BDzXupwufMmem1CpgXhr
6oo9UT1B5oBfQtMNG6rOu5TwAu3Uh8xdOU/StCFbwVV+7MQpQobuFPl1HGlnEjW+Z6/hoDiZKwCf
KKJ9f2n9HT/LMLXw5b/ha41FIC6vEKjX7pOonyQv2sd4gNEoVBMPykoLOVzr080cdyL4MYIUVnJa
s7Ax8NZTOtWgGP6eAB7YfSQFRxhWlzbTrDYCJ0NEvOK9SqlYhzlfn1X1XUd7nj0kITkmWRZVTf0M
HxUJ9mr2F19h7ESADZ0BQZJiXtpBR+MMlnUB29S4S0Rt9fO4ByuvoTBmLZyyzQFu2hp02+pj0ClK
uRYTLz1CXlaZ28ANF4LJoWDWIT4IOhlIeWlGmiXuO9EnUacU5TDpQ1Cpt+v2lULMVrEmgX3niaoN
e2x93LCoRcarYijZJpncGheBkkyZtIQf+drfsbPSx74v+x5SX/wZdYdTYtQysUbwZ5ElFosQbgM6
BOqpH+jye3ItCis41tdAR/FhII9IysHQuwHtWAooxh2yPgsnOqaaBQ4MjuvLL5oQ4eTc0g1VGP7Z
tBdyOPlJSQv2W5Awaqtn/q2Cig3TkR0qqNBGqer62jyXskFozpMsG3u0iWqBjm6PDYIqic9uHCWT
aHQgDtyTBGqNmR03ZdXLeIqHr8B5JxnuyRVoUxrBIRCYc9xTokadHz7UB444qLTXH1c+KzldsbWk
vczza13eGrNnWRdzApNrmGqYUjth9EfL6JNeht1FpFsp8/IcB48xlSV/+FLwevWrP50hRI5K6u86
htk6yPUJsOuMwo74Dfc5HwELyiFs21VH2j7OM6DOdSk/zoYFf/k782D1UMGNEVO55dV7dX71oHuZ
rj0vDfQ5qcKu5Jj8ISJR2RPlcsGYEcVXRSeuF+3tSt08vzes87SiDvgyX7T8ex/stI7tvkf6Ghwi
JVh4BlW7jF1Nv+c4x8VuwXcbpI8VsZFFRvoV9hDqCcrXnrgdt6FSVmrPgd7UZI541FFAhN8qoZU2
VQmBpiRw0ImLj12KIYZ4CKP1N9c4D5OUyZGVRshEm+vV3pMWQoIfYscn7MsUGjU0b7v0+oFY0870
oWVjwn8FtgBATVXE+S9Cul2/afEQJEhlZHKnwemOJ+j0MKkJ0I+MrW+7HjQjB2cRLDa5fJzF9Vlv
aL9caYGHPMrVjcx8R7hypxzxlFdN2v+46vdBhKX9BbvTTXEqMrpZUSvIUxgdw7qocDZjEfuwx0Yl
xNpmwuuxYvIYl+3SWkMDqRJuw6U0cuzbX+CT6i+r9TYg13qoUJpMutT4qD18ND4qCUjA4EhhEs05
eoYItp5sppyzJ1k3w9k1QlMZ/I1hgeJzB8yMrCBpbJA5EbcSUlrCcX3UkPD6fi0N3R0x084jvH0D
VAttqhDUTQc5p38daM7egUptip1YHOK6V+WvGqAbA8DtCH0cFobs+4Mccd98Jr+7pauricbX08zP
l5qpvbUHZamjKcnkruFvH4IQvRJmTrt+uUouHfhBd/op+BYf8cvXJaWCHFRc8x4mTJWjo21zJ6FS
gUjwkYny2O2f8pV9a3acjvpg1DD7ubXwBZtY184J4NyXQ1yeaxZ6bAR0D0ZBVRi8d71tBpgNEKiw
YXRlTBm+GHFE1nOHuHZVC9N1GPaBeyPq1/fyx8Z2pUeEr4mwQNLNHR7UMjrLoXKcQD6zhkoj20tx
DgKU6OslSlymtGNErWdr+srjJy7QMxLYTxJoWWmQlP3haF5/WZula4LkUALd3kIof4+g+H5YY/WA
TlKpt8enH7UTnFgX7m3HpVdXpMThBPfbGxbOPF8RByegepT7xmAAtUbuMfHXAoMXnZ/ZsFjCaHXj
F9pJH+ByT7OutyuR7582QETnNDzallIILQbejbhNQMl30gfqHH1edOK8dWQ8x7bo4GlMG4umr1BF
Eiz0mkGKZPxCYGVic2fbt2WGdleuKhRYabAfoQqr1/Zt87uoqkHpCQCM4NPKrbEcPZtUTD4nm7L7
PDDgQOuiqWN95P9z2kLUnWL9acm+pCNgnCsqRepNL2GLf/E0g83GyQsSQf95UyLui5m6hQ1q/+5U
9Gn/nEQyJql7a0m6yl8mvePc0GtMQWszfRt8s5aoBlGXBUk6PNxpiQIwh4Hw5mfluOKmGz58VyaF
haaXn17I3toQ7hjb1Fp0ObezSXW8CWxsLpDxGYPJeK9TOrvDrooRRNxN9Yraya+SF8rG1uWLDJK0
C24FXA2XxQc+jojMomnmWIQ9z7CnIrgn+dwRtvsnc2g0WON/peAS2/NfqF2CFq3s+EcFrhQsOGOS
fdigWef66EAcJDDzJL2QZBsv5zz0UdhG8R7xkiQ5PquYcmCB8+yYD5e2/ZxcEtYmPeKfpW1Du2eb
HU3b9Z4tAUu/SEe+81H5DOxekGdLA428xsYMIhPnjcGxoTvGUsfIkOfmA6dO4Kz8m3fDNFilLwdt
R9z294rHCWYKwht4KtH/HqIwDVyL45fT7L61IJnVHV7rm1zIp0QP58tCbyJviZ0HfabssFO1qq3w
C0O6LoLdFBFE+BWZOBLmAcu9AT2G8NEZZXIT1s0P9GoQhUa286MXGkyfHuBffF7jsJqn5u5iwQd/
z9d5Fv39SpDOsW5AiizXRLyxeyMOEejeWBoEcAulwuokoIYBwmUr7PQYuJTVcc979bMohq3JlBR+
jokAzsVAyxoNuz5aDDK3LkrnvOqsOwbMGkdL/efy/zt5r99rI8RvlRbOCfJJrd993YLyKaL2QIm3
gOluOC+ciDoJAV7QdYFV4C3VuzusAE8+3ciYO4c0hpO2ghpZ9cXt0ZyJWveTYvEZJ/jRFET1mXtb
wMXXfD5x3MwufB/CsTeu7tqdrHrbiN816G1ui3xlRg+TtTciqmAt9SYWix/hl6MNilU4I+hDcLy5
lIlqbTnqG5KkXXXgdTg++eKYsDLNMu62Q82lQse6zGBtaN+2VOL99DAJCS4AgaxntGXs6F2PqW6V
cuE6AHp3O1gBHokTv/2+ACpvRISu+xdjKtMG1CgIHRx3Xs+CtR0IoaRZu+jxFwxjJOx8vqs7gHOy
EoHRign6gpEOCMU3gIz267niZhuEQB2hnj/zoV+tBMk344SDRdZkNcPVVABCAr9o8NtEO6wC52LK
s3PLWsD/YYC7+tI1DX+P3SxCl6+4LVM/QNkfsDmwUDCTaAaprItzksJtLKifJaEPCDnJVjddme2o
JAVB3234nHBpwgTfdm5buiqJxR44BBLr4MQY7hrjb+QxUzq1PZGyjtOXfaFQXWu5FfmlNIafouvP
1faUATzSyGdWKSq0l+7ck+uFprFjEitknrszz7wnJzbG7vpp5vFfpUvqDKD/MdjSTcSaNm+GOKOH
1pHAGX4mZyIuFa4NDyhumM8QaguSPkr0pddcDmv6F3W3jMokYC7gH3jJy5mfHT/xVNVqknusw5wV
9NLfRa1dOF/SaibQIvfkGdHcWLWNf4wIX1Ie3yR27LcC2rxdq4bP53P87lDl3xg6puzt4plKPYOd
Fsu3uLOwhDAR5s7MMi6EEsdcICU8NVmWBu3pZswKl/sFcwP8wwk9FVKhYrDhikIEVAAvvgCN+JLJ
P13jOiY05QIx7MVi/Onbjr7xnO3HdJBJSvMbkWPXJhVgYHbxgrS63oc8KYigtUzETx/pVLfsya/i
fAgFkQDc3I065y0IWZEoRFvAw2hPfBlUHpI/aBOWc0IfmWPeNuDhM6YqAdRrmE7Pk9efnR2/ZUaG
eE5CIOTH99QloZNicqbs/3vHw6JIL31XP1L9mC+2uTEkCkqGVrDVSKtXzLWHkerKf+h6Zn1RgS5T
UgTT6xd1c7cmm0KXUFcMukBZnRQtwhzrWGVcPQnt2vCf6UdJTKY7NTuc26RW0zX+JRd3Hf+Fy5A+
LulxD/vvByYYe5+qkTrXZ+VtHM05nalKz3nrWIk4EBXdpctQ0R1ikOn3KR1zYQRqHQZPpYYqJQf+
43VsUvpbc5lOr8R1S0GNtR70thoG7mwJ3rLbLwAAqmNQsVNYKcxBDTWDSivOkQqjyquS7ARzyz0l
8bFxUvM/VwACPw1HVrVj/lw2Cfkshml4l8NcjzPrmY8N+9i0fEyUhplaiPK1/utpePHfDxNQ9jQv
+chxuHe8cB+REm3k62pjvtimeoI+NtdeOhKEtA39mvXJbPKG8vMrPCOs2oTJAJwTQS8N139I2qq7
RysPsOsqBk8Kxen8IPIYUOTKgyhAqdV6npGqzexlomHXRYp+tDHxe+NYQsGcwhUxbcPnLojkCRzh
rjVBbbj5ysb3zLHlRPgo/9X+RVzjwntJU9wWlnRxd3E1dUQB7xPkGW3cmQMWHBLV/aDlLoaJy9Cu
9eL76wolc7mZGw9VrB83OqkoECqNTMAOYicPjGK8SrACt+RJnwDl6R+IItAePXPnHq6Fk2bS9T7V
JhAjyEutHfZSA104eWUBsUC9kwwQGr0eToXdprt7BJPjpyz5MapcEcrlPWfdkoI3usTAGoTxTNlG
jwlYQx+JgxIgK0jIoNMOFSDsoj9Na0vOULsidsEZhqs1EWcWh4c1s53LMYth5idj677f1HXunU5L
kwsNmijnK9vyxKwgXzwuZhxKzfTcme7G9wA++2wa6UdjGR4VW3eUYAx5EPaGimPsMQYDVPZdlfA9
1hsM+UoiQNFR/ZhMUf/sbuCjpyf6Pyi/o73z8SwUH8uJeK4VD4FqPtndk/k4fIg39kxlI2r/tro4
7Jdpi2tLff4BIQN5O44rlmjPCfBsv3nUJAIq1+1Viy8wgQbGy5LESCFOT3izh4Ie4hn4U5S6Mh5Z
44D34STSEj7imdNZu1cabziE7jSzZBDA/34G+lQQgDnxeG6c7qqMu/Iv1SxbHsP6EfXHFmAgByV7
gaG7sgjRJ0tOeyAf3DnY0X/7HVt1N8CCLJ7nUdgBN9StuSIhkvh2AUMnnTjpAqGaAinobIjx3dm+
pVKy72gHxoQFxV+Ufa1fR4F/0FH4DsCn0ETkY9s/laBgfSHaKC3OU56xm9Ufqbg/Wk4co1o97PTO
megEX8Mr5mR5Xtgn34aWNe33f55HIf8W8/tAwdRuoMmARawlE0woIMWMm1k3ZvHRrNYQkIkIQEL8
T0BMHekYJL1sA27DyFGA9rGnb99HRVLu9bwrB3V1THicZe/VZjC/HlZbNIlHZ6FVJaLFwGIW30aM
iz2WNxMjZ8vkSuGjFAekukqcD1/SQ/NtCeHyTOxhvcobWkyruBmAQ6OfPPImRbOSm9n3XXi0d6mG
HnNptFSYJyD/Q/14/rtBf9sySNODU1f5WurB9wvJJtVse1kWG3jKh70IWJQTO+qBC7MSnZnTKVvJ
3VgaHrpR4RsyGOE4pKTNU2DU+nk/31IlPtMARLDP/q5n4LEYvydT/ZhrTXUvMb3a6T1Y+5eH7UAv
KTZOQjcI+KpHiKqjwCSmmJY6f14bfW1txUcz4PNcMRMTKGqOVl+4bl6jt1FfLXIYpjyTArufR4bc
ief3SRnLP0nYRqfMD48zzBNkOEJAvm5YBFfcfmsTtBxWDHMFSX0K5k75VLn/ZRqFse0XsS3ud+JA
80vK5UM+v0MOwWMljWWKSorXKhee3j/7EaTGHP8mN1nw3z8IczCtkvFWlJewpkSd4M25LqoHE1qe
hFPtHop6dpSgqw8P5N63HCynJOBA225tfM9aFXi1DT5Pb2QpdACre6ooB5JdpcJPaCD7j5E/C4hv
v8Q//hxcdV6hDT3X3SpNsLVIISIXN3fl6AmIVcGP4SybgVgMzcrAs6/12ulbKqY//El9ZV0bBT18
aTsU7eaOBzuajbplcC+oUuNUTJ8FBhNCNynaXROtU0N/Et80LGkK5EeuiVWEi4ivclD15ExcTC4F
Y3cHcjhnucqFRbYO8wIdaodCEvYC6u2v1CdA3WHGPg5tlBsnuZa3kwYkQrIRclhqeiovNYUQetEb
LtMW4rmqHBGuXMtxFXeN3iPnW5WIk8nS4Fg3Qo6aj4WcZKbrsn5eTNZXs+frg00+vGSso3fk37kB
SP+22tVXPvEQ8WFh8r6+5ZFt8anHGezV+mbIBb3QOGM37aSXpvHez3tvVNsfmzysV7HgTu0xsJTK
YDjUdEKcWmcQaOH6xYItcCgnpBG7S1yLAfPuHIkxziFaMTso18XvoVlOvhbHDghS8klJBCy6MoLr
p4ootAKuKCaRSVZaQHPKW+xtRXGxVdC//bbz4Ga+a6LHWDrn+OzCmN1ADFNZZOO2cWH0mEQDqPSg
NKn07Qg1r6JJ+dr/Q3XAk7MFMTFIrqsego54fQ8kWtmDHJoxXXL5Tgyo4XJs/YDVUujKgxlSBcaM
AqorrG1BYAbp50o0kZeiCLMfv/O/u19qGLjVuESsv7aHryIo4dYfe2dPyC/ylbA1M4HB+uuZyVwm
ZUrnlFXW8KvbDIBsB3AiqFtpvfNuglkQvtplVnaavDyTUKh7q9fAAz7y2e8tDeF2IklxIyS9biVH
DB9hiQlZ9Nhk2GP951eCvr9q/fLGYsCKOK1mnHTHqGfgCeQWgeJYdZuQwQXjH3SN9rnJwqj/XcJ7
rnMcQCET4xl6p3wXmryefVDfmWEdvWVFYAeZ6ygAhf/3DVUqojH0dyD+juGitdMgF4pGbGUAfh21
G7sAt0unNOtWANIs0vRkPhdvDMgkKXg0Ht9ErEqDu537ErNl2dGWblX5IRDjJTf+oAMyodccYOVP
beoVy3BJrBTukz0ptDTrlBVq3UmKjiFczMMsmg0jcc0nvG0VjGxLd4dseg9cAAa3BcG6+7Ck670a
PdyEkAUfqDHNWG/p4EcHjuLgBJe1b0Lmqomhx8yqpaO6Djo41TVLbbs/xgCzrEHDWpPcWXCoG6SR
ScCOZpehWFpvS34osH4fxmeqA4Jm7CVvhO1cbDQJI4CAgE75Nyy600xmC7rsooayL+okznOh4k1X
TxOhXPgxd4igl/jZzQkRgPyaajB8Hrrj/XxOuCAm7JdSQthS+26VF2vXn/cUsA8KPQBT6c+YR4W5
gNhix3b2jJbxoSZmLLEF3eWMIi/5wFfp3l/zahRFAHAjYxp/l7ibg7soMxBbVCxpmHwN2g2DNr7m
53AiUsq2SvwbJm/trcHbtR6BG1XxiPU4T/dF6yFctjhI7yp/FEQGl2wjeirXjZKJhSyZf2ezbqDT
RJ99+rXUcBVT18NDQ5h2iaUffdsrFxCvTXo7iz9vamQb8QQmFyl3ILsLc5j0Gx4JENguc0g1QiaE
3LVmY8JYVRhxeTGiIwAD3jzVmEHDena6tcJGALbUhtBgwnGqgIsgqqBjPGbfsx8Cl8f7O8KO7jAe
ijGnpZ/DH2KkE1LxJYIhsW77ZY5nFSRvtuAGD+g0l2IcgqDf3SyJSG08FAkYQ8w3ag8XsPzXGw7z
cMQUG4MrYC/QKA3M2ASLoA5hjDpkrH1Yv8Pkra5Vkxe853VSbhgx0idpIUePD80vXSX6R8KXdWRM
jYF6GmYRbvFAZPEw32fxobJfVYfugu4Lf8exwWqqZO8z5324cDSMdKkd97+PcuL0N1AQKuVve0SC
ueJ+PuTA2RLXU4674bKb51bWm56m4FXqMat5hBu5soVFRD8MEJHMPHFNkHIsb2WMsGUv5d/dCDQd
dGf+BoPCNM3rhu7D9PhRPLDocjC5pbtRGOVNfhX4/dzEhibM8VwHnSA+4VNtgnaLwqs4t3Qu/m6I
6NXB8+eaxnkIiOJoiibBNxB2JFTExvHT+gRk4/69cEntzdAttx4DdqsUkLxvpcwakaKMosNjboVo
7xRF5FAunMsiWXiEwcx74bqzA8RVTh82IsZr2MssnHDAugiJ+hpB47ss9LbTEhy+RAv/3rQyR5Cg
usMHzPp1O6hTTl0j+LNcfShWYSN1KD9K0ZbBYMIQ5Le0wcu+cWwNOPx7ifXolMnMFp/D18htP9ud
KFBnx66ErLAq1fcA+pujij3RK+TkmFmwAfWkpYczBSzYqdm/xByFtN9l3EJf8LJQGbM6oVgeoTys
XrTofyER9W9okzQG+ixMzWLrqWi+lQx9EGC+wdRW2K7dQ5FwcbcSCvd3YgmS2FieIXTQv0YUH8R5
p6kbp+2hPo6umc95v+zpnuKXPorsTbsRBkzux6WdALqR4LOl8ux5pGtFLnTAoHOxaclz6txEQBH8
ty4Z60INp4UnF9rH4tB5mHMu0EOQRfPgo10wx6av4QxpSjQrPAyVYNHr5WYu3PqHfcbaZDmhX034
9hko/Zb75VMrAdJm6c33rmuxE+Z15zuJ3vrQYpyKOW5OHjNNSDfYMdlh+xlTN3gzJqYEMBjPpw5p
HYdb+mv8lHYyZF374Z/lfahhXaWcc1LMvDe5MeIDHnYmT1lEnywq9rSORO/EgopQbZSOfBSkgau9
4Y1WLGjk46Ml7lbbhQKfVsZsDsuxUAIdWPWz1gJ7inJAoqNNzksu9m0nvcO8jmeXsZEp6MBNbz+1
gGxS3vtqPA7unCflriKFeaktlCArX/gpZQ6t88GKf6TaDORrXl2YFFqJbIst0NQ+P3GIVW+UTXWw
sq27/ej0T0U2fb/YxXHNJWL7HEmaJQ3p++zgj0qiVF2XYKzQp5LBuKpCeV+zIpM7er1MWJdigWGr
uehW1OcdZoZmLlZ7ksNo4aBMFs4tPbNdoWDm0ogoI5loLQL4XMqobAL6C7t5rJjvvcfZzZ+K7rUK
8JU/eHzlvDn8xzBiD0uv4E6LlGy6IZAlETJEK8+ABB+SDwGkce0d5MnqTyuXV0DM/mDY74pr+OFj
2r+XIN8nqeZhZxXCrN301I4HXauAoeBLZ4z6hH7BfQgE1O9LQnqw+oh3a8s+80bwF/FezoV82ETx
Y5l1JP8VqE+2P0mVUVLcUz79ynBIOPRVXrmGbkrsR5funRVZjb+8nMmfgQmki5mvdBO24exmMaYK
k/ArguGnHgCtgN6OOfaL/m977+Z0lv5uSVJgB5WMFNwpz6ibiRRQ/iCf1Q+TW/t5oqtdC+/qIytn
iyQHl9795c1yXvdXp2VaWkvNqsGGxPiBpqCPySxd5oBA5sas1xdYAzEipcgBOv9RJyRTh27K190H
Frd+h4DT6Ga4yGWm8G1Vxhdh7zM//v0XppoPuujnjeQ5YSaxfxFSn0F5CAo6v6zSt0MJMAPg72on
5QY26VD77Ofq+fVcOdTbwCt/NbFXcdTWITo6Dj+Niks5AIcMdMu2I4Td3tuoWjRk17LHzim+AtyD
wDLfqRxDF/PMGIjyYpcZEPJu4uPL0pWCt1V28l6YgwqoKvlz/eoLa0ykEcSwZOaog+A958NdyPLr
V/wmYjkUhf+gERvVf7L30s8gjHUqn/YZpgwI2Ty/ZxGGMhCOXKTx/00UfbbbDW6lUPwaTmi3q6jI
U7KbL/zKwCNwk/yfQZXbWCFRwIiEhVOvyWeTyaHFchciWw4v6g8XuBvPP+ByC68TeylGGgkOYrQ3
ctinH7dIsUO3sE5pHoY2kTqc21YkWAljtKCjzsKBFLwGTyN/syQkwSMZsalyIP/ubCBhq3aYGq7B
hgwNy5NpKDacKEUFGHT+3PHoHff0Z6/yyJLOTHwWyGXHEi6vqfvxOq3PTyOW7RLkDNfMTzB1vinT
lC8wqBs+ZNIfutpqBPS1g+7QM+CaDBKq3jfdA0mc4Jd2iLEqH+XrXj9OJ4MxBwKe2i32ym8TPLqo
3f5/bWIRGkllvESOjLSalfKy3CZgs3OIsk8g2/OOGbh+bNmY73J+sQvsx6hkSH38L56NWEYaNHS8
dmiP1okPSC9dh2edjhVyJazLw+nJVo53tjpJXnRtZcDpccPaZFnSgk+5T8MEBT308hrgimmByIQL
K32Q3QxkiAJEmyWseQAFxnhl1G0ZR1NTD594f2bMoSVbZ4TNX4HAKr4nd/5WslqIIVsfiHJ4JsNw
o+enGX6Lkjc3+0UqEM/PXUhCvEdz34ZR/b+aD8/8nqhBg+Q+Es/4d1QVODjnEulBgA78giD/JYET
b67ihCjwTF/ZuCYb0I9r38ozylM0rslwiSMtTL3JZB+itHq2jLxJLIFuK2m9Imoei7CKF++jIW5/
vGdEfkB3wd7tpCEZbuRunFqFDveMRMf82PIMFo4krkwcTEFwlKQdUYNhrdtwFxdU5OvH/Ze+4NgP
RBShVRVyehgl/PlyE8tWk0AxdfJpaAnLjkAHkiX0IdNM/+L8kJIPFByaVRJwGSZmCnzVvR4zIo2w
JpnwC2N5D5fdhP98MQc7VabOBxvFC3xVziz+J6JkQR+zHtpQo9+wPdP7reYRHhPhrG72cMOnIAz6
48aaWze6hTXBVEXr6TmG1SOqFQYEfCZsA4lgJJTRtWijFw1sXPjZLyF/nUjSl1R7wtOnyqHn09dV
d4e0DOtCvXloVqs6PDbaSG89kWl75r4Su/5wPloz2VYRuAogx8ZZU9vKqisiek4MGd+eh2CpT8BY
AMGE+X7GUefFOrGqN2ySF/5uyxR5McPNcn0AWaMdpA62BCjFZhUDCopMxexHRXshe1fGO8SussUB
2jL1qZp5dgddgk1o2JtEUP4kSjQQ2jsmn6vT/JgYVMVEi31/nfG9S0z3vtkRcUXAz93eH7m7uqM9
ha3cyFmYl17S4XaHnPxLttEdhnatZiU9V+s8aTuVbU1ObGRH63ARetYaudnm4bycqTiS/ANU7tGZ
VNOQROclNw6nb4T7ulLZ8LscTqZaHJC+ExMG7pRy877i8vkQn4Bp9xd3k98Id9RBHMafimKxYdZl
pKHFY/ODZs5cJYHDPm+ce1CTOjU8JRaMm/fhkPabDukb71Or60jk1icBSllWIVfztVacQHEFvMYW
QeSxXFsVG0eeChXogylvK0WTHGZe3JZYQ9bdRWvfeXz3SlTtr++OoTwIiWlXGdWJncXNraLvz8ut
wZtgM4lyvdRIdHR48bnWUrhAYwafyPD6UKIeQsvGbbxdpPoYybKCjkzLTWUSkZFS8QOYEiI4zgo1
+sKpijJR96u2BcbI1ekMLivzJRGyrafI3R3ju4wuyPt7fJsYlHsE4a6kHDlcpLfYcBww/ZeTfAkO
IOLAAZJFWkCNlu2YcvE0Ht4547xCpJCxxMkIgR29FaxLN+dbqKp7IkSFVmD1WIMcgj+OzJRfHt7J
XwC1EauKdbDHkuJzgndMGAIHXW+xAQ9AT/wWoTQ+ISVirwku1403hfYzazkmX2LIvsxcSmFbgqhM
K1Wc2ktc8CrGh349j28RyOlGuFErE+DMG10N7p7AR4+QdxBriJGBqCm0ob4jDuPQ4Yb0SaoHkeJk
SwqVnKY37mTRQCKNWl7N77ETaKvvhXGO3WOhnBW6sEQcLI1PKiFCoNE6nu1lvfw2CuERzJDQjNg5
EIzhDyUrIFzaBrBIbJG2VNT1LvcQNTkH1bq29qP259AyWhrq2CB2PXwXnOzA41uK/0IaRH9kUZWx
cLj0wn6Z0Qugx5I8ZK0bCzzlDW+snh7oN0h3Hk8umxl5JIdAwREa7JchhGqiiYxKYZflUADL++E2
Kjcf2yPyQBuhvqpaRGuZ6h4uDeEE8eymokNn77e2I0t0sT00ciAI/n5UK4gs5XjROmvidjurPmKf
QwyqM2j7Kh8KPOOMFrC4kNEXB0oWfM6+FvRHV2q8IjjcKXhp4Ff7XGXocf354UttUooCBMHd+R2s
6GW7FlP2jIs3a/jnqWAYlbZy8bxb9h8eKzXXDtVJrFSDhvD56snojyYCdvd1CvmCS/WAZt13+7qi
MqkZ8bL8cDPYzoWtnA6AxUd1mLd3SZvVvdS43PEt31srEwQFLC7PRWmC81W2RgX0xAxpZOaBsYka
XCp6dkMjFjDkhbFkQsc2o8Jq0ilVsuPLatith8ufdzo3ErFt4qiR1+j7CGFR27rUaofUfN3DAmig
k77wifFtCFuKpJLa/qq4u1K0Az88nLIOskoUJmjCd3+K+d8g+s5Uor5u3UbiWH5SqHKGiNmH+XZw
9rLth+Bj/uGSX4M35SpOM6Czoh1D7COxBrNieK1AfIp/QanOe9+MenFiYiQZlwfr/mfC6ZLcF4r4
jvoViaS7vfMpPKI8o/fdjzd9ivUYIaXahOd1S0bu+FUr3ey6mH5/6fyMeqANYkUfht6zNoohzsqa
KMWfgiQtx0f6usH0ijfiEGiMfyd+AgJTF8Rv7TWk42pJIQo/8WbvU4u/BckDSe4eZdsQnbNR1FzB
Tq+qPHtjJ8vgc21paeZlNZmw0gtl85/jc9ALId3z3fUUmLSPuMWo/g/97Nn9xz6uo5yY/2bL5cAC
SAzqA3TFu5qIOwjEWpVs3FfX4lGrO5qjUM+3HfKnGZASB5nOzvxPaqFmPV5VVIxeOoWOQrFRbTkJ
8jffXpmBAvNVokq9jZW4qkHd0AMiFWII6cDn5n7JHH46ctRx/uEzlCAyIpRh6IWPN12AusiaNikJ
fhX+Nnz7uqvEyDb6qcyfA5z9lZGsJsirn4WHOEK2ZiyHcgBQd079tBPMq+b9564+TxSY2BvRNOod
p9NCduNdvD9uY/G16cjbEyE1i6IpKMoVJEpV8WToWc8JU4BvhZtFM9fD+OwcxIVMiYLE3G4MCSf7
L5cEkC9g5M/ehtO+E80bunFVc19JMorHOllXLy370b6LOqk5BocESHF5Vo0JFBWu38X4+Lrvu1aK
Ra9FKiQAKvSlZyqqsUrHiMWg5GUEAtXtW50yhSD1bbEe+O/Pnwq7C6cy7EOyqo18jlW9MNEByvgk
EoX3AMAPHtyDcr1HnqPwL3pgTmQxdRE8qdx7Fvq521HyalY8ebZ1dxE9KeU/NdN6BD2v+i5U2M6o
qidig6tF/PYha7eey82G9wxR085ysbL7khlzY931bqek9NIRmlXijKvIyhWphtKfJU0xH3ywOHHZ
dQV3UNCFBnAelF3tiHj9CdRK1FNHikfWdhC9f98CcasWLpc8ZMr+Rxe0RJuQADqa3QkkejJG9gOt
5lyRWe1HK4JpbzQpFEztnPhJ7+yPUpssjqEzZb+7uQ/y+aJ6vlcpCT3tvV5XOET+g5gVvKpakGg4
yMrImgCESEaz9fIY3ZdKVvLxlHdvVUDBBWypWLkr8CZqeGCaLq4V2D1HTyS1BA4T4aCupXtn2l0w
QiN7bxhw6Er/P9ZOef5QQs4uDLPKKBVfi2N8/6GqrIse9rQSTXwnERV76t5OF68SI6J7+KdS6qxL
j9irUjuZm5xrBXzLNMBxbv3wRQHH4WJa6IRZkHuQP+WeLzqjQph3zqHr1x6oAq1OMWpY5Vha8TgN
/Bn4tUOmrRoVe+Fc+mGmKfm06lw/+hAKhSlflW+K3qB9kqzVpxbL7CRdqWtSLrTHNllRRPIaiCOa
3nU3QGsV7ZGDrxOjLJZjxUkhOMf/oq4wEbPpuxt4PiIM6G/YRGmgVdL0Vn8rnIEzGoJi68nm1U41
RdxrSmBqrOytZhz9clKhTJbdbXtdckN6C+IJ75L+7OaxzPuy7yAJY0Vw++9CrsrJ96tJo2+04fdw
GIfvJQafbx6MMS5iG9trvWAzRZo3wUjGfaXrgdJRgVuIJZkg9KnGP7FjwezjPo6y7sc2nSbMCyLj
7FZyXdedK9Ppvqy5g1li5mZRswTG01pN+jc2uIN33J2Qp7eV1sonLek0Um+nu0EyshWoF0VJtLwn
kYFym8gcZgUvSF9XWakWxFz6wYGgWccc0V6CBckplnqj6wwC2Yy4+S8ZZhERulSCrpQETbDshXnO
nLPxQ/9tnnmABWh+9Ro0h8hbfsTVKDMWGDTN8x7eF2Qd+aCuc0fzt0nvoZTkEpAV7HfGNyJr0EOO
1K2w7Tox08ZcO7TZnWwDJLAOQtx2GWpGQZ1yqX6BGaX3pl35oFbPOCsITHG8FLC+0hwDRQGGfQOx
Lnp3wExKSdCOWBHUk55KAgo/iIiz/v0/uKX33/djb8k4KomXLd0ZCWWDsGYXobYo7velAKz5Fg/q
s7zH/3BBPeLlNRfOwriCgjph92ARhtYkJ+vQTMdZ+ADJ6xH8rojoyyULREBGS4NwPTXZk1C2GIhf
pHfgsiEUYVTSSjCIhustSKa8jvgSFeRfDqChduWlQ2EyTMXHgQ5He1AikBbEOlossMFSs+hdbOF+
xmx5TpQDCz7rsHQS8Cz66mEgn79D5S45K/5vuqnp5EMLnJ2GJaDMxoM8cOQ8C9dpcW7m1AUgjsxz
R9cWC3TebxIzHUntlxcPapEyx08FaaFo22dCAm8vZHNXsgzod7uZon9LQsgLiUVIBW10vdUNbqx0
rvAS/19wGwiRdlQDhm4fhZ8gbQ05snyWiFfgXuPqx7Yt7WjFQz86woBlhIMPDjTq79zWdFRq1xZT
vbFndayegoz39bDlArSSdWuQp0UwGUXZuWtTEB7RAU3xE9BjFtcqEvrGWLmNMtpJ923MPFKmlc2X
ceBGrKTl7rxVjtX8TMG75lZFFJxMYTC1AzQ7yLLKJ/svOT3CG4xBK1wg7p/DJ/755HAQr8CRN/nu
ue0MQnIfoG7WQph0dftQ8YvOrJ5gT/rSEYpoycReycPbOlt2fTpJ66mqci8xSEwLqaVdoNdkAOsQ
Ug2RL2jnV2Yu/MmmbWX0GnAPtiCKZLaLRUO0QWGlmLeUBalWYoHUGuzEn1el6qNvLjj4sKhTWXYN
xOP2hGLZxLxT62Awbrl+dPrvA7qkz3B5/0DNOgK0/LWX42u4YLaQaCdRwxB9x6mOTvczPbmOsNTz
4nU5Jm2vKSl7XNC22IxAr9naBAwe+eyO6arcrjCrGZQk0KlK+sca3yovDitVN+z0gWn+9jvrQPuH
kahABV8s6z+FEU5iGAsajL+/k1t2KyacWC/uKJDQ/iRW+FlZwgjRq/C8DjbzVSzlBLbF5X4Bj2vn
BA9c4I4lB3grYUpL7dNWnNgG46TAWwxFayN4xDIJ7bUkG3XGHro+avFFFHwCInI8wh1nmp8fsdNg
cNekrUi3Jj8H3j958VlvZQdYwCEjQdS9TKoJAwZZMK2TPwEHQMkc26HV6g84AsDRzeF5nV1PS0cd
JXQBAO+KbCs/fWM5zDQzUfG8A9TJJu7yMS8jQb+S+VXRjuVXp8fN5RKAA9Q42Q2T+M9PY7DBSFr5
rZ50kYThjrEW/C8VopeAeq7cmzbasiD3UdlQj2ccJDIlGtPtAZHeVNnV+CoZXQK+LXyzVg6NTFN1
Tbr+33r6zAlUmtaus/WUj5RDViCmk9Qi9M7cE8wvnImVAUegD+wjpEzsw5obBs+XKLVFhNid5oJ6
6iZnaY4zadzQ94kOqyrBIZV36t8mJr2o6zB3xZDK6hWNzbrxxdu2nZM0UeMekD9juVosheOi5I10
+zWRHWWnrIIOldYI63fVLhsBIbtIhOwkEAWqC7qAxFcO20tLhLNcXXxxE/SDXzUbfco8ciYK0k0Q
q/suJ2oojBL8Sq8WP+dK4Q8r6DWU0fedDL+BsT/F8ebNWBbSyzvJrDjaGXuWqyMM8QtveWsH6xZ0
p0+iBS7Or34Wcq5uGREivzUwvX8p3pJQWYGyUYr7ZB3SysgU6zn/GmiFi74FDKdL0D6GM8M3r8SP
OhavtG1vyWPaBoin5Zt4QBTrSfG48HqwhreDj49I1T58MRfivVyNnUTV+qw9ciHffT0c0zrBmqh/
ZqPlSfiy778U3/2Yp4wYauNLhNx+pLtJR+h/W6f35d7/OE84RO5BALxsIaO1pVTujZ1o+LCOuvKB
AcvJ0y27zBycB4zj4ejY8rKVJopf6HWoxdiVM3gt9xFdoCv9b1zglBOQsWFWjPyis8fDUYghHnrr
ekjJnkzKnD9wVfDKJEQn8K3e8VYRxpb9RE12t3tP+F8dZYNj8az1TA1r2nn8iepHW/NFAVSTgWVQ
bTlS1Cmx1A5GduWaf3/2w5GEpe7hRMBgmhK+/GgGPibuN9hry8i/SWhHob6tKc4EMe6J7b7zPLf+
C8Z1i1O0FBhHr6qVJGjCq8UukCjUm99JHwW/y9exRIK3GX0wvPXa4BFyyT71sVsuR2pyXnJh0WiE
tCbY+9H+NHFLAs9FWT4u08Y95eTC2psBy2PpUPUfH3mfxilkGwa86tm3gDC7wzC84tn7ErC6pnI0
MjXVelMPFLCXKQQE4tyuHkrSbS/M9evvW5XAEi9QrYyMeDnXjU9GIiRWhzZrhP1toZpgCNe6TIi3
JGbX6PV0jfThGUN5uEJjtXPtcMlAgRQ1r0mGvT4wq089+m8SPbeaXjPskkpkOGe0Y6MN4rPNRoKL
4DiCbwesqyej1e5qI9wpCuOxP9JgwCAJeztg2JuBq77F0Ew0jeh7wJfs/FQin3HQgT2WFRq49BtZ
Fv0Vrh60dEJQBpxKZvxvo9pNGMRFhVwo0g8uce6TnYAU0m+pWwk2e2SFAoTdSmQAmlGuiHGqSf1P
2QV/KyD9lvyKXY9uYzCyEI43lea+Q4X9F+E9asuT0EG+187OHWoDxqVeeXCuzr7cOB3PEf1zYhlJ
7sIa+wn7CvkSWgDLGeGfLW79+bfBgcbWAEjepPbmHzAK3TVlfoC7sb3txtNbvCeRb290yUj/eaE3
Icao9l3fdMTFPTJ2jahYJ/ZuK5H/eZylrW8Kgrxjw1fqU8Yoe600MGQP4xw0bONT8zlmxpaAhi0D
6WN+eMKW3dhENEr0S8jW3XH7PoHlh02/oix6qdMtnwhJkpQzOJtoOnsYyaTCyR8yzq4cldLjvPS9
/r5QTnwMWe88MpvBLknXy2lODh/apkLKIslUL1AfYiUmEOC4paSUrDlqLtxNXOEOtuqcybnDJX2C
G6ESb+5f5niRBQbtoqOWV6rJT7JmAAoKWrJVPh38IfH+/o3bKqi1QqWxM1A03R8hWwvLL+AH7W/H
OsvXkAnpliKIbHOBNNF/5luZBEWSBIizOQsjbeC/egNNn3fAsyesFyBCniBhs2EbyqHpKP6shesd
VWEG+2oo2kfZXjrOVnAGYXPfXNlQ0HwdD6FMiZcdPaG1WtQUUPeiSezCS4XBEUWuyfSkh+K3lOTL
YMtZUOwrmloTVBFZOtmXOCTJzMZV2wUJ4LK+sghNdwTmcrio+GFXLPcxbti2X1r3ZNkmHfQwOmuE
koMMZK6j4a4VQD3bJmMhwATmu60yzrYqydPVZNRnfES/+uDyDoHOPFpniSbZ1MHljRsldwYMdkES
0XAZRlJaErbA3pDKjT7Z89GDI4D2LE0sP7o4EpkSswLgNXvDzkcMtWK35xfQ0bj2g+CIlrhZtc31
pUS393kLIBPBarwEJ+IhL2frq6tcVRLIcj+4IDbbD7lX66pXJqbmFtBcAwFKEKPmYFAfRbfmBrB6
+Sz+b4zO9yxcRLuIDwGZCxj5jFgGO2NLyEFVaNj5+hoi9Q57DNylm/rhkS35tQkVIvDYvWXY2o3B
h2Z3KtfsYkc2n+OHR6VrRTD2rkPUu5rLjncx3z0CuItjWh2ozf5Vzq4/zJo9KMzsQFz4SrZGF7ao
P49Vj8xdUvYdyp5IA1jKHKpFOLC3h0q5MFblx020MDyyBY8tenIL6fleVb5Ihm2KoGYvDeJSOCaZ
UyYIbqgOyFt8e1cmJehuqTxXJtBqJ3kDzAXkrC8NmHQFh1ok6mWM7QPchHuEixFTrsEIv3L9rVBY
wwAMTkMu3up+JrAUfK1OmWpQZYJVat5TZwooMmESlzwbrATNxIOO3LTzUKcKrTsR+WMHgJVmisko
s4izAJKL3jVo8w58VRK0+M3nUCWXL/5KqbVvXReKkQmkgReKgxFMHjyvhkwkqQzQNpA3qZXUo+h7
vkVjj06krkLy7LzksZJpo8ddDwFdvqRY3nATJsE6ddkWQnJhaN3gUxU6xfv6WUMePJeqD58vB5jq
C06cATg2J9e5tVwkTCOAAB7a0sK9mj3jT39ix6gzwSHPuAF16BgX91uyTjQnqnAYbYfxFziPSTkS
WNsHEpCmWwJb8QJ03XKpQHHbnu4qF/cXYmbFS1SqUAGm1IbwMeJVzQsH3SMOqAVyRPXIPy4e8mTL
PnVVaNRfktmrAe2O56xvLzecK59BJGR3m2XcjaMSvd8ujfE97oOcDW+3brYUn0dOC9jD7LHXY4yd
Sdyg7AyneaS4n6bKd3rfuf/loDJ8y1aqje0bxxboM4NhSct06EGJpkLMtMOQQR6v3Atenr94UCqZ
eAxcbmo4bGOkTTLY2nCj/4Zx3Has3/N9t01rgduWRAd/S4ZhPYW5FWuIwj3A53eQ8d1Y+scECkZy
HgWXxdMqRlaL/YofmRYHBnY1D2/7ojhN7+e2TMQ6YwUWJn/q+HjH8yge+PtkNkKYRbHr1h1YkXER
sOuw/K+RNUmno4lW9Gn1E2X/DCe8YYsSdYW2GCB+MarOEmSHWsUE+RYaNjPxOTa3Xp4GugRInK+G
6w1nJ/BvzM3lsKOx+w7hVwnKxM/lEhkCAKJ57YMOBUa28OlLDMYAKJushmS8alZZM7x/TCDOOTvC
Okx1x0lxNhKFtLQyTGBQpWGCnFjA9EmVWRFsbkzABlFF1h3f9Us4EzZP/HSkqf7KA869xhB6njLN
gWRSQVSF9+YqXpEhOwwsoFmzolcx8hLbn0TnHbGtcrC8W69VRRM4B7pnihvuMkdgJ5Jycw4vG0i0
1XAYeCftQYN+NJX0tZaxZkBN1uscuOEkzGoOtvpIuumzxJO4pw10x/1wLYLBVqLT6+QRXaKZMXsy
PUy/tW7W5ozPoSeVgXqE0eYe3za4yAefAoGfB3S8ZoXDloORzXceKM+CbhQyK38TIEIwZhgbcNS6
WlEDqCa5sdNGmCsSAlHvEv1haxHpbCx/TiNQExRSVhwoMRYvBDbvLf+0F0W2zFtjiQUgXSi/zeHA
mBgEYtLuyHjCrqOk8N/ltQr37A8/9poI/9uQNfomWHIp+20rHzQapwB9CSibk5BOtA3Ks63j1Mb3
qdJ4Zbu5bFyV/GeJKXUiHOqmHaH6oErcOlmytu3lJa+pq7NhEoTbJ2dLHzy0BzsZCiXhLJ0I1xp8
Y/i8Q+p/XKwJ0RzDR22aMmL1Tqm+1P5IejLl7xx07+8neKImple3rr3YlgjKjXaajsZRa4wbRb86
FlhxpBHXWAvBZQy1+y7rMTF01cbWSBx3aGwqU8Np1pxCBNul/75Brs0L+PDV4l5jlKCl4eDer+tx
BWVsPLHFDUn7fb4dNeKH8c8uwURg/vaNXVzWG+2UBnceH0wZrLTn8/7iAA7jmTtJABAnHxXZicQM
fLVySM3FAww82E07DZteub4ss2y4BMDBL1wTB+snXV09q3eYbJk2bk/vff8Ek9P/I3b4BFbm2Jnh
dXRrbYhNmDhNr7o7++vuKHEYXYu8tGxkg+B4ZeCrbILgMOehgpQ8ZqNh09E87FArEfTvTWf3qq+Z
4cW1vaoEcwEg36/0eLbCGl2KvbXTKviEwwrnfEj6BCSdUyGtubCdMdID/Za1ow6cTzYtQNnk03DU
jOivGZCaTtDK0ko5VV7XoTrvGTgLiJ6I7qGnCw3Zc/o547lEfZLmm8VNH6svYTUgb5d6o0tZS6A/
sDfbs7DBuSMXitfsr4iY5JnG56MbprhrDal1udWUpHRAv0lHdhGvnaFrrHkJLJI0NoxBPVvGOirp
5d3AAqvJ7rbSRq1RyiunE9UUwXNXxEBPsGzLcVAhNk/H862dcjxr5aiH4sfNcuLIkr3Cb2NLgfqp
hktzgFWx+bNys9l6vl8rKnfc4A2fnHrxBRhDdrZUZnPy/4gtW0snoXmAsCuBw9avomTqr3ZUj+2I
1rEC2uNfLCiRsVvw9SmQMKZSYoR5tJR69TAHONFCRYltEXHXWhWZbJF67Ixw5BrpBd6QiESJKa0D
cXN6O7G/0cCtG8cfb5Y6Oj3AyQrqci4slxt1InjJ526l9CN90YUpRHSXjbt7bObZABsvlIt27Bm8
f/pnWVVJ8sgw7mEo/eEysKy3FCEpJQ5NVz0J2Y5y6+Chx+JG01YkgqIzSbOshe62SjzQ3Npt3jin
5q7Kutb1sOHXLJzuGpFdnzE45nmkRJ3KA0sGbPtakoxyzAvlFjPQaZA2GSA36IZGuJi2MAejv/Wg
KON25H+HTR5rylOuDxLmpzqzJpksSjcPfbCIRRo2BnxKrA40izobQshSd+x0i7qnmkUW5jFQwjpR
uHkSO5ulKJJQ5iobPvMKZ1IWKe8Yrnyp+mMyhUTgcp8XZc5josuOkxvb6NgkmwwYRoLginq1VIzb
nyq/Fow79HbgW7pZiXBJFZgGDKggOO4B5TnRSgiA0mQ6xvl3vmZOERw30yIIMvTJ8kOVdWlAcuh8
t5qReaSHvA8rqeb4nAqiSVHGaiVbVdojhWmyBRrcmaLQoacL77U8O2UWLn37UplTjxuctH/knqfa
uAKlgUh8wjdxZ89Z4qk2k4xjX1hNUx5Hh843cxV2ydyrSFktaowznkP+Q1N7T+vhu4Re6nZXxyCE
w9mV48un5TM8+P4QZ4cOWV8Zy9Hz/XzKsNPFJAnLB3Y/G+3s2/dJd94Ho7imW3BKQPfv1YjbULeM
yiO8KqFqgo/hPWvxAMPxAmjirhuE4yz+VWZvoD8mdba2X/MhWgjJlwpcqkrmqTSlduuqvTC3Wdr2
Y7zYsnsy6YIL3ptTulRoF2IvVqwuWVbsmwKT8C5cCJ8eVS9UZhBH0NIyZ7/Fpqxowcgkvkq2xeTz
7yqJkSi5JqaxxYbS3ny4AzGo3x8yTVUxZb6o7jj02GXe7Vh8rL/yla8qw8teWVXeq9vMe6z7edyi
CpDRG67OeZXE5IsvuTqE+3GxxftAWchjavzVDJzBQkqEXfW6G9YBwhbKs8JHQxilPk2k6+yECcdn
bJIC75jmTLVB2fA9MReNuotjR2dto31pig6H+DxWF9Eq1YLMkLKw5uFJzdKLFlHCVWrS6fy58QIo
Ns0KCuewB8pWuEwrk42ZDnMs4UMGuyHLz5l5wNe8itE2agxTsN9nC3ZXuRMXo7TyhnXqyGp4VB9T
My+mLYkmEhIwdBTJCoA9i395jPTcw0nNqwiGDnH7Ylnn/AjiZnhEd8usCMFrrCah90LPcwUn1sBx
b7QSlvapxm6JoHcnMLJSD0n4ZZMuNVqNr/SUAcgrhJAtl/JNcwSs+xkCxvDlQ/s9Mum1K2gZTr2m
G4qODFSINRgD3P+oysN0ubHuGSDJpPYJhumah/xiO0LXhiJH8FShpXvG2vRMI8SlT/p3jlwa3QOa
0U2MUxKwhXd0HPrZZamOpzH6sLr+kZEQVogE/EBZdWX+R6Nw031ezR7g/TpTHHB5RuFfZoGKuKX2
C6pqTtSdiE8WVUhR3M+XJqYT9xVmF9HQA69OlkZ7/5dTRsoYsDAMIIHgrQNuohraPY2zsGc5SGiH
AlXPAMCPaDe8z0ZFyNZU1t4EYLPR9dYq5ukYEtczRTaeIJg+Srn15sBBNNSN3YzsEep+MYdtmdw/
cTMcIc/5bQR/GhFYCz23UtcRqo8cV1zncV5xdg1y8be7GWwJvJ4yI7CupV+peymU3j09ryPKLfjP
SZlFpJ3zjKhyD2T0gZZ6p5Is07krYYBaf3qZby2II88geZx0K2xBJ8EeZHEpKln4SyugXJVYkRP5
EB2Y/KgZqxFYJB+k15D5XnGWFDdMD35uC19rDLRiOFCLP5G/N4QfHNFdVEG+RhM+IumraZrdYnIs
cxS/JfEaOhZAi4axu//mMdcVeVAUfNJ1Q6f6JNICUmRhqUCtgE9iUJCShtwfpDr8OCZ7GlDjh7j7
ryIhjgRZRa+b8keZaBADIIxOOKwvMQSDXKBrRRCItS45Vi8GVFsgJpDPM9mG+oz4Ho/35A7hwr3x
rcpCtRiHsLHaXsId5p7udsbRaj0/5TN0QkuYv8Y+u3MDtwg3XqcgW5JHfzQOfXM3nllTaQz7wPyi
eUEh2ofRg+oVflZ3Tdk53IjH33l7I4CVE/3fUWWPcBhRfH0kVYAxeeiHO6p51kL9R63MVGPfSlQx
R4a5a1YT0FozbT83mpsZhHY80UoFqecPWrBt7xbc4l6qOZaI/LmBFKzFBBF7Xm3IDH5pHv0buJ8w
34Q2WpRnYmQBg+fAUsrajOCFVcNuXOM+xPh5P7JEDmVYPUO27MowjgdQjlRvccScLVAMsfiY2e7T
ezCLNjBYnmBDWMW7fLzWg1I4raiwzv4I4DO2ez7zBjwOEtbDmMkLBbkqbe8uZaHDomPHbRxdSO+U
SJlt70ANX1oQ2tTuF2QuWaYsFCgYY4ezILA4pqB02qHWYbH4UR+2dGx5ikLuG2gEZvPZVyYvvOrC
Ti6pYvVmczv9R8+EBF/5TdjWFqG/5Rpi829hx8KtiLN8yeCDVHUG/vqA1gMc7qiLeckgWVtt/dkB
pT9tUjrO169SAwbCIyIQRR+G8r7UrGQVSXqGYzvnPzvMGGv831XfkSSNgYBxDxAbk5SkXLuwuzz/
tYuxuLXgHe9wwviC6AlE7Fl4GfkK0r6L5Q1pd9FxhdZD88Ojlhd5SsU4NAUe4puJh6Pi9BJAmZoG
TGoGvLhn4DY8UCPuuhA7UP/dNUeshZ6QNw4JQXmqovuYvL/UyPY8/60RNiVnZmmWKlZyYeq8pOgN
IdZMcbhD4kbgKdrxsOHGLNtqLGqjO0gf+sWN/OUifTIEe17Nr6gY8MGa4LemBG5YsKmwCT3Kz5Xx
+/XTBQ3HYPUgX415sr4n0XLPh1MRrWCYGYlYD2M7f0iyAll7BXoaq3D1RVvcTDXNrsECNv9/ZBSQ
bmGM7760G3CtclbHIEcUW4urN7Wky7QFwziHetbCGJrkPfoEd4hvIT7q4FZCKh+l3pku1uJoYLq3
k1flMLEwjFAcMzY5uC7mvKBTNbPdwU9YeN1/K9yXWWbgrqW4GsJABLDGt/DKoiEH+ik8DGnlZybQ
2FWhuxi4lXacfvIbpoW+zMkuljIsm5MPMsIFJ1bRKw0f4SLWLvAicTHcRerIM95db+veoLb++/gm
8Rb/clFsBDCT1YKsbs00hAGcgSYSPTaP1cu9jO9mrvEEAsq4BPaguDVQ44HEeWD6ojR3xrzN+szi
4TtIffPHhrP43yFBqLrp9c3rD1fhobppk0FMhkx9ZaOftW+oVp47C8VXeJ3hOsa+8nK5KXA345qL
OAwcWd8/Y/CsLoPKuzQ55oExywqBZ4VlzC8+N+j7VCEqgXbodkA+j5uufRnU9DAi/sDdnvVgVaOy
OMWnaR7j+idP0Pgw2CDNSBZwc4vpnPH38oHiANyNL3/jCGXULU+NUBWxDz9uvMNEJexEB3jYb391
zO0VlyvMYPHjP0GXyEx1lBodpwh2w5ExtxVIsGZGuIPwfDXMvjdSwyNkOAskWO6/1C8RdBssD/Cv
u/Uz9Ucn257ZQHvTD//Qd+HRayi4fqPov1ycLoYSmm/goHpNafjzl/im6M3+5J/Xhv3ngVSaCyEY
2pvWDa5Po2YpVHh98mGGhQOelNMeKRj9paVoWIwga+5+59ckY8IOJZ+bXX/MKncp5inf0WmiQwjc
S3VccXcOas8+MH9JcdiM8x4pUVNF2XTuDIlJMkHXRWE3cUr0TXNNS7PUJibTeQSPM4muRYlQQanl
1uBUhcC7C4AG0V+biQ6LRzxtG0j/S53HYzKY9I3h0je0nWrGOuxLKYkuNDG232/sBvAIw8jS0OM7
urZY4hBmo03n2+FVitfXe7qr/PUJ4veKhYNNGSxVL0lSvzz6Xhi/mVzwOy8nR8pAuYffvVemFJwP
E28d+DnVUmstQEGduz4TegaeVWHZoOPguS3a8H2IFdUgDi/GXYMlcd+ECHx8i4/BBOvnRst00mta
FPwy3D8IjdPhzfn6lmAqlmtvQuLDoFOq+8PhTN2vAQZsspw8xN+VnmRca2NHaWeFQIZW7rx99O0O
yPUbmE2IIYkwMIfmsm6U16Wv7yAgn09vDf3DQAMvDFD8gkDqtjgl2bkUPIVKjMyrJKgd2Uou88P1
ijbNqk/7hjgw+Nq5JG7U/PPLqLdIP6JL2/l+wdB43gFs9WtEhLWxntAFgNYqm4bmVj4rJPA8jeek
Z0wVDeUiWYIhuHHfXk9WEboTO5HpptQNMiUL4bAKhoRSc0ZpfDmTprbMgPCMlMs2959QjVK3OZPs
hAlX6CWh4VtBF3N5a6xT+f+5ffj8Wioc7rneHcRvCtZCOPWlTPCeB05UEksL4FIv7HB/w/vG8Ben
7kReoG0qL9BIodG6gDEyWosW9QC9lhngE7QnK+XeMzcOytAjW5aGPWESH35elMNTS71FBUx5kcRv
4KUhiOYelrzA1ED/HVUzUynIiW+XVGXRAm7xQe9NpCkSY6w9iff6QaSM3fdnC4M5xZORMNAIUAXU
u2F6xsszpIwnFjdAGBUMI0oXJiumLB9HbbNpZrFVGb+0o5jNJ/iY3ZorsZ/ynGmVuIu0hm8/XAuU
wybWQe8hb8R3hGb51FQee2SiK8siDmlPxlWd35bEyLWm0ZJrm7ujx3XRWcWem8X91L4BEOg6+1LJ
tTZ1/k6pNxjmuYPsGwUXrDm7qJfcuuFH7VH4sakOYdxMaoMZfUSzCQQqiEbeemUYdrR+aM5LfuW9
bNY788jQ7PqMATtZnK30oqI0ycA74d0PCHcfIG9OBr70eGXdi0QAbGy6ky9OefnmiFawEGYSxkzJ
licQKGKh+SdIylAx4lGXXb6ylOrlMwzrE2SAGS7aIS9MXkneFyb+40oMPjpp97KbgFIBGpPPEJay
uvx0C4f6YZHxQ1qNKYZ4VblWkqH5MTUW2JV8e473YdxbzlzAr9/mx+p347NTdWFUZGmP9bXIJUxG
6+pZEu05VbNHIbcVsBhpT/Z6HdkVMdgzRApC8AVBHeIt8h3zLr5CgI6drcyb4G7SsRCmAtChLXa7
CMRvoC2KAkVWY3/QE/0XZMQuMUmbP8BPyG8+D6VaLZTqnR2dq8A6Cc1K9je8pd9NOgZA8+F1/Q3l
34+VJKMv3xy7w7aIH00fmWj4Puj+H+Sjd/iHVR8cRx9PncRZNSNmfKKdk000jHzbscv/hrDNsi+O
cPam8rf9aWLuq3lkSwz+EySDPCb6UH7U1V6DPW4EjB5HbZpjLafo+7ntB0pgd2cSREbANx28D5rF
6SqkejcD3+svpFyoDSJ9sQPDDnidolH275KQYhkokfimtO62lqSjD/brMyLj/FClekLm31ig9X5z
/vbsF0UysDXEhiGyE7LBRcYaHW4cvo6ueam8Mt/EM6OCD57tQYijvZp0PVVE9oWnh+U8nbFXdU8M
12kVbWy38CY5VIUgD8/gopcGteZ9qXdxxsypWnTIm4QTA6DH3glpFu/AmmfJRzWIF1/CoBi4HfBq
IWu4RBYWuHsEZnvihnrlwJC0e05XYWnDthEK6DKWqvsA2Dkk1ZQHFofOWLrIQlf8lNLI6lRSKhxd
KSx0KkDVdKCgEPhFAaICCIsdzHvftJT4z4gUDEtIC5HQLmsKATy1mHcQ8VyvDnxlO92xBAtgKSk5
+7VD2M3r17rBDb6JirxIq+nSZxmY/OU2MSPyvRSU2XqU+eDnKS+IdWbp6z0QLkU9N9vuDBSMSq7J
76c7GS+zMbjXjQAyg4zF5y0H85qltGTn1873kUYNexYkcoD/beEHh5LTOkOWlS4XDg7sRyy03kHq
h5Jm/A0CyVBnodVwHT3M2tcwkj/llz+Goo/MCxqyUMvFoAcfGzAtkleqTt+RUpNBl4biK1Wr1Q5z
xdzHXG1qdoXboeT2BO+3WBV6YlsC1znXNUkDdTk8bcJjcY9SFAL2TXwA7HMdjhgJMLyrra5yGBfq
JGyFNix8Ek6TZ+njHhNd9Ea/S3Iku6nuvXkCUJ/IXbNt8Z7e9PLVheDVWlm3m3+REj+VtOkhljC4
1n3mmSzG8Pc4yvHUCXkSoUqfVsK/Ana45JgTQkxyOnCgNbjjskPvdwcZquZZoWQRGdrAP070CM5y
V3bNQziANFTDVN1He/mWpIaPp22QnVqKYksIRpoxp6sfFUUUWOGI+njjvz51Z4qnALEsJRsjNQAr
erww7iUnHiadKv1CTtlSrqy+R8VQSYe6IqY2W5Z0Mex4lW5ZwqRnpRiF74SteedRNetD6kUhY8vI
UA9tGpF6wrWKo5l1W//iEa0sVSzg5RLtZV3FbWUy1pnt2nSvSY9qpacj52A0y6FtdEJBxN8gpyP+
IX4zX3N330Qys7ztcr0QzIUfuD0fGHeY1OVkVwuu6+hEJ/fAbPhq447on5oJh5vHyDvZMdBc600X
XxfZ8PNYEQCl4qjF0hTmEuGMkFvxLZ5XHzv+5v9ipz+RpPZsbs4yG/iyVDQ5pUxkR+1WA/ZsOLk8
9gh0dFhAcnSJ+/5uMVoW9dFPVY6QHT/2v70Vvu0NvbhEOCw0Oq9vA4RfPuFjO94CJiPSYlfnMQvF
nC5VbWaxHXimcTopexNq6omrtJKKAvwOvgFxdKDmOeGg7X+0lllfvsg/ECf8YYbr1lP3riXMbZxw
Dyl1NDeQX9oYUaphIZWfHTECy+uvRuTi+3GnjHopJe6+4vjZr2khKzdrO96+8p5drRroxOIeZ7K5
l28Yvz73ZSDKdJbc4UkoGEYsSDEmT5UdlhvkHyQW7L1HhprVJKPYqJZJbKtfaXii/W+h1jhSG7s8
KBxd3Hno3Sg37jmcl9hEucBj3MnTCvlZj7tUEkmvU5oEfHDaiBu52uISyWJ0HjEryFV+aCm/hO0I
m3/Ssruwr2vlzCfsFHzdQoJubmQoEtnkLXvKpj4DylXHJysa1EUoBxCgiKJq7/dV3O4I7p/W3je1
VuGx/30peTNY+ODzE/SDVC7BJdF0iuzzoWKjfDQpPRmRik9pNnqfRUJifDJJ6D1myh1LCGxFt0QT
E4N/6a972P5ws4nrAZ/cnDYnnwCF2VGlLcSXhvIzlLwYAWprDOS77aCano+FsMze94yVrnhxwaLA
eFEaxCcMLpERc9YzyFZjCxKgf7/l5Nc3233Cgwg6aORlbw9y4/1MgVCA5koZuqZHPBErUZQUDIc0
OIrNRs+7wUgbbQ8fJbqGxhCsZhq2DSdcpooIR+iEJwXqwQRlb38AXbqsUIBBtuHXnk8Q99SENa0h
we3Wr5jI0kKAP1aRfqGyQSQHo1DEoo+lEB1QlJEWdWLayjCNynnJeevTwnmY6kno84ysEp9qorod
8oF1f9wCzKqk6PQb5BFuivUU7BPNdIURiGKqXGweL8eCiiu3pwUV9vRzo+e6T1RadxzhduJpizMl
P/jlJhGtLmAsJYy8FgRUhT10CiWLppDDphPamsGhlY5daYA5JDfQYUR29a4A5hcCz1LLnAfLTpk5
5eVeqH9GH9LsWV0EcDtN9hp8y1it86rRK/AVNLb8I/Qszo5cGkOWlIiRbvF/1FMYSnS6EZjfWGik
tQVViBGx29SWG+gmv4cyZbVFhVjhOve7qkSnJBvkrIewudatSLXxeeKjihHM6wSDzIF/X6BsOf4w
es7RgA3QEreNNUrjQZsIiaxaA6/FCV8wWDgxsSHFBcpBEZWfAla40MboBXnZi+yAbxT+6m0UDKiD
C0I9tTm/kVRSaScpzaB9VApcCI7aYRWETNOqJy4blqgj6SDAzKysI/Nm8ZSpEyDpKodj5cdL3SUJ
lV86hzFRXcm5LoPFJxzf6XIY3+4jK7ZgsYicJCVuymkgG1RIRS7jIVfKPOF7maoIorwZq9eUEm06
bb714sP0Fy2QTau8s/nmmh2DLAPHLXNm4GZO0nEQgJNsq9Vm4vOb+IL5h5uqFlwAme9KE1DrBp+j
509FYyL4SpbrLeAxxfT9rp5UKdZrgR3I/AwWJzK5B06Y20YenPptjgJC13lNbSxlmH0IzZ7UR1H3
LhoIVhi7RjFjyOAuKR8K80/GpL2T/S4g43+wxmMYS8G8hUuYTo0WQ6i0ek67NWvYMPh0fr+eI5V8
QrHNHnZoR8phEYz08QkCU2Slf/vYRXbKxqc/X01bTbZlPfefHDRt55yOq8UzVpgaGGJVXzCjDNHf
g6kWNRnyhB7F7wv1OeY6q+AF931rpze7kz/MXvk3F6WbgNUrUtuMZlg7rRiTDzzQZong3yml5rp6
5zUbE28faF4X32EQvP4JZOt+sokRb9yCEtGA/0MQe7vhv08gXCyk/36+fKlYBiTdC8UQBuz/YYsk
twX1RuIlLbdHfCJPLa1s11hW3nc0ffnKu5YB6oeMZXMSp49HN9ba5UsV+2dANr+6acbofDJgjvmd
AyqsUAJkl6IFPE5+Go7MOIHh22+tPoRRsmr67+P+OyMSpDg8+jSgLv2nLd5RUKJfqpsj3bYshp9i
PMdzGrLkLqJdpwxzNCXFADwCahunjYaEbcHBdMHDUr2FwNiaWByNhrC4rtKb8Osmi15rNOKORTWs
Gz2ZiTpSpMOnmypcikYNaGiu7MkMytA8/PKOda0DUPbMHjzGUR/dWLcN4dQZlHoHZt7yBn7AtMie
1mUKSN9bJiVd5OouzS/+ID5kqAnH6xBbupYxZ5ZvStYIWREgDBEQKJITpQdjrJXaRW27F/dIvcBc
n0hUp8aWQfrargouzcZakBSEVQacEHeYhk5NFXwjdB2OVhl1xZMZjESQ1r9rT4lkQdQgqGggP9wJ
4974sUAVZTyQ8P7Y7JeGeY7uQT9xhhuf5MTkOfX6DasVjxKY5B3WycKKoFRzGR7pzRXXqkJ9Nf45
x1bDkHaLogH0892t7fDu+7B/BTunwveE7UOEbpvmPabQa14ALkmR0TZ2A+mI8msKfg8EEhS5dBDL
DFOMvSkEGGerl796hNnp6R4Ge4N2cuTY+UwaLT+XVgzh6jL/hhzV6Mk+4VqOwHUc2dPLAjgixx0e
2FvRZ9D03idF39jZ6gxOa434ug+7RNQDJM6IvhgAG3u5hx2c1C32kzEewTZyTu41K9x2HYrpjqZC
UCFNvHr69PNu0dLhDfJzfHLsO4YxGVB4isL0p9jzmwSRMBq/KU5iuR/HXcY4S3keMrMvyvZl3Swv
1RknbLillGi5yXHSaV7DAJCryr5dEiE5Q/bNVM3wcroR4rGx3wMVfbNnpm8YBcXxDjPdgxREOdAy
+EX0fM+wIZZUGX6LaYTY4qiZNBc9Cp7wWYRgpPqrPLleR5XxozR4uVhCXz9np5LCWmrzWxWn4a5V
cDK9+5rNiF9tvkI+eMithQmq84ICNXqpQUPFREsd0vKa0+A8Ro0ncVrb4wgQZO6/lWrBv1HTTiQi
opOukhrLHT6a4IQnHoI4jPfATjqlMcTlNd/nmi7yqs6EK4O3mKQJX2rFfQNVNrTMeW2xvwSgCqAR
GNa4GRI4I9OssKmaaZbcBpZTyI6eJKb4ZUTECnJ0LmhZBAXeXc8na1wzhoPhH2froolxHa8DIpNO
wc1dT+DTN/t/VRafyk3rqHEpP8Sni8vIrytbSL+d1lpTkoIqEdStk/hyC0m5NhWzj3LOlKUKupyR
Q7tHm3HtIFboMIuE6U/PJMx7iMCRxINrzgeH8qlgO1q1A2huguX3VhRmC472XQaRyIBNzT4r6LjQ
Ql+wRWAXfnGShMVMGBoHN/vYeE00KGXb8pfZys+bQhB8+UgT/TMu2vp5LmifVyPlllsfTh7lI8Uy
MPl11vj1MSchCF3ciT83a62wuHdXijUYzPldimK6cjfqvnQzKx7rb5Lp3TW1OAk5zQJFlwwC3Nqd
bDjLOyVRui9MHSQeWY+N4je2RI5ow4pVYjBfJ+O9uveUgC+z4bFGLv9qb4ePwFacS8FMPkbP6Um4
cbzSy68N/aGneZNeQKoH7/ydPQRQikUugzQLtZcD7FGwvSF7eW1c0nPmjLzim1xgNHLg1UCKMZHG
qQM1Y7bEwQIrkXt04ZaBCE0NmUGiJ/EJHenncJbZmzDqnPF4CRS003kyy+9qmZ4F4OE+nhxGJPx6
p0Sh1QgOlQkQV/1EgEwkbob8oLhPQuHU9/F7dxRF8LoQSDhNuDwCVcCXPgLBZzVnf78H44BTCOu0
LLaVa5VOnSBsHLKxe6cs5wm/9wYRODIAGQNjLenu/FmpNjsKK1TV+EttIKXFdKdZ7ojyMsAGNr6z
eQeb8riSn11u7MwQb9AcXRcBMJQHedX95cTcihldjrtfcuTLdSN05S/5jeknwLJeUeUeTv5wwESa
cYIpA5C8fC2VvPNu2eMHPcD3qotjCQ38Xp3OskfLnV9uucvyoWFirDQFSo7k4hfmSlQ700Uvt0jQ
pVbE4Kg4siiltKgVFuvl8B19fkDxZG7+vx6GIAhv0X9sVE1INISfSbyT2EIUcvSb3XmHXf+v/VHB
i8sY4Yo/vStIwLbBpSd6AklS49TZMytmUVdpvlMv3I/EqYgsAyIvh10uTOizdRBEzU/F6hHD8LZn
XfklRy89BU57P11TouycQx7IgjIiTeoznMT9kFvyCODROeGNKz/tk7D+feNovcGaBFv+w2Wnu25P
yMYZN2PM+rNqacufQolkeQWaVViMiWXNqvGnqNkbDNVLtaT1s+P4828bVWsoPw9MZqA9NPb1K30U
8i6iyAYkFKSbsdAWgdO7UOJ5x69gJr/Cq/2dprT7CXHOjVmqspF+ig8PgzP6Eofcv9OUQZjsJ4QB
L41SkP0zyxeD8oCze7MzRBWdIxZcAm88N1t2MBzxfwp+l7dKo4bs8QVkfv91xM2+F6rMvJ3EVvwR
cUtkjvAfJGYEO9whKHTt5vc8SxW7QyNNKikjdhn3F1K/2uia21pyfsGmt2IE7Zh6oN68yrexB5B5
zRcoYJp3I4xpXuWu8ycfwiDy3YZ0f8WQezXdWg0VtsRKGYJNn9R6/mlvXEv1ym6MqueqST3NxlA2
7qWnFydxzcTl5R5kHz2iGf9IVLsGcv41/f0iT0VMhaLZX3phFn7ZMrzZgIOYHaCVOMPzWW0ABTi8
N/OxhcyEAfRrm6kkfDU7rykMjBcFAaGUGpyG6x2/DWFCBupFOyOQDIn0OaQs7Auw18QIa/jtylP6
h1zv9oKwIbLJuxQ8I54hWiYu6G76H9MIYBqsvMGVDYEO8vzwTTGoTTE/NzArtAjKR2r3lDYizzNc
v4VD7LxzY/VPTb92smU+FBXp7cZaPMS4PGsfne9Vww3L4ui5cot8/c+HlfwQNHNr034/llUVtpr+
DHJ+DGNsD9eDKyTtzsUzkLjKnkeGtSqUjuA+291GhSJWIiJt3wEtLFderlKLDUAfiMacu0MocYjY
wreGrUeEhsBtjFXyrOjRVaSxNe2HsJA9cbSTOaCJa+aUO4uKqj4ONQIxHrMDr29A6kk4sbcbpmVv
rwdXG9VbXqSolf7EWucAMOrDXauhWpGg25LsODi1HPc2XQHoZajWycEKigG9p8Fi/wBFFnq4TGJR
my3nOW1ifUWVZ/jTGt9jYFJqrxkBYbWF9VxfZI1bYcPI5h1X3Ye479zqH0puOOqbv1oia8TU+ZfR
zZekVvlBTPfiVefW/JS8txwTYOpuFV7yi+inFQ+IZCaUhFiYIH9+FyAKBPYI/wf2STC73P1W2eaX
Hl2jh7NShPyln+grnM7pL1XN/P2SrYfyCZGKZzTVCrgg48dPNx+2fSf5wcvQQ+9JZq9XhAEgxynW
Pp1g+Vw07klwdXixygQnoUe4HRRkqNPJzfdT/o+kd+kUMtQ5e8kKf2pWH3BYGIjQH3RHm7J64Z6t
xVRoaQKI5P0Hwa5Tzoxv2faLYFHZM2LDhmW7woZ49M3YWt/Bb1VYxQwXuhriFag0jt/U6iI3Hl7C
fTGzxvpIdYuUPImmcbxon+PguEdQVGTaZdOqZQiO7qnh0rdiN/+FLT1NeaUywQNqf9zZT7N2beqW
MoXmQMGtYBdOZ/8gjFGRs/W7vxaayMryOCUL/pS9XBQjin3U5Y3eq9yrGThx6s6ZUH60bkDqlcA2
eKqpP3LWH8Fq3mBIsp31BtLxV88IwG3508E7dnYwIqVM+HUEX4R5cSG07FcxF79zoH0kjB8bpj16
ecJUExJVZV4HUvBBKIa1ykWqDCnQKuPQNpz6iHwq53rs7qINlfvdIHZYUsKVU52T6JHDAo6Ex17+
uZc45mXX4c37Nfi3UTEkJ7jypmGAg91EKBZu1BLzwrSq/UYmpvi/Ws2GCt0khGzt8kgH4VClna4W
pP5SiWwYYkoxYnGeHpZkLVfyCxVsTuByAnI90DiKAbllb7iIAI2dX61vkvHhl9IXcqPNYznM2sA6
/FjUg4CpJBF9ojwXe4PLKDrvdS/gitW7VmlVUpFq3KbNJO2XeG9ma2Gu9aV5Fp/0Ct3yzP5a8r1g
+NKQI6ISAzrjvP8lDiX21Ugt54R4ih5fKzUdG8FfrYDiAA8snWR9SvhhXi9Nvlzwsxsz1Vz69uQ2
/6vJJhzHDJlvQlPrsl5iDEPbE6r4017do7EsPzYgN5ezTuwh7U6GbVQ4Ks4Lq9E+oJEsT8EGRczI
VwiiM5ZQVDHR5L4tDKNoeuQo5ndYyGPsR3lEzbUP05pi3kQ7b7Zspzlj97X4tMmbe9EvyHA1dfvo
h0tSh14mmTuGxOdHjBo7zYqOSxORrWj1mt475Cez1TI/gChUebTjHZlppg2slumVTQsdmVqrW0tM
QHl4o10RWPn0Lpxgb5AHcRYSszI+8KJM4BJ+Bi4xt86CJvjvohs4BM6EKmtCb7pVgB065djbpNGv
phNFsMYhIn3ldONkGdCV3tG1IlOuieJphbI7+uz36v27mZxYsKY8N3V4oIxnxGxPrxIotjpWnHZy
N48mcKbW4ZUWQLbk00HfGyXYs18Fp3C6xlO9w0xgkTUABcR2a9JLWtItjyrBG7EGXv+TBdVwR1FO
+K6HhLDNlBcpUJMHxC9odqGKgQCMcb1Zom7dWD6OPEoja3T73+MosPE28OyD/M8tC0qqoeiHVpSc
FaP4ia/ilY4xEuIA94DT5wt/S1Upxy8d//Zrg0ZmeNyLu6u4Fd8yznBA5XpzGz3cQMyNRkG2HIgA
KbzytJy445qne++95eYetZdcL9Fqw5g6Jj7wRQBiv/n7x0pWlBG7n6sgAzNCFWEawOA+O0IWQAhE
1HZpDKAyOU0xhIMZguT82v+VWZZPXrj2gOnl6XLc42SBq13NpkvIvEWx64AST2f8aHYJgjw24r+g
YCCYcIQCRerWc0y9OeepkTeFhWYAMmVhU+WfOxUWmDeKC6ec9rBFPRJnQ7k6ihTMo6cLC/9gx/Tt
LCaD7UJf8EM5YACBjTkXVrxdpp3na1hahrmxS2i1PYU+2Iw8otOIfEkrZ/GYpUXP/6F8mBCzutrD
BLP2DKCoG1PE+ndY9ZdCjR+Rf8rC9Ywwn7Ea1HBDZ12WfK9N1ms+ooOUDpZBDafPZhsItaepuh7p
jvLUV4RMbgPaxhcJPGzxsUUpJiLzvR4qEyTPgITLQuceHtP40Z6kUlKGvlrfbcmFQdml6hW2poMk
fYv7yhT8vBE6JZxQPdBTo3IjzjzEygt8gzOafM/I5HMQGcObxk8C+nBrElWFHNZnegDwUSSWxMCV
Nby4PP6ioqaPldlUC9gKlIFrBYDmFPSC8CaeFoKHPISToPuitN36x7rT8ialHdlM0n5Th92+VSWQ
dm3OyEqp1P1XaFBY6S0pFt/QH2VUXCZougCsX9B9Jy8XsoNFvxs3ZtnJ/HgkIEmoAwqa0+0n4ce0
LhXDuGajlxP/kIDLScvwDXXFE+M1uDgfThg4X7uaIoGmvNFmn4xWS9QLIBoy5lIcWPD16psqDkW1
hNoN3pebbMRmPmEPoydOerg0H0fobJgE0idZl7nPIfBTkBr4ihzyn4ppmahxwuxAqxfTM1be044G
e6OrsjpXiACJZpqhf6kGHXMYoVO86Hdhs3ICRGXQUdz54yP6oohqpaY0Q+ApEGtuH6Ay0FwvFXDT
knGObAPfrVXbRo/lXU4GF6MqoPJcC5PK1A3HGWmbCBrvjfaDWIDcC83nvtWfz0xF69Jh9tWwjNUC
zTQIDCTkmugZpqlo5YZd3yIKzM0eWpT2jHSwJbf8w5WBrzA3MEx2YAf39JzxI2cAMNSyv4jdySzG
doCQBJInt0e/gv/DjSBjYB/zYcCntzRaQaF62fOhe0frkcq0a77UH87US0DoshaNl1YqwabqEVCY
eNL4JawrK22cKWOGAaTFwUeMSL1vxyYaJlv7st1E7H8DGH6/8CDEhMkwtv3vw3QMzGQAY7CCoZRX
Y5KRHYM6/wpvwlNUZ2TlVhD6v6iaeJWfuFFu9uGQ8lGzqVZW0LKVLcYNHi34NzscF+5IlnQIov6f
mIMvL8rKPdG8hg4kSFz+Jj3oycjaJztdNyqG81YuwYFGA/eN01qXChIi3Cfse6dibQNJ+WX9O41q
yS/NmqQaiNbzGL5RgD+GwJipkheAnQkicngZ2MDHekjqhdhpA0E8mqC9dOyhzOWdstmJAbT3lRPq
ea896AhJeDixlAy3+AWz3YvF/BBgN6wov9x/cwGm6cpFjv3Naiv5+WFEyvoLpzfQl5s7q/BxQDtq
RaMlwISqgzor4B2HXBKnmZV0QSKLUYHIFL7LAFnkB6cyuRBvb1eZpxtcqbepBJEQ9DU8H4cOCAFV
UQ+3OGGQixiqCIrctGQIG9L2flAPgBtrZqD/w+YJ7Qc8I3Dd70r6ErvDZB8WhgE0KBStXwU5+1kT
QU9xjZWwL1hc62P1r7YrYnQYTsinvXDbY+Lq/ZEOVC+9666Vg2WHp31UnMXcpLtUTbhpHC8yobF5
cUGR+82BaM5kSuXgOvXiaQVkGzdAg3DNsvoS1ij80Ctt+gA35HKNnWCTy3ygjm328TE167WjQtnn
T1yMRlc7uy7Be8ecfRBFEQvEbmyULeINMqSZchk7WUkaRrg7ApOHuZR3g9WnnQ4NGquNVM7XdDXG
hcORR/qcOaTlG9j4tPLpQnnNuT3kYEz1VwF32JIXvDcoX6ZUBJveCODKnL8G+4/lHF+7omklofhx
3xNvkpf10GmUQlBfoYSt0MHRhXuPydLqsX6QniGQm4bW3z9Uwfbd476weBXG8t6d6XSjjlPyRGKq
pvaVde/yYaWxh1jpC2YFFNU91aGZuCmimzhb8FVVtVisUOjPNcyDZTkpNWak8BGeixgNKFcS6PTu
sVlmDp8MK/Y9UFtNwQjL5/p08qUUFaCVBf9+1KLouG0w297I4zEAn5r4ZX0LCA4PiDyqsZAICzNX
SNZxhLGTHrhpFjZnMOkFUU/HbU59wHOvZ2/aP9AFM5RgiE0NtxJSgdsEIr9BaGwFYgcCcCfvxuwL
LHswOu/g7aeDWdINTtq9NnWkFwtPBf5ahQqsFfxZ0jLCE3B6p9597BMqelBIWA18p0kQOZ3ePrGf
ixoqLxuQWDrCDferYj0rTQkzaPgsXX60qfRoDcvqas9Ho8tP3QKLbxduXB6iQdNe/gMcz2L0uxLN
+9KWMeDTR9EmuCifEHGJAcci2AchtSJ/kFnlPERn/yPkpVxsn6UZ0YXMNosK7LBlTHurcDK7PqVE
cLCYNv4LBjCOWVzsXXCaeEXmlYt+QXBk+QDG164Ioa0AUInFY+FJ742/+6R9P0dtiHwRBkcZilMU
wiGZ1JG72U6INykDtDlvKF8ZM143lSQLSqJR1gWlj5l0KjCLkS0aOfXtNr/aj9uE/dFPz70PPXz7
Ap6Dd8lRkk2yNqoLxR7SvjpTTaMAB6jGcwvvGLooPJEUOTKTIYoiMN4sm6PKgD14doU90WIaOzhP
rULfhhmpNe+pSzFDq+w3eK2mjaveVlKK8drBAAPoncPmDxH4N83NojPhXYeGIFe4L6E3qkPlQ+PQ
dlf9LGB0gAlpusqS1YZZWDrcw31h29DTpAj0pQ08BKlu9P8MHQ7GSn9hItRWmZy1cy1/bZROZLAq
lEUIq5F8rbMPdr/qoocP+zZd8uHGt8tRSbZDdXxZ3KZzrPbh/LiXrdae29quYljR3iMgnj3LHaUT
fqjaANlIU82Xjbp4d9UyizOyX+XzTr/4djzGHS9MahzDKioW/K8ue7Al8+exbwbY22PIINYB+Q5B
kbUcWtyMRQWKfEJ3CnoROYtR5ZvtnlahZhuNe5kV6OV+11cCprxsDFXFtP4MZcb+wRPbd8I3x3dF
sI4+ZeQYFgBV7ldrtEYl/t486kETZAW8KIUBIN/lq62ryBiORYSzbYB3kX8PlUwPJaA852YtOKSe
svCyNRnbOSn5aojUUGFBvK0/1MA6iAVV7C+uCQUVQcAyPB/10t3+lyHTMUM4m31PzkGPVoaL08kB
NqrK/WDqlJK3C8ADpbOPunYluMFve4X2RaX5a5h7laKuCEXWgWtzTdd6s70d5WrnBycGohpZGYIv
2GwzChJ1Za65Xtoh0fkJpMjn2nj22NSPaHG4gbJ3daeZ/JvdCpO+cWn0CN6a9fnEYGSlnLwQNMks
moSyRKwFckm5/QR4Xdt58OAJ4HQsEroXCkuhI+GIFrQkIhT26/D6RjCaTW2enZteXXwVpMUcvHJF
P6lpixUXQ7Wm5f2UNLgXWsATdVTJJAE/EJZAa8eG5dz9gE/klUgr6M6IsWIBVV0SEZRQX4ySfqYS
FB2+635rRdstPKFdOt1wu+nMMNugsp0qjixxF6CTpbEM5yzI0ktMwlGLxsOGXhMMDpTOa4KUnfqe
LiMQvBx3AX9UTLpXsvmylgQT2nQhD6zv8HLcfkG/SCkn+k96F1Arm+XnXHWOh/Oa2XBm4NzrXbu1
trOFDnTF5tvr6DF7/yOzCrlHxlWDrnb4aQ3vJ39nqbHwz7wWVoKPHWFkPKf/zBY8J490nBeFLh3w
CCACElQweVsiPVMnyTfxJ0X6oaUs1V9dUWvftXLoQLFjTyW/jWSOacmvnDsLPFQAGWdbpkyk+qwL
jPtTjq9vtEiUDEt5nI+qUTKCkVxZ1MMtaA76lspjuUz3ZuiFykvLPUqjSL+bTA9jawy3cYSNbxI/
pGkuA54TzhrLWBvzC4o2sSzFL19JqinM24ghpMSqJo7VPfx4gpITjB4FbwUJEbkPUet3tVRq3kg2
CJMSmHoBKjP8ChLdfhlrRofnwxTUotGWZ5/32FPxrHZeK2DkYk5QVYXB8h7McyfJDgLRzvpf28z3
33Uwbw9kaN+/A37zWCt5j7Pv+p905UbLiSM5gOzB669zYSrFTKtMeHurMK/VyTkibsKKMK0mH7K0
V0gpXQqOk5jSr8nbassENizs6bhTmAkRWvwwxOkW64vn1vSSTAyOW2iHBCH8H8fdHmRoqzSMpG7I
UJVyS3ipFMcAoBVY+45youht2Z4aOcdGx84Xkg6Eo6+UuWPZ34ywZUAYBBCrSu8HAxMoLu2aD9IC
7ypEj8tvs9aX85fDzHaXLYH5XgAPosvRRwgJowIGQMgRq9LaWQ5rngAO3McCH0eedXzMlE871WNK
+dthYuI/KIW8LiINXXg+EwwDXhPWXjjCjsvsA457qAYwOJTeOg2Lq8rJpqa4nIuvxEmmRsXM6yGl
wSGdvWVbkMhXYXopmIzsn60rqiUJ0Mpqw2mpT03ZB28HHHSRi3My3ABUyaLq179uyQrsmp2WzcdH
6LsQLJyqhwW0RfZMufhqEFk4tl/AUOIhaDm9ryfWbN2EmRVurlH+NBZcq2zy7Uxu7MJ/tZgb7B8N
Uc+mnt+4F0zW2P6S0J4BFDB6zvDwxLpTTxoTzY+EZejRtJtY/vgq4cMxJS/QoW7FBiCf1bLSqsa1
h0nO9q0HQpHkTRE7NPbwcfnCNG5ZjEuimiX0e8iH/UPxgyYVm+cjZXkI3r9QFkaKHFqCdEJyY0Yv
BFet8xDb7oeqqwuYTXfo4OoS4vrWRJmUzIOf4rWPKtSy+UetUL5CUAWwmmnIwPp1tzLDGV6YZygB
qaGSdEAhYGXjvEJejz6NeD9mzen7rZQANq1WHnOgcjFRTLPCZnrPGoVOfAVXc/tKVVZwymFgJ5iI
fjb23G5Tc4gzRpogNftj/tXGK+K5FYdJVqz7/09HwjE5/13bmkLYkguD0EfBEfVCNsWb7Ofxmr6g
5BzXY52o75SdKtuD+RHdOJ+sC8RLRzSGj2Mz5QVfxQ5e8eqmxB55BMzp0gwptBY5F4H5R2pPiWUB
7m8bb8qYuCP9wm4iOD2ZRLu23M0qqNQ28GeFmXGgYxWgOVMAxZzK42I5M1GWvEX5p2FpvH+XzXj9
jt0ZYiQgOP5vQSfIRE4Hc2wVYpcPPnKu1KUtXNAonuy6OveFRL4Gewcn83AcoTL6RkACjmWcUY9G
mhhpKwGBsTt6GWgtcokRbNQp7guUv0S2FcObBxNdT6drFPfnK7Lued/j1pVZD4P20hq1HSVS+VoA
GD7KE/C2n0Vc1AkDD2KsyvE33bAVYBhECsrzkNOa0zrBgxWdI+DJO05vrqrMbmFIlo240qcE1wce
IrWk6r25MgELWBPfOcJBbe2+Gs+sebwt1fVkwYW444fgsOkHMIquJ+utHgbRZqk/RTv9LIuHj5p3
ru64pPUYnpVaMPUvFzGXSNX/jmz58w138pZLX1LNa9WPaVvWOxXgWUtbK/NFTEnuBWmjY9EtUfEj
Lcl2lghkSb6kQmE9jto474Uswimj7kcNcuuoDUYemfYj5Eg1TXF7gclsAaYfok4GlVMcrofk/o+S
ksC4rBsDrr1rGXNCdndZYqEZ4SVa8065Qhx+ZqBJ9wBaH13XGlyJuOCZX0kb1gdhG7Z0O8TEeXeb
lbwQt+/eMpLt8Bpt5O9Ub/z39qODsMBmkiWMSvjhy6tkPVbyXzuWYw7l2ZjiRlpaSjCowbRn9ODV
ZtVHjrzC8VuaLjlwfPfbQ8jqIlCTcnHynXOEKsMT+gZRrVSmRJVua95mTJ8IcHxfKsHbnFTdRVsO
1++cmotqHpHFuGhivo731elBLCrtXp734p0YV+HI3No07eZ+mNJnSClbPiTTt2x5KKZP00Ki7LG7
u4yNFsy34VTvMVwZhOHm+M18ci9omcMCkL9IM97Ue5oMFyrNybn1KtEn/UKNBuJmeoJwBJ4Os9w3
NPRCPqBZ+cE6s/AA7FSeJBqWOUXfxM+FQoXZdL5EwxTSVTQsOJIdP1iLTENJO+vz+bMzKX2YY7qf
pfBi5YoZnRFllgT3ywCbR1dMITy3jvhaA+kAWmPGhyyCvbvw1KXJl2qMvM4AmMlsLLNY2vVu0bOh
xHOAwN1UiPZ393hclwJvb3+RG4gbu5flHSe3aalj13n8ch5KWyGAoZL4Z5AWnPVlIfBWy2j8q0qp
BLF+M1RgVQyOcjXL9euJJkWnY36mrgHyRtcMl+gv1js6hYEBNuhBnEYEilGRD0z1hMTYBijuNb/p
V3oTX94V+CbDv1ioNEg/AjaHP8dQ5LUP4Sm1lo5SwCAzQu2XXiKU3rVmsrEBO9Gfo8g5XZG6DMob
wWK5LCSvhaU9RYIqBbHAKvckdqpManG3upDv8xQAjk8/E5iH+O3Q2OUPimzUNGWZBX45NsU/vbWA
AdeNa8D7FORWBl5tvNjaYaUjIOEZEM3EtLKdAeExqLFW/LIVPiKquwPYaWUpoW4rQzXwOXKPKN5X
1t7l26pX/+LvvOuSVrrvOj4lJy5LtN5I0gOxHG6jVWIQISL5R3hVn/ZASWUyt9/efhWFpvInUMDW
eOfSaZR8W32dj8WVTMA7gkMr1dZvyepJb35+fjhJguzt8GApr04VROETyr155YAbAHDPb7p3CaqT
JG7IB76BkKZ5mZwYo7EYP2OZWwdh/y7GpqFn59OHCBxlGfbdV31rXA1fEf81zBDQdiNh86I4NHj1
Ui/T0dxjhJjDYMhSvvfLSs1918vTWwdthIClUBCp2rusnBAvoYRedfM5ZJvAWPG+KKdkBsMiAbDt
gMG+qR2XHK9jIu7jPlxmCpTkPYrW4maaws4EHbE1gwF7Y8oR5SRzzOLzwjLZlTFIpi37OUM2UWCv
plL6KTR3alp+Qr6bFqnE51BqngM6T4tx17VA+uKdDV73/aFvOMnZeMRIqSvbyVNMAXVzHtKnFZSq
RFLx9siFneNv7BXdLGFMnBZtI3XxrER1jAB9ZiO7hicFDob1L6EqlyAObK6+OGWJDxloI2I71KBX
9T9U2pkYzjVkPUJl6NvSV3FShFb2DO2lskPICBUFXVr+cMdBwzygppi0LgUQ/38A1sO9Do1So95e
WDkp37FDjMjcYq2wEawWvft+EL3WR0LRRbnjKYlX0vOjWxc+LlS5NWXn7jN390q/swVAfLXLZJ9N
3ozYyCh/L50jN7xAG7TdHxI0IyzW6ZYlwBMJUcuD7Hajm/30eqsof2xahlo56lrST//2O/mkRB9r
O/UEuQHC0Cjjwd4a3W3SdfQMyqaO9G/nGPZ8tDNfe6q2epxDWdaF/yBjab3ogC+DTjGVqRckRboK
FC9wNdYjla5iHPc5p7MdH0pKIo8ZUq1dGwTA4hQ+y6FZIKHUz3OYlm9MWxwTCl3tO+Na2oOx+byQ
vi3n2yWGKfVnfu7gN2q24wbqsQ8XZ4v8ZIc9rGliDQR+AUAMnLmUqxTpKQqSoR2R+DrPvjbNi8O3
THBzec9k9D5m7UiypAz8/W3z2hlg/56rsaP18bkPGZ41u7ZxEkBNshjF0Cb4xTz52cys+868WmGg
3E1lfqDvb8InJ2wKTpFMcywxbkTBJRWsIv+c62DgO1va43GqJc9G6b1D/nVA+mPLs1XzakkJekR8
y6JshU9ojps9GfUhdO1g7g1iEuwa0PfQh6cXRWJIBcZ1DcQXZ2FhTjbUV+bcemUZfko6BoebZHCc
gJrl6EbzTw1UAtcnNdpSmCnBHliowupX8n3sBNjVNwWbCyrLwFFPFciEpI/9xMPZNA9Idf2qViMt
PDWsy3DuoRpEbGnJz8olM9IcxKVAyHWfstBLCQqNXfplW8dJxB8ckv9Lm9HhlOv4j3t3FtM3sD6r
TLMkiHbeSL4NgsZuTJJiVYSzCgDGPxsOAZD0q5oNL+Jw7rEy9uF2MQBZivMlcH/FQxB6lGaCGHa+
VL3Iq1hpV2l4VND4NJk/jnXxbVNUEJtDXJ5a5TvX0w4fuaU4pG0iMd8KRVs422LC6HCW7CjQSrRZ
AzHTwtnuWDo5ZP5zMolTpwoTVGFS45/HBmduyUlSUbj1EBPjc14KRKlsYeoeT27rqBR6THRibMLG
8KCSwEBFcyzfXRXUNJdaeg8thq8lsj5OtzavXYfnrsC6oYvou7zicXkffSxoMKKIzrpZfAj2/E1O
cIq3SqIPmvV23FHeSPmZuV00D2g0u/qGqbDdM7uZNI1QAVA9JQH+nogyaNhBTfYmQdFJ6xUPH/Il
unR4AztpDB3h522OTZQPOu3iMHxhNBrWyvwKJBslxzT7Iq8tljGX8VupV2Bg31lpr0JNz7jAgDIl
UG0SDO7GXH0L0cgdIcQGReEpmEJ1mPudzEXeEqeOBH1ywLTAU/tdgt+JWxV2VaHWmoCO7Q5n9Rz4
pCtxzglLdlZhRW1rz3rD6XQnmfIgOYf/OPmXdLKAS7phzv1CqO4yFKWNl0f0anq7AElej04AEbHY
Hf3wvQMutN6MhNYfWDbI5I8j/WRyv8L5d7SFCnO7cTkDCFz5ofmr/9va79hdD7fHn7oDz8zNdyra
oSFg5MD0aU25s/wFY3PIry/KFPxN7X6bgpYIwU0MnN9a+pJHH/GjT0qQCXZioePgR+MV/gnxjII2
xdfr7amGSli9TALTpn7bbc772NvsOBhxeJmt5j+OiDFC8oQs2Z1Rb3UalDIkCQnb9pz8zX8xPdSB
DzwmAlE+uiG4K4uLEmaNmAAzwzQ8Dp7nbdxeRlU8Trvq+k0TFUP3Ms+3km37Nz7UPhnvMomnlZzK
JCMflzpBK+0dtfyiE8X9O79UyfkCTu63hqqxEXr2zt58VFYQgKDhO75YKpC3GyTPgWdftb2I0TVd
RwtDDrXLVmlHmxPUat6ArCAD5MQs1p7FEvuYjFURJ+K/S0f6JTr1VNus+Ae7M2PUtZvca8e/3yxB
wGC+x1/anKxLT7oZr162/6g4nUFxI4hKGB2HliBBNvUkCo89EmLSnnsd4h5v9MUPTLvWLstcWMLx
xeoUjCfOP/lZ1exCrcqH2eJXczXr9oDV0KeJwMB7pssICj3zq0KosiaP7AsnMotj7ygbqBnUxD2Y
6tiMvyoFBSKHr1W8ijrwwjnHHSpAk+OL2QSK5/jR13zLW+y/I1sQGb4BVNXTQ4/h5zCx2OCp1soN
yfSJBFRnaNFrKBAbPg3LQZ2TGCkXxWvmx+LZN90Ie5q1J71KQOakfUT+SfcyI+VLMWsAJ1L+YQ/Y
f/UGk4Pm3MnWxhm08VvUH/1kzXJEoEZ6WOuZeBtgYtV/pivjbmORWSiJ0EFG3Eh6SSZXLCntMcVv
l8E84LUpw1QbUpltZZPZ+thMuat2Omz1RxG21D++9J/ugpoFCUk0huteOPZXO7fVZi189M7gLZQM
g+LK6+6dlXakQ2bBxKD3slCGd+ABG+MBhEj9+9yank/4JxSB85QbUDjd1/KWzhv86YXyV1aN5cCF
frh0SseIZ6OhMHgOPAphsJ8sOZZN23JHXqWp2oQfaqGHMADEWKnSxHz61jEh/nIaLYFWtb8prnKY
MBeuiwp5wAiFZteMOVsUQueM5cl9sIPncqEGIuHYnq9isy4ztd0TK6o3DLahWsC68LCScZaJGW4s
8XBhe2LS8vivFBHO1MOz6oX/SmVAEi3RKtGdRH/W4D2B2MdRxErukLdspgeK4y4yH7J1jJDj0XYR
1lwYgrjDfAATXb2daSyr0A7HWnTH82h9C1Mtswowxm2ptnkApfOHoh2mIsOXdVfM//l0p6xOvrO4
zhyCk7by+JJXzT5eYHgow5s+WdGD/zdhZohlt8CbtbgPpqSDlJKlfs3m/MScKmG4k1MNbAimW75b
X4Zn/5tqcVULdtQXv4jZAC7OyYULWu5iFvjLDZjNT6F7dit/S9bbPyYAzldrvRY8VkSK0zH0ZQGn
8m59wbZr3qWhySy4GRtOTD+iPyKufL4TQA1HfBGD7KtuxVqPHOHCo3cGfOWfe4nhR2BmG9cr7hB4
7k8I3hGeJpPIvbyg06OFaSrY5mnkGAJ+G+K55UNLpuXENdsB9dKrYwuticE6p/wWQPrf8hB7aVgj
LRyUMVlo+WD2285i538QzSp89TvHnH3AbePKv28Ppc3vEek9mBWsJXkljem+hHkypCjCz6VzgF8o
62Mhhb3tnsrY+quvFS8TF8ZlDd4ipZyV5IxMzw+DefaU4IRI7H2CUdBGk8i8IEbm56NK9oXljARR
ZXuB1Kss7eAYOdwJNSb58J5FrtiPuT02OfdNlmUj6wwoSlUsGUZQFZrZ4awgCqbBouBipf3Ocn2H
cpgz1On2AZlitTZYrKaYMGqVJv/AgRa5mWzjPlbtyJqsfkd2gqQXg4xCfNCmJOhzN4Wbe+fxINt8
w3QFkzSJ/zuA8dFPtPvVxfYvofeWZ3qT/k5oV8grSfmOhmgPMbYTFWxmcjGjuq1X9pY+1G3tr6J5
BQoCNb1XDFmxSp/yUoUVFoADQpeSIXkUX8oIeUxyDHOYk9caChPABJmqQMpVWF+Rq1Gxgi+Hd7hJ
Vo1lYkO+2ZWjDyX8XfQejie7RDfucAioO9jkNnIICmNJAg6wbcVlyqdW0YV4rAuJRIwiXJxI2Ya3
7QKq4Cnen/53CIOU+9+qEOrA89dnhxE8s4kmIBuoyf6K0mwjDYnggT/RAzdKV9x7KDdmOPixLXB/
rvXt04w4CkMXI4Z7Dnu8veBtBpPNmMAo6lEi49v7GVAUCnYDJaHVvIxNTR1tqgBR8mUWxsN9nLVI
3/eZM0I0K6bXGQ6JmD3US49yKmoD/rg9zpzu8v/IWb0kWepci76FPCUzIJVKd8IUGY+SWdJgJHaJ
2tT/6iEyu7jmP4WrzGwjIpuVUFeg+PHxtSDiuEdf7MHMpZXskWw+mcAmbhRBBvSrEas+QitA5Rey
nMgEC8yW5CpQ9Z8oQVpypIcp4TNiK7YSCLcvwsLRwQj9L+4OQ8WemQxKFuUUbrWXT1RBoPfrt2U/
uWoY3wBgKg25ktTh29zSxcfE6TAmpm/DR1zpyAf498aufIIE3ttvCacRVJm6F5GtKdzheDM6dil4
2Q1YIpwFAJge+KPvBrEWFKUUIvIix2z0hKyVfvvs8Q3PtO68D0+CZktXJwYErv289pYwjuuf4pTN
R1vX1etMASBPK6eegjKS813SDd6s/0IPyjpGliSCUadKNHBbdfXk6f5Fcebgde0mfjVQVOdYB9n2
Lz3e8DPvLvsT6hlUQKLXwky8MY30OohE/rMoFFr0qa1XTsGq2pivgrINb1cig3CNbH4PGDmpxTl2
eAZ4ehYD2jwF8scoR670aSGvCANFsCjI5OehqmUAdGdkYUeLHGO9zVYAneLIcgX/HriIubZaDbgv
qw0LShSL1PXJm5r4AYk+RRZjbNoGbuoTkRbc0Ab4vMuPUZadZ54xTcnBaMw6jQoJA2RXAxs5hw4n
CJ2GVRJ5SrKZW93TqAroqXqhmYTlpJg24LgynDHxQzxQRaGv+LemZsyTVWQjZT1dc3iCnppJq3Ch
XUx4JxCCrWtcIWAhrxX+HEFh2OtI5yywRJWcL6FHmm1pxXB/vI+tgVG0bnv6pX8bTWyJX6CwfVj0
BKcSwoszJ4kgTH71LFkgH8qOZSmvabV+stVRhpxLHZQrCFnyVOeJqtzMpLjLvY3Tgmuf1iT88H98
vsGwbdxnnweIuDmnsgW+pCIXtXQRfBIYVosmilhhRz6gYZO91fhhzlSH9XAkAhIiv/TN6Feiliu/
NqdZ66T6R45yHOzc9DdZr3iKqCmu56Yi7ZpW4ZmlC1QdQ4Z8qdkCRpboDJkdPJ7p9thZscDLGFkj
r/tiZNxuLyRO5HkJhN8EhlcbHZ1eKAkxUbGBBusGVE6IUeOSISwRayWb2GFaGH8GnL3A8Zvqaz94
jBojz4mB3XLTdcFvwCAYPBmRnth+rW2Ueal3dlBVGiuTX5cce5h6xNJHzQqhsynKXhdr5l6gIDUk
rDhZPEVBdl5V/inFMbaZVk9H8TxX0oI1jTMHCe87NWOZc7ocHUyGs4CPPFOBc6+MsA5qC9g+0uE+
mntHJowgpQcYmzc8WOLUO5rIjwOFdV8L1W5ucGxgj3WSIvWaL9aX5LZ5omvwhGJTHs4rs4ry2klz
oKJAAOLNae/5JOEcoh1N/1Up3yJSfZcT/RKhdf4GUfmJmq02LxNLFMKQ+NyLzyiIMG0mdtqNmksi
RoZXihxFmt9mOqBLXsBG0BvAfQfku5SUuiT7lCAQPbLMN5jeP6Hyon51wLLMTBKlB70hP+HSD5rW
76/D6ROSuyIVIMfvdkCbmSMigeHIpd/lHgOxNNdAEQROJCf8/NVUPP6GGPxbiAoNs86rC6ccD87T
M1gmGXVxvTPwxVn+bn0R/Kr1pexXy+PcXuvcUHN9OlAroevHqX5zeRPSGOsIpoPRvvkRH8aORBh8
yjrXjEPVugTkqOHzhWqUkvkG4/HzElgu9SDMUeorEgZjZdLRuNkURK+X888jdeZg2CGYaFxHhdQz
4whoh17SVT6rAuPzvdnlzihJ3d8CbMPu5uRl8yg524NnHo9Gxfh0c/AGRMG0uvG7rY7mlnraXgsm
t8DxvI+fLjCX54XmRSFcABEbsXciXBt3obW05QW7TFFBHyvqEO0NxhyxvOB59vP6M2PDQdsMobtM
D5YWu9D3IqKAq8/Tz2B0pWSGXYKuqdX4khgooj3hHfCmAtIrjV/0p44rM3fmAfCVnoVWNNUumubh
w1X2nkvtMiXyS9FUNXJAL2CbsqaOCqMtvOGe/SKUWnh386hvVLosXBSN9a+cOMiZqeIVnsMVAAlY
QIQYg22HCv5xT8AOkUsb11D7ZsHTdpydda6gI7hAepqcIxtQZ5y+GEfMNEEvPRlSbsd3ASH6r2nJ
QppRz+m64RO1squ18AOisXZUH0JyL9edelizJLAGB1voG9Mxp/c9aolmiLuI5nxyTO8sSsh2Gke5
JiWAE8IoHruWQiou43h/llQpvhFO22jkmvKOziIc5F6sIsCFiEDPDXEm+lYZDom/fVhnQcLGz/7A
f2EpCmMK+S6FSYzHKJf2wF6D9tLJC02UKb9LBq5kLdTXc8dxjLRA4I4hi/mVedLWUVVhBfn9213y
UYM2hx864v71WC3FcUc5jLtssYC3g2xobXO7um5Frb5nwhgXIsjJCedhBhgU5B1dLLJ3beU0y+f9
Voyy625u2RC+eiH3ukLOWrnB88cZamMgOVXyCzw0h0SOT/YGL6rqh9QQbHN4LmIBuDuOt8dSGQZj
8vmvgkafFGxEKyNPUK9bsEToKbnadPVsV2mUk3YcMH2sYsZYi2KYWNMPKHkBsfEUho+vW6f5PvQF
KMVtZIU51dTCRdWTx26c8hVefdeAPrmciKxgB8ztvxOomBwdHhKWJxMYlcj32eTXUIRh8NMttEzH
HCnm05znFiWKfQ00lqryv08UjEhK8lggndOGVHBpVss3/LLm/2ZyPetzpK4CvlwvgsGS55cGZr4X
pHyeuPLeNBNaM9IOQNW4uvjcowQbHoAcmSs99iNPudo0YR9aowJr9AkzmRXWM2EGKAG6EK8gk5rR
XkI3wzKURosfBE8ijIG0OCa9DHMUFU59KmbHdyrJavzZEsXDX05qVcGhBCrZz7xxscno4kRI35td
Fqy4rwCa0Mi2OP5jJNLbsQbodWL8rVWO2MZeIFMcb/XxuQ8pt3wzwQ5gOh/4YYJ3vtjYbK6N5ZU7
TPomW0Hs5kRtl1RQAXhBhUAP134MiQwlgBP6zb5K1UhzMyw2zqv61+nvk56qPolqFMttV0Q2mGu6
mgJAptjw75VWUF0FuRHvOvFFEY7KwyFCAjtwgF+lgg0F7g9709uSLeySP8Z7OGhXV+plgtF8jol0
WZZ+mgAgn76D0pdyJGwXeXvlcO/ufEZJ/g8GQfSwgOBNIZdKfe+tBn/ulNyqrR1/oV4osuh95XTE
m57oChLbew6vjSnEXP6ounU/ZCbH6b+XTnTLRqCQxxZDy9btIYk+goRMggjyUCiP9TlpUXG9I4nA
2jgRwF8x+qkf/BhA6mJZ9czo8EuWcVe9Dt3dKtDDIECDk9Q9SK5q3VV0b/a+rJ0NVkh4WIKh1htY
/4xesU5HtPLvJYHCiVB+rWFWUtNQs6mLQ3fNZUDdL6JJgVktNB8o1AA1QSXI6vUdqsyuT7jxl5it
vnnjZX47uSn58vhEqzYg2Lp9MV/DWLT0Ipma9ypkFzy1jixRNyTBakte45Tc5Hb8wwsc0AinLFDQ
cIRqJy167Rtpq+mfyHaREkGeO71ybFHNln95RzNsh5zehDdW8oetkqCo2+gRBZEa2Pxhm35spS1p
MsRPzmH8YGyOP7jhTEF0oVMnW8rcVjQwbBxpYKeQo8XVcYnUaGYg2CkE5ZyGyh4fPNUuGYYQ/ha8
J5h2hdOO9FzvQ7VyikZ7PfkpokH4/GKfooyMkRPYKY1dQrCN0ppnuyjFclF2dlTkNbzTRYfJpF4I
g3P+CofNF7kUyqz7IdtYzrXoVPxupe8LPKXtQlMRK42DVJWHgZwILDmUyXCHdfp/OnpPnWyy9ILj
/UVwnDugUlBnwHS9fwIlR1qXmxbE8zpO1mDqBdq5sI+7LM7wnCyRAJSF20Du6T3EGsNrq2ADMxZJ
flQqArkgiH4sudt4kQJOUuQiSOAPwa0mtAG1L0+WQzplPFDc8jZ+199iBybyzFGBhCGkHG/wLz+6
9xypg9gAzAp87iA8HX3Yq5NfxJGrM2gmrLsUt8d10ZJbO137bSb9L9MG2hFBDyo2lR2F9/xUKULd
THPWqwoA5iTjCq9Z9n/BTNug6P/KRkujiSIZE++OIg8rIinY6/XjIU1yt/ccXsNjV6u5sCDSHo5s
7osoiND6Cx9Xh0/4uEBga0v0JwHXDbcuMspQZ107EJG2gexudn7T80e69CMW7O3OSvaig8hHKwyL
IqHucYPh5iZc1C5Ny50dtGRAPsftSXYxUHblH/gUTOwqhk7f0/tHk0MeXiUqAtB9LvTKrCfxer4b
B+0geO9Z6O/xsJt3ybvfcgJTzLwJLvhhpTUuw3WvHznXK6QGTPEkyfmCpK+wr8upRtJS0/Gjf/kD
CmVQsfjnaRpON6JaqXJdqOEf+1blzbqlgIrVpxAahFUbheSrcmj9R+YN4jUg0PkN8goQlEND8Z8H
nDN9NuXGQO7+dz/IDWIenOFF0EbVgpfdPu5vsshyytiK7ymsfXG/dkSFTz0rs0B4f1XTvBA3VQVE
VtBsn88hV7fkMkfJKi4V1w8V97Qss5zBKopT7Mx3al3Mjii4yU7IXATQdXx+UPylK8qn3/mcP1gr
Yn/bGTmdZhzYK8LGg1U8SBjxIke42/BGIB/NVLFuES+0pyNjHGpeoGrPRu5MSwGRfqdZzSEgfWhW
2QfA2nlYmPVHV3tVpy0u08GzbZ/aX9x/0KOFp9wVZtkpEJ8E51JosoHLPnGZ9gsWouJK45ckgO7o
+NvCfzKxbKBaaHQCrn8ssgvMZxNusXlWtdR5z7gWujm73nbymM6csnsyUjojqAPOWXxozTZ87UEG
jiGWD0qRQgSN3Ex3TYAs/3nMKyFM5D2OscrsM6BtzGUlfFiPacXeRIvPW71ieqW+1sOa4hLqKTd8
TGCNjoZ90qJkvKcxLaHqxN+EN8JkKkxqf0OhVyrehY0PSifTHk6cB+Ex25YNDZXM0Q0DeBKGAYkh
bwRV7Us9IkDDHQQMoSjhidR6dci4mUfLjBDWCwE5sxB1yhUbSMImFoec67faw0LGv/av75Ko+/Cs
27U5gywYlUYsc0T0JzhV3E3eWmpPWGMJ8CCtszkNTN+1Do6ekwkRF/w8tPYzN2GiySM3JuAVtXl4
LUPe8kFgrrn5+sPcEPQeI+QAIYoijKgFvyliXAxzV3VHdyKTbWV/fDz7WMUJNVnPmIqWMweuDKzw
uGn6feTzILMQc+cXf/Qh/8kA84JXA/WkvzMaE4P8pCKi/TvoqxIn3Yqa8XZ47AFSZyqO8gHsXCVj
5QnFWaidFDUoWDv+3wxwkcnQgkRdT0+hs6RAoxiEwEhnMcTpC157qZQ7T9yBqvIXaeiCWIRHoiv0
VRbgQLUSFQZxMJy8wsu7lYXqsQk30XsdP8YDAfK3Hcnz98HxqFmwghofThwOkdOnGtX4E3D9rDF5
OQDmhrl1AvJYTbo0LeDZi2VGyD1Ft1SOSukDgCibM2ZhR/gByU0OOv5ph6XmnPrf165RN1pqiUqh
1gGdWA70FGZh9kuRW2nXSIrLbEA5Yf+tZrfKPJ+K5+cgQol09phkLIJUGLbhd9e9Pwnu9S8jZA6X
VF0TbEKwbrSzoS6NHzLsORKLwm/AixBPwZAet0gs/LxDCkQRxCCfTvs/JAAwisJrvkfzyK6mD3WT
NGzabobqkeNRWThbWL5bYd+b9BjaKznNVvUi7Vv8k24SAc0NPapZzvv7nc73byrkJs5seek4g+7c
JA/wQyx/NBtzyOakKdbveQsaBGMu1pbclMLNs7hArY02AG40WfvIV28t4R1TSEHunogKJbYN18yv
nIHi5mkkOhgckwfXWot8Gpt4BjU7Ar+7yNIHesmBL9LE9zUNwGabE8+WuDvVv0MX/s3MtiVM2Ces
PQX8q1cQ5i9+iWHEcendyOhabZ2OYkJRmeWt9JMc1FfAyHjUob0IysZyaOpXx+7bdGWHCLWv6q1p
kslEzrgMEB6gvLQwRKc1PmBDA6zlk5sHF6dN2x7g0ajzHxyQsGjDvUpbrWBHbxbOdkUWnr08cSJc
rhMfvkmPhtSWMMc+asB9k8CrqSFJJzTf8Fi0DaX9RCl3w/XkqNQ2pHF8iG0K2KDUpabNJURQLrDH
zr3+RpVW7Nf0yBlcCPORGML4g2TXuEB0jSiUz5H76FujOh/cN7WKKKQja7L+JAo2esBHRpDD4DOt
hWDsuAmcwpdcM+8d1WsNNFJeSjHe4XIidfLkrYxKpkJl00yaByw+HA4pL4FthYZma8XbhpCX0swP
Paua7Cs9e1vhooAhVlmpzVd587134ZLIpC9fv8LltozFaOyRbgTStPE+P3cZGJr18NsV+0dS/MjW
hI7kydPJZC1LNst59M8oGyeiPTiUgtO/EDy/p3KVwYF5NwjaWnazplg1KBviRbgKHsFahGW6Zyez
EOpWN4jgkQTaaqcrdT0/of4GiUYQ1YtG8of8UbJQcaOK7+Zox17W4C+rZA8Q12++AAAIAzRyO7bO
2F5fY4O6biEYFh3CWhbDc01b/CCTEARsMcuB3oEnhD4mOnjSrrykIFS8QuUeVdMBee6gvGIwivLq
O0G5LM4j8XkJ0YnKV8fxlnUaEsjDp3rf+3DfMH2JubJVlgqs/n7N9quErmy6B5mgLDqnf9NlQI6n
wEc0TBYUEapCUh07hhRLKKt408LbOxddYMMO995L/gbjwBaUX50Q75lP0MpcdRva/wd1g6BWYkAv
8ccKeZ/l/xbG0FIgo1yotBktdMpYHwAVYL4hV71w8zXmWbYjjiIxFXHEXj+e+heBHOcwAMKd7TlB
1QMSCSYR+EGmIVJlfV4LGH+hnxWV7WFWsJol1lKQIIIrYXhR909NapKT4mCD+5FHhOCRPR9lnIyF
B68k61yNlQk1RvQKNBlq7nkz//Yy+TYO3/Ihal9L83VNGbxpU4UqgrD74Ox9QhcymyPM/crXhDri
OrBmzbY+bTjGoaQfWTBQsjlHIHv1tb7HHRibgFS2JNxUCgssQlmAl7pTFIX/uPH1eZljEa4ofTWU
gdnFH64Xlw4gLJsEcxylUQCmHxLjomj0tdJkOLbTVURfznQFhmAM/FUcor1RhtqJ3gwccI4h75ve
FsmVKLDU+TRda+Rl8KFZ+5X09q54CmRf3JMbOBjFqWzjitlW784H2vHnHEmCIf/51C8SLehXxTkM
nSY1eGOsBZJxRAJy69dutMZXTiFZtobCLxMu6X1te176xpsNOYCwJLuPp2NKYbRXLL9Rv1ZHnlzl
q11+aYdLdBhrkqgsW159x4BEmG9lyL+2UMUMoACttEj13fYK2SYrwMXYyeSV15aekOZvMYxOW+KP
pGYAUuqDXm1Jv2UmcS1zxQvm/zcod4RPnjWSB2guDz85oVCEGnjNADnNZyqXrIXtKkowkWvNczUF
EplG/8fd9ARBSXLABk289yAlQLAvEYh4OmNi89p4Wq/RBckZv/IkIfa5AAnVmM2baIpp7Fv2Xpdf
1kJKo+cBD/vhwFnsx75xN/4VJ4aWhLQk9+B/oWOOFRPOVVmeTHMiH6yz4h6LVdD741BWMbuIiCj1
1VpH+duUtjyx1W4iwNyUrLDmrCfQRxLMC/le+h4xWQzw2olIg6bQvNl2p5GpIxotyBudPYeNnm3C
1zxygEoiJXyoMQGaP0R9OpY0ntrWljVs/mIaCwFdDVAcRxGQlQWpVEGteRFX1ecMG+FjC1EyQUgU
ERLWvNn3Nfa1PhjFU/lnmWzPz7onvRnpVlbDanqVTaQKiNwuLgMA8RJMCUXrmgp2nliWwTYoBPwJ
s+vKIDAuZsqv1H8B8O6mdsq9z6PsTc2Xhxx8PD/osUdvVIUB3EnSSVznIfTEK6RRw9S5uMccqkPS
v3uNqzXntj+UtBQNUog5XQXF8FP0ViEt1UXBfbdumGlk/+mxRExgYla8zsoduSNYqS64j3EpG0dR
MMEJEZvF9nfTGUKMEUHb8yziYfYutHcKYZWDBw6PaR6jDE0AHasH6SYZK6rkBAoPReCkP4SWhy9e
JxNTMcwOWZPmwiEJMmo0aPZ4KpfcsqWRh2cQ6jCvlV2H2ckF2SDnJrAawjDmAIuGmoTth1D9em8t
Vn+5o7EjjnVxEFaQk+iawldRAO9+ceKazoX93brLXNEjPMnLVTucU2oHhMy1OfGBu4eixvnblrj9
j1vfUCEC5qD+XQg58cS++DTZANJrNxKb1pax/nmpssx+smkv9Hdmp+i1sYt1L+vIji3myVRztzQx
TwQufXUcNlcL3VVyWxn3PheS2sQHe5CCILKhRUoceGvUGVi3cL5cE6oUfTlQ6LGjsbLHMFLbwHKY
qfVZE2iRSfmSJ2vKW/A4Byoo8ej3mbUim1yblJ85a67jiz5WMsYA4trrZONgea32+Hk+1MDb6CAz
GXBu3rD/fqyGbP/Jqae9eVfFHa7+8PerVusds9L1x/bDYnnvy0c7s5ivHLCshdGpDuExnfS2PX00
cZNmgg6yF60AMS2Ba8gicIsW9GUO81FuI3scskK8sJnAjB9bGo0WOzkYlGjWS14cYdog+nux6IMX
ZalKTBG8dm7l6cQIjELBXzb0CNCDhA42y63wVD95mBB3hnSwz48LLg5qRee/siGz852o3t99inVR
pczINrjJuQh56B4ympobBwSeUodPtOotM4Mo3V+08EDJ/z4ES4/d8nsi+4jqLqoKIeTSz4P+sclY
jQr2VbATZg4wn9xW7t3Y6Q6RyZ5Jq1BCFwyc+FcK0zVsqvD7HcoX2qkVCJIrZ4yyIG6q6X8WKh/4
bgjZZrAwBAFVGUQTLGbUW6NgSRkP09/YKu1U1VOheboPKqPk5kDkasD+ZpSloRCIT60x8PD/OxVr
4RULjiMSOGhhXgRm4xiEYj9IcvtU/yYs2ggIXy1wmYSjEXMZnx/W6lfKIwXAQSeiio/5jpDdVxfh
nci9duysnGmKE6/073+/Ce3DzZLKzcaL0GBJ1GX+ukPFe4c9S1fevt7Qf+8+cncW7HkAgzj9fQ5r
9Wz273mc1ZeqMXZorFtg+SkMzz7dgGPjn4yiJLGWX1S8NXleYwcZBPCUhaqS+wxfoOFltoCcb023
9MfXjw1Gr21PHemBCDwIebXNH2HYIzJ4Ka0zD9FSwhO6AB2FyelDGH7mvQcQ1IUV/pTa/em/wpMr
BLPN7QVmpBkUeC/rhJ/chMXgpKu3zkJMOAisrhz+AX161rD32nQ/Yym4/yQ+xjrFyyPkdBwYO6ji
4dH9SoVAiSjIHDmufzThFmhdK+Ijoac/b6O84YkgImeotmOJOQ92acYdIdfWf9G/FKqueYziyvqA
mk54TysQz9PKpV/NZ7vcY7krKKd/eStut6/FxlpohN2ip31bC/Pxd4HQgGZfqbSm5eRbwifjaxNU
pDkG6kLIksmm6bGlS7VA1mQmPbgeipUfKP9sM2YkjV8Xz2Mw/u1pfzYu3OT80mLD3F7c1LxbQ7Z2
2lt90Azs9p/5WaFREStZZlkEtt6KlUSHfU4Sr+/dcOTT9wnFuJSse2pX/HaHq0dHiZiqVqSsQL4f
wj3UooifNR1NGX8K7X1OY/wsJTiwAc4oqqB3AeaeqgTbIijn0O+A3vMw5fxC1zSXekKMt/BfgNcx
3U8TLGm2rM6Gc3CBlNqJEJVDWxrU+ghZqLCKhHKggCyfIC/kNqtjOW8+5eaZa5rS4lUwpcwfFGFH
pO773DXaXRMvgrNOKkb4qekO9T2lRdPNOoSavCO4aRM5f1qFJdTJjWyHgc03sKgEtAFe8fu1mIym
hbFT8cBq/rrrUYqLS12YwovJa7FZjFBDA6Rbc5L25X6ucQj1kWjsDca50PsyMOLPOmGAJiO0yFwa
k1CA1yzYrtH+KpubjcG89vtH2TxwhPys5nP0MI5LWlbdv2BpuLexo7NVLKY0jeQ9Er/2FnieBMrH
5aEsyWq72ROUwDfGyz02YUwsy6Q2ZKpTPmL2M0adTEyiAy0b1HFnrav24iPH4eOk4n2M8dtfBQV4
lB3EjtFAn1lVsqU0hPa4iCikoAzd1MDS7NgsvsAfJaJGRPLKl4txutYNIZaBt1OublApAlrZqE5Z
rLmIAtsuxyBQwHp5MUdmA0G+xPxhp/T34pmeHuwDx7Is66CN8s+5UdsDIWjyOjqcdUHtLhRH1frc
YvupmMWt7BKpVjqgHl7UrqOzXJZ4xfzuY62h/zt+nZsA3yPhqo286bKsmKyUadUb31H3Fam5XX7V
hBpdKhAqqPfqGXchIuhp36hCf4Rzm2ofveCS1TNRe0jQnkcSzYri43zALQ61Xtxyogjr6EoEKSo2
LgcASPkw6Rr1LYcpmezg+VOd+/zl9R5zAO6bmogVpQkhBLMBPWgq+gg8JyzIkVIKKicKavwCTBw+
GOjAPcnZjGqRzCVCfLfJwhHzDySxingNm0ptpY/I2z5YGMNw7L0ad9j88vv7+nRMReWZaLxzr4fY
UCWCVbwSaDNjUtkBFdyOM1Ji44RblevuEyX8z+DVf3l53E3xCJ9sZySg58wV6pAjb0LROb80EZSE
P9iHBe+pN1lucK6ro1PheMfD/24sChfWmprBTruwvVisdVy2pm6wCYaj0rJC+M/eYMu9cig2OOPP
XHopbBAHv/Q7wALXiX3qELp2ZB25Svw1qrhpahpU6keT2U2SVf3kvjYAFd7AB4HbkbcrYm8BckqG
wRBCIsPja09D2AFlCvXwQcFbvVJnYYR9D0EqCPWBz4NNKXA1wEnExMqtRvwK/cx/DACAjfrQKn74
ra6ovGCL6ikDb//cAV3jdGDeGX3O8QTT1FfMF7qfvUoWak8wlWLFQhMyFVnppRWsEuJgY3sOMbnv
47G7eHdLEgiHJVj6bGM5Az2fcG+5V6Ek2GnybCKmaI9xY3IzEzzOAvB3skAlq9NhrfZhUqFsGz5v
mqIjSOMYp4S+akTBK+lxKDEGFJjtigmE0Ne4AfMVj3OYmoBNRESRTwkcjoPWlP9Hpmna3EJuQZeZ
hZG4CClb2SIvDMdCG71W6aEee4HPUH204k2c1HUh+VFs5RADVGor47I807/Suj5fk3xKuaQBa/H/
fzxiq8pRziq60yEgq+wFSe11pEhZAc1PygMNWOKVMcTXTTcSdlIeN6HTA/a+rfyzjI/t4ZjENH+I
ESVc0R6dCF4qxyg/50nSQHKzzPiPd1OA5mqwq5ql3C+fw6SBNsZQyneyTcEhx7OtBxUXjReeC7G6
1QbT9rToBdYkGGtw1+W8Vq9KdZ/Q7nuoWteHkTH1+aLouKVgD75+NOayYu7nylGJ8l3/aNaDTiI1
FYWmGYxHy6TVRjFqo1XxbP2M/ww6P+C+E1DxHBK6dvb6zqz7qOt0lMTfvet6igOi71l/zVQnPmFr
udrvlwhudPfJd5r2yzdJcJk1x3xBbXnFDUg6Ussmk8O29vyBytclyQVM4z9Cnq6FLRu1Gy6uO92b
fITgBVKotlZlvkm7E5tWb/S44wCdXWJcY9EIFSS1ZL36/JwQrpJljPJZjH+ICVdDQHxwWsE9RfsO
wgwhRpeAaJOFYtOLo7WnKONJSpw22tlJSpnJyhYH/+NM1c1vgCMafVbLHWk0QvV5Ve/d0kXOWJMN
7+ytuXmFJX5WwxLFgzHIxyvAL3KtQafvj+igQTadYFm4KSk7OD05kuXDaDkRjO9mXWC2uAqCEpZ2
vSszl9ksD8ZjFALr7lGNGpI1JnPbN+fNn4kC8CPT9ANq13zHGnSPlc+Hlzw6yYGTSLPPsYZnWrQN
OwqWXrhxRF3VRiAoUgZ6MMiaoUNv8MPhloPP9jbHAXps00FoDKZHVPYo0KoDdJq27qqGlEaOx5LA
90PRTfDgWdTb2Fq6V6Q9ssrREmLUtaxOEtTqs8NQj95zfEYobO6WwdKpSp82RBoKSPOBAeyxna6Z
dvaREMammugclR8p3NzN2Xddc2IxaUQevd54kFSuAkeJm8xgE1JGsyMtKvUqj0Peyeaypr0u2Q+i
gaQidYZog70iNogaAGGTnGgw7OFC75fdlmmBZYNgHtGP/wHcARkSYPfZltz2TTpJnqvgKT/NdYJw
JY+S4Vpb0bNOM8M8P7y9Cf6YBUFDoGndnx7ERDqg9ZnGrwTcIEymSJR6alvT3RPPw29OQ0x7mm22
yyZU2sH37DFRkFircPvCoB9NcRL1FrhHClEtRayI/D5+JnBJBZKRsKaAr2twY6EadeyNuMmM19rh
5dVPIRp0XI+mGPttFra06WAISsMo/TMd69VHpFwlICRxSwwy7kaiBH1FPUFZu908tO7Dr41iyt3O
UgDbDyLorolGt6tTYVqjxv4gTDbg0+yPQbBN/v6HsKc6Wga1CXqlTOwh18S80FXrqNdr+quB4DgF
cqsdfJdRgOsZCrUGL7t/+e6J82s73WRgHs4aMPamM+Zjlikhy2axCu/cwww6pBwU5dALSEoJy99j
Qes8L6ScrjTEFyY+D5Gv4NTNHQNhDT7x/deLLZ7NIV5RYyxtsHleM68y3UaDLmuh9rlWwm/v5QZI
exCGC9c8BNEs0od43YILB4eVGMR7hUlsua7egP5pJB2teJHP0ujSEAKldBTjcKK7bT4AOZ9QfN2o
kqxjXM6qJxdadMMCQ52NXMKkTQQMoZ6hHM987xlqvD5YSUof//7waIPTbzUj5xMiMi0jMHOZp9rs
eQpZn0bo0nPM14ZzsheheU87qW+tLtYqcf/I/OQ24JG/u2r8ZE5h8XTYCZa2b9VdIVwvAAJUsnQa
GpUz6TJe/S1No4myIHPwfsC/G4kxJ1LIPIqVb9vMJnt+RBeJgcYnRHBTnq/Z9mRzLzZvwr/fMPeb
MXzoAH2IKTDU9CwScRnbP4jJegIrZgbQ3Xx1k46h1UVI6NOTxRmET8Jq66+ALf5l/QvwesOvlUSK
3uLgXG82n1JbfWhREWYY58WiiGUYhPHQoIqgyXBo1ODFM61a+KyHWW/m7VCyPG0nCogUYVcXs4jT
kkOxF58oi9q67tGOLgzE20C1551T72Z+BPLHkZT8/ENV1gY+5+uIoic+EBtnfJ5BlshfH8QWJrTQ
jSwST6ikwLXOKKsJ9JPxHTJ0X1lTxvV78zkKQOgncIW+59hyYFO814sfhc1LXy2mKbiBefuV0Fv5
8ZTayGNW0qCiP46NStdT6QkepjkbBDYVVzzPfBwRFf22sa1Qsl79G1rrTkEFch6TMMrNR4kCT6Pd
066spAXNDt51FRwmzbCiq1/KRuXui7WGSF6uxRBbHE5Ovu2VGs88u4DN6pgf8fll0fAcxL7iFKt/
rMO97iBOOgRmUrdMUqO5KgWfkdQ24DV1/ScqZgUR+7q/otubWHTuSLcNwkHD6X8SSQfejKRaNg/D
ZdF2cP3EIpsAcukVJp1buf76MAz9BftD8B9Xw7Pfh0Hy/3wNvPYZC7+xhVeiyEICoqPwKnhf5LkZ
q6kig26bpScnuCb4+bnsqwLGbCBoTd5TGaB5lENbk2urhpotPhvpdnQ36fyybpNXGyGXBpmwGcuA
l8bPldS7L1uFQT5ogXPIEysWSaHLOU5sjj+I3WrculI1UKJ90+dotiNM8EpGfcKE//kJVdfnwvGt
CGy/cmLJlXshxjSDwY6KXO8hJpn/8QwfJQfXRV3EfcVZklBD5jAudHCzuWx4S60TUryvkMGK3dlK
vIK0nutMIyloHEHgRdoIayfl78u5/upN06nuoFI9I/3aVBR6Ob0gnDuM00zpog7yGy2fF59KOAV0
zCmm57gWpO+a1MwhBnA25eyd8d5wllMXU48xVJ+StRHAWaeaGyMHCcxpM6rwrnQKjHaQOSUpsTG/
jfjRGsOnoo54gTW3Ucwh90baaT32WA8ghTBH5DvWgKN4S99qywEyL4JCmz/RLExhzN9SiwnzWFKS
3/LzqiHRPcC+BWtXlG2F7QV/N0BE9hbXMofvKqcYV4IXG9Munl+ZP5g2UQ4NzcobFyyrPkykmebL
R3fYncCU1OGzQzg2CznXpVt8J7gEq/4QyPdXY/6KoonompG1XF94PN59FHrYcwlJ0FjdJFllGUJr
gMiYBj6BRNnvDYd1LrJ/aAsj+wCidP54UKL5iXsQokgZQtw0dqcQ0mFVdm4CaeQ4/3HGJruAMszj
KBOjvPlo7yR59Eg9BgZ1MtN7AVMlq5w4mpyYDlckjq+01gshhwGGPBeAmIGGtx+zkdQIEc7qJrlA
+OARGw8r+z/H32vNRG5lY5UXZ3UEiDbYjDjrMP3RG2jqHymxRmQfSyEkatWbg0Ap7x2TbpyQZnzx
Ka6/Wd6uW/klcAv8y47riYaEJTedpl2TbhnXUUKKb8osBhmjOQoJzNlRCIxJDzbqyc4yElN4MSxZ
uhOVwwD0pOxiVNvozYiMgPpdCJjVkx1g+l4YvdRUjploxU7GwxYWyJAIyLsPCXpfGf6yX9vs+2sb
CW6KWcuefBa6n0zfoL/QXY815cnejnTOTaguONgOP3G54WJzB1MCS9YoPneB336tkZP7Q0+LuQ53
AZt7Lps1/nexNGLWRGFjlK/K/r5JZtJAAS5yjooalijzM+58Wq+8/6rsUtt1tEqphTTnSBryfVkN
2gb756RnuJpKcL+EkO0doUYtoVDzO8CWXKGpJnJaRDHe7BQGjG6TFgOPUG8t3beHiPfDWNWhr1V9
N0Yzyn0V1dneyG+OmqkHrwWYRDDtC2pOqympDJKtxCMLf3PNIhTgnVtCjr8HY4GBxxVPW0DonlOc
dXZj+av8x2CsGDWJ5hzZFscoFJelPDiz+JLlHuwuXWFH2RZaBd/JKfZRrQl3Tv1Zsm8g+Yu9hpt6
wQksy+k18+j3mqVzQ7geJ1bEbAWi7edQa8wQETTx9tjRwH/K8aeCLai6ft60QwXnSeiWtL5sZwal
En5Q9BdYjM+Mzh6gGqfz3dlwDrNJm4efRM3qSh3COg5LpniwBbel4sKD7JXRYntJKqOo2gprQtRt
qsCOzZwDx+XBTu8PSqErepYwD/vo4iE5PsHpX1v3rG3HWoh9IjTLQ1c4KVh5Unmb4AoGF86SngIi
T31FFXrIQxrQbHiLi9b9VPjoj0m/sg6WIPie3iqJx4X1mkGhQ7gMf+VdUygeyB5yXIk1OX6mFGTz
frV71kOR6PE+6hY2nYcTNUkyZib1MvYXi3QEJikl9e2xJTytCAEjZgtBfGDWV1Fwzk7cPeCSDKCh
mDCmz8LKt8n6mJt5F1p6ieJf27elHF1wNd59bUZhdcXWra8Xa4be+w6041567qk00G1VftO6pRHj
xTMStU28J1/rqoznMFbwwU1b1d5HLCmHx/oG+cBQ9zoyhZl0G/ijviXlq9syRU6lENMtByP+24G2
e74WwASv0UtH3QjCGXMDPSY6jhfQwLJeCOvwCGo1nR+z9llApoWOF9W1dgZkXedgkPZ/vHayze8/
YfPiwZ/omeU9wdFc24bKh8C8On+WKLkT7qL1QdlnPkzP/q6wlcCV3mo3cMwlHFFuHdmIGseVtd39
Q9c5QC9uQ8eVEzI54EwpdaDMfp7q+VyyJSP8pr//h0VnD5s7RdvUdmzJykJwLwgaINXKG1ePQgx9
Fu94JHIAaRCLbB8MrOtX4Sm8lFoAuS7jbthWphn+Y5XLeJ6ltl1jJmDX5yk1+OTzXZ1/WpYxzNqo
Oi0dGssAy9i6tJD0xJkPeZaO6UpkxkbhrFJzjaUx7XJSIMyieSUNt94BC12tgvDrwxT2pw246EgD
fAShtf2CTXALTrK+Z4JTzNP8EG7PCPUk60sVYV/rrZjQr83v570CMvDUbowuAPN82u6z5IM/mYGL
bNMXbsbPT1mK4RP1mOCwVrDLClxbdr39t2vejx9ZsAooCrSDr2ffZo39ha8Qc8N9UaI9COimKJve
9vsOrktWsy1GSPPUqdzHDhogb4d9X0b/VABX4/rJ1DX02R+bzl2T8rKsg5xja95NKhBm+bMhDgE5
n71EzFjMdvuvOdIx3sq9BsinjatqJ63sunwoVhPi4c+Y57a2QmPPV+QcHsnSztMtHMGPB2x4g4B4
9LYI9krr5j/bo3B5EiWFvIehxb2IpT0udt00x96njjvlbw2BPlmkv9uSmwgyqC0PuOWHD3D8u6Pk
97g/1lyTeowEvhRy0axditVyZewAiUyyd8ymutpg/Qr0MeUR4RHiQl4lGaL2iUENBRvw+Uw0x29W
fUzaB3JYwkATIUGOtONRo26s+jbixj53JseDu1EFK59VdexpjlXiiBVISPzACF4TXGKOg6p5kGdV
pzqTKVz7xaHAI/+FZWwVfPWJu1buySlAoUmzJFqoiGD+SuuNauHcbnOmhdS6vosRNI0nhU89d4bb
mk+HLcwwzo8MH7pMQvUMicacPjsKmKHi5WmGZc//ZUNmDia8EjEGWhz2h302IhdfcK/cuxcYt+b4
yY71wWtDkt2jqNMipc5Skl8frH3kTeyOUVsKjNPdzVgT2L3wG6eB4TxylY4chImcKKteA/Q4SzFD
j6AgW+QmBYhQGGI8ANk+1l2U+rfg+CZCe1N1fVUUKLfPoAdPa74HJ0mmiXI82E3BHdNQEGdj0jL1
KajfJMjw5kE0/YlJrYEL4SVVGuRc81Mog/+3BkUViA3yRuCgOuPQe05/ATSZEZSv1wloeIx/4K+p
w5xFU/96gDPnyb2IrYL33kTUg62QkGI/dzbDUOUEXZFBnUyiMKaerMTplJvQM47UpFmePiOWMp/v
mwbva8Th6Vdaewp6BMP4OAgsoHh7HVxlUP7mITUhZbSqayXkM9Tw9DLYS0rqVk9XWsykUVEjKDF2
qDNLqmwfg+f7mJdlSsmGbGA0ZqOz5qk7UK39eFKt8pQOuqQJ+DxA2VMnQ/FjvXxz0xFdB2n5nkrU
Bg3veUHCJLBymMOeDdArPwYnrftwbwGUQhWdkqqJD21FRJK4gOQt4xb6MmHQssGnXHAs6Ci8Sosl
j1krdMEfIisYdq7LOQHFwiTZRocEu3+Bka5WuUt0cWM0DhxDd1vTXkf1hiYam3A7cx2vnfajCflu
gArElDtVg8yk/G2WpeIIq2/K3guATaMXa+7GEo3JsxVlZjgv5hDXS1Ku8Dh9sP0taZeTzS49DJYh
gI8RtVrSIpgbfWSD+cP1+Il+LcEP6tm5J3j0o5EQMs0KQegAgrav+G+vGP8iKRafycmc6/VTRg2s
MgCypOP5vqE1bDpIGCHslaohxcSMVmoyOMx46DGcigE1C86g7h8+3c/Hi0NQ26Qx6u4a5Fbfd1eM
fluPA+7Sv5KghsJQlSmziWB5kIuJ95nT6R6ZLvF8e0+1ULHC64/l8WZRELMVzJkovqU/Ma3y3XQX
56sD6frNXTIjur7Wq3B6OU7X5H0+VjxvS17sjYgzjPlbY8JYDnm75LXeTQ10IZhcAaVqliT9fbng
91CthOWcRS6gVJNstWyhcYlkkmqKzn8mDbyWUAEAT8MX5CtMq9qbxZHHko3TwnjsEbh6/rcAwqM5
AtFtOFpoKgTTdJTkMI7Z9993ItTm4QdZlGdRa9wdKOYPMAf3JRQoBpuRNNGk6xSrPlcc/gxPpBc/
N6ApNow7kewdJ2ShVlecdqBDQ6Y0o6rr09dPwFmq9B+E6QTzw8yI3k+506ulSe4mGEPeZAK5R0Kr
pSC/+6jyke5G9ntwr3Hu5AShFunvrkhY7zUt1saA37iKbHEgsM+WOHiIpHZFR2tBRFRn7EHftx5t
r71MtyRI8MY10xNOBDGF6ges8qiMdOXbvaNMPMgeopGywkmWUsrFFPH/SmjHcROLksYjtg2xI2o/
pKz0FdMiu+mKxm9RJv6gcAnwbpaGtJkX0wNMfI8TBT66M9kkbUWKWeP0n9iBHIRSttrnao4Mt3yX
XSKiGUQfepX+bPohFe+wakeB7tVgsS6rm0WDcnSKNXKWzToUSmd+kIAKLUEXdhvPMBxAvJFbgtkD
D0nAvNBpKKoaiZ6oNwPdCSyv5HOsJ9zpzChaZBbpjRsbXDFdhq0PkuXYZtBxAORbiPSyXjfq7nzL
E5PcDKJYgyYOqhFPeYpKe695y/Ts5BIi4IE6ONKRHop5vHIBXE8fMf9O+vxeJyG6Hs92OQ0qOG0T
jJKhfAKYzekhKyRV1aN+Q32N9mcox/qj0PzYo/5eeLJD3G/6heHeBJ/2ZK6JXdmul+8d21sUbvhj
4Nidao9EwPbIIGr41j140GaX00r3Yq8OB85I3lENeGtREYgbCUaoAUjr67Py3VMxA3A0R4UFRUv+
XOekqGw7bJoMh02hDvlQUMy7vJcNOdc+QokgpE+Wo08cDBtyyssLPTGkqr4SnVwt6YeAeWuPKwtI
XfPe2Jleq2kM86wPPO1MIjAEkjerwyRPnvP4MnWncaHc4vUKNfz1UwezklB9jSUnuDOlHFpmcQFq
YOh1kSRh6yQjsMirCxvOYaZXyhDg3L+nTI90HyYIiolz22MVcibvQl8BEqFr8JEWE04xqkXDqz+A
KWr+8+AWYhfMnH8tPjFCxoPufZjZTVrdG8PXDTfWSCKKhZYh9ixbtG3Mb+QwJQLG/raiOY2Zlz/B
roS6lhaBAdqqDZl6eh2RsJzJoecUhQeNkMCzFBSdhg5tFluw20OY82yD4hB/V0bvulCdstaQfWVu
qQVS+xDgWqD72VNCQJA7gnydS5TVoO5lHOMHaNVv9cGKmVDFhhsFVkOEfflC17dJYTt3aC/gi1sG
HrbYXArHPBUHS97jgwgfzZPFYKgjih5uLabJcBgXjMP04DXKy6j54P3aueqPmux2NZF96F0gp5+0
91FaEjjmoxjPXCPrPKQM65MHbbKYvyeRcYrToFo3akbaYPwIbacvTWtnYxc4GUroopPpwXqBK6kM
l3hXsbp8BSWrKhsG1vjSvRZYE1yM7QnKEpXNeDbosVj2N/v7vETI8jye/PPDq2IJ6bqynbZHoxj+
N41pq+fbseHs0sK824YCBlHXzXWcxfe6RlCpWNOR2g48mBA6GVQiV746auL/YIB+iyibvsyovoul
zYLqzbmbFxg9gKIrZAlJef0FL4wgajxlJovFChhCcbdX2+0o5ypAzG0EMa899AkcZcW6rmGa4yAe
eaXiaQ7PAgxTe+wjgfh3HQaW+iw4PVR29zEjhTQ0broz0Ys2zZ20pgyEQnG4n/IlYiCpMWD6Ty7p
QaHkbqNd2zHXJ14N2upQK/Rji0G9/gmyBYh+ZDwispzsNRcNbXsroo7MVj5PhYHmat3HcmC4ccCV
i2ipglRwdF4kJSE1L6AnrgSnCbULHa3cEEqZK6o/jHcfvG0twymYDdm3ofPJ3Jb4z8SEuSucUMnX
Ekc+3LLGfN7CNPTPJFQr5kZVlSjc0IqK5GInLhfYKcexNmoz/BDp4+KmoHEHqTST/vYJw0hkVdMT
0xXb/EeP9N/6yAdqsrDm28SYhGSeLtt99oqv/Ffsaj8U7yq8Q45h8A5Mn01zyrZKCXPznciKOO3g
lMPQCX23bdVrCFx5PMLreyBf2KBTDnxwhB+JBWd8BkECO8nt9j1H1+vz8Y/47U3cnUNBoEZwyrOs
PT8t7oNpT7rPPyWUdJpAy6LNRJrRJZsVRshc10xNtf4Jai0sIokenDW29OK5u9CfSuT0wAJppMvJ
DwComZ7+vzqMTGMulBsZ1IKm4y6Wz8OCPO0KMPQpuDASFZeIbpEHfbrN4xAMPVI8nuz7aw0f2w07
Ai780kke99K43otYUBMuA1caGRNiVGLCftiyiax0gg5ufbtMu9DQlmVu38uZeJz9me/kFFKgBkBN
L2J1xTQEIpAPGq4/P7SVO61HDyCK85J3qWj6qtAIcmOsrIZbA33kSfNCynOlWhqbyGJePQwmbyAw
1XLEoUNUDpFQvz2YR515YXH3xrh/diK8irOQqO3N34+bmqCG4gq7f+b6qa+BDndYZRMcbDhF/vY9
Xg/ePjVQ7v5vmegW3TC8bDPOUCNmnZLCm7tJmKY2WHQz4f+cFxl904ji8KSV+LKlhSvidvwq4nMp
cJw6KWAO/gG1xGatSuWQFVTh7BZMNpA3RusnDbxAKa+VXtYjpRoATLO9x7+ZwvOpO8DojsBtXfHH
joVEqB18EJKCg0imcGIX7p1PCyFAG1zUp3SrYsRwtCzVHSuM1Rf81eIQhdVdZp17HLR2PzyVyKgN
rBn7RN6drnN/WVGKw78UZNPzKTePrYBhIW9XVgBCuZTiOoKSP+4Xtw/Ui/37u6YFMtoJjl4JkS6v
JEM/cTmrvdK2Ud/CfV8EHeIiRtmQVCdWw7/O1jWFaBPeMhGFdylAFf6zPBQdh+T9QYupJmiJ2l7Y
upnGdD15HcgKSoiT4JzcDbFa4KkhvlFQTUcef/cGc0GkFyYIpnrf9m0cQHXdhnWyP4eNdILrO8Eb
KeQljbMiLvu/2lMqe1pcM49CJ0w/HlzyM09u1SaEw9QByPP+BxtgkqrNz/w03hRSn6YrcX/Suy15
4qCht/HkvR6nab4syWi0lyVIG5bc1XRn3hyy+gIe/DzyjL2XrcnC9eOkFI0NcDwP6RdyV5QvGf3w
O33FIvAIpopEsfRjOIo9UN1rcKva6NvaUO42n+mhEmyojXs2ixRZQ2pRniIconVB0vojrt4u0SvY
ZxCxOoZTvmSi4/o4o15DqLFTmrHABPO4ejKl6s2piIHPhiwGxIWpUeWi5h4etwvwmHcP39Qb5fZK
CIi+tDv7v1kE1y6ZGYzMNpuaxdH4AgQcCtYen38BBwh6kvhGhsVwPP1mV+V31pNELUGvZPFWwu14
ecRJPP2K5SFcIRbwNLBoCTcPkGVxp+3R9HcJ+y71nCOtNLaN7a8MpZMCdbXCXIL6OG8Sy0aLROky
j59vUkmPsnsEZeDJZpVDvTqpP0eqN5hbuJld+oNUeSpf6pNJXf9HICGNoOTaE745cbwGxqmLblpy
KnYgi29PC3LLjjQ4FFJXU9PHwDpE4n/f6WBsqw6cAZYTDvkCdCgUV9+6Lx91se7Z5txyUnbO0cF0
aMy3t5G8w2zS7STFfeImqnJ7r/OdM6CIm/GN2PMuskOsKJPqDBePO/bgxcVRId9MyQUVM36Ekzkj
ni22lnRw25atJQfBirDTLIbpX3KjpM5gCsSbxCAqvResxgK1Ik1PyUsYI8KXVaMVckEDOKNEllTH
c0D1UUsfInmR2/B6MH46DbkucBoO7dPnXYQOQUIe61ZxMQxhJePnXO33sQ7mzG/ptdy2W86d0zzv
aVHfISNLzkk/T0eRpeoUPLz+doGIqsn2hwGwlEiU0p1FVRYWq6aN1vlMUMeVSLxlC2yKt/xKECIT
+2oC/hskQL46GFa6TOUbjL/QKVWhIFm2k4G0U8NUS2bTT4HjopujEpNF0PDjWAvBrCwWqPMMQHfi
CgBKkRpgYyTUR1vmtCN3jiF61uiW2LYNukcqIYLkq2WwdDJ8Nm+2/vjo7zcktyoOMwvE0xuexEJb
hyzA10TFvmBCadsxw9HKDDUlYC5GDFgnpJ/YCJ5L+aIgarWS4KgdwydbpvCRy1MGJGenYrNQR/bB
4K0xuoTzU2w8u2TV1yBLNt7q4IgjZwNDF2HqNMOSIwfhISAz4vaUbRP3leJSMkSqluHBaADCRXcM
6oiCEcund0NXIJH4vzdGnqU+Zam7vYIFL0I2O30TRT49LdjFNculP6PJD2NcT+RfGtK1+VLIH5kp
lmiw8M6+FROAGMJDb5a6tqudMAM8V7TkA95LDfAeaBRbfwPze3KFd9jhX8aI7g46lRnSoulUmvrW
i2OQIhuSWQYeJOU8MqQlWpymGypQMLEq7pVw8aEenMfDyHDJYazZ6+EEj4gb5ZaxDyub/R2SIOoe
DGWCkEU91tJT8emH4WIoboAVTkPTZs2jHSDiHgbx4XlbUfuNXduDIcHU4yht7Dj1ko0W6mBmRUro
i/w0AO27lqWTGJZSnSxHJMl9p2KYUQlyrVsh4SOvccAtx7SFHrDJp7gEIgKg2E+cY4iEMnqbY5xN
xT9kjSZIXTQ2s8EcqDRfTKHQD5X8Pw==
%%% protect end_protected
