
module lfsr_tb;

endmodule
