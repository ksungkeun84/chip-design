%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
SH3vnqV+2XAHk7nrFZRM3gP4uCcqXDfaZp0ZIPt/cGfd5+p0FeyNs2vmyE6Q2wZLiR6koRTemzWA
Q8lczcSoIZKa4uWmWbtd6f37WXHha149Cg8F4JfkgNPmZ7gQYkiM2a9TvJrN4s8M9rFOlBRSp+yi
eN+X5RhJW+yC6kBrXIqhdl1pFHpNrGfgoI9w9CSNlclIdyRNSiyyYxemNBxyvuwlxyfdnJl4Biox
rnXQe3qDSpE0aCV/2KsYdCWUqY1cDl65NOAv2wLeyxJ2wDg7tU48z0+R/m4RrbQ8BmK2AmnYMksi
GDFjOVTsfnYYpPgSj2Mme3o+mwP06srqdtUcbA==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
PoOzlekESpROZdVRX92fF46XtwnprYSC+3B1pkDIs4aDJdLDZnH0qZnbQUN+/gQFAAfh7ItrM1+m
0wwcAlf/ZZdbUpaWfmShQxliAk3z29/eELGzRs0WkiHt3F0U6eX8gvVLoWLZU+4r1qRHYf+2GmhJ
vyX6bVTsEad7wGNqvcOFi7scOh8KsJfIKdvwQfwBvVEoLJJYaDtRXLqPn39AjZK7sJvC1mFRqMKp
3cAzj1Lg40tuRBmrJ8z1hLBTiMrK/7vNyFiAxW2uV6f59VPuouTIB6f0aZ5UiRF2g+Lgb+tnqhCk
d3dHqgcduJbCqaYyp9brhjz9cb26BsnH8NDR4bQLWF9u8IQtrOgo+ZLmWeV6i69/JRYoROiOIxd0
vltKkRvceBqEdI7zXhj7TNN+u9WIKM0H1MhrRHH/VGkKJtMeZxL73SZ5vbM1lW5Zb9OqkBNSM8fj
yPxCTsO9yq+DPL70usuK+P3zSNZooHbHjXSdYZvl0KpYewvfM34H8nDg/OJN4329NF1PBSRHn/R3
FoQIsGrV8gIwxuMcep+XEtb847FQs/OTgmPtemP6SL6BeEFJBgKQLgZozMW4/f2K7PLWVU8Ziqoi
l2NfomKsaI9RGls8zUuHGfj6FtwZ+shvvYEdFKElF6YFohCiNhkhvE5wjmRrTI5FVzO+i/h9E7ii
S9vPGflVSeGY/VSKvWkD5TagowbKclAGHWAo7USACbhMQz02MzRKmQKpkeRughG397/eo1Sqqcez
kmdpoG7XZbMQYvXBQcjn65XBqVutzTg9k3eS4uCp9OCilb01Sq5nuEg1CCrkhWFyB0R3cxm2ChVc
0Urls/oK9GwtISUrivpIOnf6dHMBKdv+EXZ58oC38eQnd36zt39sv7OEllvV2UXZQKRTNS5rzugi
0uIZGFR+fJSuadqvil6jRmk+5lfkZ4oOkz5fpYsUtZbFIzCaSAEYh/gcdn5WeIf+/emxW+A7ccHi
U+1zCKBNFDB6JOlLe+TohbSI/oPPgNYPVAy3PXoFZMt3T9iZKjyA5hOtHdbj6ulQ07DjkWNvctaz
GQNN/81NhdYXuFb88XlEaUP1M+DMEi2/bfcYI23Qij1Juq03ePD8FekzWemQNgxWiyVCmPoczYAq
Y55ykoFtEDTQoiTDe3aRnXPD6EWV7XDbEMMlo264HT3WjppaPUTfkL22pO3bk7F4DsNg8zDMlmqW
Iayal5Or8RM4iSlMB6HRs/38XLftggl/5TdeOA4z7+unrwdpmUH3VaA0aZ1tO5gVSScfXLYN170O
ycrdgwNNjGFlrx5yG9Z3qgavbNBI3Rt1ZYdUUJn3VOnuZKjcW4jRlqwLISf9RMhHPSz4KDWSNi6u
vKlifjx5ug/RklJSXO41SoxpL35Fb9apwlxLzsS/hj7U743OwJV1OvlXgqMemm1hCIm11hcfsj3V
y2bA6elnjhoYZzSHRA0a4iNlFm2TyR2ojsVz8maxg3/TnYF4qpZB26o6Xa5V6pWF2ngyf2vDp/sx
2tM/8COmyLse4lk0mdG+0BxAzRsNe5K+KlpdJTj/hmPdsjT+LckETLN2mUYC+B9gaOiaeVY4qB2G
LbxdKa+7Xblg3ID/lt64ijYwqy+F/VFeWgAAHSSPJingw6f2+o9olvpEqgnV1BVhox1hN5Vb/NuB
yaicOYIA+DR5/yyDsx+N9AQ4ykDJlAJJa+9+mxdYxyejoQaj9EwXLTSzGPT9Tv+ejex7i/ADv5Sl
2mq91TXr2UsQwDhm9l1Iu/xqu29TWXQjDNQ1KQNEWjeUFEaUw0N5Q2uLvfRes/OPjf87U5ohYJ1V
/qbQH3hcPeZZgF0mHAI0mg0ypbiV/ZTS+8yOtFLy1Gz9yEaoqvXF1NPto6Is5WhqlL8h8E6WSkH4
rq+zkQy13YNTsCrqgj26zgQbGXU/nS0l8VC98xejTYmH6O1h3luQdI8b+GmXVfkMmPWQD0re00fw
bQ9XsXHLFI9TSpvxok8r1XkXerrE5Ev/Ih/kCQqSplC8DJs7yg2pA01L0kps1bwMXKeBtMSQl9W2
eD0FLVSBnDp0MhD8QREyXCckM2VjrGK4hx5R3j1K6/AtIpk/Q+pmw5AklmESYCIxNPDU2ztgQawc
fBbgBqtfi87/Ulxl6Sv114GmnQCUeVWkHjVUtmEOoBu7bFPlDWpeU/d2G8SOJn7v72BzOz90Yo/7
d1QgXf6cCR42fHXBWVFYeOQG3YZFMRQmwGKersTBVlEvYmjDi03ojPKDFkVCbhBkOGhq72fXeVhd
bpBvXnZV/VTVg4guJW5oS/V7u1heoGut/aqnoue9uJyfPGl0ttCEuavOQi6rXtY2Ep/8r2yKbgsm
p+0XgK7srzwi4PNk7zpcjymJXUjjl3xzyJ24sevIXvqXpqyS+yiv+Lb+taj+M3k9oEMlJ29swtTc
5GK6fYj/aAS2/P/0FO8pgIyF/0HF01ZBrdd1DbQKFBXX3ZjwmVbNq3Ke9nvRkugLR4nNIIKciPqb
svuRw6q7ByFyzjkuA0TyQoo2ZU9pIRUMW+vjQb3vXyMEvJ/4ybgW6M1+8TTKYePAR/IOxxyOx9j0
FgI0xG5c5QNB8pyaX2bsZO1xj/ttFWy/vbqIKKFYCDnuU8PEraP7ZNp6H7hKfhFjALWJ2ixZDEKB
s0q+LLL9C6/g53stUl11c/oLQCsXtRNd/K9nRtDp9M9pkYzyvQYX3n/qDbEQD/m0bG8EjtdgkHLR
djZDyyw/H4w9FY3MRYYmNllmlQijNbil86eAs8zg3WrFKeuPk2QdgnuIYYf4zZm4BpRp+7i2KSc/
24xmcsPq+tq6kJPjsvbqgAO3R/dj9NutYn+vhp0x0DoNX1o8lyTX1aS6CyUS+1RJ/OHB7u1GhEcU
JuqZDCqz0LrVZPYT0Uc+Ay924SJzNUg6ssbNKvHAX1JIuDHER6dDOF6s0UydE9CcO7YUajLiPUII
xG41NCkwfWOIYSQbCTm8Mtc4qKDXc7UOoOBojq5+oaO9GM2HBrDRUW9/rjNMFs8HwnHsOBqY0pY4
ah47ies2jN/7OynGoewBJ0iwhUHnCOPKyZQFBy4y6ZEcjwJHH7WwYYJ3G5eQwCMx2HqrZzPcRT5r
LRwthkvnGGRkEAjtWN7d6/5WUqpr+mQK5cwns20M4QfwrbTN2lcOOv+VSWgKRfK5KpR4Xm+P4GPq
t794JxGS+o8xg+mEnB4agHmvcXOAOa5606JcM2x2YdtxWx0l8KNUbMzywfTqu7B9IxJVBm9vrHAt
PNIsov5jX89SSZktAni0Oc2DjIyCpdGiEaxwSVgdRkvSb30976UFhEtx0cBZn1AG63OjsDil0pcK
YDPaqH+0iyjzPn64LJd9E0EKo9tyOcWafp1DJ62UuwrYzNnAhHw1+jscMXzMAZFB7SMKfl4Q5UWJ
/2blsneuN0zBVRy3oc+x+XoJWkuX5WjTyTJbJLbYZA3XNDqMdiWa4jQ7toJmORrLhFD2lX/yLgOX
x+jLBXy8FxVDa/pqfRdJO5OvcBJaoxgCbANryetttBBseGxOKMWBq4SnN6tu0L9weYxHf7SeEa0/
EE0vnvwRF5fi6ConinQ7wKf7XCyj2mzri/4Uy7/1sh/kbBahDV6pIqSxbdya2m5ywwUBNqQ2816e
p3i7ustHUvzTjBaVEEneyEtdk1ePSigIHt26gG0VOrKPT/xbFQ6s1AZixRp2+pMePNijcew7VNyi
5PQu2dqYsym/iqsQBmXovzuvLKhNXRItOEaavrofX5JO5pVyh8bHX3zeMQBFjnRefwOnSmFdarn8
4hx0kqRWgrjAgiAou+isjAYQ5YOfdTd7CHFvtSUfRlKplpfB5gmn9mSOm213EN532+5Ac44RnnNo
WEPyY++ru6M3Cu/D0QgbFUvDGoFEIzKkpdDxSOLKLyGGXEQ9SFYa0tHgqrwO095rrBwMZcfowcJq
RbyhzEcs+T+/jE23SeU1BFKU+RpGW3KYCmdQS8AsmXk7SKWqHeAVt/7F6XYqYkpEnRdvSbIRVYJ8
F0dlzC2KHLwHodQzdO21KqaOWvsXcCg8w6L1lc4GziJRUmj9fN2vORXM1/bWWFbcJoYdjrWQwkiX
YT8sPn0/qlccainVMeta7QmBL/UJjKMcnAsdBbkNF9aJ4PNDmJ7wltbEJHZ+w3NzM0k48v4czoQn
GKdfp7UjM5ap7kurNcQCpMQLFMYcWPy9M/3Fp/yv2jhpQ6yw+tpQ2eVU323M1VWxHsYUjPU23c2h
8y0hHFilsZeG42RtKfPykj6posPO3M4zFy2/0pHXDl4vhcKPsugS6nkBGC3MvpMJxBdSO8ewQncY
dm6LNJA5LXT+QNwQB62YXMihCZ5qBGMM0XJ+0Ddmr7sj/SOQRxYCdEYFyf4izxuT4XLqTj2qnN/W
fUxqnc+/lg8uNZogfEQETsKVM+SFriprRE0jRsHwnj8z0ozEJzkIyR6KngJgz4rwL//5DHmJSgRr
VR0hxS8sHOwdNiluadWnKkGj/bB9XipYem8ID4swRq2/3FIzK42GDOUiKkznBjyncYYxW1mwWqkW
NW52+ipiMtePfZ/onLSUgyaHbCxHgCOng7nIc+Z28WMUml1+/sE9v5q89FhDsv3im/oJymnc5ppP
wAsqxYNTdYqgeY+E2DBpPZw9F6fZJQE34/UezHsVcvvF3U3oY/WYO8Ng749B9O0u7vsgIl5qEsT0
1FRpvGC8Ik45rcDUHSPQFJRR/MMK7aNzaU1JrJdsFhdeMJQ6FgKgm3KcIFL2DDSmszfm2UYxfB0/
ZCx7d54euFfkgskn1oZTpR3lUYOyPQqVStQqUGC6+lI814uzgagcY03DOv6RqFBHmj00EJ44/Swp
IoKEzTp6iM9Y9ng4+JFlVrW7dT15WTgO9E+T288ltfPuf3b/qFMDpTxBe69qJGL6FAmPQQy+g3dF
D5aMO3y7larF/FwsLMd16ifNBgeiRXwfIy3DJv4OAw3rEptc/tlGjR/4bjZtfqJqNAFFsI1QP0rp
9FJgkA4XDrKO5ZkYwbWQa21rOovNacZCgGaZgKVCO9+DL5NFOrwdxjaVB4/IdrZ5mMlE5VttXMRy
lk6n0NUlIr9dM5OwWoBJNCZy127v5ki/S7WLYJNR2kcocZV9zhOVigMbPsJsYygvt7h/HdAAa09a
Y+SsICKD/lJ6vu2zG8VojYAzFofhlO32Q5gyw7IuPOR41sOwXC1gEHI7aSA5lWf/rYcK38rYFGEK
HFWBaDAMQJF/yeotMEPxG3PQ3wWuLj7OmFIoPPmKsKSEA2i4NdqDSYficz/H8VA6U75xkybcxK9d
UKpkdeG38Wnz37Y4N9UJBC5uHuDtRckqeEKK+7kK7UeVmcrJqiZOX+9jUm718OPQ1x0qyWCMcebh
8inGBKjlG/maDqUOpSCDZSg8JLmf405ObdnGKnJrdsL7t8L7Q4hzmQaRXfXX5DH/BU7uB1jKvuUt
mjAq1+zoK4J5v6ixSJtsk09zwej9mitDlyFAlXdMoTDr3G2ZTjNzo4wTNAqSg4zlNitVh/gw/m+t
K77jfhYGMyEhRlUdIMvpF+gIOgNIuPO0fpmXgd1dpogHiXfj8AqXfivy+XRW0jKY3XsjxAlUEe6s
npRDs2ykCF4drUayTXVpIa5yq96r4lBNqSDksgaueECqM7ZICxKyo10bVjDwJiKV3CmKMFuMmOrJ
PP3s9Gh+zzM6jvjceA+OPPDs4d+LdP8mBiqAYL2QZyRFo1Uo5CCAhsm2QpJhDI1vY9dblFqBUH2G
DHpIWh/LZ0wb+Hsk6g+CA1PdxU/ZDoT5n96vA0tES0VCtR16nbiaGx6DFP40rMSIsDdvB0Y2Hk+r
jZ6VXU5C/kjpn2krdbdezHQeBoFzy+WBZe68umNORf4Ls3TSjfJsZfL/B3U0YMjn29b+WFzioX8W
mPg0hv19xl0Am6+axyTAiCyJgIEqcxVE3hGuvZt3Nz7+VuHJkcRKvaViWED4c8L+uHJKLBnW61T7
Ifqy4l8RKZTXrJuZRk2fc+BgnWVZk34kGHlFE3IDO1go/gJEvVkvTMqbcoNDZh9Du3BQ/cCw+Qqm
2JgNrKOgwOQJskFq4Q1MtB2UH8Yxvwkg6D/FBD97D/xuMGnF1WTHRhwkfRsXcH79f1ES3RX0JCYi
/mHhyYai7YN4YU9JbrDgVZuN2q29JL8Wf4d7JSV8+HTPA4tN4flFuiT/TG1sqinJGsA3PH7osRMm
frFDbXjpyACwS3JTADGSFIGWUKomXlYxpIsOew6PpSuAPbFlRKdoEgQ8p3XSHP9J3iMQGErNzZ6R
Kde6mItAwCPLmMpvx1ZCZJGWB8jBXnfaHyCLMuJTxKNUNfrtW/GsAFp9JDVVE0fJRMV1XJ6qs72Z
2UZAQ+C8iysQ8vumb2bI9eJBnCRfhJfEroxri/1xWEwg4hebCRKLY3yhsDHYP6y1zaNmTr0WVajP
xfSF6VLW+BK0TJwJRfSlidk2FprRl6fXDd4z0DXy49uCNI4h+y0GzCdUrCNkrp/gitbB+7i6+sQa
QI7qv2ZclY2/kujI9Zqq4ZMsK993rXiBdnAL6o/N1nkCfNVG277Zz4w4uVq0DSi1BAOVdjzrS8SJ
da1ChO03LITdindYaXvSiQJEuB9l03h8gZTzG7kTzU9V3rjP6tO0ifrn+GinBUJEFVBEEMQoiE7e
l9y7VXPrymPL0hK7ssRTSgWjg7QX/cWEP/oNEk2cseis1UCGwtYKghLDLX2AG3WIYrbMayHh4S/z
nH0Ntf/msVQxXk4o/IqCZSiuC4UxRKbtuUgvLDyOdKjtQ2JWLrdIuwkjHvoPLhsAn/qzI5BC8E5Z
wXfpW4PX2rgb4MdTSbwpNko8cAhSCFDFaAJoxCRchbN0IzfjKRViPRb1QMRVzET9TofgEz9UWVgF
kMz33DArJ4AnsVK5kERZfHMOFEsRsQhbVhBtsTdsancSzn7lAVYyoxoYpUNX7UfkWEe41aV5dh5k
lOKkE3002FVFQQOPW3eDWbZrPgL4H9YH3STtEjkqp2iEHuM1Hy0h7RhAx6ipKFjITXoPpA5aAmIW
G56JP7QQ4hjuEfU7lX5BZ8tsFObel0bBjovr6r53qg6Pvi2ZJH6FWRYsZrDpBFeCm9p9Hyw8pETi
hT8QVP71IukIgt/XJGw5SMlZ5BO84hx8Hdad/aF4ELJYmE55CRVYtH6CT6GqZxiihWU8KKvVa+cz
tG8C4BIEyPNXxcgn6rZ9IW2J4GaReOkzU2aBOZ/YEFEfGwhbc8X3Oc8UPVwvsXd29H35xaXx8fMB
TTpx+dg6JadKrMWEt+QQ2doaO/agq+n4P2yErAkG7EYXj6YG+NCWkQMF4bNIUzhPHjrJ238962NW
rzBI/EfPoldVAAk2mlKsaZatcMVu4Utj01jy7X5s5QcqvMKWGk65+SqvCt1B+M+MkrB2PCbT37kR
7nHs8nQHGbv4f4OQ2HZ8GnhcK/q6RfxVtMmK/Ej0D0t38BAAcNF0EjmLBmKR5dFnstT6oi6ZNIzA
4Wwa7Tmw+MOM7xQSmquhEUfLf5Q9zq6lwHkzChLrNPuOaMBsPWNIRW50UmGo7TllG5nQlc9MV722
IdgZT0TodY50aUsaXfOhcN/LQId/FAYTDTa/CXxe3hss9wJz7z0nyKCydPO67W/QwX5NCq2Vrvb+
ZaG+59INjRBvaON3fCTNfEFIUMvESPIWaGRT6CfcGxF10fLaRne2c8WZRNesqEA0RUt11hm40eO2
Ypqjk7Dmvw2pq2Q9wYhiRLjgPiZ7oI8JD6PXW1dFQOV0DbsItohNy6/l2hOmfse44jIl67LzIjgf
U4bPcJ77LYQOnSEoB3srBE9M2urL4ssBHH0fUn0wNVvP+ojDI0FiNW6WT+Z83geuqPfgVvgrlbyV
/ngIq6FIJTWjA0YxcLwCNMuVOSFzIDLux65B8Z9+iRgK8aqrZLYWGSBHMzZvlsBYGHwDh1K/u35B
LnDqScu7UO4GAQdTRs2gL9YimbVNJURGv8hDF07458BC9keRnxduayGYsJAzvqf5O5Cj4AScJY3z
XxQ3hWW6q/Bp7+YCzoiQ32Cax3oK0rGJNYFXuhMd+M3s5LBlEocoDLGpV9Q6srXtWsyolgCzhht5
Tr7frscnEBq8RGKbjf3ZBxrBleTS8IxoDH33/Yc1hgruV7rTl7VfIkxw4BBPbygIECTWGZNWx2Lw
abdTXOVsMA82/77WpO2KG+ZFk+119uOLBW2ofl7SMM8cvYgByt6Npdu2+3I1eK+/UmD1zVSb4Ajb
w+EnIByqQyLo+fKtQaUrEa47kyxyTetEcPM0TJvMSYEKQPGyHYK+bACxujK07BQVWRo4X+vqEJXg
3HO+3d7gXBa+5SE/YddKaf/jqyetUPPeJxUcCX03YFNLCXIrcEZ2Wu1OxzQq+GQx3bE2fIw1mWjv
vVcEgpAK9sOY9LKkgcaWcN1mx+qFLebPOn25TfHO6lWvo/ujbW8l85ie5BMuh5Xp1nadsAisYwlv
HZMHCMQ/P75rXjfMsuMOuVKIE4nODukpRoHn9Lk4fscyZBHi0UKxUAntdxd1oKbRtef6NM4/VqI3
1O3cDT8zWPsOW78UahCr05UGngr/CzhaQGVYYcfE5xybpAZ5HCcas3f1acnJGrOL8Tg9TpyW7k9S
1PB4CRZm0csuJZT6EFAt6gd5lVNP56klob7OJBzPovT/jxyQfN8u4su+Ygj8LVSsutN7hRYDa4PO
8FrHrhTaabm1Q8DENetnycN+Xwi7uipEFv1DevqzQ+LhuKZIcEVppmviZJ4zrF3o3amRd/EOb7B5
rgztNBAwmxZZQFNaiYmZ3g3n20aZ/HvDiToYMfi2QfrtExlIE55qXR3jARnkBnmTl4OLEzf9ggM7
OWiephkLa6sMM8/OF660QIhqD+8L9Dq91S/rQRo8/LwEYjIPcltsM5OtqOhxBy9eTpzA4N+mrAP4
uhXu0YNvO8P/87NiBy0bK1xbbpzyXb8J0TydaKbCYXqTZ4hV1xwTL9uo2hzTpx0Yqv47Tox0avLW
0DcLj1CVCdVMFlN/WmMQN5dO7Axg3Q6cua4R7L010kWssYT+B0zj8DI1Rn0RG+54pUWX/6WHIoqk
GIXD2ztnqIEkAsiBkRMkAViMnzURps8kq8GJqa53xUWTQSv3JvbkI8VerVbn3h4p4avKQxz6wCfU
0rK1lk+IVnzl+/uj7wcOqebx9IAZvjBy3UOCtEPh5lCJ9uA5U2pqVmaz7sBMirdcelZcbNC4DUV+
lpslvUZaKzvVGCxV6T5vJfEBSRJvn0t26KkexX9y+gL2kqLQ4w2gFLc7WUuHuXh8ng5YCqpxtLKz
kyOEMM7AV7+Wp4vicUfR9NzW1kTkzEZSjiEUdSXOFWI8BKk2hj6kBAZua3NGrZ31Lj+oyBnIAKh5
AZ/G78tGfhX2jR1Hs6qhTfS7/Yu7LevcvKJg/+64UTlOcmeSP3a44JqUq9pZ1W/Dv6d1UIeMhM/T
tHSll7JF44A7q4KJoHc9SuMM3sY4V8DOD/sjt9iaNzcY6SzgNolkV9dmnEE8FCeVqFF2OJYduBSi
gSWE5g0d03Ig1UpUMKh/Fw4jma/GlTiiDY+/sgqm5dKepQ97ufbkJho9nw7i5sjkaDBBGwggrqu7
N3xqxVktyhRpD+cjtC1pdGrEhECZnoiAY9ZBdZ1O+3o+l8AyExlxx/0hZN4fYgJBshx5oGY5qn8D
Uln9wFiFahLjGjM9PfAhKY1aoYai13QrmmOq91sUbvQa/BsdJNNkocU+UaQQqqqa1jEBqtIsSjGY
oC6CzyuJ80uLkmgScbp5JLH8MmC2YGEOWHUkpdyOpEXspRCeAXpRJB/Rk9cPLLeNr9LAV8tzmWhJ
jfRbOSbfBnjQh5t/cYiX064uJ3E1SDySPbiUVmITbS7jlTcpNGRhKSgz2qDvritQCS5K7CC3C6ii
AZ/vqd8fcG41RpTr9uLLIERBiEywaCTaTK1QQoVXCC67ThJLfPzi8nTJNaEFF8yj8Sz9wd9u1I2E
mUIBsy+o7VsTgPV8mvTrwz43p/Yh4lAMtuaXqpOxq4E+jWbLU4zuTQWtpn5Pjtdcpj29R2Lo9cU1
MEME+KGx2NzbziuX5vebN4j6Yg/EGBhaa8OsrIwphIcph5P5nbj3RoyHCvNn7afpCbK6tVMtNWSi
UoaUcriMkyGX8tlJf9IexB+jKtOBFvTEtEGx6Vfeei1B8UJmuYSiD2OjIbrTam69MkcuDQ6QAF4L
Xh8IGbUgOxbxhSecDxFYcXsAPLWCzNs56e2XiyrW5EVQzJZwTER2rlAk0wr+VJDKJsRII17X9qIg
zA7hIZt5Z0RQXssWCHQye/tAPfyUqx1OKkR+bznL+CLKKmWd715KN7ZiaPC6lHrel4S+GTsJcmeb
effm6V8Zk2kbour848Hrj5KP7QSmJVQoHhXX0wDmVb9ufq/ejPZPJ3fkRgwjWcW8U8ie+GF+wLH2
zwS3r/Bat7MH651zAVMthMnz2qSvzCVesH7uRGt3VOmLHVj//a+yCpLGSaMp1qS0gdh3/v1JKwmD
5m9SCBKflDazfeOM22TUiLOf5O8fnqM0vWRJ5RFTz1A8Cw5AaPcTr9xsp9+dIk+OF3mhekvw5Vbz
frl88dhFx+1Y7aVQeYiaGuQz+87df12GTwKQJ05FSPGeOzJxjymKEs9QFFv3jsvXKxac5zsLHVAF
gBOj4PpzWILjtSgg8zZTVyB79ymZdJIhVJjryQjeONApUwkuJaM/IZvLPL6zH9vYdnuy8J52+skZ
AByXINsJdDjRGoVcn2SV03Y33LMnMCQS8RzVgGExXs3i6AEhueZKHZpN44qkSb+d/guV5mnNsZ6R
7s2ASfN82heyOJnkrhGCDh/7+6gnbywdqZ9pp9vpVj5FIAYR+RwKy0GAnpSROFylXjAT0TCk8tx5
e+NTKmyi29GWmA15v12IxP6JUQC/sZFRdyCBzWTVrgKFrhxYegZsuh3Rm2SHVjrxJIrKXviTpxTi
MZezPXJE/KSIZn0etuzcg2COr2bdWQm1uma+ZYSa2dlIhGmqHsAO29Jp6c6PMUXDMbAV4IoDXCEx
AnWxEXaCkNU6kxThp0WjXAr+coRNiJQicpVdDrro6jYcZCMn5KimvSaDv9OtdLG2B/iBwZT2d3WY
BEQ+G+lJbqQn8hg0eIXmO3GTUXCEqlL104lXJIxtze+rQo87oEMUYczFZbHf3cQp4YbBiNWX+2z0
uE75YoJE6eNys91/sz7iO8mwvrIWWVsj2xXxDf/hCliwDzztE8tb5G3qyxku4L1nso88LrHHelW0
k7HF2z+9tr/r+YNL3R8/sSZsQgQBdGYlqq2itIJhQ7QOlP3/9HVNX3TMm0Tv9TERX6tEzC3+iG/a
TMqkto0kv1b/u7tthRGPpfW6oPHGDxK0JFlFcFkXvMdteWO1zw2p4L6IDYY2h82HkXplYTyxbDP7
ydXHSu4XxFz1Qj2TMrntIGtPIwHhQH5RvmYvF4jNLoTBEwl7zwCXfpd6nyyJ/7d4702ckQb3Ia7e
NZRTYr7twAbR5EyUEFJ5UvBiSZ9ZGKhdoEzkF30HTGe4F85vYr3+VtuLWt25gg9MIqfcPqpIcQ/T
nEdtNpZ8nawa8PCH/rJDwEeB30Lx9S+Lg4ODxCY7GjSm9tB0o3WkctkrUxTj10u+lkudsGJKAnPB
N+f4Er2KG726cHtErdW2GvZhhZ9Q54d1CXFKJ+/LaVltNkKZIRR5dYRSf+1fjpqCZX/Xk54kGwJw
oSHyKRMtOAGMog+YOHZFJ5nYwj0yudKywStwJzQhG+KKjEyr7jLE3vZipRDiWydxJIBTydRi0x66
PKz9yAAnnr+nt8Lk4EKTQw8UgLqwJDiy50OIyjRyqvFebOA99N5BjbKmg0J2lobEmOfzIR9uPX2s
nokmZfxpoeSdu+ouE6vQQ5PqAHA2Ac0SwJ8wV8rBSVcfYtS67hkPqAtovjiDomyjfpYseY5Z+/4p
Oikg/h1BcrgHWcmCp6tTINO1vuDwdsrjq4Pn4YmbhofslRxLOKTPEbYp4qRl/R3Rs6+FVukI6/wI
4Vgp/WEsKtS6di5U5I9Hnjgn8z/LVhxC2Mni6B0pzX/kzRMPppOtKwFye5rk9G1c/WV+qaHHcnkD
l3P/rc+g1HK8lgHG9jU2XvXetDJXZyn8z04CznFpmH2Zh+kkDoOhEpo9lxflCFHsQSBFs0mPJMCc
siH1A7+CqhNLldvL1qVXvb93vwYz6jL0gZVCnSGDPFBf/RdypLx96/Gh2/mySCcoh6nURp2qchRM
4bLB/IYYBRC5lga87l1lqSjeXiGnsbLUnYG4O0YCfXMkI6kN5ZuByM8qJ8ddBk2f82MtqZtyBJIZ
hIw8ExAk1tTcVUvqTr1mluLG/vdz2gjgCt479DT/RgzMZjY5JQdheAYjcb2EfbPHXX1r6VYD9pl1
c54RwZvwMMzWaiftkzii63waI/RmbaIScZk9f/BaRfqfjT4VmI1dALsWVlGnfOJoD2qmMMbYtAiz
L8TyG1ZYU2r/KSzfhKljQj6Npeflig6ryRDBQlzEftdZDT0LollfKTqOSSB4X0pi7UWP7Xd4/6h0
5iJa/iguz6+vDCDRDkysl+NJDsXnMnNOmnXs5I69pvE487U0PQptERHgz9i5tYTgZj3eXhtcyFNs
xTOL0AWXbGoDk6JLsbfQWz11q8eIydGVURQxj4NTbYPBCTVEoFoLkmLQ+I3yRC4S4ACJZsytXZBz
iJrtSHI0wlIcJjBNY5cKIt1/EwQdGmcit2HQpSM/lmpG9llNiofxx79L7jXuUZPG3Fn7heIqjdBe
oh8RB4QnNiqWjaa6g/uoo8bA4009ywXJhH5codT260+uusycuZcRgyoA6Ij2wPk410Xs3fxs3/95
TVtrr/Ay4XYxOoz2KEdJ1+5gpE7wnuP01vCSSviAfL0TiTlPuwPOwWOtnZ7kXkMfKv+5uVKNyqbe
9KdQIaTUWW4WPO9+CeZm/v+3SJKUYiPIq42GG/goX5SgpGNPHDPDgtOySH/4m+fRH+vw27IRclaS
0rPopZX15M2yZuEarNlt5Qull3TKa5xptc91wTtcBpDkRlRqlGfLSNjS3nz6fo40Mi7S2q4OfFTi
jPoQtyCW5r3xom0+U8LdZVaXb+HVIIQTnognykXa7P5EHBDfutZuHSpri6YjTv3J8XUuw047JugS
T9zjfbrXTVFGGWhxrtm8S4Lw9wEZJc5Ixi5PmqhJeakAbhsW/v3Uh3HbR0IAWPDg/jkt4d/RCOd+
/OE/gpw5j1nIqE76YJqr0rDKrpBoxsXL2/iTZ5Z9XxT77nkFHifSsKtvfwpoFqultOphNw4zN4e2
WYGsDWy1kfBHKoq9IdFe77AKp+sndEbUycplb0Wb3esO3Mn9ptXjrXBmIzyglYCnQgbguQRAE4an
Ww9S5x3zjtnT3YjGXNE5Mc5k5GRdqsYuPSJpAELw6Q4dL5hHWIDGcE45omliAhCkuFzKIbkqoC5I
Mugvc3Q5A5xMv6hQsqPrTEvjBVqBU6IGW42RtBO/wbfTLe/Om7+NIRlhLGtsrkip6sAarYcZF7BW
Lxx4uxPx8KLZZLmHenxVYxDPgrRqtT5v3gf4CIjVvAlEHTMfThn/yXxIHa3rX7FhEGCzo6+LmhhO
k5fjmKmTuHcVhy25FJh4H1vfxAnXe4np0Tc9azv3kUpH55WiiLkdx4EpsQlGSGQut5qim1jkNJMG
z6uRw6Vq9tUmAbFEiULoU6v+JAV5BXZAkbXmYHmGZimBaAgsu/VjVgnPqpoOcj0sJZdAhrxgMka1
3+OUsrvJmBJt0D28IrYWuAUQ3QJFrVb14pkKAvHTav0NPwEBrv1rrkKKlyFW+5MmWQcKBoZsWPOi
On9wcX8SCDKx4BcLiV//pVh83/R4dvo3nVDcKmPXz0mq3BqbzslZD3/nQrNVggmJxECe4Yj4tAXD
S8uImIhKsNeMaAPKyLjqT8FhwxOxSAB9Yje3NvDUKV6wyMEbcGL7TkkgKMvcJcbBWCGNVOmkjHCr
kGqSe8SXjkhFW2fqtA3ZWaofVwLYSfBtNnwnc1pWVarJuuURZrnuno3/RRo45YaKtNz5AV4dGPTE
GPONuA72AYbFYmxubqRm5Ps6cAp1eR3cDcyN+j61hLDnfh3FuvuZ3KCPxCVzqhuCPORTuiZJaWE6
NrmQxmhn5CaWhPmTRIUUEVMgPAmTUEkSf36J/Kk8g8gi0NUPNZePLRDwg/maZ1imBmMWK3BS+A6H
3yNJekp+UMv0WsjptIWXxs/72FqDGM12xmZllX35H0849iqP+Skb0eM5+0z7qePjDXkns3CWtAQ0
WS8uzSWYhK7xlixLnoPdni/adnM1p12zHfDYXOieip20Lp/iSSJEE1N5mN0impIvCFmapWHrG9qJ
48t6MyvsSa4vrdViR93xah5aQMmemcUFMsHZZI+d9mjtdaWZpoNjs2LttoruYs9d3ovn96zU6kSJ
e/ALeRQZQq8sVL7PevfGSr1tDFbjrt1Q7JoN8jOF1MRZJvL1BM1j9MiXuY5CELbRSx46H+RD4zz5
5646O0tOwh2H/HRPvPtE35i7n9XCA/Q8Xgqj2A8nI/YfZjUUGYPgYlkJIFmSIzWzm3Fu3aQASK+D
ee2IReH3grzMf1WjjyVpt5u//XrrjhAJfH0m24QQRURDstnII60d8VcHKcznHjvt70TsXoVkif0R
jxoS0k4F7vwzsSAzljrb8DRjv1ustJ1T4flQTKVMRXYS+6f6Y4CL6TO/+2rawIqeipWFfaomwGJW
baRSXlbJeaL5fkWYCof1SBpAgK+pBQDGLoBYdBac8teVCDHq8XWIbUzKBk87OS9iyh+QsOyjj3dz
RlamyjKAyiRTqRhal5RxA7gB4bZZpfw4bcX1bSt1BrsljnpM/11ZJClxlA9qlrz8kbqQRWnEpyPg
1JBfyyMN3Yfk1hnX4T7SuftK/a/evkcv5QbG1GR0ZS1AttRiyFkbEHDWmkKBrTCE3b4CURQgXx3L
Z4NQOg8XMhCatQyH1oB/AHRND5L2XdEm4EnBxBcgW3p97WJy/7CpJcf3cDLSqPsAQmCQDbCKbaNG
5xLAcKz9HLEfYF+h7EX07bgR9yDbGAK6ppZBSV6Tn8jPdB13AvfIDZpIJydPFzIOu7TrgE4Aea8Q
3R5pIIfvHgo8o9p7APFofys07cQxnghMMVxld5DCPUYalEq7n7V1e1+BLGc4M0SK9pYb9IPu+gUn
CVqu7JIdtdsWPJVh++SwSZUol6TCXuysLOIc0p4h1R2sSZ0JYZb4Vlx2Scz13myXZt5itWJqVI9/
RLbn80R7lsS92idqUuAUlEN3dxv+0lzmE1q8pQ0eOKBTlEmJ3jLC5oCBfjrLl0qZYR7tzWFT99ny
DFRgyE33zzkQbmcaf+woGF8fxKi8TzTVvaWU8wjlN2ET1qLZ1HMWY30IDC+hT1xONRUNowYpFztz
wpTLhTrGGLPkiggmQPfe1fKEeixT1dBWfCFBot1yJqsx3l0h2CM0ap8Nb0wtiGnHzKGhLor8gR7y
5kt4oV9FHIxBhdG/xKH4s29JPD7EfIGzMv5ZN+hBOIUIkcak9NACyfWm4C0Eks8HRdZF3wPshYO9
ORZWZz5/kTy9BAB8o2sFnsVSKVDm0bN1PgK+BCuTjJzOvfwYQKxjT6EMd9uUa1svUBYBHeHxHdC2
8cIrurbp4jqmzekkfOGbyqyzlwdaYQI8gGEj+dggfcQlsLeGJN/1Law2m5TKg0Ox+r0jZ4puxgfU
Kg34PVa+sM5eyjUQ9jD64QAxIkuhxrz1Egdq3rTHyJMuKavk4xb1yfsOqzI35xWqU8y0j+7IeXEC
dAbRed9pjNl1RVmhZ1MaEC3hz6Mt2EFfHm2c/y5wLNzsInIJ0d6+Mok1uFgxmI88A70nHGc2DNTc
Pmoja9C2QO3gWSgPhK46L4/Iers+YUQTN2lgyHiu/2FPotD8PcT+vH2tkc6LLOxSyyFLBSBQPhMV
csZMPRw1VIgSNAzbOUYF6VXD5vS9kafHO5d5YhcEgrSBE83Nxf9x+DmAnDd7mXCxprr9jA1+wAAV
so2YWZ4O/LnkdHuzcC7g5BLvBwkjtyJLDgQEnmpQnYc8xERBdJodpK1ZmoYkb0vrlc6drtFMkgCp
MXvdvrEcBU33xzlLk+tGqLMEcQnmLUUYxXGTBZAtVvtXoIAn9DoZ4n4nRh7KKuHeUIQ38BsQ75zU
8FppXCn9BKk1PLspdRC8PdwXzMY0XG1e+Mc3nHyFXrT8WZepSDBKFaVXkwL4rj3Oq46U+F1YTGcN
kDXysOG2Yz/vfKbGnlF2ox9qzT0Zoas2QGfRM0UnmQ8c2d3PwTJSWo4271HaDvmoChcxIAFzlryb
KVd/Y0Le7Edn3DlbEASnyUQt7Ocar8mCModb8pvnoPOz3mODtX2gtyIB7ah/7xzP7c69kRwPB+KQ
TLg7lDg50za7TYo0RnrBTUt8g74POure5uI7laM+CyDCymjs4ouvQ7wyBzKL7XYlo5SUUuylsBFs
imTA/6mhuhKVf588u+TOlipqSyOP1kcVw7ylv81o3e5h5qbneX4uT0Zl6Fvm90xWCZDh1uE9snlP
/4GfmqnNIywN/KgEOOJ6nGNdeAC/cE/vZEydIFaptrx9NkqB2TuIpKk9MXWgAmqe8s3iLSAVYv9B
IEnK8jEX6BknHUqI2uAkaEkZ7jdpuMp6hpUesqbecyagCpCkdaxSM5D6xLzms3OGIsrnPNYSyJQ2
X6qmhtY7WjndJRARzOpXKmXlJtYj0HgYcYa9xbOKl5e8Mh6DSlwrItMT3DCkUeDz32DdAMQxirA9
jYdv8WVHE1DByAGwU2UrQQ4Xa/NBU8I89JayqZV1LGsr3nqbCQsuXkk9Ypyy2ulSOUuUbIpJmfqy
qOut7CnRzwMwVSeiuBdsC9iO/dOSVSGiK9bi6s6nZ4WijXteFf5AiIVAj5xMfDT0uwEXDlsN8DWZ
OwkOPL+5Be8abAEw882AFaLuvx0mScVeNkmH+zW2wLPsm561AZZvQUKrxTsv2Sy7x1w9fcLyRedl
T624D7RVi1MjzdpTb64UhtZCACDbv1lHZv6xDc4SCg2aSiVYe1xeNmvAa+etfFNWO6bhJa6OZm5i
es4D3ZsEZgvOjXx3faq4H5RYZd1CPqKCERK4Ky4HLZo4AXLotpnbqKlOXmP90kPQAA9IkODO+D07
b4xfJQb9sYu4K2AfvHoQ2Z++xanOXjznoF0PNZVmEYSRvstTKTqBVL+n8k5xFzgG6ZdqltuDlqON
rxfYnCOe+FavpdJuaUblNhh9FSUY7neobrmln6efsDf3MdS1NaRjeTivEKsbcMI5hMWvicsKc09O
yrA+ohSM0u6V6TfL0b5EECDjh9BVmkgIwjiPMED6XDZf/cqQzQT1yGTd9B+NyTyq8zDGH6xikwYF
pIn8HcQuPBSxoOi4TBSBviGTm1UEXbLT9bJ5zOZoLLcSZtSejuHHYgtysPBh4KsLKw7WtWvH3mSy
cgKgDgP2yZk2iEul3sUICJ5wyXkQuQEUcFl/Z3RNtw/cn9swuWwimFv3syb3eYiwfMffbJWZ+qEk
qBggTRzRxj+mr2kfLQc7XtZ7PaVXBxrLOHD+104u9PEKM6QkNLKzqrS/uGoGhzOUREXVCVBDhHLX
sV3bz+U/cjeHVOTWL+jxcKZIpF0ENonPq8fLFfJ0WbzC0i5+LWD1nH4cVIlRehouXPWdG1289dNW
lUNQkkvfLamKRHfbu5lrQ+IFfIqwiQ1OgU4R8EOwtzmVnDRyMq5tbaGCu4rNttacOuVWgWKCn9lb
Zu6LfFViGtOEm8lSEUDKgj5mEfpZlA0OXpDJvtuvpsJ062c1HhJ9Rd6Ve92fsJ2YzWd+3xSY4F/W
Bc0cmDNIFlQOSV72O8dCy4GVoQnrCojmwz63jkgNOB6dCLsCD8riQI3RnuhiaqQoei8CE9ycK79h
JAJjGyd8AFndYMt1uKPHLhwj3pIKXFH0CNtJfoLcpDmj0bGwtl9mi/4zu76kAlF0SzyI4AH8cIqv
MN19AGiw2BejG2NaHQDxXV9zHHYpQwbsZZ2/sgpI66hi5GV5CnapyzwoKq68Lg7tXCnk+zNA5u8D
E5NwoLNDPCyQwFKGT1ghaFoLeNfXmJngRE9INcp6ChegCDk0dWiU8DpEGgESVosnz3BETzltLker
KNQj75es+nbY8RqhGomSY++39ilLFTv/QgeSu/FO1zcVZZmKMNb8J+NE0Z/1MbJxmKfdyggG6YLk
6qHNCcGLmQtOw6VLygX4sxvwCxvGoDttY/w3CWkQqaCccFIUjwddlHj7VvZ73C0FoxgB2N+rNSD7
cn33ASnBhNa5de0gmMmEENXFTgmvxXQ4zudydoIU2Q5JlTbRTlt/RCLHBZY6S5xJliETafaT7kw9
Dp1le7ezRWyBPEVrv0uFPfyRi9ZcW2fjQYw9zxDEG4c+DOIg+enaldhahV94VEj71YKSQSag8FpZ
pFVCcMYWhAK94BIofl/AQKSbCArvE15O2W8LNBRr2chcY0GEdtNSxCpAnlO70ithaaP9VeWWId2i
0JWElUhO2ud1wyDIkyOpOSN6n+vKVZJwQWuUNxmpnUsTY2EnzsqQHE7iN6puPMXFNVLtHKDSutfB
gqy640IhYqzOa0PXLyixjoTCCZmtBUA/PyebH827LsWarSDtOmCoWUFdKY6CVao+5C282LlAMpaq
kI/pv/i9hNkz8uyl392TuvfsGNstMxEKOLMevlOSFePMSI3JihTl+qqhyrPHCbmYurxKPaykCMrL
iBR45vEk/gpTnbmqGG+IlbjVprr1Rv98oXP6NXt0vHrLK9E4X267bcD6eLvdGHaRKAjAGRZ3/Zsl
ODSwJyBE/OY83k8tq/Wn6jV7Uo+tUdonvAq2YIkDIUecsrWYpoKVuMHEj8qATEJ55pR+iC9MdryX
ir0LPi/xzmdCT8wwWNaRzJGIsbFYL2cLTsLidPDfNqydRHywdjJGVan+dm6Ib7zxl9PDQ1ZCM6wL
FJnxpQQvTYzjnxSYPtxcd+Sk1B9LpAA9bUK//JQM9TDGBEJQ7GDAFgosEErZuD2XMqMOr00Qfs4M
EOLJMUTJAg4SZm1UvXX13a9uZKR6epcZKhMkD6P1THJy/MYkjzgIDL9/qQyXff0sDbf2zHyVZtFe
QmIJfCsK1YZA/bIkPiH0H59sYw0GzVkwEkHKs9yuFjmhNlDaagwF1aBH0qpjAu4T6O/53VVxj4d9
gG9Fat9zAFnYGQRj2IDCAQOaXQ3uhCgRdcPGpfFF7L1dTsK+9jlGdvUyCQ2NhQKvbb+aSD4vaMvr
1t5AnwZddvyTSR648uys73xzPom6/GRFAVVWSCTIeALiKKR+4d58qJ5/k265aWtk7RO/h2xjmYUg
L7FKfq47SA5mmg7Y0junFW/7ug52PJU5d+bfrQFEihe1BI4lBusacSTLWGOVb0rarDnWASe+8z6b
GB8ChrlM/0IULZOoadnTBi8rBDkqdF/eB4SfQANQ4Dv/Cp7gu8wuypc15mgCgZDu+0chmFWOC+Xb
raMD2subaYu5Z5vynrejKOQEDkFja+SeOSBV6p9fgqe+AXbG/SbXQHjE8Vp+V9COeCKHIRhJSIVx
ZBUUXYNLRdQ+7VmzQiNwuguyrzG2CiXBgUSS/CQ836BINru8YpqgiikWpfrhm1gZYqdHxknE3mB1
yFN8r1zxnoQgen6HxVCoaJS3lPqj9xJ+s7jC7LyZH+LKtTVBVowpok0zs5KAzrlnhZF6x+APRgAB
nH1n7c4iv9mCYZgeejbU2riiWt8cSjBpAbKhJirt8iREoLxckCXhZf+4tz94OrbW0ka5fBjsf9nb
u9U4zW7Aa5o17qdUfMtkiVSzpV4e4DlgD7fZcmQ3Apm4fCv2b183yodFikycsHJfBaWvU380QSqR
k11t20Vj2tzBYZ9giV+xdz2e+evLU0SLRUD7lvEVHYCRvxZoR4wPrORGrXxNZHpnWw0Rilwf5O7o
LT6suyBEuqYgamte/pibLQ4TOPLZE5pqwqzedDfN3u+Xi3Qmqu9x2CXHeecdKvWKAdfgxqqJX7ak
gJ+DUOYV85YpUE9zXWhIRTQ0Vf9neq5tR+1zvMgJ1dq4y1W2h+RWLwsaWP59Kh3BVGNx9MLdFXWr
S9lOVka8cN8O1OF1IhguL6ocdTu/5jtDFatVxzL13w9000S3UV0y+Vb8vsPcfg1VDM4wTzsp+ayw
14sqXQWdmV/+GhEyiUUBSqwHzbD/Z+RMjDn09w/qFlfsVbuCgO478Nj2jPIqeEhnBFe+Gz/IRh6y
PoDeVHGIz/9gONyaEDMM0m2M4mg/3YtMh8p2NFUQJMrvRQcqbqWXlW6Rt0K0A1DkXINI2pM6JpSI
vbD8Mo9DW9x7FhEq8ukDwENXc3GfrDPjyyLjvJDV6WCP9pxF7eO/zPdtgDIb/oIBl/s4w2CrN9xz
uaf/ns699Lzo+p4SdkhIzDAjpAyadzOZIUj96aTSiB7HZF5UhZ7O2vRiF0T8JPUYkz5uU2TMPPVA
MrfR3RtBdG4vfdD5gDu0EuOxbwzxsDMeDcjSnXbbOd1SveFS3YOOAiADPS53xY6KNrI+md2I2vhx
iMgaRxrobNR1a5s5hxp7runNUxA/5nSLau02O6X3QaUTh0tggE2T59E3mDRXK2WSDHveL2ZbMf8D
qDzkGUyq7OlyqjXnQBEWb9J/pfScJpLxI1LPotnRtVhwpq42eNVO9S+Co6J1SWbMr4qfnxOCftO2
dsCcysczQl25ZbqEfjxp3+zCw25L7OL+ta96krfWM/sXg2wLd/N/gGIJL95UB3wd7TfIzUzXlTF/
SkAprKi5YPZmkJ+Q6rWDs07EnAqMh0Nh2ScE6Y8o10PxS2Eq2ltNzCo6TiLdwYltZJw2UJGnGREZ
4zhHnttKk2CbXf1hJBtEkSBqb36U+51VJCm7fyt+d3xq9waIc0nWwh8FggOFf8hkVjNQBio8bVxW
O5QgWUvBN5yZqzLSwfUHPKIZyb4pbhJbBOMQza67vedh1VnDm8ZEelAORRvTWZloAdvWYXnQeKCg
As1PiiuYX8lMlTr2zIFKbH5c6GUS+PlesOZAkhItvOq6yMsZ7iZs+UulWmHM/4IggCdfi//E44w5
owd8VkqRVbxTp8YW0AKOQD4g+Seb5bP7IHyLHI5VISR7YHYF9AjzMtNNqXDVAWQVnd2Fb7mBnQH4
/DSEHshkYY6WvTt358xVdy37mkkhHPZOJqdb01y1Y2trFnjzwHycYCExKQ1GSQbCaEzuAcPr/5lV
iYtWBi8CpVrHbTdxLaSSCtT6WosERX5XiSYj3r2eSQsM6zLfeKcmhgLnvgiLYFb/gnwoaF6gxme9
/29paXEuZ5xe6L+XFLlEK1n8m5I3TaF265wlPBsVOKVked0qYkElkGE5LpVOS4WoWrA/WbUFwBeO
i2ME1l+OijSxnT9zgYQAHOvOrFtv546tDmfB1gDTYkXj8qzhyzQtPSgTEr9XEbC3LJ09lAjlXI+/
t9znoemCMhNzhwuqPEW+Gjbsg7liJ1QestBXPG0CV3pD0tSE1fam9Gm5aPSwdQo2dOftis/HqaZY
8bEktvcWGcRWfP2u6NSwQY/1tgT+P/Nz4tVgWdPhcVVr/bdIPdR82W4PlDe8IcsQJPfD5mHmtSjh
ZLGy2W3+WLN6gGhlETdtMNPOPeHBvTWj+Vye+9d0tU7Xe1breNVRxwLa8QRhVxpSZkv46RcMqSdU
FR5J8w6a+zWc++tTPLukIXULjb/XKi81OdVjECXihCyPj7sculJDG0Whc6cdO2kAtWMs6F9QqgHb
obfC/gHc7/TJdANRn2dPfWpegAP8K9vTZNAZ1BTiwk1i6QEsSPD1nTiM1rz0o4ywmL4628WYlMOE
z2pQMz8ywv3s9MSZlbi/E1372Vkzwj/f7m+OUHldfCyhPMoRgcSgbvOsw1QK5OG21NzktQElKe3I
pWGvH2Oq0eYVXny1Jm8ZOnfbjjY0YxODQGoXW/JlHAzen5bymMZwynNCE4qCh2a27+m4vJdR4Y5O
fXQV+QiL0Z/pH4nPeUXqDurZAGplAVVI3bU5OhHK1dZKsYjbllUBktvsgqjRQTdhhqo2DBcLQhav
F14gs2qAx7wIdYXaJ40CV/vw738EivMlOeBrEdJSfFEOCgx4cse2Ko9/Y68CJFJKb16oemB0xZEc
MtCvO3YXTL6HT+UF5JMifwsamGIqe6vbaTFJSDbkMZgdRJJtmPVBIN9rwWDWWOMIR3TZK1RlK3wA
rVfT0v6LPuCtpOm5rS+xAKmRMRGil7YXBcj7+PudrjpkWHd0U+P5fxO1kfg4ls+nO4+g8o55Nh7n
AjV5JQQbq2+1d5/WsYdXiWtRUI55meh8NLMtzpRbtVcJqWxMn08ugLbE7oyeZ060pBdLQr+QqxQD
UsjRpyy6jh0O/PrOWtq2QxFhOtd0FQuLT13WllLjGWBjFaXw4zaAhCObptfom6WkS2x1sr/qWOxa
OUUK+TTyk3TWusUxt3TkCTK4sKAQuaCcnCTWWbUJ/52dZFhZq9jsruldU5uRh8AwUT+fLH44D0de
VMnRzcyKagcIggKCRVyZ50j0uisLi1xZnJA9x2BUzUpbh4dt6vn51N3WBgUa4cJB3VHkYiE2wPB0
2i3mVis1ALBTyI9mjUJjhpEpxSJO0wc1eRjHT6Ha+BBpsQ0Oy29ry4LzKmJsFl7v6crFEreSZHH1
+3Sw/UqCuQZnbvGdbp/6xj7i/xE9FLrVUY1AL1K1Nd83sJokyhbuJa1l11UJ1v9lTESH0s4BgK+Z
DDaAXhscz4sR9fkLajWFNKvq3qrvYMuv4EREkCGCXOF0B1PVa5NxQwVh3CRuQ3MmXJNsN815mUzM
VsJcuo4Cz1IAG8fObistweq6yFKXVPlcy0LjCHHcTvVl2x/Ff4HEH4sIzXBk21Yeo+T3DTtRuYBW
9nByu/sc9L7sCzozKUkRliip8q3g/YcBeGr4H1v5ahXvEfjIc1iWf/SJbEsyeMS/j7Q9C0mrhz7A
xepVOvjYsi0iQnY4/MwV4m3LKgdNJrvo08DSTu1ygnUaiNBzGj4GFVQrPah20QFMAp8sExmwUMQi
jiV4tTU5yDyaWaxGWTgVwHzyBi2KWda8nFoS4v1TmWOvNR6KK+Ix1l2by1IjiEX212TyIWNVOhYO
xfek58ARbaGcb820g9Mq65q8HzbCJiAkowldWKwBy0i+UtIgphjtLrikF2heme0Ib+2ufOuzvykU
fAWOP2qooAg0iOWPL1CqBArp89tzgJf8s7IWLO+5DOwysMb7du2UU0SrleT+PHx751PUXsghyso4
jdz6VjVOWixDFlYgd/VyLHGbtTN9pXfxy02HDoQNiNt8f1eFDbAy4n9X4p9HiQi7TXgMRAusqMYu
N0WCXuDmxDF84gUusTowvBLyfRQSmjTnV/ciZGAd4izdk0WCyii5/uxRZ4Yu+wbfz4kQUu4t8dbo
9P/imEWeC8Lwd5+sR2HVE2vrE/x5UwYw9NR3b4/JuojRSou13W2VkWeBeJNXdSwrVf8jO/wPKqsb
KPeQ6aAGZXgaf5bKsZ3AYugCsAq++gjQ+A+14ZaUZs9b67RSm3Q03ejCv/L0RuSgdPAuuxujiNkS
//+JDkO5y/RPap4bxWFyvzfs3wHq+OvJSSZs71D6wovz12ZosywDQQU5eKRIwpW+E6OK5MGNi8fF
W5NUN8KoF3MunEig0h1Zi44lBu1s1ud4E6z3Lm/ziyG9u1cV+T3tdSYziDdC+s2XYmzK8xhakNtF
fNiar5GHjJk7ssR6xcp6dPL4qhiuByZuN9wvsBgxYebUrHwVZwxRH6XROtdjqbwMle5Aa8GZZ6ZV
McGI10J6QhroMNtsdYM227qs/o5kBW/Nc0Z97Prq5wx1EnZa9GfRMquDGCcCxP4zI5X69RKvRqOO
nc3FuHUl1dUMjvTgM8Mr1xkJ1YiECp7F3691iQGnlveqwxURT1X4+8Xrm9mKtcBo+Tkofc5+tZWe
oPcht/3dghPgXUOGW09XIZHkzkQrs4gDMMQWfHubX4IWK7HWgXiHSUOMBu1FJw2ysLI8bcNf6akK
niGim/jX+LMDyN9HGoGSdplTwywE900Bo69QBW0xTb/KQw8wqTp/5807CDz1zhqiM0qBAj5f3v9n
4Y2Pt8A56bMwtLX6ssUCt3FjMH/zvBjTtqIbJ/0ko/bieyST3bbV/Xc+zyoF3NozRa2TeNsKMXMF
vEHtZJvX03Qq3VQw1JWC8g7TA+JkA2c97i9pyM9hX8XHhhkdbbyeiYetAr7cxQ4Z7wD5zzOXe9bX
h5PIr73pDMyIEfdzvT9MmmsKKOFmdTIrmB10P/YNYpDv7AaKhDENIQeIvbb9c1nf7h6n9YqVlMvz
vtNd+iJZxjPRXc/ySQjn12KMt/MR3fijcyPjZ+RRP4GmW13cPxfAKBeBsq+uUksxaP9m7kqLrVmG
2nKJFpuEAmaiaqw5FMjqu7/AIxvhK6BtZ9xu31bzNEB8lsinIesW7SYB6t16SEmXBzQiHwz60d2J
6/gax7nOJL59JQMSa0Toitk23JHfH3R5j32Y74oRV6Db/gsZMDBieyO5JLs+ndFCMuA8XJl+PTI6
e5DIAvkoq+08BMeyAyc6wke+R5xyNQyayQr7FVpVNSNlg7WSO6sLgoqW2+AGIqUIByC/ejAOqIoI
rjDuxkNXN924EZ4ziy8b1VmVxdurMgugeF+cJ9/6UBaCoMX85hvbcdUCqLRniCeAYlS50nfpUz4b
Hgp2d6Pr8P9IgAHvFuedzfvVD5XZFqcpKq5TdqAUCMDIrIMWukdITZ5wa+A2UKpP9/LfkN2J3a2R
NAiHX0SMAIlMh23OCm7sWfyrQNnayf1Yi1DI4v2MruV5ZF9iE9kjJ4IqvHbUZjv6CiiIXQDL8T9v
gOwm5PYJP9M9N/PRFtxEsVVp/Dk03yxuygNl3solZltls9rjM5qVchP0ZAgm0+/zAOSaN8kPSlMJ
n/m+brp03wpREnJyNJ5+nFpdXMksW5LbMZXSWpJ9Vt8YzmUVo+GDbAvMwsYxApedYUJ8/7bWq1fm
NMjtIJQht3rIRp/VWoUmHj4BDn5Ibc+7UqMQ3vDzzgUUOJ2V2gdHjqPdenCp30hydt6VyX8v9Pvb
m/zEywmAXcx4V/HsFB+XVX/b7zCXMzo4gzz37OYKXYxBqOYPLOQmiMg7SowleVqz0nmBVatJ/I1S
xknaBhkOLNmGZmMYanI9jqHRPHkezYffi/sPt0D5fztis5U35v385RsNRtnpm9NT4GcAKD8gneJn
O9H6RBEzb+/kYdd1KfJJXCwq32gDJucRLJ3kAB8+0yuCbmF0xDs7degxC88iQ9gsPpsskyX0c2Nj
1jWKJCIqxawaua2MFmvW+DLjUBLsRGxs/EUXmFoamPSZszNEyd0zjw0BSq1arCWMdTAC7HoxR+aF
Qbmqv3aim5OkUTbjq2I2IQrKA+OobU0OTXeBCvpdko+IwHx0I7y0PNq/7wu3OXHLtARApzCn2FHh
zqa/gnDw3W41acZb/XohBqfbLWGBNlM8uF0xRYlrPPIvlg0i+4TZEyDVlbfL6rhlZ/+ZfqdF7iOp
QdSS5whqSlBpo+UsSPmkPne10zmtFGK0WFwLKF/LPO54C/wJo/FCHS0xa24JEHCUsFzFMzOcxQRZ
XbWn5Z1mbZ5yklhbqcalQkudXlnwGZnFApORMPZdbtbEQrveQqwv/i+8pgTcQ2dbIRJEYv/Cay9P
WYFqQqWMCHGFGALD80Ss/wbaxKpiaSRNZzxf24iY6e61NqlAcYBmJQEsor1sCoP15SnNvHn4c/fX
6W8iMh1Cxt5m1yEXx2Escgo3QoZC+hoNHx4ObZOVBaWNk0Fw5OYvj2gDmrcwstNuuVD9aUqkuNeY
mb/7D0/8wnBDjPyIESncFRbsnCnpbU51zg+RoGQlesWKXtI6W0nI8opELF0CFaDLhRdzv1GuJW0u
AY8I1NQVbBJ0atXip2r265azB+j5h933gRIRYru+UEqrPkbTMkQ1w3plgGv4pN008r8Kqvx+4kQB
YVOIRTDJ07tDnExIxlb3MOmvd2kNsYIg/bynYlWq1RldjFGyC5MtATX0VkALkDnFnSe7KIqLtEH8
i9S5HA7abQXGofvvIDOxKDRwoB3WgKDJT+K5XIe9kjrkN5u7strxWkwaq8DodGDnDymA8afF0Ujf
ViZUYEEvWUhTX+Df9NjTi6L8gjK80F4CtCsyl/buokRPFFJZ+qQSnCk5zjg+sPXShIJz53X8Socm
ff0gO5NaoApC9B8EhHIQWzFBJZgJBWvIEjcMuyHLVp28m3b2yHMIr1qx4T0jbDT6UVqh3aHy2Iye
i10uEXWh/Bu1KY8IzQv4FG623WdZJ1mq3/t5TxD3hvcB/eDWJtVEQHZW97M50PdeT3ZV7Wv7aJnx
BEYsH60UHSNnE8cTCS+WBm8dxoVCbApX30zxPGpwed+o1oO9PzPbJF9DKg2zAR4VjWzFky0XIdPe
6bgBU8z5S51VG6AW4jaoeM9+eMpKN70c32+6kSl+vgYZON9F2uE5O12azMTKe9nULRPZCaq3x3zo
nFVVyy8j+fTKYWBmpHf39rpolBdrs2bnuoqomJrpSbuKsd3wWtX43erw2Vd3UhOCKUrflNPmHVmX
oSpRMsKIjgu9d0OSZS8h+QyIx7KHud67+1CqhwY/wr8/mz6ASfgSIVQ0dpuXPLINS38448qiqhtE
TO/UNXqQGFoeHEkkZqcm/n1gMfb4lu/Vh1DgPIzoVwDqsUv6Ur0XT+77NGP5IAa145t/zufHFCjn
16XY3JugW+hDygc9nN5bgaslrZToBAO0ynVYAClbp58GCsLz1wFZu3dPqUsVHl3cRscwLTHM6K3a
A7uC+HvpRLkq9EbefikKh4V/4ZJGhKo04j11LD8dVRv3fkypSIFEn/Nwt8EBuFs3mbzARtFZsVNn
bs5C4/HeWDNJG6VYibcS7061716OFnp4SHIX2bAAxlvcnmgMZY/Jtm8CKEQAZtAFwkc6216kuNS6
6dwY1NSMdlF/XBzv0KBgsw2x9tGfDvQQMk0a/z1g/sikJiyLJd7Dn97se5LbbwpGTdPlrM1btaN4
mifar2f54ZC11ZzubT7FwuvSePIitnJV56iNo7VHfreKIQqo4Dm3cO6i3UhJUDrXZGVyRUPT+T+J
dEO4cuHsHyrb8eWnwBBR2sOT/sg3JFtVUJtgAw2znY5ZaXg9NWHbNzW8yx/X6M+C4ctsB46OZUbm
2n7J4wFh8+EBi1nFK701if9RzgniWpFL1yWr+JmfK6l1zDlzjzKk+L1f1SxF6UakLP1fUPwVRvB7
JocAIuCSP9UXbqh9rn+A92wvVfN6z1tQciDr2qpx2FNnl70qQjhVvNSOE2fnuRwNdLKHHKjEu5iv
9N4LuxFu7voGvJ58/inYe/6T90L3koQoaIuYpZTcU1uqe2AiWY7e+QUHBfrUfPxF2JnauILxghfj
coLyf1jYJUCmlhffS9jkTdGmZ5stS09FP73GLtJWu1ubw3lRhmqFx4kgOCg0dZT4Fk2E/JXWJSpe
KtuV/REApM9iKIFV6xcLxOoxN5pRYDNdXJD8GrIiMtrT6S+MPfsCH70P0+ENi20AuzqhBrSG4z4E
8LtheQt4sUgLaIb0Is/zlvLUoXms/n3dTqnEcZZAyswWIpOA7sLC4+JtlF74dCmvZ4MejiriwNqA
FOPj4vjts8uhQfK7btTtrZ9SjKDPpoclM9Mg+ndU6pIhMqLfW47zZiwDArlH+9E/geq3WHl9av3b
Fy6kAs+moNbODMywJoZ56AO1RJB0kZwdME4DDJUitcjZB2dGb/iJgNRk4ZNvB2t9BWUnrfunE3BM
MPrGDkFsTOHTaFKHkNzLIpA+wHN2YrqzJxPKJOXGB1mIQ1o/lvlSXXvEHmnfhsdmLH1EVu+seWTd
HlPik6pxHE0icaWHq+zG20dARJATq7WJJjeWqVqFNSU57G5HprfBXI5E8qv0oBcnmp5rZ9GPgd0T
Ft9/zxf3teSsQ1/YOKgROOfHvnWDGflP4H0qRS0PlKvOuwubVXZUj/1xp7jkBzyu9biyB0lWoPp9
Q2QvWhj4ByCwNmL0tGg2nEMsOASpayG+rmPQTR2dZ8zckazi9gmi14lU0jCaX/6weHAId0F7MVXq
/dvBmfCstx0p5MKhW6wo3PxdDDjMmR6M4QwwLBnJwd7uDt7yPlYP3HU3/qhOOEcfz13CKLo0BQLj
yrKLWXoEj7j3JPKNlrmiqTnQaRSEmnrxKZyzcdoiQvgGvQb5ZD2e3Dl178f15WH9NBj+koEF51kZ
Z4dwN+MWMKu2/2QdbGnSdc/u2q4rr7qR4I909qDVBrd4Hk1+U3wwLgV3CAfLvEvEgcNbaXB/dHVD
xnHJMuRNWAseASNm8PA4P7zFO75IHo8xeydPnJ3DTyG+v4McvMWEefOLK91n0igdH6iCX+V49SEt
RE1DqnMV4zdsUomcpszMgJwMP6k0k/iq5Z/Ahm7MwYlcl63s2fZL8P/5/Oa8MLwJ765qeeLXsFJS
bVxJhiMQwhKHXGLiWb+Bx8iZ2TBoh02u1eLnJrnXK7pVmI/S5cOp7UwtD8vDkYPW2r3D2ZdqbJ0l
xxF4+ecYNs7bOToE0O8D2U7L0wYX+tISC556FxnRo7NbGSO5CGwt8d5n66vsiebJQGhgfWxeO3CB
/hSkrvsGNQ7o+Y0e+1h/w33ZeaDpEF1CH7uSaCZ3sUJ0kSb6A8KNjpQSdwkLczix/7qfnLnY7laS
wYhqbeVmsJGlwIUfqsSakTNz7wyE3Gm26FjfnitAWhAmVFF8esYSp4zVGs8+aOxno/jV7EsrSRUG
zNVDoVtZHeh6zFhHyj+KPC8dBGyUxfPDCrjobNUaxYL1shO5FtUEamgT/jEgXpkOsaTU263QyvIQ
O4x0T+e85tcbKaU8YVb4kapVwvP0E8fkgjwrZjmr1VsRmgF7p3IoRJOT0qKVeIfhotEwXAeGLzmr
34Ymqrk3GfjPVWUzwrA/z5dp7XFUaKSBnq0XTVCz7hfwEG38pLpN65ZFlKLXuXjRhzBLz1dDvjQ5
gu7x02KEE3lbk+IHXDdfhzfTPEkX927h8gdoKNpN2sDxp8GQS0MCBPjwFG/28T4qf8ZIDfeuv18M
3BmkycdX3nbyyOaQlGOq08sKT7atenxSx0STL/f+2eXa+25Pxt70CYmwX7ez2JGTtKuTNk+gnuvf
htyIydyIxyYsPN9thwTBqSzgS3hbVFKkzgJQnbiheKRCvaJEdPakRz2P/ZzoEnv6LExkdhBpenVZ
guSGef1q7KqJQ2o5SiaBz10gDmPyuERbZbeZIFwqYzlg2Iu+JeosOE38xmu3C7F6QYY6avhHGLLp
p8Vyv5xPMXBMo0LyYJk5v7S6iUr4pEcmRCA1MwuSMBGN3MAcErz2ty6SpWvauNRZDQU4ID84ohee
RFIATuA/VVlnYIp95mH9UmFsYctaxsBeoMm0lNKq513AJZ90B3XRZERMeuVMHcCvzgYURixoizMy
uQyLVD3ER5lEleSbatFPLYzBYpuB+ssdqL2Byp2+q7YLedul+uW9p4dFtugsRKX1X8xpmrggh7QR
gidwqssw5NMZ8iyeZnTSyHr3t0quXHFRAGomK1qBJOPtNRU9qzx8cH31XCsCygM8gZb322fx2AaE
f+3lwIV3XWUjZrgtO0ngSg0SEJWBltnIfnw2DdGBNNEILY69iJOuyyfT8Q7fUEIg+IHBmlylSKeK
ZTRVRkXnXH1D/p8qDIZ8+HIjuHYE2w4ScShRel0/Jw9obCrpgnLSjCo6twNYtpgJQXEDnX0lJx33
/5cxB0TJH5AzjwhxCdfOWAoZBSaeCzsCU2e2LqjfFbsPYdWDakEkTWSC00Hu58WctGWXuOFNcIee
hlf/yopYe5RNJAzKQOO9FsXvVZ4eVlXGeqDX3rtJ9xtitujBmcWic/a1A1zA4neTPSlSPC4nUtTe
9wJv5EWWsMpdEtvJh086iHcjHlblFRkUUTwmMlb9C3jGpy+2feWWLDu3LoEiZh20zRVsV91AjXlf
DjTzAsyO/Ro5w8gtkew5vhsEhzKyPO4rCxAxQfiB6TwtvKgLlBlo/+p4A6NA01KbqZ1s5aH9skic
TEsu8gETzDLScd9pgqhSRrcmXHYXe7jK5AgGJQ3AWhLiR/Hy1wq106bA4+udoMS06b9ixeJkbP1U
5awMN1fV4kVYZ7/CTwErJTjkPbGrGH+01zYOSky1AALl0li1cZu1wjMVyghFiyI/mu96Gu7//eWC
jZi5/olI+f2VDJh4RXx87CdWAnlAa/or6j7QXWzmBFS7FHJXyZF4JOGbIhgCAisK5csQLqXVVO04
wJFDxgB5mAFUIQwos5bmLtzQyC/Jmlgqb9FnFfq9jWcEbr4yUIQguzZ4560ttgR5J89B9y40t9SX
E/b280mtDChzyQGUZn+lWrba+/PgGBWJhm4//+EATnk5V+GaMTipZHzmHqs16nUdHcC5xjrzIxsN
iHER0ivLjxX/bVa7xu01YnPFF/MyCCfE564wSNcqfKp9TkKPpocnZsEzyZoTdYt2wAMgaFqgfE8p
dfy2rMzKNHTfjcJNLeF7XdWcFEj4trD9vW8swgqXxJQmbrAkUHUB58MRvGZWHB+SP9viUrbTYZLJ
VqqlRhZs4+ARNR4OA+bZ6UuNvXaq4yr5HmzapH+sdVuNxR6EQbDnF6JNWchaQCmRZ7sXfaxMFlz/
hSfWSo5h0TV45uwJ+25oLLrF2StRMO0YEvM1q/4KhyXd8d76JJ0apRdiWq/MdZ2t1yfguX3gy+43
5jLWMzQyb+FHP5II7fudv56LRW+WuuksYuLXQWbQ4ME65t6sLNnP4bDVCTuOGL+MTII4Z6G5GO7O
tC7k94gIzUlH7WXDRHW1aoXY/C+soELtKxZJkh8zc2S3KoZm+Yp0/qiu58D4WgzXgbKw6pKznCXW
itK07jc7tSoGouVEIQ2sqR0ylbiFO02KPLbMTrClhz3v7m5sX88crp4HShLklIIJRR2H7k/Fn2bn
RkCOu+0B1c7b57uhSXNtzhKfCCSAFSH/0qKC6lrjprggAMAFBuAVG4FYi84tNkvWPlVELKWEbhd3
U0ePZx/D3nikEJV3pbyNzM1vUiEWH05bUCtY4TU54mLYyruzErPWELnW9OWSJIvYrjzQeZEgg4pI
gtsll+8DJeB6Iw8og85T1d0n5drB08d6At2h2mVQSE9jDijpV5yIxBXcoNySgMDixo9WopT2Vfg5
V47LOA/GdaGAWx78sCqDYEkGDnRgT/XmQwrLax9KRNWShYAtdk7uEvVTOq2UaZaLsfzDPwOD1/IS
CQFT5qKI6oAd+nqHfmxqeFogZpYUahehML8fuxGfqs0i50FvCV90813y6EV0awepn5PgPe0aRIeB
GfKhnoSEVPMLWsWo7yWwTX7Sn1TIRnOV8Ultqf3729QDgUgWK3ZsUw5QPM1Hfx+fpNSixUrLtfCH
UE7VRs+eJ1svAvZX6pdAgSMS84gYGNpGz9S7hbZmbD/K1PJk0Ein36zMv/HMcHmOBqUXBHm+QTiX
GcNmsacboEkiVyFxCLoItgW4dkQv1aIl5GBhw5HYg4UDOcUBCv6/c8RKFSz+G89C1BYJ5sFButes
awcPzB/Iq9tQhMI4bgOLTD35Wo01yO9Skp8Ttq9e4IDrR7l7rtP+htSRHgwg5cXdZN9H+JEj6Icl
Kyp9GWYlmmjf8L6ap9PhM9ZGreh+xtz1xP2uYQuvmM3zGCuIsqXPNjVcWQOMxClMZsMiodFVpbq0
/vdZZrGtk9QFIE21z1QPvnbPUDo9a6BlhDIrJ5gciW+o9Ra4/71y3u3ZoToRXhxGY/hELfSdMLj9
88zVKkECHvA75L8YZW3tIJObgk3Hg+rXGhwS1pJZ80MBNqBdMu3HNM9RTvaYK5DE0SNQPwb5jMec
H7yNmm7998URS920VIvdcxjyc4mxVYRBUhj6aLa2Otl49ed0CJYAOqXB3dCUjw7VHS2zUuvBzkc1
zMtKSe3/WAJkmQRImpyVeAqHmpJRG3u/5TP0sDZTWHZFto1+4A8gRtCfaU87lNWpZfJVME3mP+jV
qZd2LkJdu5PqlQQ8bpDGI4Xz2oWUo65hh1HDevZ0tgOWUcCPiMShXyAuE8PynE00YYWEkO4SUhed
obM9lTjcRNm91dZTF/M8p9+orxV0gTSiRPy4/GgSt77YL3B6X9EM/kFh6gqtoH97nWRtpo0a/Ub6
iQznwOSsWipasgWNlyWB0wb4DyBOQT3ihCs57mcDoz+acE2gbcsrMxI7HYU0dvVug2i0lD4aNich
233GvNaIjnhw6H1RJDVFaU+/t7o72XKlF0/M1lbGarcairc9Sk6Zf0n6CH9QieAc/kIUbjG5d5Pf
wI0Keop0u2L1sAMKE/YGLbvr020H28WP1zwNvpb3WJGfw6IHI1n6VmgjJ5RQhmXzJlisBsZiFbFP
syahzp3MRfnL62aWA+wo3mJTedsUi0iMKi0qH0I+12ZZKfn037BpoVted9hdl6FZLNNo7XMMIzxe
f3UAg8AVKJoukMwGaPKJeHqVblQS5mATNWKPnYnvtyJilKLCR+qVBA1E8eTZs3aFUW4+cBQBaQzR
qov8787AffqdtGqsV4B/wQyiFb2l6U4qI29nlDW1I1rpmI8bpvBBwohvVPNpTdihPDTJxElf6m6z
ZGOACbuSRsgJY89gesa1wfATYGfKzoKY57n9XxrEsLCQJOUvGl9rdHBP8AK85tw9V0TUUBwPs2Au
7ce2kaPCv9xNXgHv1aE9aiDbc3IjzjxyccmFzpoKAE7A054qtncVh9F25U5qN0v4/tvbMJHlrVVO
rfWk3G6/AKTE2kFamHJhLtrVfry66c9zjbkrGRLAK45Y7ukJUSSWpY9RmQxyA4b/iGfsrycScVhR
rPmZX1iRAYvvqjhLfxyS3IXyTo7B0LCVuIJqqK9ZZSX/ScQmDj9o0lGGNn4K+1zQbpZxhnkafmuV
eOQoql93C5NwfYqcVJAI2GEyM1r2hNm0tsCZO35z9AU7Mxk0BH8Pq7Gsj06XuPzwKBXH4pgKRuEw
4BxkOpMm13koFcJGrZgXk9Eje5K9ce0838nm9cpvFGFzeDd8tCfJm05VTdfyCWecKRMvPtHxiMDp
hTye3MR3oZ2a88cLMoFNvhDiQAIKkTyPKr9rS8Qwt1PsmsVg5utA3LXuv1NOhRLfpo7sAP7XutYE
YFPvGvvBZwfyGFxbL6TLS2zjogBUznQaSGzESsKqhBD7fo0Li0ZYYR8bMi0llJO1eYoc+XPVuqIB
5JxZ8qdgp1Jf2bDpu7VB7icqtexsDHeLEnhZgPimm+mcy/AxqcNoatd60DQxBjcrO+gq+yZHvdvl
xiaNX78/mTOddTYbucoyuboQCavQJ1W4yWroZPr7hCWQ5ty1RaISYTBdDXASKEqB9fJGuY9Ui6XX
Zso37b3x3opxaFVm/gDsZuVY2w3khS2yxw+NXjd5inIKhk68oiyx027K38YKZgW2Y9NQ4L/y9AF0
KdmzZTpaR20PtISZsW4t1fpmfAEcip0N6e5vgGhHpv0zV3g2+yx0gbD9QNFigaf8tOVA/aJzFsl3
KVKGwnd1wHmKJ9knbtAqsrV93wxnfDzFGIXmfHSqM7bywDPfJbGx2alMO93Dz1gSyul0Adzm9pig
D5zqqe767OC/duETMFfVghLTAYlokbWYzur2SyEKhmrrn+6UhBmKlZ6BVbyhSUOu4R5dOYhLiYi9
PjLelA/48eCn/icGw4epXF8bmqjNNC6DCdFAXeriQ26o2T12Aa0m4UKOzS5NKlJmGWWDHVJPro5C
1+zoS/4Ez+2sB0l4v0z2xUeHMjY8ArXIt9KbS6PsDEqJ8C13OPw9QvgHvDEpkVdFqANJvXxAilef
B9I9kHdXUKGMCnwmbIYfSa7JWyW1ri3n8/+7HPAyyR+Nqd5qJCraPkGn72NM0fDsuuT8dW6A4nDA
hAw+AJIldSBAAXjyVHFjzW4ze9kXncECNBCIlKrygRQ9pH8fo/BqhKM8AQnKnUncLCi1FN/dmyr6
+FwWP7iOFrqqshTA1611fyL6xYl4/OfJxOhK0bGufPX5sHNF9kI+xchd1sW0PZJG/zY5uUfG6I7X
IHmi3shyN1d+wyX8Z7DJtZhYcCdTJmsVdlycUfUMnS3OyJJ+7+WDkvGAHQRvZ0ineMO7PPrnbqt2
9JaGFXG6DG3rhQQZEHupCRHNIQ1lXLffiV4Lozc2UGwrrr/XV9WRTfmvRdTJ7HY7dhbEpA0QFB13
fT79/50aw3SHg44h8QsKqGL0uA3aZR0zUjjZXs1TXnAr0islDDOeMnVeYs9LImJIQKle3e3nTqlb
IRdoUSNkXTt8uSByZ4s4Z9CNngo1QOQTgaW0/FmF5Q80mj4GNdZSNwlaG+OVsncOfGY9vUAqM3Ro
bGYzFmnOPUjPh2yZkI9LxYXLr3l13H54NoWL9BNb4Hm3YFEeW+ZGoHp83Ctzl9P/l0E5ev37Pf1f
k6lH1skky9hr/JfnusznC8rl0Rj7RfUVDLoUFJnvcvGxwqp7NloTDuKaOK+UXLzoHTLG7iIag7WQ
j7y5ITKGAa97TOKlrtVzJim4DM/7t0xZeslDpXMP1QhqQxvZNw+/2Xv1NrZ3W3BpXy3kSZN5I2jW
V/SHlUA38lAoTp9RQrA0N7O+r8VxTeEWqA+cjU6d3qjWLCTmrk4PRshXVe3BpFvztDsb1KnegzE4
kuPwELlyVB3mMD2szAIKWrDCoZHJveVMNiWxyeG9pF04M04Jo8ELtbIDTZpJ7jXp5Yci3sAdpaRm
d/EvO3+w22yWENdd57wucUfw7RJBpdJBKG+kakgIKnflDb7GcWQtFgeYTlReSLPlY+yh6O4Z3utI
NshUHXRg0N+SgawI3duuJPxEXO/i4E3tEuOXfPoMxMVJ8Y0aZhHFdelVlHbIlV2yNNFOoU430wpO
I4CdU8z9UyYDbHG1Q6mRUzDUeIwzKhbKopA91/InUYYz/+nMSsDr2/alCcK5qRRRIpLkdaHE7dWq
QALv48WtiTfgBB4XZ/jCkdoNQAZ0GBksyKvmIwGYUQlwWOhU9GxOTyf3FtYEtJzZ+ej6J8YDotdH
zjAP5SAnZC7Jiv8aq6+660QlF7WWKLWmtJuZ6YUbC5+dbSlOGjumXdS98MdqjvoXtNjGjJ1+TLLT
v3HfjHtstNqHuvoh73xKYmzMa9JnaCXsAne3oZxEc/RJW/CTW+7KJEG06MBpJmPLCLmzebkZUh3l
0XHNm1crTl0Ob+YMrT0O3bI1iyG7MauuPVbs186JIunXSgYiiYcpPcX1cDu9pw5dncQhetLKMBFX
F0uu0jHuVOfjKoxkHm3b3QeJW/7C3U7tpdmcMrmwhUIt/7Sv+FxwkLGKb2jN+E4+kOhX2m+SEveC
m8n4FQ5mmrmdfhBW2m4JM76VKMmAjwTK/rWVlygyifxVfj/U3Ue0JWunAp1XwK4Io13OhDIESAYC
nA5T62cotk+bljoVzKktBzYUMfYZDtOwYDCVTbos/khYsYBQoT+goH3dcOYPiVDt+Qio872GqyeR
gdlxc81/utoTpIODnfImUXV76s2sVGRJfJHlPEmsDTgYazMIjUbqyt+HRswBz99pg1FU0diprySZ
UXwRpfwIbUcBkus7n/lEVnthelpE5Lh9AwCt0Twfpnrc5M5mV316F6QedDZiLrwXjzmIhWkwFi8U
Bv2oVtx4oCDRTza44dGEgmEfWV2TEuBgZmCCY+B2WoAADhbqkL1LF3mI1R4DMBwfiSaY9Y1H4Tm5
Z5o8Kts7tLZxfrV6KsWrRg5hbFIeG5QL2VX67WmBR5ElKtn7qSYqs7I5NeSMZk8q/L3mzLXzN7Jp
m1FCkJCgSG207F/rre5JVl2fHiN8kiT4/3H7ucR/7O3PMS5EpptsbdRK4evo0eX+53HTTMjcG7ly
8tMLMAXTPnfrUFqJNHgNGK45P0/jWVnSI9NbscLghaEDxIYDCF79ThQ5qHT3CPvpgG7B31RQj2n7
+pW56Cb6nVXmso2z+AQPXbJBvx5h5Pi22P+fhFWjPxDJq4aEkXs2+S5pwGCqurlKpMyhnQbTqBpM
ix8XufRvX8hhDp7UafYEh0KkkY9nvUIciMePg3hyWCp4yLYyMXhs1ceXma8EN7h545Ln+Ckou0oU
WBBrXRaqIKEYD3iduJ05uD4oQ7DqqYhjI2NpPt9SMmJSPsg285nBHAiaGq/e0ANuxq9ciKSupCAT
CeKrdMpoEZmHse2dG4JqAXTXXs9Q4V60Tgkgode0g7IGjxxwZ4jRTBk+kMEBB2Qst7GEJbfgz6Xg
WvUgmi1MaiH0FN7P8p1FZ9z3xN/HXwL1KKTS6iEGP1LMZdzBmQg3E/J3Eg6dV9HXdtfIPxP7wL5Y
AYBQ94R67ZN0YHIEYj7BePKo6HuLS6DxDxsn270G83bzQnjZxIwbzV7/FJm4Xfcf8HlVRxmRfhPv
Ey7lHCeKRLfxKn8X508tK37mRJE/dPllREm8KOqPCii/AQMSYCQrfNRHZFY3u1EYTeg7niTIIroP
DtCtAEQjVE6n47ZfWSkyfSxudSvK6900fkm86HM/NX326crO14dPHaaLrgiYEKscEu7ixXT3AoHo
WPbYiCrIBhhtSrR8N9S/5nc+XV4Qy2TN9hFNxzC2HsB5lAIvFGto8wsZQlFZTy8BLEazjajnwrWF
0FZgNKPkBu8O6O3iuhfHuNw+6ok0zwy9qJ3AO4y2I/aVbCNgwILSQbmB1tM945XV8GY1IByqiHIN
+29aV9t/L+hoNCGSdUV29b5I9jKmR8y9PG9tVqYFecBpwJ7bAS0V2XUq7IeO11zrUoVfe8dqIUro
qDKLGSmfi25wGdwKIeCAXDD5o9oj/0UWBvN+ULv3a5aFKJAI6AidMpYRNPhLAEbB+crXQPt5dLyQ
4ggPaFnUCFSRb2sDgd3TAMTyNIX90XoTTCdCdFO+Qh/KBT4H6DH367cmODbeIxut2WHD8CfYr9mp
qJSCVyExG7bazjL+NSBKBBVuR/5KI6Tq27A9ses9u/As9KzNd/CX+u+inf90fYFlof9SSkQ6yVmV
I7DSKGiA0nTBFbcL6Ve3N5d2IsSP0ke/ouFrfgenV2OBC+Df0YUwjRvY+YuBqLNGxHwn57Xr0fOx
2gLqr/foXAK99MpQCI3y5P2DV38foFJt2OvLUwnvOnybP0pwrW8PX870NkDB6/OG+jg2PgJWr1TJ
hJowW5y41L+DLfw5dPBLDms/1MkEKc54wUPxQ1pRL1a95yDkyY0T9kriZkA60Lpr/+CrD8FGw6jq
p06ObbqDd+gGI131uUYc/KE3ISj8v7BHYn2/HH7inbRKhTmc+kBPd4a7GG6RJUUHK/tMYwD7cAaP
G74BxJQ7KkA1mUgAp259TX55W+AqE/un9dxFrIezZIPAjlZT04j5q0RJqgkgjNo0iaCslfqFVW6O
FHwt8wbytYh9MGJqajFMMpitkskq7fW7UI23OAt4mEn7Gj1Rzzq+L3ln9geIDgGzFU5cwrDdxU+N
GNYfYlzMWKZp+fm8fJgrNn3Q1ZvrIV37mJqXWwaPu8hxZOoAbNolEPDAAmr77Ily2f4m5pDFlb7F
Y66z5cGaIgzZTPXNxk77fRh6kIJczsebYDXI9TiBdHmGwKhBwpkwo+cJTPpzTL4TMZ33ClqRpUc7
QO8t4GNFHH7DR0uYKkqCswASbZt/1lMrXHXGpWx7dP/rDZ8aNAlwrpLr0oX/amvEvc0L0vUMJbLT
DGHQ5kn3tsrlVBaaLBE5tpPgLomVTfENfMC30vEQeTJvmuiz39OGFyrXzpLU3N3/K0l0HhHtRgwY
wiBUvh3bonn9SJd5bHZ34voWIrAWGtve6KjFODB80VKm7lAHZdNT58mwRRyn4Ej5dH3lkI5TlzKg
eMsFuOeL0xvbl+2yYxgiEjJFE8BbbiMy73CqYRdvrs/HD8sVtiltfMGMf7FmU3h/qJm8hLjd02OW
TkE75tfbnbBu9syaWJEWsm2qEkqa+ogJEhWhokhbVqDXRRDcw5Qxvh3L6V1UwVGXSmXNenGmU2EY
atrlYCYzmGg0Pdeqpcmniui8AjaGVitCY514HY4D6Yb+jIoMcnKWXD9Xqyfodwrqzwi6oC+WEKzI
CVvHQ5xU2iVGwhiyr+oAXn3kzXiB6EeGUmkeNX8IV2lkkutphkUYpL69BSic5U1jeH6OdSEH0DiY
FQBHm6rHW3dfjfiRFiMTf/tGIJVaKJMIZekqFvF1SUo4erW+bgZuZXd3co2JlX5kxzeY2i2pv6yi
fR8r3JPUeXqCv4J7JVH7cirK/OnJFEDpIe8jaOZAcNcMdllKbs65R7L8R9WMl2JNb5fgzfhq+ibO
g1/wFf3TXTF/e6g3+l+p03cUPJ5YiabVLIAb90bMiJAIPmmYuCuhxWmgDB/I9B/VkVavJUGPU+up
E0cffaiTltNIXlFJhE0m7DZPcnibDAIKZZwcbgzB3wRP/nkSY83ot3gej7m0/GypGAcGMJAabHJv
2af2n3Q+Q1NFtrUGJEDOZKIn7WV+cO3RlfzafrTlsSOJ7GKeT/BREnCHoJudYq85xT5dCJhBuIlP
6IYihljlMOYxm+Ya0M/y0ddgmQZ3cgESkpePXL+afYe6w5g++iwaz4814dm1OWHhYqhih/TsgbmH
Qoh/vO0oR8q8CYhgMAnMmhXWZ214Vux3CJldUeo8XR9Sp3j35jrYVqSyF8zMobp+HD7H2x9KeBJb
GMBt6LTrWzO4wOiFWmVGurFXWw1A8/ifWgIB1v1LyQu/FXxZa2O4l6Tz0J+gveYMwzhyrOlh6s0i
W4Rlcn4D8UnXxe8Ag95ICCE2n2Hkkp0tRMX5kYVB6v8inPydXmr/bcvwKpxYmpKFTxnAdq4aqazP
zGuRZd7sUH2MFhkxFaY/NkbzwvLrTyVdiUUnLCDbsRbcPCQbqaxk6D5tpPHCP3Yk+Ro0vTqia9tr
p3qLV7dvl07y5f8fIfin7VKgGrDwiPxFkHsLP3aSs/ZzngZETeCHXW7uIydN2HcVByGuAL3cmErr
KMGNVSi/mpzIDv/tH9y5PnnoShRJwOSrfg7UxZohIQtCnuk8A/4jHAaWteF//YJxYLwEt/3Agm/M
nVBxxW6aJS0FuLODjs/+VAcVzkkgnp4umWiOf6Z40p1Au6n1XBU1ryVdrNNfXppbVTqlv9i00wjh
nPmYO+jVsbuTzQckXTtp/NlosA8vFPcdJdsILYSLWnNqGAZNqS9BpEF1/3nN40KoPYa/aoGboT3S
kWxSvwsVNXTzcaEBspVFITRE5pUnBmX5TnNguY6IGJ1V/LC+CcLb1nRqW2aXJfHFatxVkusTzxaa
runcTY4Fn+QhK5WnTHwCYRFurTkjoBMegYyNil+SwyUwN9oadrgIgQa7Pc8n3TrreZrUqVjGStbF
sVLY1rXLj9B/Mr6au2m2L3riF2Nu4sb0IPiOO4OaFmWV9PrCeASXZNmnC85EwOGZF94DLRVPqjbz
tejar46ykvJyxXXwEz65EdbkRmQZAgOQMUeZVqV8b/byIOb0NTApmVgXHVJoz73cG1tvpfueyDae
fsnjrSISSkH4HHUcrEwUW2KBzv8FORUYSWi5iIlWb9/VOwPJrGTQNiIRWDyiy/HNVhSqdhAywFf5
dYnjBHLYH3fGnw66UAW7FBTTcPcpSOT+ZcY85QAdTreoMyE0hpAvS8U3wqbskp8stGicQpt898wU
xxE7d944epZtcQZFxLYgD8iypkQaru8XB8fqQiswizXxzYs7bpSD3gziyVFu9iPvT/lBaOmtZXB2
uTfwqXLyXziTWX+Plj5gZELvzfB7A37WTD89L2HOeY8ric69KzJy/U5a6rQkXbrfJVuNZxE1xpd2
L/ImKxsr9DGG1AVCdHVowQrQHHcnc49V97F5DOTfec7IROniRQmSbCKlLEiK1lkg9If2hS1+zII8
yFAaedFyZ3rpo5jEqfUnkMD8L6kamBVkzBQE3FlTzspwQbAi22IbSe/JFa0i5KdnNYecpB9bu44w
95eag0ftrPEBYrGhEC1/eGTihFizigxH4IeHzTHSA9Gyx4tF91UizfJi/R0kOfMWhrb2oPX35hqa
11ZFFgYsKbA1HFk2apyg84JmEkSku3rhtc1UIVxbSPIxsRVuLsHxoou6GL8K+aPJCV5xo+NNmu06
SohrIRogALh2FAEOSy6Jj1vD0qrLS4LBwS0uXLukanysDkjdaoFU+OwEDaFzd2dgolar9SFfOEkY
PBv7sn1JOZbwSMVXmxdvW0WWxW/PSnCNrSy5xRJQd/8fA56EAFgGEdjxFTnAyrcNpWueYayqpte8
q73YOrormhUWg05ZsNVrtscwvsTpXp2rtWxWEVoG3yn6L7w/KStHpNyjcuihdfzb0B/V3mG0Kdc3
Y5LmK2WqYClCunTTV4gTtqP5Q3xxyzlMOoMI9l5CAl9pxxv/YHRnA+O+8dGJLikWF2fnM8QB5Lry
ajpibUAIeajJJ5ZhlzBs00FPMvBIMXoCULE6WkTBeDqvlCEq14medYPBnSGLllpR4FAogqWOCBGB
odejaAJadMDfJxHJ9TBbHktzK00b5P7SRLBpnH5fFmfbDMO7ebwAF+2VveMcKdzrVGfmdw9A3RrK
mE8Z1BjVaQVmnaeA6SY+DZhUiFqa+shfm1aBJyGAwVBwtKfLstIjufF9vfkvqSC8fyAwPrvEiFGL
zeYVS/5sOP3bJHN6HwXOxibXNnoVcpTO0h+/WUqXSPRHUDxn06tukaz7mzuaqsR1ZUBfBx/lTCwY
Iwsp1eKdd6EhcUZTB8YVTq2rS1Sl0aO4b+Xz/1TO/yLH91VzADLrOSffW1+gHlohrRM23EBY0RX+
dfKKNPlJlVSLqAukQDrQZc5QpusW0ZDin+x5YwJ2Bi4MFg98qFd+ZmaEgSNPrwcihOgmUFEAl6eI
J67MNcbheJ3Bqg148Ts50Tw0jkl129NBJkWSt+cFsXITXvg+L/AW3h7yHNn1gdTbbt0b+kBHEASs
mQCApSCT2Oa9HgTnLl7MyTdcTcrjm/99XRuIfUAkJoWWfNYqqBzQ3zjdXwyM46TA5DzupCzSvaSa
BvBjJ6W8SWkDab92YQCGY+I+HHrIWE+SrSoe7NgGOsXRRfNHuwgLocCKnS3W9XU0M/lBI9loGKvt
yZ1vyvLRxiVqnWJzCuj0ADxR7cwy1UrY2/BEz1IPmlWjBuD2hznDvKkWAIqZywD6ctj+oQ+lWWbl
reu5H9PdnmRRna9oWDeCSd79wXgpUrvtVawkuoGCi10Zum7S5CW7fQMAn2dKS9dsd1YvQgwhoouP
WcvbGsxhDoVK5g3JxyESbCjvanrm+5Cwakl0urvQFWpTyXm4mx3qlhZRYoUUBo2rNnQvgguwCJ3C
+/lOX6P3nsezYLzlPzUB7kQ+Bduj3rpTwtZhmfwNNjEqrlbK7k4STJYFnWOyyBt56gPgqa86H5pE
50/nKprm8UTAlQRucxTWVw4OliZDtTn4+prJlY0ERqxkWDBvt6lBE+M7XKaek5GXN+C9dI3T4lZ3
BG6IPDND8lZs2GQaQPLFFlJG8edZCxllnkSAwSFz/u4ciuB6E3jvxqCkr2sg14O+KB6TXhvOMCMG
GuIIckCXzPx4VnthdKt37D0CqBANqz8/RN92g8jEEl8ZtapSqQIYkng5ZJTmZ3c9LTUX7CqHXU29
rWwj71BlelktpubocmYmpGo/3k8TEg9L9DQQRaUpCnx066IdDmaHFs2/eifTySaJBxABwCDZM5Wx
i6LSO9FPwg54VFhyDTRHIKQYg1lA6v6KuIS2g5s4SQQseksWqdj1fo2dWarhBAobP/ZSyCI2nJSz
KU1erC4xjGDDYY5pIt0Nq+Ig4/V0oy7+6tLjQM8X4c+0zFiFsXhC+EbjDJb8Dz6yN2YCVeUvaxBN
6ffScXtr/p3DLAaR0K1xa/+9U9WJbqHez/7sKpgqJ4opJUstl+nk2xDcYa2W3MJRmNDbp93R3iKn
MrGSzjfVAZrh6uI+u9+oTU7kVZVbQYdFZfVqaTR9CmiRuJ8fHBa0MZHmq4DIUp6zoCHgKUkc3IoS
9MW7MzJ5xnk5lx2Wz7tbRhe9Q3bbAmVnWY3hqwz+8Yf/g7PmznSnJOXYXcBVv750R8W9n9+7oS0I
YtWzOA+urxc5pTzMH0uhqngxV3lmMrkxQlWIFuxZFR3xmo7xtoi6GRR0KYMa8tGvRO7to44w46sl
vhrdi3P+MdGsaKoPc258v9oT0rn3q78wDgQ3LrlxxJywhOyOZTfd66NTSzSnF647t0wCECa/CmqP
QtMU0FIkumiI6mIyLumy12QRTrXSRx/a7Qebg3h9JBSxjhjgs3m2RYnUmEUsuq9gpbv6DKLE3ejI
saMzW9akyytKyV7I0Kp/DwS69t8L60vd828P+Ga2ohMdAxWqkdGwcZZ4sSYsE0J90DiKRy5LsyWe
s4Cgiyd0JgV44bq4pGgCCCvabBkpslneIBRksWcRxsysMGwUUuWJI7RP5/qOzHnkrG0KVXpvSkf7
5EleeeYmHp8pjFXGTvf6jbWQEYmaltlFON5tfiM1XQ5NSiuev7DbCjbIy/tRTY3jpOSOu7o30iiH
uTVOrvpxuuha+/IlYep4KsI9U3tmRRIk8SMi2bqlbNoB5TT96cDLVQgNqfEPjX3ndi5yhD4QUKi+
BRFES2fIrqxZH9J14qVorP/mpNtdpOfB1jjPIkqR2EMajpOXSR6yQimIAhPpPdh4A/457eTjw87s
R22s7FDCublZ97DNlNuDkRxM1SqO+xPqGC3rrnN1nVCtN06TQSkjq4YnSef3erydkevWNa06pY8A
y1QDkP5uvJE2WbiXGtqTfTWpX6I7xq9/VplfioG1VzqgItj1wjrQOpP7aNfSwb5cLh5WkFqt9OYy
TDOxJ3K/Yuf94X4Ihv7Dk+1ujiFnp6krrG5FKzOxio0InkETIt+Uq/bS9oPXD1zzmEpdK6ekv8fe
XQEZKD4aSD0ZpBR/qGRGYTPAmlsk4U3PvC7KP75n971dxMdyog1GD84dnSuNr8izT1T5HDjFOWkH
xlkftnlaI+tvMd0v1JGjFkdw0AWklF2dntJu3V+e/vnOlkU4VijobkWNnS3udroflPKyr1HVjcdn
fLGRK+4KYlSicpUjw1YAp2Y0mAnwdWyZEezx9Y4K7FoXNUsd9oXAQDa1ZSNRjHd9F1TZZTTwsJKI
5MmEs/Hba4axogMkARVDwB6tssYulo1CTNX4SrarN4YsXfUHX1z3BWYxqrNZza+EQ/4/ngDzQO0S
3A0W7GR3Kvr/LHn5v74uRP1GyTd2F91+O7VjuhNq6Jn17rdHmhh7G5o9ffUhsy+pDGRBscDc7zDE
0QbIQCQGjgXBdE4u4tlXysodQLPtrpYRb936VHknDBQWVZpfjfMS7jR8vNeFi0R87Usi0dEbql97
E8bcDPq2v1cg2DQzljEbqq4ZcW/72Rl7sReUkYBwTcW3LKoc/moZYUSTmCFgWKHK5dYSx9wsizgq
VM+vWTEGiajd7ZeGwvNDYk+Qj8Fi58W9d/Grm0GwkibEFRSGRFP6fiZUfxXC+BDNoda2KkNjf0so
U+ZYJ0sOW6y7EsWpJpx8hm+fSWQKyfsWT6cXpvccurp6ZDM5ITU5DUfiZReekDQCUMtgb82G8vZP
vGA5OKjFx0Dz9ImKHBoA8rZp1vDG6uJM/+k8BRWk8WPFrv8xhGiVSvqajVPt0TEtI8+JKm+8Yl/q
XR9uutMsyp8hz7cZaZmmDfDLxeaLZ0GX6nZ5tjMX9VTvRZ3qKSPVfro8U2wleI9QXkUyVzCuEmgf
IiXUtf/+cZsRwBZQHyogG77N99qS9DET3AhcaBAJ+N9GeT5ZXX9tiltCnhygwdVKuyn5XKdOq3g6
lyTNOf4lzoSD5BeBv78yhlg9vMpx08cWYjKWFGYnJR0yZhT7q/jZ09v7T1gupHkVBHOtAskPUPhF
dwijYqBayPKqi4qrjYhyZOgS63KMxkmsZ1UA0U5/Uh8taM2Ds90Ew4/cavSo2oN/gETXE4mRFl/C
zG/PGrES4tQcUAKPimfTxk2QqF009ZasbGoBBNK8t6f/J0n/IFiv83ZbVQw5mpUf1lTYhHPYhzIw
UQ01x0Elf1wtpJsSM+f+DYgbKy4zk0blam50ykizF+0Geta9MdeyZS9ZuAv/FZWnzDxP6n2Qbv7U
T9YB85N3LxUYgPRYogWbToa8rjRo3woCxTVzOgpokM6u7smxc3mkLDof65DBBV4QnUT35ne3YVhF
jHwKVxxHLb2mY9CT72fYPW5kf+HzhTUKZ8NlCmECJe0680R2zhcLK9Br7RU1I1SE1yZD+6Kivmbu
n8UXgB2jjjElPo5AO/tTzzSJIlPeHIe0zjljGd5dm33O4bnUOX6UQoHX00lkU8Suhn7Gzvi7o/CT
IxhMe+oLVRHYQ1Bp5WNWPCPjRRoiaGnuDBojCiOGTsaZ5BkhgyTOxkGwQaA8KMuGdFrgBjR9VtB7
RBWJoFdaEKK9n93ys91XzRFA6qwQ3+rUizYte3wZinyi8hSfHwEkpHfQVAL2kP2f1Xn0fa1KsIza
oO2wNT+Mo1gH/6LRSvrrDK07LzpMR/IrH+ZgtON3JjcIYBh8dcTXJ5Lzg2kFp1SBdgk7iWMH2qGL
vGAZT+tEZFK8H/Ic/fTghhPc1b22W3q+9MQrBWYIgRBKPLgamoDXHVtxQtI4i7JXjNP5DEXKntYv
KBt4+92QcyWhcGC3KDkvR9qxOxW7HwbmTGHqjqzMIWRuOJ65HvzvfqnXN8SI4Fc3HUPE9gzMAJcP
37nHpkasbOiwlXL4kFbpNZHyUqATJ6Wdjt31+YkdiVW4Dp5MQ8x80Ovf+ivlvN69g/h67FrShMNg
HlzjShNc6gsLiH867u8Uy8jyLnEU8l8JBjhL4aAItol/qIjFMl+ccGJVZtJJx0IxnNnsy38NUoRM
s7ZoXM2XEovB99sRkT0OG1xhtNZrAUoPEH5s3BcwN8IKMraMoFJLuPLDsbL3NsCLPev5Cf+SYrYO
jXBdHUAAPxf+wWhiDLcvkxplwdMTvtEWLkc3+heyNwb/+wJN/5MwaQLliOLaz35sLePeJxz+zbEP
u66dD8sYiJ8Gf5S3ewoKVUB+mCLoUkjXsx/QcHSTllaXaFmBduOjxLfxPAzflsddjpZWqsQFKhII
dTvqpFsXeWRuluL7K/xVriIGkqekA5mNLkzbO8LbvDIWop/vXYIUHxe6CVdq3dybPeeGHrrUFNNX
bwXFZ0HOMMNdFW5KjgMQ3Cr6yxm13leWV5+rtaFefCdEGeOUPQlqluWLBXNnr/L+PoFbnFZW1Xqn
LL/MZWIp4LM2FzCPww9i8ygeUeHmNok3xnWloWdXbu5GIZ9P6+TzCGapNW0BJXyr4RvTMDcAwKDP
MdXHwjAlBhBdltev77lzs0TV35wb9M/chiRxMjEOwwYFCGur2D/UN9RbIUv0m+2lWZTFtEOpe3vB
zzZLEMqXbi51IKfL3n9IMO97PnPQQHMWdtLlDxw7b9PUi7TUQBP6ZDhCfrP8HZHeFyDh43Ku6x7B
NwHB5gKT3yniLitiMVtucwCaTlxPjCKpB3I8EJs11GSlyZAESd+lckBAbr2l0O5nT1+ovx+aNUl4
FnXOQdMjYJLRbNNWRzhpsvfpg+x0jc+ogFLDn9FNEcjkDnbRjscCOWIE5aYjnJLeV1qT5Yr2DhjD
I0MCXimCVpQNpjcWFKe1x1ZOBF3tTFSI14fxK1H8PPinDclPKqp9RgIURRCBchCcTU6AI7I6B6wU
gP1rEwc88nmLtjslgFMTiiIYGcBpWdh0yzS/pMZ/wK739O/xb90ze5cwSWx5qIQAdbXwpwYYnej3
JNPYFyWC3GWUiLXDNZ1vQ91ePCMy9lYtEAeNlqno57F/kdDPLpBDCb2CH57fa9bBjgHnU1qh6dzT
3F8suA1NisM75KisqQVWgDKfoPoO6icAXvPKneFykq9SmvdZnMJgpDbyOIGYyLlkmem3mWgoVVDO
AkyY1NQQGa0DyWYWFAs4jANa7LVsjq/HHchLJgSFX743lutY+V3a3CJOUSseRZJo/miCSuY5NLci
CJHiN/ezcIKW9RNbA89EcwsxbuH6SmPvFzs+2uh66gHj+eARcFQrpDQIjo3MaUK95d+/kpd37QWI
448V/UeLy5iyRYHrslX0VGrO9x65nLnf0QvS5H/fn13XyDbsw8CmxaMgso7hJXf6plcSq/mKXEmC
flHofI2R25x8Q7sLN6NUKnyoRPDrOQzrZupE777l7prUshsJxFPBEoaBNGsE1KrW89M9JD74UK7A
FUfT4wJ/otxLWv4CH+HiBEX/LHXSZMUrOqBzDBP+omEDFW1Pmzbn1DJFak/LIBnGffk0KOFOZvJ6
19apGlyAPxdgS8+y9Oaxxc1qSrg/LzUs5kPmpsi5wnoOzcHbJc4sh4K4a8pY0sGYoq6zDLDW+E+4
xTct11wn+scZMq/4zAyTM7ukvfI0ggGNDuKTHEejBa3kKIyYusx3JIsGk03WcpTPwjNTMs5ia4ZI
bCO9FnlEJN9iXz60J2H9nXXjcRcEUyeFKOefamuYxrzAqrx9L5xql61Vaxeq+RwDyfiITFmYNc7p
WQUJnjmv63FcagTvXtaeZUSdLWioqarMbmtGcdPG6IIsQYXzsw4ey8795bGT12cIcdYjgVfwVr2v
6dYci+CX1O+f/2pqWETJi6DlVILTbqeqMqX45YrylrZGzv+84M7xkpUl//2yb01JXeYW2IijWVgq
3LNZhz/TrCdMj33RyIsMkFJSXNud+fJPc9aMlx0to2qgXrh5Jvl4FaOQ6I+j3REef/l2fIAMwUBV
uHJSVAIkBmD8X6BUoxMmgdyPB6bdaBENMn0mKCGB+sHN/Dwf4xt4npdj3cvGRoIqMzjvfRHo1NKk
WvDZfbzxQaS23LFqsG6gUN8Gk3NBn//9MCCoSig+l2hK5HyxWwbAaazQX6r/akvhFGDqLlITdUX4
trAKm5y1I+0aLBERZeEIjs2uWwU2N2uFYIU90xlCZgl5q0jML5AQhf3ImuLHG/WL//uuMxmMOA1j
AMdQV/lkF76oWV5ckhBQ6YYUJmDaPK+Vlxp2Vp7JTLTzlu+BXQVBG4k3GSypmmq7rTKrBprpof6H
OPERGzZdgmTmhrlAWakq0vU/LXhIHVOA13dMmaqjWhTA76lg2T9wDW9/4rACGWhqlwd62nA5b2Hb
5tGsFjJtJf0GFs5tTxZzgLUo3EBXW2DEHi1AVFKoXDfaWLZd7vZ5bbkbBX4p18tdp8704bv7ldPW
oBZmPoyFk0wGNVRMHaymxHXHgg7Ym0p7ortEQWTzbHGLAeyu4jRX9/ajOuRGD2p0vnLYBS6m+i32
MEAss4MhUHhkP7TQ7ZApR/t+gRkN/SlnHp40UaN1d4Vbq2vVTBGs3VFqfdglz5g49W2c8PfIuTKC
VCNrdDJr/aWu2NDa5erslF8/5L7FukrHojnck2lvibVmUA03LYRCzyaJCQcm9a8XzUS1Axa/70DO
qTdi7v1eDx+bq4lcfcy75eb05qN0cFHCodkaoBpp9egSC70w1wfZzsIIbHMr7uBdN5nI4DUFXZrS
7zLK0RjgRVjRZLLGgY2AS6v/doXWZ6vOw9a5Ao1+iOL1HGJNZ7HQxu4PZ78r2tRcED3AvWSBXfC6
5oNy7wMuF3HtI5OdhElN3AyYIaF85OTWCiir3u+f7AYo9tHyJjyDAK9JcjTQEPW/ti0SecggOoSF
Tv10fGrT3kfHwH9T6NzTi0aU/oZa6ipV/yyYRlB/Kz6/6O7mIjMK8nYhtvslbsYrvUctmk1OuRPX
G1TBHbsDiqqUfrEjTRWdmJPU7zeNlC5i6e/EnhmWOHTM2vGfMSG8FJxE7zeYxsVHlWl64opCYTFF
VFDU9Obs/IrKyETAwlWkSmpPYQLHIPs7swKxaEUtBLSmjivei/C2u9ID4XYvmv3Qjm7HjiJcJ9HM
jiblJ4EUcy03S92q+Q8Ep7/eErO/2Rg4/nX0vfcNwZaBQW2/3BIk497a4BmFRA4gLYsOK55H2GjN
20JfGAF9mo8QNW/CHr5/Zk7rU3XGUnkJkJQQSRn4MOysNSMl4nW6jHH2Mv4hOCVZKkUSf5rdYVHq
9IHxoQuTeINH7v8SwFGKaz544g6YU9wN9gpT21RzyfmooQ0wYoMSZ8NJjoG02+ylbpAQZKjTvZxO
HZsuVt2Np1wuR98QBSfXh87KgwiCuc89IqtVBNn5PXRdj0txGvDqhC1LXihUIOpBOXBfI+Qk3mpl
1WFt7Y3BcnsgLuMnhn36ztT65nobxZsc24aHyRGgrhr/1yVNuqn/vpb3VebPxpHQPtdmNIjeg4N7
sIbEQdUb9pwt654BDx92qfeb8r1e44mRXBYIF3EfoZSouhAZly43/BUIdZ62c8AG9kHMr+4V97UZ
G98efJChIB64mCYV4JP3p5ZA2Q3r/Xs/zaSVZcCX9HITuHfbAvR2TFxt6UmR8IZelKI8Biyjen3y
3osJDufe2ZcAogcFsvrJYdOE7InLgxEeKvqp2apLPeP+IV/FjkE5u1JJsK0AI2G3j8rN11p4nsyk
CbDkSAkd20ueSXmFUUVbgD7IwvPkKz6LC3CDYtjtuh5zkDzwJ5a6FovAOGdNZXe6qji/RPXi/+sr
VfBRziyzFGLErItETh/B4VZ5XMksPB9vYcTcntAIMB+H2NtB7Ix9T2EKzRle0a4wgHVr1wEAyx/4
fowVCiq0EPfx1RXTAue/wFsIIa/Z2zaNnUwXWdcowF112lfs3rEAAWI1DbAX7K6Psxc0DQmdsWTl
vgv3fWcqvIRd0xI1KqoWvWsXz05x22DtqnOBcNCMcW+U8DDF7qY7dNmz9wVE26nGAZbAr7KdzZEB
JeFwZ9/tiW2DWrCOkRoHfyf/KWTaN3CJIXtmrXexBIz6aqII/8UIFEobOI976LxE4jjNBK91xe//
KxkWy9Vk9nOD/cGXHBJxpe+nKubCNtRog4mynpH16UZSKfsoj5+XE5RAm69pvZYp4NlFzzDWmwLb
oRrHc5aVgF4k6Zq4u7SIPIQnUo3xj8kF1cJWYkqqg8PD+oBgsiugLZtxTJ2Sum6soikwNXOuLgRg
zJAWkZzSdZ6zj9smSe2o5y9yiUPrtdSzgfmUwvG2NfntrRLak7epaXPtDSwyN0Ezj7fA2D/8lNNP
ukS3aaEISkLXLrEP1mEdA2Q1cLMDRXN3C1POL7mAaMFx2t9KlR7nm78Fn/Voix9+8IM7qgmY1UcL
9K9Bnc/xCuyslBC6n47Qg7GfcXjhxVgBkKqT/mtXiZRxoN7bqvpF7Er7tsGSBsqlJISsLsRTr6QA
P5aN60wVteZ3Liw/OYlHtpWEawLGI41jGIGl62ryWBTmhLXvFGFUiehV2kxK1MexquYhnGtvWmeM
dc8Csw3j+CohwVfoz5b4MUHTQWWDzEHNCLsSNGTqXeM58+vNdj2jlVi2rnH2ogB5H/ENbDXzMnJD
DDdbDHsXqLKMMxUy9x77GHbteaqLhEaIhnwc9pRX0FnSIK++rB+uVJjI5wC4aykxP+Gkdcsh0RRm
q7WjM22s0R/As3fbyXhEw5GCwcYhob0bujdMkGoY+KKMVfdKYs5Cpn6XcJhQuaL5HFIqxJKezO9x
PPpFIpnT/26r/uM4sYD2SxPaOZhnRGYIAqS1j1fpF+rjQ6+XcoO1BiN+GvAQPIcPyVXSpVtL2cjZ
NvgzRzmLL4rS8+wXoWUonLyIS1xbA5r1JzSDd0cEFW+M2nHI368OqLxw7ww3yOrcjTrnWjtB+/+J
sa7IzWkvuUI2oWfxntfp3TnYraAl/WsLTlOqzIe5sfk05HP9rHVTTE3OmL5lMuEABx8GvsJCFmK/
jViTOaM+XJGfKTfMQ6p2yVuC4QdTW+jArw3VEwzHZfvL3dfWuhijGnr1WCSKmmqRSCIR6meUYgr6
+Oy6Ly9Modf26UBaLLE5pS1y2oMhGK2Q0ZU45vWB1KZQZBOtOM/o/GTecaY01tvSHMLtgtmLPnM2
ggxUL3kIZrY4si+/AmBslSOXadcRiS+yKHfj3qAppDP+k3r7Vh7ZU+/70iju+c25aRgq2/EISe9f
SYBHZeo0hHO7rIDDa6r0niZnNW6I8nxaHtA27cftC2re0pGA2liPdM/xV6XIQMD0i566Zn5634bU
vQ9NFsu6s16SAvB2+Yef3O8fBgHLnLJV4ohuUNusXAJFwswfpsDHWzftl4XQsb98FOYNLf/BFtbn
oDoSPbb+JbLsGRBIKKqXxybxCJZU7KfscNzT6H+iCmHA2JNxSMVQh20G1cXHLuPa3hUaOIAymp89
MtpwmZ4Ldp8F9/uB3b0iBmOBPY4RaAh5RpzV7XQEYQ7eGaFFUhpZbaoqIKZOjAmEgIgfCmHzTiF8
7QfDAEltnMJSRfelu9eGHzLvpRr19qeMHzDn3prL8PufJs+RV6NdThOG0JugNBq0HXAVz3DUPJJd
B9S3Vqy/lFwtL54et+O1R1gwov9FJIlEwd+Y8VddxCbfO8VKZAyBPEfCG4/fhrgA+i3Z7NL26uIg
iAZoWNVrnwDRBA5QqiEA/qWpYrwMCuWwoDYYqndBXDhsPNxSVqEKawDMupWVGds67zdZAljWITGm
wtRJu5fmAUiS1QH8lZ0SI4LuIjCfQVEmxwYYhVMHNifhTg3Md7Sl0Mej3JBInAAOfReKNAr9gjxQ
TmV68svctyjpybMk7ApOH8IhTrtWk3idqu9Y0vRX+nDa14uX/w01ZGmmEQrHaHEyqbXb9L6McTrF
L0YMZyLoL2bSobD+yDms5r5n2UMt46D+PopUFTYpD2xGfCJCQEHLsMH25AcuuylbeP0WPtTimq00
1R2FLG5QNvX0Y+6O2oE8nZ7pn2DwOt8H12FhOe9lM8vJTEnSdJhdcv6Rj4oLgxbV492GYOM+hkZu
SWR02aIPgZNfN8IygkJThUVaBT3uoKc7hoxUiwiS0lq5yNZEty3RGMmE5sP5edpZY87m7ezv9Vro
PBjkv5FkafqG8A7V9ci7CqLC59oh0fQH2qgotpzU0+jyxztOr5gNWzDkHnT6jaDkvVbSCXHfaRag
/vkJZnirpH35pn9AFAf6hnilaUFbQR4klMI9XuEW0GKrcxW4O3mNDUvum2Rc3+FbKm+zmG+/73fH
qu8G7zYuDXCVYilSpM6GmuxwdTasb+iariP64V5YgvmHvjsq3+y0oSa5V8oyiW0l1GVzcQAvZWh6
lWKELvTNfDjxGnmJsE6P2HTsfHhPR3KxJEnIqMbEogiw1sSdGO1uXTmh732CEbiQZmaPFk/0hMWc
CRw0PTe9FKlWsdnplsEchNNEKD930HaWKVAE2pI2v1wesx7UN5yVS7TPzWAJGaRrS7hszyt5lmZh
8naLRYnCewa2mndRgkkySwZVZvs61d4k6iZfgyaaxBHNoF8lLM24iXLZPRrfoOazKCpl2QHimSMH
4cDjNNPLporfZrG+LWLvUQ1WNKp4wTaMOjykv+8US+KKW3Jfz9HLhKE5eulgv7cyXbyQUHF5TfUt
KQHHrS7sG59Ku/b1q1Dv41DZwqLh9KlEIG7FxEU8zhPVK/HDBj+w9UM40rxzE47e9qnZTmNknPmh
xfLf9UKuv0UtDFeSd8j3oMuI5J65JiE/dO+E6SAQmHGHOIl4xEjjS5xW0imh+uVtmLc6PoEG0HuP
Nrjtum0x/uMP8CHMMvrJnVMInu4cPRtwo4xlRLb+wkItzKpKlANhiNQ0/TJAlXAbDzXIlkNr+1Kh
nwvHQ/Eh0sH+sZkXiDSU9+UTXaojcfwLzd+8K42K5S/38BA3sST9rEWSNSD/lQdgoYIWWtkcxtl9
e0uroO6HR35Fzg61yY9iWpyZGmxK8m7tlSQ+1nzqs94RJ7Tu1XdLJt4SceLLOuM8OoqM3ndhSerj
0pPKBpw7iMguLU55DJzJmw0P1RMPXcb46MEAKFW7r/a+wqjVTcEH2cBVcUFVsLTrvRc5DSDHRoJm
DvwjvyJCOrATQIY0sFnGTVWuNB9owWD09WCHSngL1HHsGDdfNuiyeQTOwUCO6GK3jPtUp7m1+7ba
PcGhiwqbvRp3Ou9/SCXVBayJiVurv4HP+DXb328T+xVmPX2KU57wDfjFoggD9KnW6iplBv8lOv7h
9RzsnCHO8CZydytaY/8PybTMUl1Bfri9FBkpMstpY+iXgTNAx5KH1MNSVdAYrZbVjgcsoztMkyUw
58kcsvPTcGBdEuo1lk2/xj/53IwqZr4U2gafQzFLZBMBZOO3Hdr0G+GTjYr4itqVge2H8HyK6N+4
GyAFAyglPZr28CjgKU8H2t9NSZdGT6b/uJo55LYjAgljO7U8nL+uhled+xpxsK9YzS47Ptu8O76T
3EXXScrWdEUrsHsC6rKxKJd1mvxEsXzW592QXy4ct3EHhDDggUXaULlwCH5GZ0Q2Lcbxea1uTgaS
pW+TRkjJ6G0ODsiWVeGGuSBdg5emJ5NwfkF9QPJLYi5AA+omwAubro2zECpKgfbwGbx6y7x2J9m+
EuEtClfhrUighHthMa6gi0m+3vF6JatOA2B7deaihOx3I6/DCr33Muf7uyF/HhOBdHNPmtDMd6Ms
uZ4ZrWKABB9kX5TE0usf7cRF2IU6ol5XSRjbp1AU5qVYXZk/fT8UpSYYl59OIcRh4ADb/dNXj1pZ
Q5t7/5JJCdsCVC0nOQFkL80iqjxOmh9MDo62gU/CATh3tfrJSttm0TTzjPO+Cbtt3AQFrO9KuQwZ
KOcBf7IH2ArA7NmMFAyGxmDTNP/+9iHJeUjhWz7mMyL8TqkoRpSvXBfMEQegjW25hvCVCL4YDmBV
gbhvf8ZK52mUlQoLEGGy0jKVfB92WzmZQRUmcseNhit/OTKknezHziL4LLMlo7HUk+vnOOiiUtvH
evpXqiFAJBEp2r8IMumQGCwFJQnn7ma1dKkDsbAkrJnRbKwydDiB6Q3nu6vdMczP9YlUVrBE0Pio
4JcIz6Exk307hVAxPtRkr3nepojsbQIwJORygMGNt2cJsWzf/hj28NPjsTUxbsbQ6MJKROFcE7mi
1vMN/WRbv4+ufLH1KYysqDQskcXxi4U/gXAXsXVuD0/qnv3q7NuBPDpn7Fw2tnbM7KBSRFsCIqYW
Fl/JJtejPmt6fgTmZ8OO9f3iyvzFGNchSRPP3A3CNIV2G6QD6SmvlXQqazd+KPozFPMpXGgZ8PSS
kboK/U5rLk08NHsV2eQGdp3Zo5i1nm1pMWcWDC/SCmvZ8wS/Ei351kQj7qhjBk6vFB5u1p926rT0
fGJWi6spFboqRp1Qv103H2ObImCw4AHQs+IuvNS4g1qgu4vxJkTHStPG51pBbgIkAFVmKWNd4Kll
MWy0WkN6QDgnWO+NU56NxKZm4G2GhYZLHL8mS7GyPjX9FpwVJpc/ICTcl3jRXBHFd7h1onOAi60d
bA81XhdFFOg+YrmlimZ/t9k7c4HkEMghpmKjyv9jsNf5TMBw/rTN/zbnnYbveNymipEikagni1qD
Os64wVqd1n+euIh/phdDkrmIvoxIB0Xm94WaNfFcKg6/lypjidbs23ldQi8Jfp1KXnLMVUCxfELZ
QyBI5ifMUd18HOpWTuuXbsTQnCBX8UjYjNwtqbNAfYcJ/o+kH0EMUZCE48aidK0kQPumw+RUzqFt
/OYi//gl3KrbHNKB8rYOR0Eh+AwOEVbkuK96qleaSHPYrWEXXlgZhSDq9AMDNR2YkItOlZV9iz9V
iWYinV5Uw4noSCWN6ZNwT6VwacgyfPEwpRBo0N0i1fTPi1Rjy1PK3sc9cAHIHA7A43t4AI6+wd53
i2eofLQeCO9Do6tY0W4VS+++L1Gt7rolh6csp0U7DMKo0I2J1JmwWjnXeNWWNY+9GuMfm2EBVjb4
ltUqonSo4uR+G+yjOKQzfkSAm9wCEzPZD4Zec02b9a9pSZLMSD7YodOjFs8Fb9JOrAA02KuymyGO
nCmhktlEcy9jev2w0GmPoSyTfLbjafc6WL51aXzC8d9bctJ31NRdyinB10GOxydobDftVf5FcRXo
E5xD69jrNz66RhMHj0VRBM9Euhf4Y95C2dn9dDWmTaV/zLPi7n5CmEOMKUY8GAF3syE38HS359P1
nekjPXKKFBCiZQq6u5sNpp+E3fgkPFXolq2qIjFjzdOfv70uVOyZ/QP+D1GKeAZFEadZO2vi5yEM
oMx0U5B7xLX9/TNRAu2VXLRRgdb1VBrp39Ci8JIs3Y2RytyrugnPSN/aEnqeHnMeBjwKXdf3plsb
xCjCLY/cThoONwYtE8lJMs2fLz24Fex52otzhAIriZZULLW0DjmImiS+6Hd6XAIRfzNmupJ/vWL6
DT9vinYrrySVy/tLlK7SKc9CjezmIPvhg7LDgpaHN9hnBWcrwuPH4Nd0V1in9mRc8ptjSOzdOJ4w
JWmzxEAR0sFxBlzN1REnjRnTtNyd6fOyvnZtoJh8Kn1hDOvkW1JFa1cknGKIEmJ1r3452C6EIznG
yFwPSBNY/u+nj3v7efFCjJC6yYBPnI68MPqcxKep0kkafF7RvDoO4vh7Qx4ry6T7cE7qTQRyBwsT
ywTOcn2sSfbIj3He2sp88NK9J54k+fZ4wHR9gANtBEPkVelpbZ3S5YZo4NJL04uPRfCyQVUwu2nb
+cJgb/MRx5mAasXx6IXX8ZdgviMDtTYC/X3/+MNhy+jklH3IL6ltJp2xq4Ip6/AhV7aiRxfmTzpd
CsShtyQADB2D1ilUBOI6HgNtOLNIaBNm/WHpIixlJLtiogNuOVw4/9ckjDRyrxb8q7LS0OPW7DwG
/T6KdfgEvE5dhi/0/jO91E09fu3GTr7X185v8kkszjeOkHOMJh3KFuQ9omuhE+lxJk1wED8T8A0j
uZLFwqb9XRVXguvwxiRBLPzpYyZw/Ls093KTmvQOPGiQHJZb1yhLO2McB8soxMFS0j2rPN8qmYN1
CJVCmP5Pvyo20EXIv7JJL7+8iaPajlnjD+UXsqqfwMFDkmKtP0Dltp1Qw1qJVo/8YhY8Oyv6tNoA
Z9SIsFZM3OTovqUx1fedLIMutayWjgrCEYDcYJAppv1iVQUc/nrvvNttoAG7wjAXrw+F5mXP26G4
A0lfHCI8tPIfVXtuh/5IZZc00SWZJpv6v5+Tjvn8N0PjVDGMRNAVt/tL8gr867CSEiKTCHJlfocf
FjtXqfaUlXCnt7Hlc0R19vNJilmdOFT5EUaMjSU3hPsVc8vzS8b//fAaV4YzyruBNvfl0UlCo2nV
b1TXcEodS/aOf3qEOY+Bd6c3c1tukwOyqtVF0/skOEl6Cn+3qt+bHgdFjrKNNVCt4yFFinDztbjZ
9ek5UAH/x6oOYUGx5JT+kjK+SsXyBE3XhF5vGMxIYDskA6z0sTfYlsIdVDcMesM9H8VZ3ave66B5
j5lEHCMRg7qCOZF4/L9QtLzyjFxjqoDFhaHDkfWanFNDB99+6mRg49MA9bSA/3MIG+EV6J9XTlmX
e67SBH29UMR53XrVLIfZa35r5FiVSaPAWORD0qD4ljXyp7YB9VUvf/EKdMsB4BLrqW4hbjC95OQp
N+gj9Xm+S8oPMlQm2+PSSwF5o/BKbkSwimWVPfPY6YewBEL4ru3jDf6TMcFrypKM4HxNxj0UFr+U
wl+VLqwMxp94Ly/sBeQU9BqjjLrt05QnYv2gGB3jDSVxOjJ+6LPQe5U4MNGj7f7+yGhXsPs7fy4/
wydsCKQ2oIsZF5g81Ni4JG1xkuJYfOmJncdpk9AEEVQsEFkvonEFpqD9sU6o43ZzD8NkkjJfHLlP
MY1+3g1y2doumWMtqV9BHeW8WEV0CyKJvleawbvuLqn9jER0rSCkBJv+WVdiyofjpp5M1IKdGvcc
tjKieVakZ6LkC4oCthKhEQo3T94lzBRe/Gbpm+0T9esyOyUxNi/lHAotLkBJDNjD5yX1DA9fjq7/
M4xCaqgSkQAuOkksQLae2vDd8ZHpv6K8DOxViXmmEuz023Fedm8YTEULvZ4/l6KR+N3CHGSt7Mwo
bQ9zzKLrOhTdVyI98ShaUMnDLqlXYidUxAmKRUngtAsTosarKuclG5CAnj45RbB/epLobM3yxqrC
H+hl1JKi/1/axR0zSZk06oAlHcFEghzwbSySkcMb7mANZJ3b0+3ZOyCRKUKaN9QcEhulpCtMSDIC
Z4myAJJQEK1X1devMH70BCSTLB+R+eZr9Jj3eZprWQ50BtILjGZlMIbHWn7chsEmRaZjIYJBdrqV
siiLpq5f8v6iWk4ayBOc/0AsUt9tVjpSmhspCxqvdxJc+u1hhABHvgG23YlM/aKj6FjXTpRPr3xh
qGUOa3du/Tze/wIUsAa4FnYFrVcXElLZrQWf9K9+xR2tYNz3FUED8/oohWo8uj6l7tcZXjBZfHG2
3NUIXMQbudiIRBbnCvh5L4yswNNXgm3XY9UB4ppz3SvEd9wJQmEuAVZ9fihLYiG9d36ltGvJTbtS
d2bunzjW4XItmeZIK6NvQ5ED/n8UnPZDAtSHylRJk/VLH9mpVY4PcknUofW6RoPiQg4kBo17UbzT
H4D32iP77rG0ycVI3au0mZ9PxVTHtoApJcFieoYf5pdKPAOvDpQOQJJLc+z4xpmKTSx6XQFshNda
vtWi5oEhg/wDkBoBdOlgB3kYL77gTm2YlRfc3ZzjAas/SKT1sidathXNJCi80IWsKUK2GAcLrbzv
1V1dxbzfbOD8AyMLh5WELWFKftb5PTcEdxijntUbjnK1Y777vO509xROwy2djR1zKG3ht3yu7lgy
WIcnAvIcJmRreH1jVTS0LnLmjKJteD/v5rfMo/aQO79tSSzoEJ3lDo9HM9dbc1iWW8kUtrJ4D5dt
Ncth8tZImSszlHt/P7jjI6mXgsXDz97PlBNVdT5gLC1hcUEZsdEmoAZ1qmCRwyTNsvjcnNSHuiS8
oTjS59M2Wpg2/O2yNuLir8x/QtVIfZ+Nmfi0Q3nGcj1qWDMF+xzUmZvKdmwci9bZgZlvKlKIQCrS
BldK0MMGgUjkxEMCPNfkuzEFqkzl6oD5L+tPVV5gJxKgSq++eZR2PBgtPdn6xdIg7bR7J4mKD+zd
gtFxR0Gacl9WX9r4M00FOp82V+ChDXaErxGv5felwL4g7vZrnQfumlC13hjsYjm1oPogmdLJj7B2
6vwLFtUNLzfYCI2V1mTM57pIRyKhpt/qCt//ush1b8BUP5QeNllVeGp9QjIW+3t4syAex4Swn7PF
BjnaC+92AWJbDddPqtM/KNpX0iT1Js7oLDqSQGo2hmJzZfp3KWUTeIqd6qaCG32PeKVqliLA+FL3
oBbRXAxJ2F00JbwUA49lFKsFKZLFCB84evBYtxSZNgygJe9l8nD2aQ8f4vtGolSlJvHBIe4bhUu+
ej7E04lW9C4HsRjFGlJnfwPmZv2kaiuXTO0hIFVPp4epMqkLLgERsYM31oVYcKhws7WjqqmCff2B
PtnkfNfiFGpk9+YS/KSZmX0Tj3r+uja7AD7VoZk2933K6cfaNuBcGAVUhHaUN66xCBPEWvhIYMOb
WQ6BPuO/aIIbv0dVpMaS/Oy9fphB0wA4LSlo+butjoMThhZ0d6JpZ77VjsjwU29rkuGjb3Udp0cX
vL5dZIBJMCNXaxYq2N0RsCwalHLSlxBhBe+KZ0q+17i/ANFt6MYaHItcBUHRXJh8iA+7ZgEv9oxe
jCi6SOIqZAxcCpsPYkt0ph5ddicTu5RbNai+IXWtZ8yaR4B1FbikHUJODMAftfYUP+cV3eOk2C1P
sGi+V8TcXC6uKAYKEqTEgAbIiQRYq+fzT8DGIoDvsR2dW7em+ZXoAy33ZdjlkZRJvV7f5//W+9kv
mxQykDyOCIxjReLbELDJymSebAWf51hSd49QkamytMFacZvKZh8YiAzemfGjCTiZoMqg5vxIgyQS
lvr8CZv2xBzDr9KEoMAS+dmJ1WW/wSGoqY0fPUHSXYnCE1q3HRoxy/2zCQx2hGBQQiUcTkvArAql
+jBYlCrnZJwnK1AmamUtMDnUGuCYFCa0zzVEC601uTXM2Xt+QhK5CqO4GOmfPrFwI4XI8PDzDz3h
PsfWfvFbyJuRdPurypfr7WIU+O1ZHEP+gHXt7nM5oNK+r7UrC21QyvXbbsP871V8yPvfrQrdvD00
bC+6BJ2d/mEjrPz8MADtuwqq1DwDNMy4SPfh/xUSC3yjQnqq4KfQmBEW+nCNnMCjfrAOvZORnGjt
fONnz6dxrTVYmE3Aqysku/tEaFbxwCEwFYrN0CsqMreFLg+eONnt/bACc6EgxQWaFEmGCtqnFZFg
+ijbrSeDp7pn5kWDW9gzt9OWBht2YKgr7KNGicBluKaNoQGZr0vDJJb8xoPV0zauoZCr9e7FwTHx
P92h28FFJScZBwVGKioclhbURvkWfqsE4qBEYQ5xDNERNbSJGruIqctGmAyZ90U4Wpok7lLc+xuw
3R0o9Xgfj0VJRBdb6dtpNJjnDo/xviuRLY7CtCn7gcLW243yVgfqMJGjJL1gtQ+ExLnVt8jXe2su
hCCDZ1efH5+zfctnDS49IEjvyaB51w609VtIXYTQekADA7MSFjXZEsegKJXS/cUsMgRybs2mddMr
ySmnxHPQk8AvCWpXWjV8D/lg0f+lqf3Yc46uvlcH3pTN3kjE4WNbijpl5gSYQzmyb/6EL0Tpjrwg
K1SIZW/1UTGSR42OtnGhF9iRv7GLlAhBeAz7mes5ayn1tfJYEVFQtrxoqitY7jS1TaLMDhaD/xJF
EQ6fxPq6YjN5cUK0eNkTiemg3wq7Zcd4v+bAyJS5mR2XqN6jFMIpfAuhY46JvyP3dWheGo76uYdH
5nIFOuPZwTKRlgO+JiwDN/0Y+HRl3m47q1u6pGWfy8mZHRN61Cj0i/mVG1Uf6DKCsb4xan0Wo/l1
kcpt6Emm5rd4nLTlE9CrL01NzY8nv8kh3HbcV/4RIlaUB+gkpkSO2b8zyUg+FPR6YGUDCcpLMKWd
UPogph30b9ESyQBwd4MtyZ43FHZ7E5djSDzKfkFXCV7PCXOukogMM80niT7QoXftP/M5neObDxB/
Oseig9ur2S6KyhrbKNiwToqy4EnrTqrMddXVMQQMXUvPhmjZsOov951y/Xxy/BZkVqgeuWqNZdgb
K5ZsDWRgW/+TBG056kZTfZAkjsoufs5OPnEfCLPJEmo5b5L1dWvhXXfRYTYm1akFMUf858rXRgU3
VDZXLfFet6Uj0iwij3+qh4bBMduhOOtsPYqCXr2uY17a8+WFemeLuwpKYrmGm/mgENcqORe5WKkj
yZ6M4K2Mru09qQcjRFCl1/ZIM+aTGsW9YNkzhkDvfmwCloGx4iOkVMN1RHS93SkdJRrdPFxfOsw0
0mjSvtIL84CN5XX1H/2zia7/AQC08helSOmzo3I5qhzmtSy1wxfuxr6HEOnGGdV8uqhG0sSC6cuK
fqecdlLgE9lP2Gbh8UtnB9BTGpCpnpGjdGH/UCAkIuvqCCJjQyLqc1HmL+kPVcDhrBvrvhq9tyDG
KL7zh1JzUNHgSRcYh58iMlCeGw9pzwH3RaBYLMsIRoigce9MQfJsn0USvZpNAysLTd1IcXsBYlKk
jrUNgFtCJc6oGQSEg7tKZZmKQLwBB8AfROnmKNn0vkzpknrsuuSpGrFKAVgBLuj93ZHRRTbYoEid
3kZPFagO95VtlY/zEPJZ5LY+C3gwh5UP3ZuBnr5DJKzM+Uah1SnezwIt+SPvlKhvo5iNrEOFAABS
8TNoNZ10XtpMzBAA1DbqBplj+PwUJiU71QYbyN9ORODfa3isVcck3eF94tYS2oJ8UM2KWJG5OKU4
77BNKNnOWA2tDapjcpub5U0B83+0f8iLgEbNBZWDuZS/Hfu9itXINQAOhsDGtTnhGGdVbFRnyCiz
SHPv1p1pVvdAA2I1w9agXVuz2Kc/Lh46+e6orj2lc4o1AE6sOcA6sUg2IWhAKcW5D/whru9kitK9
OR3VB2IHcFBANUk4KW1zz3DDRPrYxAn4+0A4C2uxFPmZrbAPoPHEGjmqV/9L5rvWDe5715bv0DiX
WcuZbzsQJUPi8Zt9GH6Y3CXf27zP6q8NFENT8plqlseTbJTu8FMJP0pKND4h4Yr316N2PMfaZmey
SMf42FIzVQE7v2Oz3iUKLPEEuVRqzpZ9lnlt8JgEZXst7/+JhnVV/TILYSRYzQ1swvpjIQ3uJxky
8+gbYckdqYy4B82FvSeIaoB2kGbzHz4EFatcjNK2BViuGdWg7vdioRk6bSKi0R/gJs7prUnCzRti
8jNj2b9u7a1N2qK2hoKhavGHT50k8NSmLPzBDHtRI+Pnubm29y/uxH32ABNIc624aYSYzPHJtSXZ
+iWjFeGO4W4n0KYBC+vkJS1FRzFP9/F/EYQVFQHCQpNvUGt++dR9Gyr7ByS7Pof2BZS6rUUFJm0f
UD1d2oZFS37tRe+hE8T1mmw2ADd2M4jUGdLcnCNmf0LXgW9KIZzcbGkZFscZY7QF0joVC/QlDSow
IQc7p2JkShAXcstwBlMl0x5kd8oXjwWOpbjKbpzgxBhGnpXCXFMjYWlfftuOPv2NX1+vKY9kO6VL
lbuspHk+LF7No1dpgZPcanF/kG6vpGnT8FGO+aDlfV5Udk2Oe/TSPshKcx3sgTLyEPX1lC0YqMS8
iDpeo+yXIZsSNgkIbKSJ6UseYY0yqs8xAA193bCCy6g54z0GEjbzmCNkkgBgiKj2oBpWlEiwA4Oy
ZOZ9e8SB8t0j6WZs+g7fjb7Gfge5yeEPloE2GwLvUPQA9YTY4FNZNSLE2hoJHuviVvvho8UAlwSg
CkredYWG5L/1kKWTtahIac2P5jpWzbRtcuQJFaFtfsAl+t0udNkVNHXOaqPedUpSiraSMKARmWY3
q8jMjA0W4ZRAdVnmZ70UsyrIt7eqjMmYMBvb81icsiycN1ic1zTxCDGxuVMiwFPrHTSfZOUipo2o
I4GnrXfs8GDoGtQyPcXjg6a+L+LtOXVtIMqDTivH4u0wkl96qp4bsYdv65tsd87yzBDC0fQykWxj
j2vlJpcMNvggTqn0k32un5UPTos9kVflRdWk+YKYNykXKXp3Amyydn5Qchx2GDOAf1CUyLj307v6
vSQ2mxHtMbM16SrtKRRDlKs9tvf5kCrlgwF50z01iYoiRSSH3NJqL2V1qNuGdr0bHvZBBJcLwoDp
AfygsklhORO5YosykcUjzmbXt0K9HxESd51xTQtqJ+w1a1F2OLscHssNp1Vk+/+5pWMj9T3Qcol7
TqbSEZxfhJogVHzSeFCYFyECGr7k5s9wKjx/5GkYFv4F6EQdhR5g/Ty+9Re8xJhn09erNfz9iT4J
SyGyyXVzDbWHc2aGCI67nRucQArd1iK0s5QKv36n6LVyVIl28zaD6q8zsGakQ4596Th88+d1ZFT8
DOCodwx+mRcC20yYe0yV5NPE+isJXl8/iDkaYRMeuYABbYlZkgBShoSy3/FlsU/U99jHAdoU9aHG
xUvWJRAsG+eC/RXeI9fbjxJWYrgoaxcF9J1fWHo5/4dvpE8dIIW6edZuKs5jmsKN6TNZmZM9sflA
qgqF2K/cZb9h9UurGXv8iRw1Vs5K+R2Pa6rIjji5aA1VHZL2/Af2Bv40kBLg8udrJyL6Uz6jWy2e
TKidvqypEU2zxYgmbH/qhN0T7Voi3feMuVlSnDkFXa8zOpf/ufv0VTQ/99dLwNX9jn/Z8+bw7DQ5
99rdapQwuvH+XtLgeELLowUIuOhbfNTYEsTyRoZZlZTST6dErKKREG44y2aFmnVJi3L81BhcdnEq
SC3bBZ4Kwd2IWf+XKPtXIeTxIBSaIuIgogNCrzomq0ul7hxnBuVngtTxZy93JkTFlCPrcWIfy91W
ZbJDLMaH+1VaHXYt3rDHhGrMp0r5d/UkG5CmdTU3cqvEttfDkB+KrebF3PhHjSterupY8ke9gsKj
e22Wu9tKQ7SjLcp+R01iYUZ9DA3eVfFCBdrAu+T0Ouf38Pk2b/EOLnTFziCBH5cij4z10eLldu4F
DokWsULqCJ9XbQcCSn4XgpixmfnBwQSnL5g4hVJ8tb31RKru4r4A2A2DTrrua8a7s1XNtjkEL4Y5
fQNojlGUaEjrOBPjoEOlYJ2XQd8y26z+d6DMbhSDVtTjT24wJzy+HV6aK4pgxtJ4wTGQHZnoBTu2
77mcvNiwFjs613eXMZs0MsMiOWVxopEnh1R6/fbcb3E/Vcn+xGGAsLq7ONh9nBSnJRZg3y1VnB26
UygKoownQOjoe3qPZWlriByqS3bHCOgFbBs2PXWSA+LLIvuE0mrwfsWfXbUQaxwia1pZAJvSx3ji
sfq3P35Xt20D1mgqXkLWVkJ98VNAokBLDWUFmDfb1xN4JPGMPAxoqATHmw595aIuriAUn1gkwlvv
LelhjTAPPfRtRcOXsFB+wcunC1Ux4WtQv2SpLgZNIdK6QoIpGXn55k8pGP02l3hg7GrY3YK00Ouo
6H9ETqb6n6NOmfA/ILUBl/lbtaebds8KjSEOyr6SZ3Op3fCfs14oaIwql1NVjSITdPQBwCZUxIyM
Uu6w0QIVe1KK4Zo4MtN29nQlud48LbZL/XKenI6Jece7KliMtV+39SfoyTeuWJokgEwOGpQf8XBS
b4E2f4pQfpy122aE3aJXn4sg0QJuzVEiUGqcfoweqsba+oh1/mNqNeCAU6yKK6fHbZUUBRT3Dih/
ZrdMU2yzoVB0Venc5/r2qhb3xOMy4B/AaJw8o+uovqGR1HF0FC5pEd98KbeC40UQUfXOUHoKEyFQ
DHG+ynUIHZhkp8lCOnh7usjHzfWzYTNjYI3BT4AfDfiK3kHfA3PD6oFCl8hOuzyGEMH2faQgCTgh
chw4i18yAMBif5T28cQwzj70VEqgECmHsVQnCODTDYzq1dkDq0SYD/On5QDvTg43LVW2ExoyE6j9
iCZLXsw6QnIHuqkduQ557AxScsNoiK3n4utULahUYdbbbYpWXs7bIkKfGHNBFuFe1pJ85ynyaJiC
CqUZKxSdgcWYsUqCupfxO7RABYqJ+N6Wuff6w4J4wTt28tPib4hyYISY1L0m6UHGRTMc2yNnvDeu
JOJK9EZfEUzcxd8MBVmyibePoq32v7o8DXhSQXBtA9/RnCEBuyON4RfPYzeHqi1pH2oGI0U4GPq7
XeyDJ9ct4J97J6n1KbUtEtadfZ8QKhXQAEVCW0i59MqDpTLzq2mIw+aBSra0kTYanpPfWA0fDaOY
6OOSkULt8A2bqtXfcSedHUsUxQfv+QiLxPQg6EEr9KPZpYknMVwVZwi02RU2oJcwy51SJ9Qe6i7M
9gOkoNfoXJg6aU93NypGJwXTUaMZOMb6LU6fd1G54LWEkLAQtV393aRZ2dZ+7xl9cfQeK0pSLg7t
MtN0uyaB8VsmGJXHtiXLOfz3qaTLWuDLoQvwYlEUw/cybu0vzJHkIPhluH96RIy5bTknSFxteuvD
lPuflP9WdxB86gi8NDFi+9R916N8ZSHNWVRdTINFemegqVVsQ505cnqya6tC9zXrjVAwsz85G0sJ
ur++fEsUXXpN3RSZ3HT4Hhh+B3OLPXnQtJXuKKF/9zlhUswe/drAtQQLYwaX4IE+eu1SvqOIS28c
uhERmrGMVZhfxR2czl8Eyek54Gk9TyHbICCduOd5N6hBuDMXSc7bg/d1XYkvc+Um7eiGDc2ejGdL
F9IyuqhxjeMyk5RfdlMYXqn4oYefjEdu4jsmqT/11fs9sRCVf5YbjW/tbuQx9sNdlI8r1p5+UQk7
aBd7m48Yjzqh8Gd1p9aRSr2O3Z5cu+4g7OwssJ2sc37elkxfKd8BtrPVqEc+Lu3N50aN9VaE14aX
wP2ZmUyy7f0kwGWg+iWuNXMVcMkNst9LOcL2xtOsfh9mwoQkn3dDKgKRgcMq0jkQsoU3ux08QK3B
Je/3ouYbxdIVzaUUaf4Au8Gb7lCN3zAdN5/kRuq5ZZM/hbWEfFIQ2taPHBGZ5gX3reTeXB1b7aBJ
mKeMc2yG0luAhpn+5A0t+egGvpWCvSvadPWwXhIcYMWM87dzXY2j0ZS9KWUiOY6cMibnj+FpAump
vHmXo7DVVeHdkmMQiheHiYKsRpx8ksmY6SYE+ZD2BqtAFStejTr9zCGPhkeNxA1ti4NNOSDdjtFs
vugQvfWGZc1uc1OWyA7uMOvSYU3k+yIbjrv4tNTZNjtaOEFTeiVRgcC6/X42Aav36+IT0YiKcnTl
jBlgB095LERmbK4giIF04XQd9Hhb5S5y04Dnz3UzCN/mVhPRLEqQIxYF8wtHUASyJAapnW4BFGIb
G/xRHkBt4/lOVG3XbDAbnSz52f3+03P15tY4hT3C34lDRemNwTJt68zmZ9JWK3xgBmz+xy9FNNZn
5TVIl/izHcfqH8lXzFMhNjxh8DZXjCTRo+6SKhA162ldVpEWUpY0bhZbBwpeQOgs4NQFCyZm8gu8
laJS9ZnA+96xGmqGWBWh0PpWrKLVh9/O8u3P4WX/ATGcTdgXwfHQKFI8cr+tgZq2b5I2xjkCadj2
PrMeHMBZZJ5NqsscrECMGY/083/F4GESGBdJHzZJvCoj5Fw+H6Incq2gwnqeejmcSyT7mvVsWoVS
yHFd22VqjYfdqJQ5eHdXygUIJJLCrA2dbFrRJbEf8/SBcX17tx56m//4VWfvqBvQ3qbTlWhDO3VM
hSWD9o8pL1z0ZFg4VF1rpF7C0n69dN5jplOZ+5emKG0v6kJ/wM/766GPWNAvC20VCs6eAmhUIcu1
g2dPxahmr+qPf0EOjK6as2N4CPotxM041QPCxDIUVBMsKJ0xU80nd4kqZri5wzJ8ECl2NGCWvIbD
WOXHAvU3f7PG+B8iUqLeTQ0dkDoQYHQb9FxqsOeFg2jG/4LY2tWEp9VIO1C09zq3wBgEntNfpTT+
3x0tFxfj/pT41+CEnJ8+SHZQNa7KQPm0OKZFdA5ziqu9WcClQI8FV7iQpROM8UguHdIBTDXgRZos
YvGSbsUnCGxIwOKLVQu9Cp1fTftCaZiJkzTO6B8HW5fH82M+fzaDfBHeEJGPiBfBEu5Zpb4FzhiC
d8ix3GZ2XkyF4b7pMBeKC4FFXbndTHQ+Z1ku0L7/26ELGNNkGJ+jITUU1OJWmMc77Yc2bOcm4nUF
JNLa7yhLL+eTJEPyDlwtCtli5xiq44R0omPYqLTdl8iWi9NrGSrsBc0cIEeGRQ9m4+LzDbebxwlQ
LYMG9pFZSXgAS3L7It3R4axsHc/hIt13cgSqMbHcqN+FmLw4YY/GJcHraMUE3BvYKvcvRR05+o3X
yHE9js4FCPmqLwwMfQkoxHcvJDFwNky2FzpdEF1B77AT33cnlvwjEfDcy49sg/igSmRa6K8EHF5Z
W5i6X0DS5RCxf7DrKGPpgjeYq4I6J3QcJEXcTNLj6n5WEDlJXmzg3Aku2l3XbOohujSY0B/iDxWW
UHqFLWEDafpIGe2uDvFtyLFxPJbkWAM+59stRExm8govzz75n4ni0aWQr8zrwFZY+rGQfuSiEBQq
ThYcVCYvnbPXpufrXetcw//NpD+kAfiXPBS8GGatYaTxcAQsO5pt0mQ7Vup6eZAYdWrSVJgxAkNy
O7QcJfHnNIfq4MjpDsLfgnZOEyfBoJi5DIxufEv8N8JTMMyZ08DTdFXkCDZRuDmF/lAwPKAa7/R5
j81DtHoTYUQXRis+EuC1L5o2XNfNS459zaYNYPMhpnn6oHNldVko0RSoVFtpAieYnZ+LpiAZhtmJ
AXOJF82aYyEaZYtyQF7FhnRmUBp/KlCRrkKw8QS8oXGE2joxPOWku9enMG8P3/BVvEqJQ2jhXbs4
waLozgKiDHp6LxC0NaDHg8BS054EztikqqOl99XACqaNlEE4rbZdCri+R53Q51oDTz+Wk3evgdMb
ThvOEIZMvMdqty5w6EBwvjWeXf/z5hhpu5HMNZ4vICoC/GbmReWPTpqBh9qyv+RnpGDDYwqpVRTY
6Ui8cYuxxwjDEHfIjzDgJLjOaBUTvsVq26sEyFk6WS4lMziLC8au9b8Kt6+3MjyQ9NqQnrEwrlDW
v+D8SUk2Udq3ZZkdmPIFTW7/9z5IVhj+qJnviXshibxI6CSYhVVhYYfqNKkDczwiFIBUqf27RjuN
/E3XA7Jp8uMVyE5sLXh6I88l0mn7irGs57Mw+fZrElawy1CIWK7kvjJ7OO+MWCTWkPxUNuy30FtI
KLpjZwTl9JnS4uqccxP5vMCymYLKlC2jCnzNIwtO9GiRscnt7Awby98BNfhoxWeGTbmV/bAr93sG
iP47EJR9n7lDg5jEq3cUwBZPWq0eU4deyYQyCIziVeYWlo8p2undw3memgyeDKXTephp/o/2ougL
eeP/rARxpaxubsNX5v0nT4mgpyDD6Y54Cs0+W/UqCaczXzwN6IhhF5OJzAwO7MaADjVnmlkXJFKw
ChTqIVl/G2tqmLI9TcOHP/4fhDsd84EEgLvvDk2ToUgYrxzyGXT5xoyk2iCg4l6eL2NYG53GxdQ6
A6Iwy1aFlDPO0GFPqNQ/RVt2yZhM8gmKgbAKCMQ7T2PVZvwdorUxXeOzDboXYHNbimyBXbsaVy8U
yawcdQz97LRsM07VtdZcvzsI/QVOFyrybavulFRz02Z+n7aQ+DHw++7W97sfmSROQYNB/uCG2WNu
RasnPLcOTVtkftB1Xna1Ky1tMaL3W33iUywGutUHYDaPI2wUSKXHrnmKA++vOhQyxu+i2qFrSja/
GglppmWFcsAK6NJExFpWDxtikhQJUFIM2D8ZGyis4ctjyr+4LOTjJANTBwOrxNpjbVsoIIcYwMuj
yX52WSGuxurM01YkySIDRoNs03GbaQVuh+NCGYyjvGBtiN8+hMFLJhkcJWKqW7vhSwXc3ABv50fQ
HX6AR9LUTB+dclkAwqTbidlDuimP9eW1JwMaHDprNy5asqnP/s4YtC2RENmmPIrrzwhAu4lwmbiF
YaVLtunJV0Yr1xQU2bZA9BAUMhIOKWZ2DlinKnowL8NNGP4TtkjclTNqOZh5YqYIm26eLUj2tWg4
ZPpGd+fb4z/E3aeKnB2s8E+83HhFTUeMiDtVR/5fexHVAWmNMGwPeexLl+oaTvYhlc54GWUuP0eW
llfPhv7bV5d7Xq/pi8P5Nthljs3O3XqDjlWnCnWF4NdqDx97AFVuRzieICy5p/bDt/iPhDAXkdnq
cWAuPXxcBG60r6VyDV883dZ3IjM/qBO/jmKZWZdQDr2sznHx56AXUzs64BQ+v3e7iBoy8zGST+1v
KcFGWDbLNBNJY9tlo6Z2MSyJvdhih9uyDPKZ1Qw5DbnV4OVh+nqJC8RChgqOuc1iBZ8grQVd0BRA
3OsDGDmsKNrbyNZFoYDdig/Gu2JBV2s17vI2Q5LtmSyRbH7/PewTQp61E6OcJ9ZJg0VTTrBUpPyx
/CaRETH468eF3W8rVGGUIn5Vx+IFMF1627QRciMF5uKRKI4RO0b3OfV9Z1NJBDTIJ0EZDEEOjLOh
SW9MjV6KsNJ2qJa93ESl3SRAGAcA3/PZOYiNAy9B4tY08qyrHSadtr/0J0e9MPc3NXhGfILlDP5Y
f0Bvc1uCbNb49r0Wd3TvJAIoRGMFQqryLEAidzXVSfCZk5EI8byNaf7UAh1NRNo+UPErcGLKDGT8
0XvUyxj4uIOPlUbkjuOP/dfcP6pJUu+QAbniattkUnGn6kcWuJgU5/QYRsp5eIDOFFa++FviYgQX
lamo3wlL43ydORTIFF9MrbR3gJ3v0H0aImjSjfyhgGgBbC+cv/E+Y3u2msgGPlamSVzgi43K6fYf
VyZugkepXaq6+n36rHnzA/6sYmht5R5vj4d9QG8jqbvBiIykjnh/NHoWFuM6AksjhrhaW521/aeb
+G8hk3XCIAY5mM4B9rHVmtSWyku7mmWY/XbcNwPqwQ/A8Fac3u5I83qIUGVTnn48mTFAIb1G4n7I
ltTfcgsno/zMt7gft9nm2jMKQEsWmvUS3xaa6Fpn19slgX2YoB1OdjHpM4TJN05pgTWnlsdYK6wr
FVDQsLXJnXsNzzpmV+MlG6tH9HIAzE7LWsBemZ9Wpf1HWx4HFd61rMOPjJd1zLklbyX6VD2mSRrL
cctOp26rKALeLJBqKM8sMZS2KuQtYAv5TQ97VMdYvZTOtgLCc6pwAHeOyjgrbOA60KQ9nQ3DSbOQ
SBAe1+Ag3quOF/bhKMjqPJAOjJ168uXpRlSzHNwbRVX5DN1RD0oIYV+CzLUGJp0rntPBmsf0eqIw
v7BtyvszTOElXgW4L9S1G9K34phOxad6Uw/PzvhqQgE6CTnmlyGXtq5edq4FyRAEIiRMGH29vQ7+
5Ns7SQdcwkaqd5YpATXJQUWOJGL5j02GKik8uFtHpb+t+n2x7mmXTNc2712uCudWLsRIRoKatH9S
v1b0gqqlF6+XykX/1Db2tJhoNtEX4KWksu7WkjT/vzHQKt4B5La7DJnjkk0mP1xZec9Jrqz2yHYw
wEmVAX66IjfKy4gACZdRstagrl/0CNLTpxfk6o/lwnANtrukB4VUjx3W5VNl/gChhkNWgcQaXvVR
K9TZu5JHa67e/HLAM1b4/o0hHGa0AvrCDzeu9Y4jJo5NYoETjHBiZoSN2Sloic8YX3OUD73XGyBC
CFtsRroQ7ZPqFslzUaEHAsVg25MdTH26NWE4iwEIMGn2QxEKlvaWs1CAZZWBoxfye0CEmkOYRvh/
ua/oTKGVDvJC7cMzLCZn+TFnMkKx+/Fj9eR/MWjeCvf+bQ7F1Q9gPWXjEkCnVpT2melZlXXogY0O
k4jQZLuh5RVDwauoLOMgCV9q5KcV/GcKS/GqPCZwnYCHpXfIy64esuo5nrfxbskTyA2VbNQBFfu4
eT5aOIqqndwZVQr9Dhsw31wdGxSkZEn2ZzF8klH9VsURINo7/FbpLw1J46ucF6r1gYmZo5b9drMS
9V3Ht0WXGRXPBpiaBbe9bBYRdhmqYs5eUfgvaEPmAsIXyj/5y0iT0cwiRiYlWecUgU/tyB8ZRvkh
B8nQwviMl0F4v7LGVAXIeQlOlzY3HvU/VcD07Ky6GIbZI81iZrwUEtlIsnYRFdQP8f/iEegR1SiL
yD28E/kOU9H5EyEepEc4CSKL+QfJ0juIJJwKyk6CxQ0Z82X3U+Jo1z2topT8YMuJDb3t+5TEQKDz
OlFa/4Es2uagJnHnbuw+RykAzhNxlQfCeXeGrmyJb9YFWIIiRzsA9ddu+A6BnyJwf1uf29XeCq4q
DJthQ7tgn5al5fKjUdso4HqheP/06x40nkC69Rxn9OxB3WZIQ31QQKGBTdp/nAsF6o8l7xbVXHdw
CpilaYvHdEqvJOuuMiuwUP9L5OaXz6hr7HX5whKAsABZO7S7aqIe+R8lrIliRYq/uu2QeT1afoFM
Zo2J4g1UWH6tkh20bjyt3LYKIeyNPB7hJcfALAn23NRKnhzLuGasQwhcxWK3RlTdD2ZmaLf0vP8y
WO9pcYk1S53Ve3q7reMl8QFHGGOX8iNrafDhoV1t5tjLt0VfguCdqJ07WdZ+qPwxdImxRSKaB8O+
UoLnMzjgiID4ZWH2x4DImX6y95nF+AYvBiUeClSBIVbPbQ/ge9GOMoETix3LoKHL15jQwrO3WWFN
T9gLt4ct7l9NlUgPFkMgzYD7FyoK7XU7HKpZirOAHv0MhJCtAcar6Z13OXplQhxZbpX7eyXrddWn
gc5AZ1sV5g0/w7+Aw9GN0Y/Bq976YKMHqGFBHTz/hNmGUVdg0hvSbd5oq9PU4IjRVTFNW995QVp4
lNL4MhqjSU+pkI8TyS6UOE+v8MhQjqnaY6NsanSzFqGZXH294X/JzxAL+hW4hG/oNWZwhZTeDZ5L
duNy1JWeldzifNz6f8keM5OYSwJAI1pSVyiNrErx4eKbh8QDgvvEk/7fPkBCtk3IGdXI0lt3M474
CQnPsBOm8wt7zrmnrOvE2G5JvhYWziYzkUaZpqsG1o/8EwvUQEJxjGR1su91kTwiqgZ++LM52IUC
L9midviC4muOPurayZny+yKcZ1p+jXND2jJH/kX3YVDs2cGcAQg8twWwo7bDoQz+rHMB7fg9sgSR
rD+TNM3M6MQdUJil6NO48u2Tb775a162MlKdJ1ACeztzO0n2vs3jAoh9gds8U0klwbz0/Y3SwsLM
saMBoVupoCfCRPb9aXArafM3tHKB5THRQrT99mE7P9xUicaGsobde7x0QjgGC3ODHHjyvZXiButE
fiOEBA31E+5OmYQIrKnF266qVls2ZRwUtAK2wyUA+QVXks7XOMkkUPyxpy+6QzZmWgtK+zDwaeBz
15k5W3f5zhiQhpbrMHmPz0hyliEnNGdhTDTUQHnnrPbcN7/q7acd7Q5rw1xAjsoUdVgXdWtC3pZq
gBY0cNGjnNaJyQhAYE13zFgHufaqjBbfDxqoUdttxop+uc2FVTVQi8RYVSXctugW8SpmkyKW7VPQ
HcdCr+5KGCQ2JMjVvnvxa90CjCCkH2NzjNi+WpUu81ibgsG0l4vRFTgzT6CEhBwHET6mdR5URC0n
fTRYYscgfh8IxW7SJ2TH2MOvnM+K/ZZyOe146q/zpshuBkjVhlde/tm6Ihs7uDC7VHgMXRCNX237
Qk/D1d2rQABM8snb8lK5o+KwAYL7eb1bIDUT64fvVuq0JLs63vw2deEgxuIVCE1mByH08rimy7pt
ZU0I6/Il01D6f4FX7hqsogfWIfTEqOrjpvQPV85sxsJjiXzzx8sZuxpYHi1uPpZIC/ePSYxEbtuN
4GcDFYtit1eCrlqGxAs4z8Uwdbh9L1v+GpdNwCzBjyClNFJZbEM3ycu4ZfWuZabDD2iQ6TD4nMEe
PA7x17O06R31lzxu1lV/v51XSc2/8QFlhm9ClZTX24HYkfC6+xlAZbsqKm+KFSE0Kswa/ZdYzfoo
A1hi5JQzW1TxmAJg0QA1Zp/srt7hgZzYjvg0z+HPiRMZE8cA7Xir5OPaS/EhUypnX+H3R7pSXF+Q
cupQg4uIvdS5dx0VgitRHOvQWST95tOCPEk1JvW6/ge6IwFIXCwffRRwZ5JORWk0v9LxBXpxlhbk
/TCr3S6XwHVy8XcVwsJO0vFAkRqejZl6/wEANEe+wabU4HWYBdZ1awQoC2bWqpXXK6+eJXbAsCL2
CVa2zAqxZdXb1HPI6duS2IWkkkgV5rChPXXd7gtUvvfslVgr4z9jfmb1mVWsvMp1GTOGResUh8EJ
j1YNgCLhvhq+wKhnex0ubicYz49agh0wei5QG69ia5H57xQe8eqoyEvFzamS7sV7FR27hS1f7lC+
bHvsiNccq4DSMAhuw7zWt2wJZWkMBQDWAaEe3xz/Uiy8wCSgGzvaRqgdzG1BQz3lC9kvpJBVpXrX
Dt27vAYZWtEiu9E2G+ApAEIiqR89bChv4lzuM3UYRDjR408beajMNp+M7JMsxIdY/Lp8qwbXHGIn
kb1IyG4aWRlFeYRpHE2lItWkjBcvAfoDvL8uE14n4Fjg6o852rvQMWaVNu1uYxAr5s/Os+04AK/L
yYsC2Gxy9URh8dAXtzSycdxIDv7QLdP7/r6E5U9Ik5Xtjh9c5xmLb8+Kn9UIK8YX1ZRSnQVY5xHH
l8SvXUwHTHApbS9/8mzobbfnRxAwX6Xb8B8fVk9VNrjYvTvv80ytTw0WDMVZEaZqQCIK26yibagg
NMzXCAsD75jmIGtilORTA3FQiHAL4ZUEemE1Vor7nNr7/aYhjSyC28M5XM00Kpd/IBU9LiIiX7gj
sw2N+17p0jIp6aCKsXcbBJQFywSR7cT4rtLDHMzJF4AXc9Zq/9QmLeC3cZVrdiPqqBYWsT1eGpeg
gGd4Byw5WnYsg/At/JkfuljQhkoY/CPxyNH41ORX7a2KG0QU4tr8u8VhnOFQH6vzZGiaeYAlmTQr
t8wVhYD+Qkg4y2D48r3RmnEUX5ClCoXAUtjhcE4TnuKwIhJrG5U5Zc6CGvD9UY0y9n+kjDIY3C/4
IJIWZEN2UpEkxLSyRInbqbzYIhWdR3Zvw5JI4yScgxfOC14MB6VhQweZuRqZ6kxCRr+6hqib4UR1
Kjy9h2PU66CR2Hn0EB1B6fh7PM3+85Mv9DN8TJkOfRCeB68alSaWrcgSddq3OmvRb90+HiIZtPIv
PiDWuk0G7qOeYPnrIUAc2lu+xbVMEA3WR3zd+uG0gAJZo3AHZUyDQv1SCsCQo/5PaW6idUc/VHpn
XA8T4OQPGM5aroD2TatLa5J3x1J9oHHdXsh7rS9QTZVap+X0xEJEVXcez9BeEnrcufrGV8OLT3M0
Drae45FYCUugAUueN0bmPYW4mKqz4qS9sSq6X+5GY/8QhBrrSO+Ge/f86ez/BbCZY03GGjPYkCDt
NUsQUxVP3LRNzJiSY/C6s8vZp3YB9QvtvV4QD4XgEDK3wE/QKNwjDK+lWnd15MAqy2WFXEVNW1/d
zWqXip+sEostC4CbA6h7HV5SaEWyTfMqP8SVzBrJqLP0o9gUNCU91asKnanHnVdbTxs0SllV1dKf
2EL83Sq9qo3ptP5LEhPCaBtITddNZ5Wg+yK4tjrQHeqvRPZ7VNdi2CDrXL+41KfkwPTbiyGtHc41
BarWqq/1/SkFzptlX+qD6/lMMWqHdT0VRxQZT1tvx/b9Z1maLBEluTearyqVy5ILmO+ZJh2Zqw8c
cRAiLXDRqivFnmwNeHvTGXSw+cORdc2RhJvFC1QQgCPC4lUZYTCcZasoOgKE3uf3p/khKKDwU/gT
ti1zUO1phM1iCk0zrU5mytPvNh8P7OTi2Nyy7NKKVDZ9Nuuz2e4ltHHJwZEfsmVqNjM3QWGhMg2G
JgSM83NFvEF+OgPdKlsCrbTj3vb3Zbu+xua79nXiuxNalbtL3wAGb+fI+mItD4jKb2w/qMFfI7yz
OuKFjigeoXuP3PJGgo0ZvscQ3orX2yLfpSPh4gxScNrc1TLJuC9nRLWmFmyhfUsep7fAixZ6LxtB
2AsfbaBBMqjfItKrd1VAsOI+AX2wnL3ezTU7eSRXQrlpvxW0HFrDIBmAqTUhtKMzJgmrC2VaF8zw
OXIzfYYALM8Y4gFSqmpg4DPSojy3FiJULXWwk842LqXBi3BnMPdyFuhObvvrPdSjMbooDMZTFP1f
3VcPbz1QPRkWsnpknE71+P1r8tKWO5ulyaffEMg8snd+AesquD8ErTAXdWa/gUd8Xp992+T+7W8W
vGYYBlP3zMX8A4iesyhFxs91FeiVmZGVQQKt2kK5dbGU0mFB7dSpyRu0KZ6010XnK00JURti+zUy
192/PqN715fVUzAZkcnfiL8QACdhfJWhE2zUQb4c1VBoZbWpXqsPpO6xnniUjRXy/ZdddaSijaRR
oPS98/D+YqEtFWGE5O23RX/Pkb/qKtXL8BzQqvz3HRIK1rsqXa4TSt4iCHAT3o5W8DfxEawnTlEU
voMRcW/bObS/5PV+ZWYanRHto23IQT/v3sfdAKkQp9MErDKnXcZmwxsOyb2UJ1liE7gxpfU14JBo
gUQb9ZC6NkftNQO9AnNeo7m4HZWL5VwkAhG2aTcw6fxjGOl6wv7h7fVfRd2mUZecGe86FBytCn72
7xPhUd29XZBbdBElfqPxrs1um7pvnyVA+OTaPnxlJOOAiHfvEYX32vBXgoUdPwpCwnY0mvX6Y40i
8KD8SzoHjrhY/fZuGUH0KaVA5FcrhBI8T/tFqzuaw0fnPNXqixJwDcl0UfcZwAxgfK8fwN5368P8
NN+stlRS5kjStBl0cbFHu6VaUQnqcVF5gUXH4uwhwL/5hnvxfDXY2udqb5qW/NSHIGz/eT+VaP++
bLIeoKR2Ax4GTUQ+DLAquwMDcdIaNRRx73a3PHM4De+x0vGYBAXXycHjKWRP4Dp0jTrzu5Vg7Q2l
3gbPyOV4e3TzZJbv66XPriq7ACyTjP6GKuUc8ub180vWK2IJk9QGlZ0XA1stY0RvOAGLpbheJ9Ls
BUNzQqT5xgNPrr8/tn/ePDcd8CmsgsPD3+7dO30pid0on0XPeqOMe+HDJp4XY0eQRyI+TovwLd/1
qV+nPPjHJSM6FDvRCH8ooSJLbA+GhUrjPDfE3GGJOdClAjzV+EdvBGXWSOQ/Chj9VHz+/QnZ6ETO
35cZByFbdfirqEwyr6Th2kUogO+DdHQJpPhwpmGrnqmHQCgTsfFoi+yXf43R6EHzgJaSMFqR2Alr
mRQKG3hGJ20VDpbCy6MnaG6eDuo3zFR/3a8MqKnzFpeGUVmHRFjvJGiK54irpl8k4senccQGnrQX
ieP2fxfcFx1/vW+i0PN6ihyI9X7d6j7dVVvQwK07VFEwbVjQrKJ0ZyYh3MnDUncsJ4CEDiJKLp1V
fpLSsPrlmypQ3x7BZahtWgqkhAV9p78blVzujNq58OcR0hG+KuqJIV2xih6BB0iqFq8TxxrT2LVt
TA8Jr2X0WGY2hs2KPCGGV9ZLoO1EIpsutFnkyvuRnDjHMTo5lHVOLpEWir+0kBca9Q75h4xxGfIs
cHBumXqTM9hgM+YIhSC2ArFBOp7dukX7u7boxr1u+DQQnFtrdH1Ydde+GbFTGmfqSgiC54PkV8KX
ZMChPnenEppy1w/Z2ioOveDLneSdXNZXvxHHb3NbUh1KhZM+omb6IusNQFInTha4z53FECgxOPbb
/C/W6iJ6UfqrOEgUKN8WVrCVpYyGDGJZw07Q1uXTihmf2DZV2rOR7XJzqqRW2I97a3Zw2FO4sL2t
r58I0WWIdgClD0LKS0/mQOrnzMdLA2EM7XB7MxZ9sVVCXX9gTeF7e/Aj6Y9Zc4knKgU9c0VfZsZ6
UnAKAgakys1UZFwPNzpAGKit61wwXhhmVdcgpxADDnef6Szlkk8be9y0EXIRPRq/JZdNQzrsDarZ
SEzn99OwvdhovE1CngoJIU310F7X++2tCMeaVcpm5PtSwjxbZv0SN6g2Sh0GyNxDv43OtJ79fcVX
lMKihxMlUpsEp2g10b/AYM7DxefqA200VKtxyFSi/pbXbQreek+MHI53cli3ym140dWV5IlI+HTs
A7BQUpnY2hdE5cALKAChIwuP3hJM+ObSe9diM7UFpnMazAguX+US8Y24gU1ToaYJ/grOhXSZEfrY
slbPfK0ay1IXyQuQIXkjmyGwC9OFsBpKsRBCLQvIv/HKF/I3LUZJrcAQ09PfE77CfXxJqdT0HDKa
jioWUeheYnFtEd6HievJ7IX5pnIj+wMxbnZjNH6guguQ66h61UFEmc/YXTSvdhnIUHOrYK0MnJgU
7H1FDx3mgPAANwXhv0Nyq8ShHyet6bWwlbtSA6AnqLN2ranP65mQRoeM4ni+ge3k9KfkroihPjHB
UEI7JEcBggsszf4VOMTCKznDCgqwvSaT8ZjIwJsAfmajj+BpuXzzIrt5gxMJbbeCoNheFDSlQhKR
PC4Ua9mrkApYGD/j/J+iALdo+5+eUQ7Fp9ZRYjaJkoVgs3Ymo5PdFuB5SiP9XzeYD59nJndZAWI4
qeUEJXYXj04oQ28TmWpVOJPlszRiWgXN6MALccPmmNlryv0D6RhBEOdEzP+y8Ql85qGzaejMYokN
YRDgvYOy+Zvd2D6+YVcLsLBbviuWreBiTpaKBm9UshIHeJ9FyYgPUNo92G7U0ENXoykS9OOcEC6n
GngWMoPfgUWL3UXDtdgaybfB4Os8hEscSEJiR9ZTRXVt4/l+gF1LarlUBOMCtS8V30x4WiWhbSKz
PFdnnLUdNkM+9UO24JjU+6wX8N7xg1jxX12RLI8nCMZchyqIGHjahug74W1hirhle6O0U/oBvmm/
Gxlz5ZdTATh9KPr+/ADmVb4AAD54Sm6c3RhVaucWSK1zG7kQrK7bVcfLqNN1ppeSoQNHTrCo9DRl
tcsGHFObhQCbPlgBw0GNagR5eo0/8G0lIaKfpOhpcKIamClUV4RXFhzRcAOyY/F+FuCxmhXRJIqA
BoKD2gzhOjZ6FXedAPhtWJc25MX3Q6drt9AShKIVbMbC7y2LQY6VsI3keaoBrbmB9GpOyhQDKxFG
ODEAKELrCT2TGnPH3fBEm9W9tklyygi/IRX9qRkzvsOdZPkKSXdAG7H9XQiVQaeBdydXCBqSq/VD
xpAgPwTozCZsLIo2kt6T6mV6z2UfgkyLIAYVVyNeU4nFbmMchUNZuwZtpPW5bMzM7iKqLHZfQX5G
jbrcJ1GHBoKMqnyRwQsPcPGKr5UDrq7wk0q9Pl82DlVAunvQ4gJvqB7xVOy/8GoubMXwm0fa580V
muGHVBII9BJQu6oNB1JxDLc52cRU1GdChhgMon+JuPvCgg+P4baSa1UydNt5E6TMqIpER9jiIwDz
qmtdjby4UdUx9wLBTHXSgRZ1z59QySj4z0roYw0Co0m9/oxWrkd3BupaLC7LI/w/Dbfdg0jlhEzR
NkssMLgqut6nj6zPmGqzh68ic4feqszrMsLH7t7jo8Lyy+0dT5SyDB/V/sfP2diAi/vXArknVrRD
gnwMNatx2xNdHRwHEHRBILIavHWC9oMSBRYNPRjDO7OccJU35hy+ia34Qyjy2gDmU6cL3NMN1g/C
vzSohARAqwg5elCg/VcTT5rxRmtFeyTHKipTTyZ4awNtJHr4Mx282pIb39sbL0d7tzuFUq6hBH6K
xjXRe+jvvN8X7pm5S9ymGLMok3/Enjnx46zKssTkLqhZ0B744CVwfOGzMJoAXG//+cssMs4YFd3f
m/J9SqVpzz+PPJKHvWRXmd3nsO9x/LA4DuWYXg+ps0W1JtLj+4fsyCsZUSnM2hCo885DM9+coFs+
tW838r+TFE9DP5W9xdDjmiSgowpkIRcXp5Fa9dmAkAqEtnUMrGnBNlZz0dlt2zEeO3mOAGQEBEk9
7Zwf4QyxvPqLhk02xpecTETaGhsY9jBo9OldcxKc3b6VibyRB/jVvOd5Ts+UgHr3MajPT7V0rHx+
1uIPdvJlRyaqfHZ1c1nuGvZh+79rDJKlqWiRXJgweGUNhKy8RsjiWUKsSs8HCUN+nHE4vYly7Tac
kKbFkqQ7cQuWpwX1meyBEekgdy5vTFdCo9nIEUmkMhEuisxxy0efHB4Jz4Xec3n4HIrraRUjp02o
Wgiu/06jLuKTMzC6BG+AROOCxwNmHTzrrv+IiAqkT3TSwHFnFMOBVKKmpeUUhv3cbrRbJQODVzyC
OOFWh4MymnVtcUcXvdljzyELoiCPD7eJoljGBzfoWXTa8nvj+6/6dBo4BYXXsERayD/8mqLLIInn
HzqgYdxC387GjV2A0bCvLXYUu1SNWKDJUtT5CWDPT1yUaFg6guHkMgyo5Z4lW5/OZcJR9SHxHm/o
y8i3UDMBInDLKE7ENBUYlGg2zp9PPAsZhtamHZhFVZSsY8MXi4A46Txqiu/Sba3yGiVT679t5dD6
kAaN5ooN4SkEjbhumU+OQ3BkYMLAWQTzVVo4LoWgwM1klu+nI1YmwjBmwe/1TwfPbCP/oFDyOxYd
DE6q3Lq1+vJqWrLLyCwkUCrXCGtsiBBDQppokLVP36lSmZHfbxJTy3lsrbahoVPq/B4QgaAvR1KS
z5ZbRjwEDdhHp3SfglYQdtjfx+B5ZJDNhxGzdkz1Q0waJwEKvSJDor3y+m91Q9nvFc4gYYAxPD2h
cAI3VQ1we9j8Hlo4+5Mt07Hn31SnhipomVcOUVl0FG4D47HyEGR7o20sKncXOmo8eZUBfinc6Iti
KxX5jtwOd5Ri5MX+Tw2ymQl34I9U7N+PjVhxjV7GKQ00j47GZfPlcg/fpmgeHeUBaiOEZPhv6Xkc
5pYHtqF8KNGLc8IoHT18fFopWAZlB3f3Yk5pUKdtw0/xPVDLx3CScCBjB4eJgRCBAUwc8v0ouWGd
ZX6oYuqkSm/cL1gzcCEcgALNoznY8LV4d67Vg/kLEs2OWI/DVs04n+5mRmrEIlqh5GXG/xzpy//R
86XWqhbSHR3Z1ypwIW4phveegS0EtUnu/cMABWvmrz+OsfRRgD9oAWvXAUVdSnlWa2knCw0u7JSj
BSXrRCF7RK0IFzf9bLfJmQb+fchGZlMZr3yAbtTk+LxR1IX84IWaFxstS1kjAJeK5S1sLdjxJ4Om
aIoBjANikbh4HlI6nHSfBGJ1leAEDzKKcEXUMHCHMd6+2iZ2eGEsRM4tZf2A6R4QxKVMCCwZXXUv
l4SxgMY8GPPAqJCmUg2oDZ1wfLRWSikJsl7XrK8LN0sby/uKeB31aYoEicLMm9f7NV2ulBvWidcP
KIjhGJHW1RbWNyDZLZ3xEuEEgu3BDexOwp1DX8049XZfupSXc/f5QxDL0iFBR1lug80v1HpsTFLO
ms0XLNNt+XveOjbnUUsJuz9jrNEYCmJjzVL3GWC6CqiZb96IGOAx00evoD5302MvXfwBTgddJFK0
OARKdo09lNCq7XuQ0SKZZYnzNEf+YMayInEIgWx4gGQ95Yx288mWYNnR4wihq4pEAErP0450bypn
doIBzkZDQErhcoV6I9y7RgNo1Hizbzfbym0HGXFROkgk3xGPPfFWaYGxAjfqQE9cVIJRmtVKM4wM
1K0J17HMfi7GV+mD58RjHyBDdq5V8d/AllRARkWdokfctQboPNCV9rX7NBBN/oxRogS0p/HYQkL/
RX77+VKFHjSfmC5duQYDUGQs3MMiimbOSa99gaZYvJDAtaneeB00LHK89y37SxZVoeE9pLLl5OWr
692LTZ2Lqnneg8jkj9NXHF3vD9y+u9MQxQWUPPXZdUctbP3GsG3s9wFUy/Oit/DUTwFoxWcFIuuJ
tiODKRXfGCOhSz2uEuyMB/9U/e82MsBwrdZFytD0pGfQNe1/tjdPE5f0RqyEIv7E+PKXk8BY9EZC
1LDWgCZn1z/y/bUiX+OYAdv8gnTbnXyI+vN0FD351H1HyugLIFtqMH4olqoyPt9OfrOVPw9Ts+5U
Ii0utMQN1nBt8HIOHiLvrJ0wsFXz1oFoWr6TnZryj3iHAmPY7dqHAFf9nyaAL68bfx01uGPsXQiv
2X6cRYUQQuI34MN7QzEQNDlIBr+QOFrtysC973bA6v9kOF3PrPRtkWTZt5Jo/nRyzcXHbaH0Pg5u
fnlz0SxHiBjOAW4kV24qrRhNVBtFFyMQRq4g1OXGywnwj67KR/vmm9T2h/J0jSe1Hslrl5T1OAZC
6wpMUc3rfHrgRNhIusPwatx/CVvl9Pafpwh7Gi+iSMnp7QySuBX8QC5Qnzs+YmiDd8bV4aM//kXF
QcX9jf4m+km73o2NqdK9OHy7iAiHDK8SgaelC+1uSI740Cz60eplMMQh1qeuTblvUJwDivXlMEZH
YMDUYk0UGHJ8cubocbS7jCTKRY3jHwRE3gDipfF8RVLJHwYEUK7MhMF/NT9WFk7Q44QbR3BuIb8S
zVVEUKf9ghQE3zoHdbq0N4YYk7FPwpoSSpZlvZT+WUshffRM2wTMYhZ2ZFsEV9f4CDEaBI1N+sdL
d5yb6egdidkR9NBbU5T9nsdpE1OFYftugWp4zUg+ghgleFOmMDKtZTewBgJW2ZgSNHedKRxCi2K6
Rpm6NSeclxxqQBlZng0zYXaP1Ss9kq4HXI1e1o5TKXAqyeRCRmfMxP/Ul6ItZlDkBw48F0+UvkuG
WU6kjlZ21UKogPGjspTDi5qTNlbCQo8H+cC0pFZmQbGeuYmJXFlsiioOEpIObGNNDgpHyc4wS2P0
2ch6tyQId3xILPV9qEYTrzUD3V1Apz/FyLFzLUPiXXuZLSrG8XoMzHCU6StcEfLWQeIdiop30sX+
pStpKat26B3H+e/oSh+EFf6Ao8yrIp9rATGR0pHuHrBXv/0ZT7lhOAYGlv//zIWWSWCh4e+emmXj
DWlVta0u6DcHst9vzD/CP9C00g6ibPN3vH7yZpi2Foa8pZJEyUmoG1Hk1Lr9SdnG8s/alICEONW1
Mj4lUL+Y86bdiTaqxH3FHPVmN0icDssYsQ+Vk2VuJd9F8+oGuVGKFnyvpuPLc8XZLRyZY9udrE1T
xJKYa8SrKiZMqMmGyMSGNWbmPUT2en/AG++XitsXrOlWJpXoooEYXKXcj1ilsHqdBXbbewHZYkGC
6kEnPlNA/ZYoTt7KcdQtof4XjKhA90kObX97qywf6+fyDB57a02kQcTHPYpIv09vNhl8ttIOFxDa
S1ekrDy/HEvONQY/r8Kp0jv2JP21SYZdrk06Jc7OOIHg1IWLhgt7fOhM03vDg8lz/COQhUWSNEWJ
cyb1mNwmBuddsz7KMW+SOCguVTqMB7g+SXJ+GMFD4iccIt393ADIx8CdbUkghnZ18NLuMJ3zRwen
VKV7i4Nv3v+jFUlUAcaTl0dE8TuKHvFsWUaALbLSXYG8rfbyZPcyfQvy0/DNkgqWWQHEQUMfgkpo
DWWi9e6Ie4iFr/6yAy36hFbZ+5tKrr3uihlBoDbf+Ii5RzaM2Cx69mJYPaWHTJbwE1e8UNePVqx0
q62ly8s6U2JIDRvPlZyBp+4+D7Go5VM6+f2Pj/HuANV38vE5Iqx7XLEMKEhJvuo31xAvCeql/3Vz
QJdzTXCcpxrxKnrMAhWPCamjnMaL2qrUKalxaRSNm6yEGSRHK+oSVXypbc/WrrcLLV7gYqHghy3t
ixVIPBISCj2/5BfMNCWeuNkaquTEgvjibUI9F+O8iVMoSb2mAfmNhWVXbOEuNdMDn83IU11hq94n
lTWcyYjWlDScY3LBfS2kK3yBN8j2G0uLNykTe4sPJk/fvJkUSUOBMh76F6bhfk/bLfnG5o1X6YbX
kDQ18Z0Q1+dasJxJshALnZEp4hyGSlnJOQE5X0eWlGkUFHtWzBLNNPETWGGQEOLvAI3N6i9p0PwI
OFNA8ZPliMs+9PaKIdROpytCDXcgKS3GT34WPWIXlhN27iUsO3HaBkEMldNsw28JoNzpMoquOcUR
GnVGsFt/AKqOUS0VqEnH97Yfb4G+B++2sIFTJHgsCn9WhqrnSBghBg/w/nbEZCv2O4mIXRjyw/sC
ECaLkjCqK3Did0WasgyCcQ8TpNgro57s0gqJhKmVg/d9r/xMH/3dMGfgQKnNDPCaJ0s49cLHqeQq
zlCzDsv71NCFXFNuJo/F6H7I0KI5pFNrShtkFDzlKP4c8yKD6wAvBtCD0OrilrmzuczWLyjTme87
hHCAouKNjhnP6in8X509gO0zbe+7twj9/W36R0yHlVYhaDS9JCFrRJKOKSfDwY9HplRcTva9JKoo
45ekHFWTFhXpy+a/r9G1zLOItIkwy7105IgNjSXoCQWaHZBFBDJay6sOXStot0rDSUq/PxPUnaMK
MdsP/p01+JR45YVSVzvPnM8N8ZmLOycIQ1gS48Pe4RxPFkYDp5HZc3Y0tDHNtfn9Wr09vGgh0MAe
s6hv3alM8UMPVbErE3IUSIdA3vkm4USEdWskhjkWVHffvRV7sgDdeQChglvD4iPORGwgP+yTBLH8
s/3usWNNp5Eu8sYH7r7kM1CbggMWe/rftQeAMn+9s0q1LAkbOo0aI7ZCk721FzwVRmDplyM8qURL
fvVdNDz7LxGwq1FPipsbwty0LpIdiFNhMlyL2dsynCWJhKF5rs3Tar7iO8MP7Ym4jZc1TsDltVCC
yVv/TnoboPIFMIualcu3kkSCk2sZ/Os094pqJ+LQwZiT6Ec9M77GYFkJC6S9QgyWFmczit0N+xqb
HgUxq4Baxlv7SfZKhSOjPh4XaF73ph6zOMPMGQXmKuPoYTstjYvu4awztaajuJzCuTDSWKpxCPew
UzavswbtkdBIQhFXbTOUOOr51jE83xl+/b+RlAv+krb2qFEPKhgkbC6piseti7mrxwU62wNHjCkS
XhUsXqO3/BpT2OL5oVVVHWXQzLHUtmInPkYAXrYug5pC1PiOIfwYmHaP8kv2gf/q1W/zebvQUGT7
ztDPq8DwkGI0GECF6ve8oqz/14mDn+TIB+Xn3RuAddnn9Qg3T1zYvIFfrRJKKxTl5rEwC1Zu3UO7
/iXakcmemaVFde/WMoz/vLj9ANlHeiud36AvvkhNYCuIjdAyQIz7dhSk6UFx2psBjqP+ADLwFH6v
bVRsGyq9+uqgo/sr8Us9uyywV5qKjMEuNDv5bnLgxG5dRb7jPL//Ra1TsHAcpJ2dbRb1jkj34hDR
JT13f642JXVT8V3rTiBg7TgPs9tqTzfPvftNe1f3h3aiLqZvuGz3W67k6qb4A4fJdV2zKrsjJ7AN
tpbZp3b5tu4lyJF4VngYjf4LescIRStHfy+JTNEiHT6tCE/49nCo8ch/xkvUXjRhXbcLe030675S
s6JT6dFTTDlr1Wv3bEAfnbyxFasx45v1hRN28mLlPR4ngFtbllJhbVWYW8mTzS4GWGOIQ0peH+Ae
5/joMfHAk1cxo+k6Ast7u1GlOVM5noNgDzm5EN4OwFLmO7qIewhJrUZONJRIrh7BAF9w6SdGHWbe
omL/vTZ8wvCRoeBPkO/d6u6+/c/Yn9dvpdc7clsDF05unD1DyHIWG0tA/z3H65XT6JX862XSm5LQ
wXufV3yBINqnzWrboj/e/8R/9Tp5AhPqcgSrpMe9UYVvhOGV2aGN3/lDWCd4GJogFiy4sTLYziU2
PwKT4B3czPpmBbOpBOaPJCg8yk9TPowPL/xuvgdylhl+WgmSzbkxtriGHc1phh3ApAGlG2zgudXU
AnMUDzKm9dJOBwumDH7H2CHC57nvqgr1scJD8hEf4wOoH/0MhPfrSdgx3DJsInHbDVhIrkSKFG55
xXaboHE5ckGvKPMwWR2TXdzeq8B3QwsUpu2CpkiWTVo8f5oMVgob6Yghms1SV60yrZ8n2RuEIwjq
9GImW8xEg6ETVRAoM5mchSbHoIsvQj5yBhc1hnTpVI0KIMCWf2w2UO7oj2BDPCzZQl9xx78UuQYA
ziWRwfQpaEK1u+4jhoiSFWGd2a5sNKH9mjFls/bu4xesIsP00/ffLU/OV2i1rY3IGkiOKhC2NfrE
NqiNEBQ0HfIKVaK4Td8wgRam+2J5NZzDOqpCWLNvyII+pKptb0HbG23p2RHa2PWvU1R7pjJTORUW
7mB3q8u9LaGYd96lRiVTuluYrDcQGq1PElpJ3vGheaG/jlHwrutUUzcMCdZb//8Mzn0UAVkVda2P
Ni6XgqbQcsb/t3fSUuK3IteqVkzI7UbVrkWO1D25K1r5vb/6TLkpcxXx3+nfeFhd6Snlc7f/5+w+
3qPrmYv+iNNVD5xbOMb/qR6FvEZ3SXHjnOIjkGMgUtDslR183E4bnNym7+RknmS5coN0b/TxsNDX
Q+QfdF1n+MkRkkeVni7bIuZELzzUIq4LrqYzwkUwW0mSxxK/lkQc9kpuUzHCdPcKoaIbEdJ4IoSm
UrlmieXAB78LBmgXIXgbsjmjwGszRwXuu3PI7wElmKSxlBLuECIzeTqUs5P6GQfzTYsB5sgu5W0w
WOTOpfWeujwdDLDl83WwZ9STd6lYAt3anUUDMzYJe5Z8J1UJZRYaTbcwcU4Cp0FUdG/KlIbfugb2
BJpgwPhlvMxFmaqHPY6yNL7tNaKko+bSzUlrIM8NRgAChs4Ak0k4hLkYak+w7DAW+IoqDK+eLFq0
oQI0ETbss+DwXMs0jSKICFyKb5edEnz+7t5R7yVt4bEX3k26OG0Qyd7RsMx+yXYknzSIp7Ks3o84
8NDbmPRyo5ghFjbJo5cfYmr512RJ89xdZYesga8JbcEVW0sUMSpTZkCfmW/EKQLQfy6koQ9JTBYl
vh9Fwj5dE+NxO/nyi6oZNfq+riw8W2BQEgK/Awi2TfcZangGCHgkFKgpayGz96VLBVgy5BLaiMO1
MJtPTb9q4hOiwcHZLnmwkUHhSSAuVuj2vpzz9xl2FlGChVfYZpEf4PUtoMPQYCvoZqzxGT4orX1o
H0H//HqEeSlx0VJXH3YlPmIcTqO6vNIamQjpxy2Oz9YL14svyCptUvWC4sxSYvojCub7O9FRRhUh
ZLCGo+pcvsmTTDciUvSrry16o6K86VfzJHTIZJ7vIP1BwOB7JHb2GfIoVa3KhA/lqrLFKXGNxrI7
AL2l9D9009j0WRB3W/aLMc8cj3Vlz2rabyq11tpw6IC/5xlLnE8O8HvKIIR7qjP4NxUtBUSL2HhD
XE2p0souqXMrYontU6Mvz+i7e3DpomQxN79mqGtmognATetT5iWB0dvqVPpieB2prNMtRddekdEN
l7hLD80J15OB5VF3XSZq6T0L/P+/nOBGakS7Jz71xQaAHqNbqG84B/jcyvCbDQUfTfGU9H0qE/bA
hHeCYNOUNoezsVjhy3ULZU9+mDyT+NTwqD/LGyQ7ggZ2TkgAETow3ex+MPgjV3qYj1hiAMndB6uK
+qYyhIgAoRDTxB5VMhAi0w0uVyhqLrcOeVv6yBI1hwGZivPbDoTFYfnsey1Lg1m8zggqUTR5RR2o
YCiPQCaUqo9mwCZAMihTBIjwh1Kdr2XmE7oqeOqkadkvZzq+iZdVaqtbZgQm6fNNFqZJW7av5FZ2
xESFl2BXlR9KEJLLJ4NELs96jm7jNpQ8imbhjjWc2sfp6PgXyz1LqJRCu8QtXNHQLkv4tGPDEcKj
4jPJ/FmIAN14jP0KjfwjY+beKnJxNq5D1wboDb4tghN1uAgOKiLDbW+sTMTQO1eVnF5jSO+EEwBA
oc7Oq1NrO7MTCyBWytxT7rTbXDLzLrYU80KhcCsGhi7zWg0LZsMY4o7ogIqMkgsq1LERNLwOakKE
UO/5GdCBuUMjj6Gm9yLrVAtLFo2M03+TIHXah/p/V5OawBshYhFOL67pHGsSfKWI6Z5SFreTqZLH
Zin4pnXV08G/X1q1eWWB8zl1rVexap7poYd478U6dMt1DcS719tBS/NVQ7gJcHGzzu1K5jiPXRJE
D1/d2eGKKHJXPEhQpJezgtfUTyAlYSlnkl+nCOQm3psg1bp9KGJOqoNHDD6f8bu/vn62IzQfleUX
8Xekk3bC7hgvDkUiu9UDrb0SLXo7qT4oEPe82Du4WSHCfuL1F8y7b1Xr9T2RrTcAqOVfZ9OnKiXM
g5qh3XeulydRmg3Sc4Rf6noYCGbetlWD0+AHmhBZNPJb2VIeUNdnBNa6VElpl0L58EAk8VKnc7rJ
MA0n/NKeL4pmnA7g0thNODKhPI4Y8Q2VZQVpi/68b3y5DJoj9CINMFu4nWlzhUSDY90A80tUnxGL
85HcO2iBrt0VHQzXc3E5KCqYSqc9Do4vap9aboO5f8jb6ESiMGFgczJoYbRSD25/6ZzP9iNwFleA
1O3xEA7zVA1ZX/Aw25+tE5BGa4mIGZmZeqiC8h+cx/7jO6I12GdvQlHjR/3SVguJC8LUUcjlMB+p
wFQj+ugMFWn9ZK1/toQ/7UGZripRgqkPuhavvrkM54ptiQROJDrm+5LbvGvZhUxCLhLkcN2wuXKD
OvESIDnG6sR0IbtgviyrGG99NjeeJveobqkxl9bf//UfVL2MaX3iHSuK5zSvqd2doHjXmXg72edw
qg/pe3LRNXnvdV3xDeUzOCz3y04uOJsYbDfx6zVxp5+uuY4JK3Q0nkexY2d24WhB1812PRKqS4tR
sNOcAGW1gJHQbeL+m9hptRQemPuhhPdv/HQSBS4Vv9fCQLcikVJ5M9QSLePvtvSMte81hlHwtag5
/tkjbG6xk5Ub0K9Y7tizA/BCsl/oDLr8LwR8FoPUEGH96Jk6nsy4CfpgGm1eahaffoQvdZAR1aUZ
8dCEiIjYQuEsDt+kmLdO4rLAZy6X+9ggSx0MkFe8gQFooWc/2Key6fK3qboWXMWEFkmvKAccxbJf
sWYZrKq1bCm70KElbpx0Xpl8pqFOue7cNFMb89M+ZtwyzyG62hoOd0MFYdFM78ZYpttggUurXr4r
ujkqBHEej6dcoCCcrggnp+R+CjXBlWv2A9jLI5XGaJtvQ2tPsBW+s6agAYH5EWrceNtH4vocPDmT
+wc9x7DpQIzIy8mD0f/PsSJmKVN0m5ZMTRWoXkL03/9d56GyUNbHEY6nmwgelRFBgf7X+wowfYTU
WzUAHYRGlP9UfHAOua+dLr82i0bod1XD0zffS/jBuPyi6le7apFeOFmaElMVHjATU5kfgwV+8tFk
54/npG9JMYknkm1kUQcy/XQG2GAzHxYusnK41J09bZSBZ16Z+iP15JmK/UoO4M1juPc0Lp77qwC+
t/ur5KDTJXbjjJdfthQTwrGr5f4T5hNBUtgiBBas02/ZqfXkfFB75uQ0cVUxbQ5rPS7kIhn400K5
O+EdZcQH6CuwODVNJrwPRvLG7k5tfZArcs+NUPLuXubx/Mf3K9iK1OkWjyh5kvHL4Alvm94IciRZ
wVjojh8SBN7SALpQafUp5v5knlZ7VSTRA2EDqv/IRPemi5DXvLX/2NNEyEh+1g/9cbLayELzTzZW
4/Bg7nKuOzD9p3vHxxvoUm+NmJ0CFxfILSDhPPOgZ6Pa+GLYW/FNYCVz5xguS7I4A7flUzpJQIgj
svln3zCLbuUUN1a3uWTAmqgjwSmKkfgHOhLhJbgaUVaQQMoN5/m9MBT972qvNQy5apC4icx2PYF/
mV1rvjx9EyKDF6iLjEVhUximiz1cF0mlp0ycNhcTxm3lrm1X6v6eDCSEv5hFWpo/FlrS2N5UABoP
1A8reHglCFkwpd0EAPTfEpau3GtTtMpAYNE7y2601g7xFm7gJE4PCJqrid+g9C/8XFZqytvZcM6F
8XFkyBidsJ4MkJbMJExe0bRzgITY8EEIh7r4lDBMXOj6CKtKfjde0+RxVuCYpCdsvpZD75ZZyCeQ
UUNnB6VCjb/TP0BohO0RQ/czAa9cTQMhXaY//bfeJ+f8ZErxv/x+RKL6wc2+R9XcXxxO5zMOshh+
4j9elDGxhd86MZhyStVQ+1xRiIw27j3Oi4i1Rc/Mk3fsADFWW+ossyg2NXLn6jrYUF0YEwYli+As
0FJdo4AvY4MVdZeCvNMHNNn0DzOXmSGcMWrnaQ6LIkacEW6OzJ8NUQ+7MokObft8ae+ktJPwqAR3
yAs5im54rKKWgv064ZGNsfYqQ4sv6MZpmaDbxO7wqjoV9huFOTtZgNoSRdFKsnyR9JiiarsXKx5W
lOU78O1g2BBr+zq+/xV9H1q4uyiuCZzXvuBWWJ9vb6xhYDzyM0zAkFvLQXkYaHH21Y/mZU0brY4a
cxqY6L6eQLyB3TpUiLz5+goliNeZvZoBgms0qDMwh3lOwSx2RzBJGrtJEt/5aRor/mh6hHSq53xz
vf+RECZo3i8rJdPjJhMhdAxNNnFles2ujXE7c7TwYthCjUzAY2lQdLNs1hggDM9K9JbyTSnF4317
FZzH+TcSabY9dGFtbJNnJq6XrErY++7oI6XuH+vz2CP0NigKE+po/H0d+UC7/2oB8aKQ9HYshwJT
8icTBhwiNJB8LGJVBhmavEkOA4De0q/Zj+pBWv/D117ThwNKXRaVrfh0afhcFO7S+xnFN7PZV3va
x2uCykA2GWSNiwfBKlvHSTkHeCOZYSoamJYMs3KTrtnLo6rZm0cxD679dQRiVxrBDSKvqVmIH5a1
OrojHvfUC8M6b28Nfa8+ehhYOX2jPFAg1MJ5lj2xXgx7w5YuIcath1R5zRQnhZPPmC5/AeEsOFfN
gg2htbY6TGHPAFxMon/PGgj+fe5FZiXxjct1gdFC/piMrnGfH+9BGSUu0iDRQniBgFoXMPV0i/XC
jh/KaHK1scF+yuIdbYEPZ3Aburqp95OVONMfIr3LNkamzAZ+NSm3wKRnc05DJq5xa6PADL+ciKQU
ftIG2qMVC0y+7OOqaWPXTWdd9NkG3+qlWah71I5N8yYjWxaaqD10QTBdD8fAXRzT1+HiCHKA/Hgp
UUsSMo5TW4RGQXqDCvkBqqCVuhLKusbPDjlcO0HgUbzTs4eeFp3EESY7mgE9P0thDU+TTZ2I2rrl
ONQIwu9Nog22aw+gv32x8SPHf2cNykgCVKg5lATQ+Vsvh/41MezpSEpH0tM2pxijB1zmtBr5tR5J
yBA3YXTGHhOE3LC2n8P5Jeb65jdzgOvJIhealqF+PjP3XzPSGFDYQsG8hRh37HNdPa/jG2+asqwP
Iv0q5QtT2Dc5KPRRd0xUCdRnXVWd9eP1Kgu4OrhkqFSjSPsod9WlqkfYsf6fR0UfX6MszavQBGl/
QFxAGsoB/cDT+mnSEWmOLz2G6SkK4mjXAoH1AueW8pl1a81NyO87jT0OJRkC9RyQAALm63GjouH5
EcVC+b8lHefPP7GYYtFzEefTN6IuXB1Ev/oH+LKaeoGFVcQsWspWeu2kTDNUuI6oDPIwj7ibcW+N
zZyLVNhKV7zZ9L9FuzZVy/8KMRtZCrj8z5Rsz5EBLPi0ow1md1d1wD5AMP1O88pWWHdA1yDh2WEL
zvv0A2TbxkKLt22lZVdSYmlsbOqlTObiL0dqIFXMf2yiKj2P1KXZios4jbr6cC+acJQC6rn8AX7o
Lv1GbGoWDCJAcUQcXtXzmPEgRmj9euKtG4pAwYl3VcJX4rHFlz1PwJWb8bZwRrxgtkkBtTE1ocIo
szOWU6MACwYa44t+xXpHYrDr3I+KrfPZV42bqEG4L7PYIskgem9Us9/ih3QRjR9WMJDmAhygJJPC
0x/Px5ypqAB62xnG04vorP4KdLfePv6pmG5XNs+LjXqNKvH/k2fZx7vLMVYojIispZx4cplW92Pu
KNg9nl716at4YTz7WRuHS64PX9TNuorjEYUGgZ2lohj5Y53geLamOeS1+HZXshHPeokW4VdTwO5P
J1cw8Y70Z26qpnn6JdGDqNjZIafTVPBxoOFW6QBJ1O4IQyPeKWbU1KV64r1DEP5kKb3xB8a7qcqn
2TbGS0XU7oGU0y2Ylh8wMmwPN+yPvOnKjXLVKg2T7MRB/9nDLa6QblCpS5HIlE9blGzB/1uKmBs3
QBJwLcYaMiZx4FHPlIaoyGW4tL94ZntyiuZnCCk9PwFnPuaD3kMVNi5wB2fTs6A6RrN/m22/6Op4
1nnetvCakTvUkwMAD6R9fZ2IZaX2BPao8NVt1bmtKfx4JkV1hVwEg/v83R3FMqIKZXJq8VvEVnxh
d+1+CxGHDl5TYr7IDcnJeQJPapfEj7l+OBYMlgFP9QElSvMSnOGV6Azz/arp4hlhkhFLGpISX0Om
CLD6LHGvkpTfmVL25eDEh5imqoB9mRMh97WH9SU0veMrWfGvbOWaLGmvLAJaSegJZ/wfv5E4/TfD
qRNmBCxfTNr5JMGtttyo8rW7y068LY5/iA4IA56jLbVfTOFu1r3tmZrnnUf5Nv+aJqEFTozwXpeD
mf4Y8OtS3i4i64YdIPSQqhtqS+mIovMvdpxcPxCbAF2ZwDkQrTB7OEi9zwLJ6acs40WjXGNwRcql
OEr4ANrRnu3WmiG3TAn8KlXoOMG0SLZIduMADlzlV6GUbgo5JbBnOX+8LXOo8EnGqtF5kkay8qxH
pyhLF6o6RH4KkCUsAbhBfANiEMPqjNWsdOd2HoQcj5T6xNbKgVa3jg5ZZCTtCXWMSjzItpHuyLty
f/H9tHUaP25wSXrqyhuaA4i2rDzbWofohin6AQ7BH8whIoLgrIQt/2+9FY+8Twr0Duspw5QkBT0a
VCyj7+SSb/qV21yWrWjp+QFPl6U2aJS4feNIwhgI/6G3aypyzKViCOdvv6GDFyPXgDsmbjhSVbNw
tIX3fqIGNvEOVzpYkNnbKZ6znbpKT2+Md1S9cQpSwGgxVl/iWkiIxgJ8b5s+EGxCOaUZgzv/4MMP
GoAJqNruMZfIPRhu05Uqtpv7ROSP7+V3epB3wXQGiRlbmGEjK1x+O08D5RaWgutEbkoFtZHH9AvS
dMHf7hQWm8peZSdR0eq9vZS+EiiHFuEfWE1t8B+EdqmhHkGFm6I0spsaR+/8zKl72kAq0jmeMezc
GnmpuviffdctjmndBobfzYA3YF3UBcECSSlxRVSU2ay1gb3MMPnK7FWAniOoH7VvLFayuVThI/aC
51NSLNgtScOk2eix8SZCANJVVyIk6B6imza1IDwlj24HUfsqIwCUv6SCBqi6MDcd9hx3csf4zl/U
0djt7lM6pRzDBDvbzqk7Wvt4FyH9TJrjls6uOAItf49+deqV+sKkjsDgAW0CWG93a91fVp/KAkzU
h16xkyK+ybDDJbSdVFcmREctfPchgGKKEcypZYaz7aUEhtUIiL8yShPaiwv2x/wkejk2S0iU1M7z
DtMn6vqNgtJtAP60KE6oBTJMH/TwueFy4/drBQXJRALOEi34OudU1DHiDlNvwMAyzVh30yvpGVZg
o2pl64ddXk+v9ZmWjhKVINJ1wmDkGCX+dEIqtUCzb2Mwzvifjq+qUw4RueC7VPNJlJJCysCoYHVX
n42A1EGMzgAyBb8CHypfRDCEuNhKiV1pTP+hClwbjrn+cqtBGTbk4+IyvHLRAbV+z7MEpQGHs8Sr
SbYQHcRsOUVZB05ZTRxgWRCySioI9A9rx0yGL+L6ngAkkcxK86KJztSgmHOs22AKiKwt4JKWFkC0
tdXMfiYKClkpCjEk+eXBoRYb7sM3Qz2HlFdDa71yehdMeSnvTgRpYCF7DVb+6e1ZHQfSMTzVvUcR
FFtfDoxmjjlFUihJxBRdgHDP8zXs3oVH1CD6scLJHD1zq3YzqUSg8Z6ze22rxtziEMz+8Z7M/vdN
7S30OphLaxH52D6Gkz/dBLvH9paWN89BiPbdQkx02CcHac2jHpEzFyDcROJEu2g5BpKsF8qOrfRb
0ThC3qUthQcRdLInPICqEsnxgIouQd+Ci1/JvkS3SySU8h0m5vmJAbkr3+9PPhnJbSiMlg9afs6K
OczZeKkRrGY5DAdmQ34ZIRqqVDNfQMwwY8mytX+7ojqA763Se8qCUpcpogG/jyeRnhGbcVYqxr0H
cZ3jDsr2B01U7+CDlEwqLMjMA+jzzvvfjC4pQxv0VhRzOVku0gWpKrFFNWFlN8qrg8mMzaxgSEuk
ka8M0q9u4q49Yfn3fODZ7HPGHDmrpwRgMD7hpI0mNeW8xl255DxgzZuU6b2YrTtL1cXoiDCv/SZz
xtvoZ/zVnet/LUtbChEnoUID0oILtM0Z4oWO5M5fF4WP73U4UCAEPVpbqPPrnCngJysrDM3DzdZl
wOaUmKYO+mimwF++vZAd1VCvNdDuA3gAI4edHj8NQOTzCItm7XaXBQpazdD5yoo5HV0DjxzpWf+H
zjXcn/r9qwwGGUnzrH1VGm1/aY52lPXJswg1fchXGpj6LbxJaJeL5Q2ZG2MRu6t82S8/gSIpZHKX
8PmkvK8fk6Kp0GpFbi75EUGYbpyqs2qQPnWateZzvOVAwhyjDJFiwxkiwXcIJlk1pKNzbII7+IBI
Zwm08Mk8k8AOA6OvmeVHdMwFCLTLiBgAp8jNzAPRE48pdoWzyigV/6wURJRlz8OxYxcfVvAyAx+R
6sEQKm8fDOj1VVIAqOmn6wkA6gNsHJzzovXCjobC29rSBYPQmLJuvEltHkQvMiHp86rHIJH0m2PI
R/LItb+OclwuVfE76zNsKoJkVvUjuY1G1ffHXzPYeYe4z6qITaESEE1JmKh02sh2ERkRYgE1l0cL
YESz/xCY+pM+AMj6ob72xXYztAIijcz3fVJT7xL3CypfZxahtXRLyqmbRe9NEiByaKXrC6AMjuSN
0F+rwCpLNeoCKpnVsP5SFQQmHZPAZIujP40BtrsTD/+24odHCFYKcy1hDgJOhq3B5moRsB6R+PEk
CQ3fYvTxo2dq0DOrgRKpB7tbWNilncvUPzKyTFt6FN+90rytu+j9kvAhG4Axxg5Gq0cYymKScP5S
Hf3SdDVYFWBE11EFI2/BVK8XmJEI7O2jEBn2KK8PejlK5vEzxVvAtvfyR35RfWO3XLGPSc5hmyhu
CeJat8PVKok63agYFjM4rMWHuJyFrED3GzMbucXYDicESuOCkAvqyOHE9mkZVvi/Rn+OuBQrxniD
sB6Pyu/8w/4LKU4GOK88hkXHYUD5pYvX9hAWzFzM9LG36n+ikJhGCV1eWkYPdmDf3Hu59PvCI9DI
HdphVy+DfXh1k68+UKx3O3gNcKuIZnuoK+fINBL+NHfKa/GubcgajAOzQxfqK2NvbDXVujKZVNr3
OanAziQsCzvRTg5BdQhM0F0qbwIa6G0FZ5QVJQQwb1BgEKzLH9RjGypiWY0+aSI4tKvBWfxfa7bJ
Fe6uAJR/TbmoUHuRMALIhhDS2c7o5jZH4lhLkmMv6CIcS+uAPHMjDpmEJHxecJzymJ6IM4v15hYt
Q5Q+i/V8aQW1mxOfmUfcLYL+E0CtRPBw8YP1bACcvbjBtqoNHRja0nmFqwsB6nFgSU7I6iSYAwDH
OAfNA5ZQRQEa7hMfDlz/DKRFfQPDz+vBZwXkygWJFSswD2SF9EHlUibuSAvJh7uIskQsC5qb8Xvh
xB5F067lcjQqD4HcGduRp8wwKYW+RMcVGYVtpbhAvas2OGUmBAxpYi9SxJ988MI5sBEtDY2JpfkK
N8daWyh2Ba4NhjE+S4bf44eD+wCa/gmF5nD8MtCsLQFEQr4/6fsUhyGrta6iEe0vsTnDZ9E29EY+
ORKAKs6WWPL5kqzpM0WZEwVLgJwhB4Tap/maRpk/MUOnoaNPAzQoNouO7212xwuS2/fuPFrrSksm
72JLa6z15MJuBK/bZw9GqGYv6YCjY/vcQz2qOE6dG8IKMLjwoPkU/hacmeQHa+MV3/CoPi3CJ58V
jPE36cTjmfb9G7NYTG+j4TVqEDUhobKsd1keJpegbsBd9F2lt5eSVB3K5d2K3T5YDmHJVGNzqoUt
sTuNvE4qqIkzJ0GQ6jYNWueXxyr6cIh/M1mUj60QjuKtm7tz9rwtAx+P70lCCYeBRu7XGPt3wd2+
OBBYVlUjoNQuKTh+xrBnJWSv9smR7UUcAEoeG7YCCCNMNAfUhCu/LJIyqisDKPm3VornV8RlyFMb
2+fuK3hh58wd6ZXQErUX5ggcw4ptMAWX2tf3hKC1tM/py5U1odXLU0tiIZw/9tyqp1PG5rq/9Zou
N2ifj2e9yekvCdEyj08zlwAns3e/MTGL1P7swGwjkR+26rK9B4P8FqgmUOFguMyTidn+o/DDd8cd
FzU0mmq3fQqcpG+Iy3wg09cv4fydE2hKjuvHwuWF7kDk8Uxfy76krAZNAO2ZmQUMO+l7JQkGcrlM
xRYS+NeMxkPUUGNLAqBWFLc5kuZUQoQzKc2LV8eRhM6iEGgdzT0WRTIZEepu9ECyCDPeiX8KGLTS
5mEjSnqz5fzz6BqlwJ+PxvzEPcaKhGDXOEZnlM6/zfmEoOajoW6/YcX1FeDmRNWjfcsPuU4EfcSs
Ub8Py5leyLMWCrMpujPbePqB8Dnw69OZbM5B7zG2dRBMBbUhnh7kCYScxEDWOC0CY5h+vWCvml3V
/Cm1siDBio7be6hmn6vv+HzcwUj5Li720egsXGbhBxgyaFwmwggsqmR1Cb+VQlGP2IR5DjPrXpVS
1V+gjIVUSan22oPaHomAmjE6mxyIsR72FC9VifW+R0yGngPaCdsbOVZH8Yqjwi2V+LlLeOyD8Us4
1ikgg56zjxCrC0ImP7dCSe7MQzsgDjHXj9f/QOQV7J1iqUc3n6XrL25wYsj926iIvYngUEaDOGl2
sQWkB7rQrBATpuEFfyask1CLt9QT7M/5fVy9o23HOnjACPBkTBl4BmJvF7t8mOKgIEfnRIeHSQH5
gYDLfyjRog82GtZi9jzKq55LDgQ3tM6XMaaxx+JYTq6fIHTRVRPkvgy7X65DKUtabrgJb2/aPqPU
/4462hn7+3HX4qZediTF66LRZtURrT5V7coW5dAoQm2TcxEdwXkITdx4uJZPlSf+yID0wsJZkvep
Gi0e8XNDxOXXV/vXdRIDpYWxl/gCwNwtqT5c4M169k12jCdHMIqDQSYTWcn6T5xRKGEkcQEhLtIa
W9wdFMhGb8wSeJZP7klEhRWCtooXHiS+AEiGb4u59PZDxUv87D3qJB6AXnj/4msUXL0+1BO0HFmW
bKrDYxcn3J8tVRUt/QWKqD4nSSYqH5czWop9h63DzKUcK83zUNbaCC8ITKWId9HFw4KkxauT4fW7
YE+jmlW6kfw8xVNwvojvFFbas66gNj+GrIev77GeE1EMjJ7qkDI9kk8Lmx9h2EYljMgkJcziAMMi
eYPvlm5QiFcwx/TbLo+ZP9YwehbI6OsukLEEJndLyEW368rr5LfdLgRVbMtUVnY5OWTf1Bgg6yg6
PTvL1pn/I/GBCxLTa2FgyXH86gg/HJsTPtaRegSzqbAzc48Uz1YGph506LPrZb23yCfMk69s/U4e
QP1M9aoss2d2v9dkfQxgcmgQK8eWg0JNJTlOZ8EKvO8pwYq42qGozU0dxxKeGo38RqqqxLHOns1u
wC67fR7ZudZbjW9UZ7JJoy15mlrazwShtz14Eo6E6//xS4s3OIx8ZWKEnFO2h+gvn3IohLc/UJT6
SKaueY9YarKXbGou4AW7NXKfogOvVj+4S+lrOdUD/byL0BQSVLwBiYH/9ToeZJz255/a5mf01acj
Swfjxd21dG92kfiLATZ1Au2fHVKIsg8kMKpmQwIp5sCcKGIWM5ezofHe50WfTiWvYRzuYT7OSjIj
pjRtji6731UZvUoqUI/olo2WOCqeJOEBJSdWLTu3Wx4TZpKKHVDrFMTFdE4ZKYYVrLxB9ADLafHM
We9INieTzYYfVlfsgvoPe5Vl7jOsEsJ4Fte7hltZhDNl8qxZU6H2REdd2mfe5UlIMrhINU88QRwU
H5YOlqhHwwhD7mtPrCzPtBhXsDwkFwU0LyiwxxBpxp6u7TiakeVLQd6nD+5mCryaqQFoPxanHkuj
rtJf/TtAH2FYaKYk751d6VrWnCkCTFNTRhmS7HKZEugQBBNpbsWEgSvvENO1tSU2NwYNk/7lP/OC
tJtL0qVCcxEK4lAOqk4D6rAiy1KTkR+Ekg937r8VP2M/hxwP3aafgWF4DMtQwMUcIuyWdmnh4T+K
PxDz/uTkaVle/LukeVjHIeDGmChn09aky2yhKyYjHagOGUX39B2C0NX24m38p0cw1XPkoM6n4XOk
pk3Fx0/ON06VPt8EK4B8AZnRPmQpX4WwCTEz4HNkVxI8lGX2qO6NH4wjBO8vYDeiLfrDHPDtaikt
MwR1NkzeOKT+2uVRHsTa16MZv1Xvroelw62Pqfxp5/u4Xey1W11Cp6FQW7nvHPqroGPoHELEop0d
TT30o3uh9TQ7Iscd1hNFPyboQExeKpWSq/9LBWr/4qH4T4F/sBoIhlysqFHlzl3f4Q+XwgS9ac4R
CsCiHCD2rDziuc6K9QC84ao9SUjMWqkELLJYN61opB7n3R+Fdu70bxz8xCEEE3Pp9/4A0GKtmGyu
QU1maqeQRpYyk5Bb6h9f6xjuFNeyij2FGcuzetRuIkmD5Dcf8c+fmrLrYABJCmFMyaoM0djUcRA2
O5HvX0LNh/Ecqxw7+w+U6F6FaQjTE9xRvYyll8Yxh9QKEgl0u1cCyo0C2ITB9DAhj18qqCRurDuU
czE/jP30W6zuilGH3Zx1wDswXOsI3gpDOQLi9p74iFd8Fien9tQ7NTof+QQwZU2KD4/6uKT9M/CV
yJ/4dZdrYA6meNMOxemjquUKvSPuiyBS+vigTBMWdjorv9WNFz9OQrM++pWuPSyG7GVYs88dtlDx
G2BWyvJqBmE8olISqBF8MF/FF6irCPcHWSThnrRj/7jSJQJcOAZdhtD2/tIfveIqYtBURZlFGiir
N+DlAQ+l98XgyI9ugprDSROHXGu1BPxwmiFnbWn3sILxfh/vYBUgGN18tZKa+Gi7Fdd2Io2hae8J
1xIqOr+jksmlFNLp6LxzAXTrnb2+uUkvzgHvc0LiV4yNu9dgNqHE0/N+81MZe7qA8s1J2OA6rKLa
BCT3cFnYUnOeVF7CuPbSRthcAPAftFlYUyWCQax1ZdhFwveD6JT3MbZuG8LHSGYIpNdJVzrR+ZMt
94FIn1RRx01feBDtvhPb1eM9jFge+4Q6So+yIxMLMmVlHxT9I/DhMyk6rA82YYbOa5ncxUfdcMNH
UpRZ+cbWOBkvCMUboBZpTdGfO0+ltBFbJNdK5aSIFEovcPVTuyPRueKeGjRLCCzCBhC4rNwfrrrj
mIHFfzGPnmUGVnntDz/eBWo6G8288PkN5EXXrdpKg7+F2OF7O6Cqa17BxjOHXRFxB3iqQSpUqf5x
1W4B6nXS0MiPXpaRVrw0b4HRPLMtY6HFtz3Ym1u3orCdBl8i+lAM6/kUt/1rvFhlvZda96Ho0efN
S8kXomMbyhkCTch1LNmfY6AL0n7N8m2hfqNrKpNLfQ05gNFsArQcvd7a5amnhobcmkCz3RMsto7L
BPS2L28In4NGWLuY3eVFW3njEwzBL0MPmrQ4WpY5chlsfZyKE7nbtzNpFe/H6AwRvslrwKgV9mvZ
A1cE/W8yM5ykG6pB+kh19QxoJFjApC78ndN71W67bfbxLA5Gb9Ub1Y8ArS22KKc8nH2uJTe82EPT
DORsOdEnhI19xIsRsqBbwpYPQd8sUMXqsZW1Uttkbhm0QxDA1ntHLmOWqi7LuZ5tQw56ZFXLuTG7
4nK3rBkt21BC2mrdl+0ZwSEM3eJvs4qwJfFCzs6KZMheeIksh5iBx7u+Js4/vZCZJEl9BuKWIMvW
EvSmoPVJqYpU9KYRWKfh3gLs3poY0+bLK78zDPDdvT19CTPniSQjY9OOHvlbQOla7IMN3Xn9QkbS
ZKk/6biLphqAMofXiPnnayCSlW+6F6RbzNK4Hwk++mIg+Sw+djwGvtsazfoKlPDYU5hV2KlflCxP
xAVlAUWRnqCNDtK8a9MBjeThixykRHAywZ/7OlNupoQk6KLoTlR9CDjEUH1PVsPnv/kuWIG+Bndf
mW8O/HIFwfDKZtQbQekdirN4SD0FTHIdMs929L4cWzoPzDsLKqYz2E36fBlJ8GTs/3H+r3JqWTvq
KD487LXRRHAPx0mm1aSqwUJ3nhkD2z1ED/byWo7bf//nnicaph8InTapShDT3CuxXf5dZ8XNdP0Z
dYY6Ml7rmBl/jc5FV/2/yowLMcGUwIRVzg9AL/aeBtY8RFSItPWsRPVnVI5r8eyvSXOCWILcJpEJ
fZb/qOfpffCYREqcaR1xoi7I6J1LPxxJ5WIOCbZBlMJMLD1q0wlClXb/DA7TyrY0ptrX7NxK/v1a
H5Gq3kc2p3O+3wUuf3vQAqnlHPZXP7/VPfh93SEKvmu6vdKJ2I06T8FSTL5BsB24tEcE+yJo2c4N
Bjc2XyJLo0n/Q2FsrFMYvbFCprXVkPYBcrcNtUAzHhWJDkSZug4qksoNCP6WiTkxv5Qiv5G3DmtL
+iDGZpz5aZo3oUR1/YbR0My1qimxwlJQyjzxcUoOr2SBTLs+uGtTH1GqizmzCXbMdzREMcqhF9wt
/I+hgAMYoxNkMBYt2j8fkZSYl3Q/rqihSP2s50rL5bXnP88+1OZqbKTwP9JWOP9eoC1N4MnLks9w
WRpgL+tiHu8GeyvZalaCtkd4T6ZxQWessR6hKK+M3Z7JUVfarBwbGlThuQEx7CCLkWZQJ8GT3m8O
02nD3hvQUPoUUO7EKOvy+yNc7PB2xURaqGHMSrS8rWdl0yNwO0tiINi5I0p5iZ8jkiXUxzBQd3Lm
lkaZW93sQzOq6ZXmz2zISRgXaWcoxmhcI3vuu6uODsDIIbwlcH1V4cQdu5EC15yN1EfYTxnctccb
L1nAu/aXa+rOpyt6DGDaZnEIZZNcijuuA7BKQRk5AMlWds43E/pYvPxuBpR35mWyVaTiXMgJKhiV
9/hLjXKvc2kVCQ9Mt/0zXBxTKGor2V2rFKzi42xwxFORuMjTmxEmaFPpqdEvhSJmrSLmlM60rr4T
ZUGSMlZAJXWIPegHqC3Y+Ok9f1TJ6zOXSQJFY4RRuyls2BrOrAWeJvgSu0dg/t9+eKdEcnqUtkY5
KtgMI25PztgIsjYtHBSSt2LPKfbgQfTr0LepyX6n/M8EBXksgI39kTC5z5gOqUP2LHigjTbtBWmJ
Vzlq16mM7sDbU1czI92zc6NstFIuh2BDN8w8r5mPjPlwgHt7894bF5b8dwfS82tGl4UrFh/KU1sf
8nyPRXJix/axguzZKI1Vt6LCHbXkVq56dznX6k0uznVRmwC0nac0E7YIQTFvpPadJgscvTWt4rV1
vPV9Rm7wcIQvp0XvfXhKnswK4MeHZJy9Z0IrnwUYO5mW/i1WXe7jR2A7X0ecb/fN0V0gq2jeLftS
ReNWt1Qm+Zwq4ui4KO2UL7tEslr8MLchgZQtFTbH55kHE277g0k2Lztt4ZVxWrnIUsFsWrDD+jUF
mmK2g2NGwfxPfL4hrxd5mfTejblJxy+x91vMGjUcBVsRd5jcmRSzmjKmQ6eM4UEP/K6Btp/Dsuf0
+b+ppkP/DoWPS24ug01mJzSFaHAUxM7Wvx6bXJxQC41c0rCIe7jQqTWO81U3TSCj7gRYxHWODaib
Los137bLsYXH0AV4moUU+1z8Ue98GQ+ncW7yscRKB5USJT7GcfJSC3ZkZN6kkE69r2z0MTsSvKOC
CVKQU/iQuDgfJrYmKmzQHUBmpT2F5fUmC0aI878wIY++QRp15TCfR00Idycr4fhxr1GL86TX2jFJ
0ZlEk7+oT4kLGGI+jUMARElcPjcKuRzP4xo4QY9afBx4hDkex5tlLymy/XNouNV9ARcJv4Nzu1D2
+PLrCF2WtRUiwy+btt5Nqpt/UKRqdWU/jlIkTqQ1gLW+TgNQA1M5XFzERPdEs5b7jnZlg0Voh+mr
2g6xOQctD8fyVLPEFp4TrKWi3kMAC5WrCSRMMUo6VryVRsDdT/Sbmj3ScXKcr3ij6NNSd2pbioLC
tXAHM7+Lb15qEq4h4ZbCpLPOr/1r0FxY2m2UQl7aE5+XUZpbiunY5asgzvlb4L3DHrARp1oM0GGO
8pEB5k1vdAXITO8Icp7JKXxQrvTrENOSmT1m7xUhTubRSQ4WM8YO3vfKMtP+/Y8r/p0SCEJukA8J
Q9Wap/DWCpfgj7ICVFB8Lh3OvHSCr4dT1fgOd0Bhyj28AF6Vv9RSYLhyVB49nLzu8tbA+EWWV9rh
IoSaBK/+X5lKd5WSYfqOo0cRFmwbKAwkq9hIRB/JWDoQIWrfNAJiBCe50gbpCRt2MIPWLalBHkZ7
plRX/vBFBYrWGboA6OK66mOPaKQ2zfryLhCwOo1VaSpdbNaTtKCltK2j9iESvYp39/0Yo92knvwj
nBR2we74MSJnLKkp7hI5YxhQ0MPVUFnf/EGyzUSOayJjTAoIv8ABeYXkjaeU62C/zilealPx57Ih
BDUOvcOrshZhzQ1N3tS6VFfNPqhTCHJIIXYufQ0nJBqU9r7DCY5BiMKOtiJ4nxAqxBU+1W8K4BZb
60UMX4o8Y98z21/X62ZcNcdS5rxasZRrk2qR/giDEqBgkyiEWSl6h9nJOmAeqoLprJQCrXWk5LhT
/B1Q6PyM7Moibg81IlPm4EJbUAkKM5Fsnt1eRMI4Ub9T3E8P2MMIRKW1HI5Ag7xW2mJBI30Y6bRB
9cUorwWO6doKQE4KSW9GT5nQeFFyeasWW1LkvEwVGuOFhnHgiZh+0sH8u2WIVkTn5VVr3DxqjHqZ
gahoWOtlfyoE82Pe+v3C70euYN/DXbdfI7yRoCQvc75iBd4SSdYLkTAuUBNdajwVt2w0yZiuDvGv
mdl5GwLFgghHXMNabYt7AQIhUBiGoc46w7NwgXgRmjSwMMFobaEOzJ08z7/XKNVjwzXY6OO5wFIt
248V9l6k2oKtnS/qlsgFEYNJtYn/5f+DAlzbRyCYD7DlSsTuKRBYnelsoO0YT+cxUR/Itpe6GYgo
FUNnmQqUrwM5oNU1oOXSJMI9w1qh43kTabcnwvOPfj+uWEH7O4PlJFzPLFuZiTHvK5LhwWtyWKNQ
h5T0axBItwfbxR4iVR/haUDNGgwBPz1CUfXvBnuLKtepqfX7t7oyDPKUxcC/bTffZgEsuJVSuFuM
rRjHpNSe4I/dMbggkqUBkBtL9rAT3N7LKe8LNWHbgz+fk4bhCy0a/iR/7WOD9Yhy5w/2ofxjhM9H
dd2BGUZBgG+oTEZbGDSkpEBjAsmRDmOmv4tE16f4BKrJN18YlbqaQStQNsvz7OgkQazMnK2b6EA5
mK4cnL//WqjApKHBsM+BzCse6i2hKSUM7ikZKybtp7dvy9XAHgSV78no5o/Rdm9HdjLBMBKoSS21
UeBHNbH9osc87jugsbEn7n48Q9nL28U4JxTpgpCllho85sIJ5sX0foBH77n93/fkmZh/BWzr8ebm
XZuzGlGCQlGKITA7aTbJzIIkr7FzSzmHEZNzcXHOtwhCsjPpYU2YkLpmM6dBF7gG2DZw48Z8heuR
dNMEuvoizgCgRqmB/1Tx6KXQYo8yUxUlhwegsAazhBYjHYnXCFYP3EakL91YYHF4QHMZQ8bReLya
hKVtoeOyvMrsYLRcsput0YrNamBjReb4v7s3QUkluNfyDYMdYIODunmfO/v/2x7zQVGlkto0zvmv
adOz7yS+dfnFZkCGeVMvgTfy1hk/DtWZIDNg+t9ZmTv+853XgTXuVrOnK1Y1q0n5WYjv7n0qjdut
FaRAnD4bgdV7QktaGLwo29e8a5bAIy6ah1Zy7QBLmPbv9mHeO5NRqaTmZ1GKs928L4vtCb3eIOES
AyyRsMQ6iYqrveD/Zzc8voYs551hgc9Xd7BZzoysFqnonB4mtA2ASzQgv08j8cLa4eaJBCVImO3a
gl26yPPCHV59H/1Xw5WEJNAOdHc8TT9rx/s7UUGShNbClMLp59Pmr8vkEeIQQUS9gNnWfm20Qj1u
L/IrvIaQeiBeps0lF39YTl+ssH+H4iPbLqYwjQiHOANwhH/JucdjFw5z0OU+EUf3qYedM3wdzI53
q2sQzSKD5Kph6BKUhXC5qgO4qm4tfyE1gZlmGbq5UIeYYmQ2ATHsyZpydQ0sBVfK3Gmu3xQS3IMh
LR206KFLq5q5wVWbDO5iJjpwIsEJB4Y0Y/iDovA+f3og4X6Kkz7PHdovPf/e7oo/sunEDEnNzsw3
Fr43v19CFxacHu3p6nEL4DkUKzAM1elcz9H2oq46pgk2aZW507E+rRxA4RlJ9JJZDIiVapORUnXL
qpVvuKxhVw0Q88Qn8HfTMMqfgEYELkdSAm/zBjeoblWYz/o+n72Iy7g3FpKHR/dl8RHPYLQyGUZw
Hqg7E3iWispUQgkGO878grppya7Eq0TdOO4gLd3HgtnvdFjPmMQOXTCPETdk/yRaphpAmwNkT67M
DZ1pPm+a4g97+l/onRHygjdW7JvREhnVbxZ96VSKvoCmneaC5tiNVuJGRt/gFPExx11zJ4dx0jje
XHRGu+2DBPhhGj1qxxmeZAnXzzQDzn68TyItX2kLlK/HVdxhBkFZ3if8HpluRxqj+E1Bn3M+7eGx
lDtVwi+phGmSJuSX5/MnNdYVLNereK2K/+maYrgcdSW8OW3rq24W7ZXQlmkkwmOVV7Vlu7b4N4fE
smImxDnguQLQx1J556dFAz2kHdfqwGINT8WdFVLQAqMmkfAx/Mcy16Xtu2cVmVyvSMNkQBapsMIB
K2Ybp53Fl6dSeP6HUtbAJrOPn7pEeBCflbDSNhgtlE782TY5Du+HsJN/LLdWL14EJUcnnlIylN24
sRI3xOCIWsPJ4FJifsKcVJStNWVyQG/mckGrFsB0Ch5oEr3uQsBPtK0Iud7uS11vSbS2VZ2TioGB
+Akog5xkL801pu5ZfTwEduESHh4/1EjkfCPYl8uw8SoZjPb+12EoQ3KUg9g7I7hKrRt/WWjidXCs
WRPouRxEe4sijhFnrHfC4CUsDnudZ2adZejz5Rbi41bIs16CiFLFUKQAAc4d2ZhkLz/eOqMrKus2
4sUBrLuTycXzuV1D0ZrZ7Hx+v5FUlZCImX2RuLBjEb0K8N5VrbcHpLb/9zGkNgXc5dZBcUeWauP2
o/4slqeRnDU3xFl/kXWIJLuQBTiH0x6Wr+LWyoapITG+8LGH0I7ZCqMw96evFnGog3Wwhzh7b2Bc
4fb0TiNoFkI0ZJaP/iWYiVigecZc1Z7yITLsxWOKhbWM05C/GrIVkRDsfXT757lGyec/7W5M+JG+
YDSWtQ1BQ53PTJ/cdYZqClC8MdpZnttI5XqeMzOG5KoRqqEC6ZM5tzHnAyq+ANw3PdN7kLTsTAIH
XcEq7AllVcwuGp3SfKCzujuEkC/iMDh28G4f/cQzVqMWWSzpCxspA//E0s3qp8RDcVuApd8JAXxu
AxMC1g/cxuNP939IyEGkhSzMbNkQYWoNURzJGtSZOuQ7vD8zdmn6RiU8yXhUsR7X5Y3SRpDbJmNc
GjM3OFWCLPuI9rHHh+pRSfRxC+PD75XTmVvx0srgZj80qlZvElceWxo5rGMSdGFtgwlaKRtELLQB
FguPDzB3t0OHj2Vnw6eeIdxfm5qjTtca/bis/11t70ez1JXSamlaG19xba723iPfE22I4Zc3Z2Ma
TTh3gRXm26mCWglaWkw4tMfVbE5uHcAuN6kQqPz6Jf5JwZHWk6Ud259Thwx7qdeXi869yTf5YDkM
4jUcoPZ+LtRYc44cLBIwPobW69O9PjwiZG/kfeQhW+YYpPCgBXYhYXx1HU1ynhBQhJf1PTzd/P+W
znt01U8PDTgIXlLMOIOFPKRIPSeaaYkcS9F6CuG1AXYma2cFnF/hq1Z89D54yOIhxK9uvJO5+QgC
kAr+8Poy9efOrsp4mAGA7/Y7jxOGnUcpD1x9dFB98GxQ4qvjS0hR6yLXJJ4I3043ZPCArNQiFYNu
0ZdCvtQLOjtnP3TWXSnwEQbFVcET5wjSgQuJTfYsPbGZbx4Eo3pTHoFw9fI+IQfK+W2Bxg4UyeZc
BQVhwGkpCsV1XUr2r4LI3ruCdBwjp+YpOIIIaBgxjPqZIzAD9K9f1SDE06Yv9O89r4ER+ymWzvaq
A2brU5GEc75buRBYdE15PtbejgR6664oTqEh/vAWN0cJgLa1KJgW+OZGtXW+W7PwN2IqgayTBnJ8
d+KAPqsXAfUY5nhuNvm0UqPfh75fxPgzfXniSFZQrXLE7KCArcl77ghOCkKh7tq3OMblhqKdWP64
YO9SXS3fhhMq1iXUh0O8cepadmqElb1KVflUwQ5Og2AjWtstObIO3D+S+Q/ETAzs0dx55zv7quhW
wyI8AYzI3mQ7ByjLzeeCC1+7v8ovsLuAzmLlbFnebso62e4lt4Qe7Ky/q1RYqJpMspzEoyuSDJhz
lS5l6VIPJIbVnJsgLB/Dc/d9WYzlonICX8THsw1YRDOBS6Q1Xpq9J3KldSwXfGCwq8nsN1e11hzy
M7cDF+Gb9HBox9ErBZ2uZ6/22n1lmosiLbmceSCuSOU8ARtqKH1jFoQcyofH3UVOKKD4R4/yXLh2
p8zH6Q7ODsmbmZ74xVOwuJGpmiHOTQOcAEXRhCj/BT5kRO0BwWn8oGZkWp3+f89iIDpx74hKkeaz
ekJnEk3AwxEMQTA4VWrz4grK+ljdxZUiunNEZSQR6Sw2Y/kaRZBVzWta8z2LoN6KBhRtQDl5uT4O
6jfoi1cqmdDA7hpe39Qhm8Ia3VwWulhEarBfg2bHCuRAqXuFoteDZkIn4YPwBayEbLPxFL/9AHim
fK/yjm8SpfJ3yyItJjOY44p/n+jcnAJ6Ya5MXyIP39FsJG7mjPeOKN1X9jR/LAN+SS4DYGbEV7Nw
1VQVz5hsU0oAFyCh+pL+NmDvJPf1irjGJRfXWZeAQovmQptIc/HZzoigDkjhM6g9u7g12TscmVB0
W2sAb1DtKJGT79KgIfNhWRCAEj8gdMOgv6/+GTb+3yobo9eUgkKYgR2r6i4ogWSQ/YPUPlvwPy4v
wz34yM6bELK4zvyTvLpq7YSgPV3bF+YuGSwxdBFJxX03nFTHbDxDgT2yr7I9EPWBvhtJBT+4p2Wt
xDUcimZDwIMeVT7ZQdR5XpRlH4m2wk6jHD0GRrUu+H5hpKUKZX/HvA0OSM86sAMYwHVoLl92PlmX
hTFr6hy54WokaOj414tujqNPp3S4STA1Up4cD6I42xGOp1vJU/DoBEZPt2muN50VEMbJa+ohfeh5
waNKqH4UQdd1tmkBJHJW4o8jKyHVqgCSj44e6yx2vOBKoWPuTPgdTzCYbgdtqmXMcbYOyfbyrQO5
+ca14SwGPrKwppUnZm80NskxPq28DvZxDXwc4++jBDskA7yoGRqhmK3PInqWAv+WM7+2DcDQDnkB
MWvZo04icN8Pbmty4UhIvuxrQUrto6O4idVJkCn59fdLDs5lJfHgrQHz170+hQQl1Te+h+Ip3uw6
n3YDcA2SwZKB4SONkFjdlvwDqIJGslikHvPhfBGFD1u7QSxBBoq5MN7Q4rkJxPFEUoa1k7/lrL0+
TrBDdosF6qJnVveV8MogxkCOb7iukX2ylhj6riM+1uaXJNM1jlQLsWrt9T7ZnR1van3PaaZ/gy+i
ebkcD/zTyjdXmm+Z/0oGMQxN/7gzOfJMmRfHDb2f31ponHejHJhCMZ8+SBAAA+8bLVujiqfdwwW3
SZt5aCKCNhVoeuN85BUuhli3kXNvfSYmwHrVX6Q9lJTRl6S3h8T+zlUrmxrzVzUXQZ1HpceQ3H3P
si0nXjygw3s2q+JFTEkF9xWuNiHxUwaySXST9NZqr3GQb14OEo6gf0Aufw8t1l+Q70qIlo2+8qTI
ve8J44Nte0jv9APDO5HzEC+qeMimnoBW40frTmM1jJpVLBlLm34Uc/qjccvDS3R387QQHZmBLQnu
a7MCKZKYp+GfhTwAKXWEpDBseGfKjchnAWLhZ3lWRnEpzt2OwlXZ4IMJSmik2QCGEETDMQPOHcka
e/aRsDJYqRJkzbPjDGDFx3/crVRhOJNts0907//AdWAeL7xpEs/9XICuwGOoJF5MGtCoGShaE/1+
jGEl7kEevnV33e/PuqawFTsYbItZcoy2VBFjbxggDhyqykK9l2PmJEPyqK2apaPwtMa3Jp05vqef
fNWGN1RXqIne4xYnDX5wgSeCWYsmz55hcUCv7jFiNKbqWZi1GfTFYl0kKwjWv0UJm9JzNNOb1lqf
lHGWDx7DomUorCwTNLJW+3blntW7T2tda1caAOLzVSnH1HOhiKoHC/B9OmQWHEJUYQfPCiOTV+9m
TGNPLHxGx/rXpqS8M3nuZofHqoCadp8vENKrpXv8ZIJwArsNSwfbN8GcBqx1ZvECEPXv5tl/DtNK
Tk1EAkKaSLHKcYmTTQarJEbTs5695/9Pg0uod9Wil12GiebdKbJrlzlH1Jwm2vZmwR85wpkJYink
Cs17yAHAfQMporhWDINLI2X+fHTjp5P2df3nnspsGY0olRbu9MdoR6ueafWJx3FnPeqHjYNZNilb
/E7l1NK9NW+lI6Fmmt1812iGV3uQuiPNpyoN6xB1ZLhj+oVhMf0uBtebGPBBaHrfsdVVLH2gv3yO
HSuIE2L82BYD/uP8kXDEUC6c5bSJlnZ2muPXBZ3X0P5DXFzg0xcxNlSy6Itcy9cQvmPXdpuF82xN
8vgNDBqCDup0Be1qX4/oZq2buyXdafG4jBce3hzoBbzWeG5GwB0JoKz8vCmO0w8kj67k5Ob4BRyj
Qzi7izJ0j6vZIWDjBXkHkfd6Nv8jWhPJXzEj2tRzjgFSoJdbXLRMXFWq+1Wvxm7jNObBh70dyt5v
HBYQhyMwJQoVBCe44p1e2dPfyDGSi1G1IJkg3RJBIfaoBbJuKoiMmOGdvq6zcdT6mNLgJpnZ1rMv
jMhubq/jNZEWsknmKrt1qcoyfwP0fEvwpsaE+BCEvkbURaEqrqYnrdcbFiEsZtfUcPyJB8Cotx0+
h1mo7HETGv4snejcWNd61jHlvZ6fNFaSYSEGHVJstoAnQLvww7rqaOE08glwdjieDzTH6id2MaSA
QD3mG8E55F87uFMz63MyessifvPwoSOi5BMGST3pjYQEN3EiTEsBDHexPMpDXe3c1Y9xDmYKjvQT
QN6yToTM7yR/HA36gr/Efsa2UsEeQdMslVPe1Sv02pNg1lUxQAQmBgTeEFlSGtTwXcPiBllFcNNH
om1kJCXr0A8Y06Es1yWxKIPJMWhLNJUglQ4N/0A0puBZ47SJw38TEaIIu9e96sQVkwjmd960pYFp
QuEXTpbCwyULsewbUE+CtaWcpMlc0f9U0uL7rdKHIxCygHBDjpjoaPztM2TEwLdfIyHxGnMMzi0D
8Ge2gyy4KN8DzhLZEKIgaNpn9myNiFEkFSFspFqGFqv8iZuE9D3KDJQJg0VK/MaZ7q7NibkvwNtR
FQyZgHVoXHnz6c2f9ZS1sLtkQ9EQhyL/GTblyot0p7/7wDG2zVhGeRytwfJpXncxZ34WTfwu7Z/e
wN196QERC/pxIQQ8TyrMTSyP4imuZbbS2tP5fGjl0R1DQ52I02VP89ilLcrSAXwtEkREQokQ0a/C
nJ2KwCBasYh3os3KwfMlQlnRpURj9k255wgBbTJWP0JaahvH4cVkupI2fQPZlWU/5XCoux9NyQ/s
yP9yx5f+yC5s0jpEaxtpx3zbVqSkaO42XFSazR2sTdTinBpee5jLQjH8Yjxhfh3j0B4P4j8HnJdl
4RMk1aEm8JX2j3GD3sCYXkCHvnzDCzBgS8Z+EyFpKZXCiOm1F3TZidjzl6nTKmCVKPFWiZ32i9eE
cLP1lNBL4WIWdWqTE6IgUGJDZMwNHbyWba/MklAZ1nAcWi44v1j/kg1KabjNAmcp7yXuFmn3OPok
yQSowCFR9bm/d+nC1liVmipJKFNX5lahEXmcEIyMS8Sb3JnfwXycmP4QBZzkNYuIbqFUIZCu1CUe
IM0s3KdaLqarRUX8zbcWwRA+hdKGceekXrBxfEaVNsclTfZ/9MycKmJQOxPu8/wVSEcsY/jE1OgK
Ofj4hgwZQrglltMdzODzZ3Gs9XTRYZmiEuWI6AUe8VH9W18EX+RX7XQndxgRE4EpYxKoMm4+hLIT
b44zA1YGYT1muIA/NsnDXvoLrkPCUzHH9FNQdg4qopJAIwp5vcDTNqVbHdsIUn/Kwlkjxy0LHKZh
tHWDoKy6rL+eDX7r+85lATF9YiG6kGCdZpCpBKquMlTNslTN6RpP2hLT2BY4/v58I17HldnpTRNa
V4850uP8AJBkFdCXvI2ilkHvwV6E2581pwf1wzcUr88oECSkMn5vsmbItiyYAqQ/b2HRzXCJvu6q
Cae9qxZOVqtbL0LQN7ox1ImiUC3NbFHm6kvZc5VR+8i4SZPya7eToMWfxtnq/XkjCBzCu+HElvx+
uW2yGF/Nm7vb8OWk/p3Q0l2R9gmqA1NMQ117ckDl376Wuv8uHnbBy5KTaywRKXn+GMz3XKgblFYE
NvBOAXYLUS7i55gbhCtMjBe/sMiA7OSJPOQ6RrV1OeZE5UWMJfhAE5c/3yqlgKtwOkqSUGCe10jf
Cx6ubeO3SzgdZlpJIWlBzlqjfO3+bVlaYPuW66/Or/jdKe3zv15YR//7UB/9i06uDWu6U7+4JmBK
zRu9PLucVpIlxkJFMzaYV5czoOGdY6XXiU/agDXQ4PDv8VuuOdZGcceeajZAJySrCS9FxR/JUrsT
gMldrEzT7F5Pt/x33JbzySOEOK7mhuiF1oijZh/tZpudntp2/f8IdDX6O3P/nq89QXNmkk5xqOTK
wIHt4lydnhMCy4RpT+VDBvc3Qj3tbfYL3bILcHcpzklG0hXAkbqHCZz/YEwB1bvvM378zF/v6vhr
NQ2pDQMecuZuXSfaW+Ck/p+zH8xfGha/hydVanz5eJa8jEVW0U+q2E+0iP3RGhFWN/Iri17PvAko
tSs0k5hUJtmxFjxFBGvLtnuRKWXTYaL9uF2OdTa9j5Vudmkslc0dgOsOOESDnGVOa8b4loMMssZ6
KekC6YAvjiaPpGOCayVro50VvTxbefNxkPDFxL8NjSlBFSlNX5Ms+06Jot9+6lnUJywBcAkb56bm
i/dNlsAVR6NB9PLXexJjafs5qCwRrhhPUu3nBTL47PekZCFL9pW0sbrS8+/kgIro9cmd4hnSIxAd
vbRQ66KaqCLrDU30iuZ1DaWP/qAKu7rLYhblGtTt7+5ZX0hA5UQmUdnER0zWW5vFmgo0WrHNJetv
6pg1hRHeVogmxVXeQUspv1y3WgVT1qOapOtZbV0GFWkCwUr8m+DLvebJAmAxyqh/d6SQ5Q/tZdOg
FHXsBFNzWLNYG4fWziQ73UqzxEDUACDZQUrzE8eILiD1GHhRpxMkrcmkaDweaEIt2QhurCl71CWI
6x6qSpSFCC/LQfNea3cScsY9FI0OuCCcaqrZI1mxl4f8zB/gHgODXP1RIlDKe8StjjSLNXHbFbkL
lk4gYfN2kJON8cQrnBGS+AYK/NdiDXxj559AgvXEjv5d+JyxZLtlt5CYd8zEbTx3qTssCI1/JywZ
B8hmmB3hOdf/5CtDQgOOgTmydAE56pnGwpqQLZLmCnifoFRG8FBj0c7lo6zyOsHQZU59MeM+JPn5
+PIGP+VZoMo7WUTK54lTwlKnexpMKpseplvc0bIiV2+R9C2YK/fKWWz5wqGFqE2VoiYaayyOWTWl
F3+dZlxascwGCTgJXJ6uBAjS/ANJVGpAoP4lL2PE1tbcq/Bs9tfE/W5g6s5+rhGuIMXSG57ttuKa
hXx49XOj9nTH81KkxuaFfrRM72OQ+CCimI7lCqhISn1/ivdDEBtLaT9rb7VuimxpAHqTuknVvJDI
qCu563zn+cLtANzk4dk23YQ0iBuaBY2Jq7444jgUywiIirF3ePbpEPzKPQ/GODJqQyWCwUc/bGOM
u6GsDMFWLYvOxr6dfcxP+eEzutw/3COlE4OZifdGnOvfUQoHFbSI5x7eqjLYEr4Ce+t6zZFNsz7f
suAFq82+7DpSzthd/KTRgssrgf5msgNVQp3Ef0zDUnn/+34ScWXO98BUdhaFCnO8O7kursKg3xt2
PgRrBAEhzI0/urKby8BwZRn7sNda46ZXuRlYWUg6NIpdNBzzcrFDiNVBc6ltcxqVeC3y9dfnAZ99
/lEHQeMfbCs9kmkueUW5WiINsb9JBkqQqdnLHykidxBf6V1SZQHFikrMOe9JW06zqeWj5MArmuGl
ZoBJ4QfCR7J5DqSKIPhnmr3QdUSezFSZzjl1HzhH5F8b5AF0z4DYtxltls7m4QZEwKMVx71yAN9p
xP95xfDAhL/rmU7AcHU/Ow8IedrFQJ87dmdhCR0UzICWsTqTR3oqg0B4AycYQ+kousVYMSmy7Lhj
cUR7nMawzRoJVY+7twzjRUMIg1v7N3kdryvt5krLYJGoUeXXEx65xiqfYW1zTBEmIJhVxHvLup6t
TbzuAzkcbwWtusVeBJFkDuAngPCehrtCJLYwjM6UsbmwqMRpYPWZwBO5HIevulG0Kkr5wargpdiD
P+BXJsP7qF6As1IWVVHfhDCch29vXdbZybDXkDk9TbV6H8pDEKJy3ls2/i7fOzqIbcT0UNoPvsUL
KRERzJ0WebPS01vteC7c493QY/nAca3u3K17ARW65SEoRhnQpHjJ5vLWOC+UvCIU3j6mnZO7Zjns
PzeqLn7JV1CG4zYsShSIV6QjomMGppPHQJoH+sVkmIa0ZwpeKwFgI8FWzUayPuFvBJYBv2VytQQq
f0Q3x8Ia9C5vkM9o7poShPqT9vRKYR5Vw45wLRcWiv7Yf+uYFeEJoKRUq2eM5UhbAMGAt8YhdkpH
gjevNT4F2yZt7SKY+DRfdp2AZLR0v1kG8ItwE3rYW9t+pM1DPTyIOpU7bRMsUAO3QNhmT4vSgjsT
PtG/NRY5S823n9zaDzslV3hXGxECqF/ep8pxNdsS+07TkCK+6A0OrowD5VReRvF2Z6/Yo2HwYkgV
ULfmyG9ZihSBIBmWozJWcWoDX0AZsVLn3Bu7/ZevSgYcbvYX3NIrYQacgiybG+N5NdkLt2SBb1Xl
0RSI53EVwwHc9fdFiM9ZoKKbvLR1bOwlbr25ugtIjMMV87XBYCfR06QkjYT6uTgKHQ51nyQr/ftC
K8tRbUJ4poK8ZA+o9qSccajNuWkZBHdSKK1F8SIncpvm7Al6F8awY+cvlzlnYMoWx9QzHFd2ni/5
fb3Jz1Wh+ZRPIiTUvlMhATQqaRO9AhoVnY6FOIvC6MCMxdG0pEtZporqz2UuY16NgEKvFmJGT6vz
0N4RuZy3aPQKy8zXC2GTVwRr0CjLFI4HTKNXUDp7AqhWRYOIXAkMRiT2OEHqCZnA8xUH8WU+aTxB
K9q//VRt7ka14AyItBOtbDstmxYErgItzsd5P+8HBrFH1klfRo+/eRpydgOwdV71dq0flwGx8Tpf
Xa0D5lUa3WoA1ZJ07Wyw65YD0DQQtzPy6Kgf7rFQJKdMrKhTbHlFajcKYrec+UmmQYOT3KKanqJX
sdy8GliJxJLoylWkBfbH3FDuoFhz6PrQje4rPvXjgAZaBFx+9xNXmfoCFOh+F5fuJshnsmNKhkpZ
RlwcifON1QES9AS3JiFUX/suq5QcNhJ3GuumFf1fFTDoU5E4Czda6qsAUu67CGdv+nuDJ1PyNUOm
Ta5bc8YwEmP90+mE5g6v6hK+Kqm8jKwcwm9Qwl4OBrh3UGYzzYwhMoD+VbUKE1e7pQTFbpV7wFA4
pHpei06pujvks5B4k/cyaBHDbGvZVIddsQmQ2Zry86nEqWyRSXU707dF4dwC6mA3UsybUekli6oP
fZySX4iXfxsMsNEZxvXdCXagx5DwrCdwjjw1cUaZL0JFzWSABeDdisCLozoP2GkRYtA+ForYTNVj
K+jEbvqYCa+mhwaxOHNz0uvt0GSgbENlxMbEFpJNWmh1fJjd/93yJylNt3hCT8xuFeITl/+VXZPE
wT8KgRexvwJKB+0b11yrU36ugBBCyS8ULyD8NNkwWc/NKvPoN3TYTQAZgxKm865siu+Yn7ieHS89
4Tl9/aNCCtZxqPOn/X22GZ2B7MZwRav20JuJXK9Ls+WZKwstprJW14Xt82W8A+Rwmy598DQ1HC9q
c1EujBrKorGgf3sif7E6+/jA5wQvwVfqwHY8eKNh5fQptH9JzLTCaXUrEqnRC0SiDBBgytt6T0Cl
f2GlCPekb7vav/CQc8OPeOslJNs9kRm9G+WhTSzXLWQlAzjveDdK5BqXoz180K5yJV867Xz56zCj
GP/vdtfLLrkVHIw4JwACdN1aazyJY4HqyB1ZlhapNEPrmkWobIV3pY4jr9ALAMUsMYpuEPCGD/hv
etAUSKAy1diXT0YcfuOD8ReUr7Ll24olViJqihjb2JIle3Ll30ycwEBE4exZLiyO64o36wv3KFeq
RCcmpunYnc/WzNPh2e7yh1ZxITwz7y6feoCZHWvaphiI6eYXveJ6WAy71EuEL7uZKt+vvSX4bf3n
nNcpjJlgopfk8QVuSzYC7qARhQkc+CrLde910R04vainVNur8Tsj1hWJlHw62HABwM5mi/lHsyD9
AEm8NjWnF6qoiwdjY8aXUGWOxf0r9Oyg/48UPChbw8rZCzEc3h0feaa4ljwJeo27zm5+PWstQ/8h
PMGT7C7+Q/u20OudPGQZ23Y5wYpWSNneYwJ9ij8OO9EP9poNlOp6ry4cMSInDo7g8foE2QjVtt8h
WIdrln7JPD4AsU5lPW3OgLvkKCjhKGZx0rN6gcC3kYMSDvArZtibJGrbsOG8NNqtxd/J45Uesx+/
5JkuV0BTYCdlj/AOCGVc1Iz/9KuemOmicQaX+qUDYwkua0m/eUHJqJZSemmoaKNfS6OJanSkq5oZ
h7tpEGOuYQgPRSeRNpwg1U7CJT2I7f0mqMFFb0ZBLLHMyAo7SJBvD9DPJWv8zQHXLGR8RlqNBiRP
9v+vKxsZE97HNyaq7SNjcYULwbgC/s9SLVoiOYWdDVNYa9SpP2f25QYfMPy+FBXdK5ejEg6+1BEK
9SIX5aN+CcL8D5QkN6NAwZthaTF73jf35uT9WYeG/2fNvIlDGTz5tx9tBNky2cPf5Q7V8oqVf3o4
cGvXEkuDM+lL+wQF22HEgR6tBsswmTjdT4V8i0PFkCOQisGZj1u5vlzE1c51yLR1Ji8/kGvEDiHT
/6fNAjiulBalRWgL/oKVSbc83lGf5kfVpfJ2wnuhHSD+USwGggvfgMtmNOC2m9DZDVNlnp+Xzh0o
5efh9AxFPp6Vq8dnXdH0x+Ul8o9s0WeUqmjiU5r6DIV8LZ6AMOOiK9zgqq1i+CtEqA8Q/C1PeyBl
R5zWroL4Euh9eYN5ZTyD57AxGb4CFpVzS1KvvKjLCan814sLy2WUMTdlTBLUCCNmxXpeLNAsZZcH
F9FXaLItcueXCmh086MAhRjIX5dUVF+XAeF4I6PN/l6MQJKaxdw+d2uU5WGIRz47Sh8W7h/7VnPo
vJkWojlrGY5nToNC9oNOLFb36QkONGwmPsv952HtJMSsyznwGVDhHjm7BtJB1V7jSN9ukFPnddQC
thBcNKtTLEAcFGSzLCgdNifGx/aV5LafZYAkrk3DDvqMVMrgL9Lrz0hPjvMl9JZ1Y/qyXHIsif7R
D5WXpDBwc+3ElYufSsuHRsvisycBGeWs2NBxb9ZgxwxEGRiZkeMFtPM9E+bsMw1H0ZdVPJTrMXIM
mAB1su6SLuyZ9CqjmIvo0fokQf9dTMjdzksbdo5qyZ2nQJOGrAJ/RBPh+72wQZhykJUgmfEZNU88
ANPHe+ln+kJWGRaY/0/7uPPEAaA0U2LKwoNrKhy7IMw2XBut1RB5RLyxWJr/Bl6o9G+CWF8kFoTW
WDhoOCFy+BqjsCHkEZOJAi4ilMHcS3e3DkIoquj3moqvvQkSarCVTwyAC406V0isY1H/5k2UtrRt
Klybj7dFP7EgGfR8/xl9jM3KNB6Lhni9sWjRlN88PU+F7WPKvJsTjAuIkTpqH/45G/T/44Nuf05A
JmEKgZxBCB1SY0e4e8tVZpX+Xp+By5yoUYea8GxmAnOvcbjbAdUjlcLYRsm1Rdbp7eVsuJCVP0gN
LCXe2gLWii+9af9G3KaUw4r9ezbbhp7AbImEcaUx/y+u24X7Qumz2aHNgnB3cN5vLqQaBWxucbzM
wgcXQeKgwc4PhRwSgeEwuJFwXWygeFZ5/CJFKkrMZSAjLh/2EL7FIm5pkYssRR3spHnBBgewRSGr
mr4TjI+p34U6KWJCDjc7kfpeclQ6ufKNyh6/Kv0hLdryJwSzUhkqcms0xTgVfR/Z8RpgjY3jLYq+
oazQNzUfEWkAxORZoqCUp44wG+z4RDovfDcZy8A3KnTJNVG1iF5+strRr1n2gMgYEEl/DMj5XiCz
qDYuhSe5duvvua3KagGEz2X09LkcE2RtGG5kH/8R/i+vBZOdbqYRwfYbVkuJuSABF8jwnUO548LS
Rc0qM/1hGKUzFgwq8Zf7+tw/YjqTnvLPLkY92tcIjmmbZzrcMN+7gtdaDBv8zRf/UAOCOgVc27ev
Yic9PsOVjVnSeEZ9T2p7B19cTt12LGRyYS5p7ZYU19Lwq03vfvhhdicPxrAUf7gzeJ/Mk+hyD+a4
f0/YGf4iOEFzszp/lT+k2xofPeFbzyFQ+bNSrs73mVPnCQwobU41Lu+nl0bSfI9TkgRaMbqBLg5j
7dSA6axA9JWjqrvrn1rEG1iqfZEKAugrcEGeaPgBCmSStEKqJlNqTMhBipIXEuHUSwY+9I6aM/Qt
Jss6X72MaGII9IRnAmxHCiOmgbgw67lBEmSl1Fp6RLM9wBe6C64FvH5ts9/t+U+1O6VexTEDhUOA
qqZ+ipaGAvykXQpe3aD8sqSlcurJfx0G9mfj0HlioxMObqJ4qgxFkXOoM6L81ifwGMFyafMZ063M
qwceJI1qCYmtmT+SGz6rElhx3SHT196B+ST5P9F09/FZEr5VQxt0hnpf/qoC5XcChMMd0Hdao5QM
bVifW+lyareuT67LhjUJFT1SEEBIGUv40Nc6wvHsGZY/zr5A1/Iuo2UzBx8HbVp779Hw3g+uYXLP
pZhsS74O2sMI/zRXA+afMq7eguu8HxIdjSsuenVYRo1IUqVuh4AkvPdhGdt12EHu9fkFMYAcyoEe
VNNDQGe9VBsu8qX7d/jzda+xjRtzqh4GNq9PJYhejxyDM3PpMSIWvY9gy6dFvRjwh8rHPi7iZYWs
wfq6a2EJp8FXSkrTZSG8Td35xFroDWA4bXlXyjBdMzzu4at5sCQw73pCNaU6lVWPDePoii0XZdb9
+JyxITHP6Frn8tk9t/nFk48ZORyhNh6sMZYwUHZ7Mp8ZO6pwR8XemjJKqY1M3h2q3opsI6+kRkfy
u02p39jdV1SSEgEI2NspOAimo+ssID4jeU1Xxd6oSyKaCYadbo7NEPmdLfOt8X5mMin3wswRVKuT
XSUw8s74w1zRZmsZUK94PIv/HaFmM/XmoNs+9TLkCwtbVRpDPB8EwAre9XTtcgLtyDbY1sI7b7Fy
r4TOt8IkTFBm4YgUkNdF0msJctU9Aq6ZAj93OT6NKjIkdN4YwnBFxVSVK8nKuewXGwC5raTgMXdE
56nqFBazJ/N7OGKF3HKYHqWhLRR1GKiCcFd92MBfLnH3fQlMp3Axx8XkaD3g6pfxa1smsDiVGcmn
kejCzwQ/yWL4zV1fwKwFZ3lpGJ9WH0IiVH571Bb0taPEnnkZDzxMec02lfHt1g/QJqeJawNR8Vfw
hGkk4bFdcUfH/lgoHWipcfTX3rpyXEemNCEZDRi2YFvYoH7hJsdSgYkSBKxmm/52uTPGS6w6UKqB
2vfO9O1cejsvqonm8vvuQ5UWPCnYRJior4QsnMcD99VmHdlpR0t47BPiAow392r0bvMcJbLWKQRv
7FcUpudxooY6qAK2pXG7oLuJf/QfhEAS+zE68cR014CmZ06U8vvJUnkAaniA2S0gGnYde2aaLJNc
jaoX5v7l+rVYxG4pJg60Zrk+K9yAWxW+WWWOVR4/cccg36Y6AcEy+sG8hi+a7lMh8pKX7oAKpOF0
46zfsDQPmI30IdxC7CBZ58e+wqoAkuotu3edzUqtwv25J5jE6N6A2y0SSjaHVipDw9KJEmP7Sft5
MpBaA/rlw++Aq1xksAZdgSLpnfrFrrzyHi1yoE73sn7ovM0Mzvnpt0yGD2nMS78qNVg2dPHMvKp6
Wh47pYMGdyrmuEl4nG74IAMJN/js3Ml7yWvSlsKzw1qJXVyIr1BjZcfJxIH0zLx8qhRNSA4QCcHn
5UzZu82tryuEQ2vIA+/o5r9imp36qTE7NijUsx5ejlmf4izWj61EmaGmx5/L+FR1l6YSQuWLvRq6
Rr3kuvrmNXYPDg0OAV04LBoay5FaSC4FOZQ9EEMI8/2twFoC7xyNpmiuw/DjMUaSa+I3fmd7LiZl
CrOQiIVZwOUvayQDkIaqKAaIFsm3MyARk0KWW/4+/R/724hyiN40Ni/PYMRIAdbRyqnOtDT2hfch
85wJIQRfMuEl1pJ4l5KGE0ZJVNzOLaTyvoyDa5GxeJYQY/6TmxoY1YTVT+tSXhtoS4yfbat+kCsE
RBZzjwDwVs0EVWnuI/5uA8/cSWEfv0Deja4baxzqOYiNksNQ8dwKc2PPL4wrnO8ve4uNZ3FRl4wA
j3VGKB3W1WQL/4xZQh5ZvPk6PjoOr4ziAidl5xb8fVbMDpPEwuxL+8eAIk73mcJDqMHMT2PdMJIG
Yp21DyVyo8ugsVlBx6n7pKfeXVM2e4IFnQ8ZXcJGJqIYQdNT+tr7GZwp8F3ot44w9bmCF0DgYWS5
7EehxeNWURxSTO8EtzGgLLpcHINPpsPxVbLISnzl8TsZvQxjLBSULLrYMCpKPS21b7aHfxWoQEb8
CA2flW0ltO0t0i1dUIvCIH4H0+BldcgHPiBKu/VQFtbpH2sf29Yvdpxd3y09xOkXW0nmp00kfBO0
FRMrROgTI5b6+zlV3wboXlwyLJkA5GTu501i6EL68KfIlI27Z2S1nTi5/aSkS6F+4B2uIwrx7UYE
7M6vBVeyWIj4rjRhEwTK7Jc0x7NvDRuorZ3KClduU6sVpBqrS+vLiDMXGhPc5E7tzJESdPB/m3zv
9wIntcLOc6h1DIjYcbqaEO7e4p1mxwPDMoDp+Njs87PraMf/Hl06NJ2dHvm1TZhdR9+RuUF5fKQn
9zjV4C17lQz3bZL4VrbH/kDz3Bdb4hA5qqPQ3dh/OtGwKOHIbHGCcAxMVa2+WWzb6e4QvCQ0YsBN
oDmYs1WCi1VutWPbMGYBwRVB8ZiBINz8xMS2MFb5WgD+yQpegSqpezo1+B7o3GiYz4z3///auf/z
H1j/Ylw842g6qBHlUS/Hj5gXtJVyPZ1chHoMKHMP6WMd2PjcPsoqgZcLqYrNHT1ua5EWk2nw+qun
v8h2hJv55Z7GFdrx3RSjUJ4ALCFD3NCpYZ1vzJXchZrLQ5JjQGzIfeXmBArAZeLmLmOOazY7V15d
1PRkQbUgzRknlKLgkxg9E08TWaJ0Ohj1JMyEi7kxBU4ZfR01QS+D2RfvnvToPC74oys6vLWqcm9t
y62QcjtEzJeT1QQx0pvimHcWPePbGL4zA1jiJWfoXLtHwBZ0j+DKXaoM+BUaacYxdVKs6GURh7eD
x1p/kVFW/REaNuXoMKC9X9TL3gqqw5Vw0Clf1C2C7IQZmnzhtArpHyz+XcwmRTla1sdDxc8KHUrq
pDDcGtBK6SKR3eY9U6gwEklZjWsTA17gbB8dQtS+iigqlELhR39u0gtdsuPHjgQ+rchaBIe+bQii
gb8hKw9FEVuqDNq08afLC7fz/BfzcEwSP3h6ZQp9ul1Vn6ujOa83Lro9YyZmG/hobiq3pN32IX7L
M/icNEXSujS8HtPSAuUFVhOJeMcKbIWNADJZzCW7yBrKBTuxTNQ1ZufOprGIgARRqnPj2DxmCIHi
lufPdlDKpSH8Z2tb8UbHvWWqPhleP+bCrLs/pEEz+gjK+y5aBzbctv5QMT+RuxXcVgyKV7KIl32d
2bRcvPiu37lEJSi8KsrgQxcEyisZC/6MWmc9fE+ZSE8ZzmarU6Ix8QhScbWpHplLSjJ0KPqhg/+y
lPGUW5tpafii1UAULkehpSbwMEw/lWCPTVuUSI00bpQJEnuBR6otyeOc4Ds8ajtuq+izNHtBEdRs
jORg44MI/2FIsnSbIWJ0vPn0xOrQCOdzIXqNO4t7ulRwsOKhwHzs6RMhgJKVUxlUAkMhvAtL0uhQ
dp3zRXclFQ4VRORCmjY4vgOFBtVlMuvcWT0bQBPeptwlfpS1uZ9o0ycClPXsw+3rHhkWqVAYn0FQ
7Ak5q8RI2TRyLKwZvVIGDVK1qIpHABnlqXvuPTRxMIkozrPDMViXspvLWnxigLW54YHyVWCpbrpB
L8NKinvyja5L4GjN6YQJQSXhw9Kc2viEAXb8hnBm/XUgR0UUxNxFoiaYQgsdBJWEamwQBB7Z8KJ5
ls4bt2n3Lae/JkGJ/tWpZi3C7kXdGOs1sipJFzWqI1s/jDU6su62axGzIwTtvzoh6T81yHIEKe+g
TVw3WCPXoqh801CSEzooqTFQk4oUzx8/NNmn9VTimBT24sSRLV5/78PLqWI8WHnQg8e2yLHqLwRB
gdjZSz6MZFgGipMzlEGBC+3a3bPS88JH8l/aXoNpgCoiJT20A3UJhXEY5DGGxpaN0AI8eckH2jLg
cipqjRO1Y34Jg3uUIncBzlKh+30IOFt6c10yJL9RsWKJ9IPFUBI7f8EAGrt/s+r6KLtnrV/Cm+AH
Vngl/hgSF8hUIJ4e717QLbWUvDPF0v42R4uvr7WS5XgzcEyc7qQum2GeeAjzZ3Q5x3Fy0bzznOxA
Q4fbT6UyfyZEwytphEZXCEdkyuZelnsqLwncWjnmkI/LkvtZe6SURyXCTITIEjHnPt9G8Bx0ttQR
sCRGvIwO1y6iROipPPBdXQ0csfrLs+W9TfdbVm3oIOB7f7W2jyz4grvWLg97BR/E5WfE7o/2ScrF
t3UFns2AVGqMU59Isp+xVwW9XWTgWFP0EVBboIb43WyJ7W4tvuKPaGdqAA8frBXdv8VzLo63Tv3e
p1FiH6qM20trLBD4FE1EGCa1Vyv5BrLQXSl3o9o5latpxI9FrhIWw11goRgMovHH9CMrECOPp+5i
s6GIehy0FtkMQKlTlIiuAdv8poNv2UERvQe4oPHTjtbH516z5JGrk4+XMNJRJg1TLhK3yMWIz8F/
X5pCeYN0yrH1H+PORcwkJN9KYbJmzFfyB3/ddZLdMDaAuZ7xX5DnY2qRF3l/bBby8mrOcY+iBMAp
CGO0xVQhNlaMLME++qkOLCYh5h6gQlXnWK0jX722H2wvjtTt6r16Hw8ng1wVbcNpvIz75gJBOIY2
ejwVwIDSVUj1uX7Qx1AmgMtmV39LqvSnWGl8NJ+Ln8yy7If5j46nTv3SSdEQo5XSyXZnst4EuHbw
OjWMAAu/txUY2ynVXBosxI7LYFHDKWrciVPfUBlnbZsGIVLcRnGUIDSHepO9gU/vYHerB9ieKJmK
c0w6ZBQZpbmPsR3k1b4JV8WQTaDb1nJtJ4dhxYGskzje5HBcmOoiaeFZdB2UdCYV2hQg2gasYcP1
P7bHIifgBep42oINC70kK3fSH011wAMbIJfIIhBsc+CHzHJGmOSn70zmQdY6VNeawOHKijiHZjIN
M/7NKN81ZmxA+ZyWauP7tJXrwCkftn8P0jahDBZq+ten3KOBGYWFzyLH3xVup8WIlErI10cI7N6I
5Gp86oFgem5557SabclsYlBGBQ7d0IB/GkahtwpZEZIB4DruvJKuJlA5nWYCHzDFz6kfiMl73IHd
JCTCSMdmZZW9jexIpoQGcxC6ohaT/NcWP5R/4hKKQxq99A9hBJqWyaQtetR7WM6IKVx9FzVNXnYR
OgrF812yII8YsVlMP/DX3rEfRyTc3TBj8ZBg/EJwW5nZm4rnDkFm6OtRo86dXNgPoB0SCbEj7x9X
/f+fc+9AcBl86TQW1t/AtqQwEyNcpvwm7YUwdGSL2uLHQx9C4E/vWX7+8dW+v35yvI3/+AbdenR+
M4wNlKnygpPhXBWCO2SFK2mOag5fRIE5tarhYqWTAf9ixB9zymvJm1leDmac9ZdjumU9WFFyEK7l
mqxNcdlsrvjgGfw+awSJmqMMa026ym28K41nvNSIOD8ulSJSC0/Gsp4g5V6Xwtm5YuFeLiIK6Rjm
vxi/9LuUKYGH3xqfMKUd90grtLaGgcMI5RhZ4eJExYJNotRZK3uucr2ADpDhMfP9KFZU8ViwxNjD
WT/VsGEcduF7Cp3E2Z84YHt7V23mxjElqv4DxZqnby7XmGdne/NjzkQD0EAmDt36DD/WZjMfVt11
Eg5ubwuIC9gYSvR17Z67XcVkjqDgfhnJb8/9E9K0TGco3Oj3Q77pp6x9wLcJpxQQkKJm7zJ+pqL4
3V0DMqpXlp4JuxO32gc5iLAPsJ4EbPpmfIorHdts8dD92yiaMD396VB8hN3K0BGuJaAg0UPCaALl
9qvSWQExm1r5ZQ6ZtycuXgCwhhKTkoIiGwv24+N6FcKahm9mskvheQYDxd2VyDR9HiDMukmCUHgA
nIVRetqEvzYpbDjG2fiC+/bLdrnfH0ZBzZBD9t4gvn4qNV9AR59CMi+Iw821PG6jvpohR65yRAAV
Rz42/BZsicseoqWG6RI3z7kGKFskzG+2mr+gY6mB+elqXVMoMcK6VVrWXZ9j2nMV8RzSlP1c+bf9
z6FNxn5g1SWxegattzrLr3jNlMGQwZukBXYQeOQEduk/4y2mza+JXLkxsAch4ZJu9Hh3HIngX7r8
5RWCPOJpe2BA1OhABL6d4xGUBBvnvz9mf7duh+uqPipjlAowQ09koBWVUuN9CiaJnuDTy2biDNyn
DfRzi8Jd5cQtpEXGEB5ztb/q/2Z1EjAiyoKRujr+fs6m4RFfWMSSwxg5TgPJ+zeaZcEhAJitWA+s
yDPDmuH9+jIaIlW9bhh1TE6LXg0ts48RUz2di3PrTey8GaOfgXJRoaua2cmlAV0rHF4LCqFxCJto
hl4+wa7yfvNU+WUGlUu++zL/CKOgeFgstv4mvFmMPQsD6Sb+X7IWp24qbSqmg224IhKQP/ZuOwOT
/a+ouGlKGu+o0QFZEaxP5ZWkbjcm9NxrYtTY0mbF5hDVPgua8VtdJMU3LGVNtWf/hS8W/JQpH1qW
JJzrS2wMqyMx97gZBmWmH6ZHcTxg/Aw6XzrUr3Zu5loQRtfEbzATFAHp6eoPL8abTQ1p4gVE1fZH
i8gJTfWoL/N12HqVcgQTnL5QC4T6f8DhMJPbWWgh4z581Joy6PjcfuC8IpttZ4mZYb62QUPUJidL
7qKSaIIAoyqDVYOgiGf4Z2W4doGChJ4ZaaifpRrOwR0tIsK82oLG/3BgCWTgPXeqha6l+LLzwZbB
xhAx9H4hXjF8M9nQ6j37gp7Farv9VTvUc5H6B8NfVc0wRlMEGzSEwHYuO5fgxkyrJItzS6+mUXiX
1f7C19A7aDyqCNJ8Qppur3ADsXk9LAR3F6DqS8CmGSs/+8/nCf5XgYNaliBDnrNhUaASYTNu4wGZ
fvL8E262eUQvwLDPHF7iBpf3dnI+7vLTIr7TgdGgO0A+YSbmHzsNk+oISvkzSzJkNXubH0F7dkGn
FXJ2kQ171QfdSpqur2LKd1dXskGA/PjzeUqOjW+McIZmcf7uIpYYcoqJWkZ8dCdpvGBfu7uv87Y4
/MzFZL47hO19YJN3S7xAbwFxHXK89LdOJXJTpMZTExfIXWPn64LJ5DUytgrw+efeO717wwlOP7i4
9NJtDwjfPM9uS9naNAccdgLw2kNqGSXOBkHOag6FGwWBXkbvZZ1bcDf4Ps1rrAEzenTmU0g7Q/FS
l4h1BlJ9E08lpblG+nIqtIDDc2L8ibnNNwioGAIP6CahnImDNF4BnUehIaEQ64A1Sk+1yS43Fj95
DmzYO3QOOwmSdTi6ZRBqnzZIQPGeyZzIfXwqQijP780B3Yn0jALubNKMFbWNeVCmrnpG/UdPw1GK
v+qyIxpsFbvINRaG9oLXsq/HzNxo56EiV+S+xl5hjkEcUV9J4iXvpGRusN1efc52idbsB409NDby
1z+6UcQtUtx4oWdKmpmgPSfYi7mImYaevOkolyO4XmhuIyjxtbtN0dM8jSY4l85brGuJn/RKAtrX
915uuXUmzUTzRnBzkWf8w/CROGVBq2t7bkGDjy2GJAyps65cx8u/TmXkA1BSEu87bKAGiXDACYPG
FyyfjMKaOQ58dOTUHzcwmUOn4x94jZDYrrg4RD4/E9Q9Z9G11T9c2vM25A48UKHkb9TvF2Wq8h8x
ja9A6+jpOeAmxXqRu28U67Yj9Ea9dsXvnqtbgy2IgM/mVxtj1fHrbh7JpJ/UNWRygy2qa1uH5CT3
trBLGTvN8MOIQxqX6YerHFR2INr17YewdDYW0YPAmy6y5+XFA2NuJRwyLAmvMHDcBF7PXDmqicXt
6dMFraZ2HgypXUXOktZgQ3D1o5x0jq3bkrVeg2szM2htIz/ysC5kCyvGjs4oLFpVXTAArGS5Okv4
toJRZj5JkPcCpKhYAS3OLjvy1k0r+Hb/P9J3vveB65llZ4N8lDBoWmKg5AO7ZPQ5g5INx+GZX8Rc
ZMHq2+UmixvMQ0AHhCPQvfmyI4x1fi2ic0/H2dCqtAgaM3H70OGfm1mKKl39ajgnZVI1/OJ5jueA
q2w/9pXyrCGq6N0qpwRDGk89+B9Tf2dG6/kqzWCCy3Xa9DtisqP8yPhCPdEXRIgXcs2UxnZQPze+
Cl5YZUwdxR/t6FUgkoKmD9OOysoUc9SMsWW4tIDAX6BQ15NyGyYfNYykccj2jSeeAEcuwGvGRMqP
XD2oQ/sXh6efx1mNkw+/HRFAO0fnSJ0vEBf0AocxEWM6VFd6MF06o/GM3BruiOr0cW8dDVN3PFja
xhiaEKYGXCs/bGLtDcd284HFpgyZ99l6+7ZlRybknXhZ6ylOBWvCZvZXEfh9Fl7xChNGBVIGVBqF
1XfZgpXAM83vR63M2ARTD8fOUpnqRT1zqmvPTSlr4kNNL1rgJbgkvGyjtIqG0KsAoqdavHvJc8Rf
raWM1qauCw/zNAZHQhr8zGVm2w+GHLNuvKUCAWx2EBeRGE+FeSXwntDR9m1dNhFJ0FG7YiHxk0AJ
jR2GV/RfTfb9nO5tRgdybUb50oKvFZEaNTUAHcgqDLd7WsZPj1F0dPCpdmRxeK4lFYstANqC7R8k
5xZ0YO9vWALqQwe8YGqquXaxHaNux8N605ZU+NqEF9gKMygiT5nfF0LYzGWW/CGHKTjD1TvMC+0e
jiJc28JYVJImvN6dih8sEd0/VaGw48meOZWlIwvd0Wxp+SFi0wRGsbsWBDFoR9Tl+RHWfp1iaPW+
+pEJVzWA1COVEM6Lsws54onDUJ1l007ZWnUmnVuXylw82ZtHeqfzQcp1eZrG3cLs1GjhNiFnJifS
sONVH+9Z/YAk/RXVgRXHyUB8vsU+TMsa+ZlooJGY5+sQt7+ugrDXxkgCOdidthX4YCELWGY3ruT+
u39s4xREvXzTno1nfJj5MxAZfP/Ze5O3lxQQifddZBTzgApfinm2ijD+Cdy+cl5wiR076lMduqhU
ZKRQGNDfzUkBCYR8yVBTd1SDvpAuZdVef1UDVatG9syThIMAY8ppaBK9u2whkK+3863xTWJDXOS/
k9H7B22UMHZjyWn8xxC3up9Ca0AkeOetiq0HwFi+rexTffqDcHJfPiMZemo86UsAnHH3I1owaULW
sJPRjn6+2RxovSUxgBPUddtCC7iRDgRP+e6O9P2QRZi3liZkvU/d88c/k5kSg2e7B8CBxsqW/UcW
GNtBa3eRKqn2v8244/R7R3a4IV5K7Oe0VUNg0dhjPrr7ujJ5zF1MQKHcehrN9YP7orMbI8s/jBTo
RxuD/ePIJKObZTll9RLVM6Jo+xyXZWMXG+4lZ6/3XE6yO3CRpOtbi8XgcjTGQY0mvZelODya8S3J
5qxDuUjQOtzX3i5Xw9ljuZgbfhG8BBFtAsk/6ZHD5G2nwgZ54vWCoTziMmLOJ+UgbbOdjb2tAFJl
YnrWqQBBqRS/phmMK0nEwa1502HyzgWJOHT/3bEp73R20m4RpevtWPpfdF+V9dm5bHdyEcDW6itl
TPqR3RAuoGWh545wrD9XvPEc+9H7k2/aUFzXjVuJDnzbkRXBcKm551akPMeGGUSmSEDZQKHiXndQ
HINgfC5e7jRQrZcJ75Wp3aRg1Uf9ao2fPjGePYDdWqy9+KuTfVRGg92pZYDIDJME4FIv65gNvIrq
4W6pnpzMQhAnbCwsCc0+flFD4LKJSG8RQ3MxpklA4FeJwVEWGfrHAtyIH1XXNdoyg14PKu4kMII0
eGW00u85Ijwg8aooajjcNt3QFQR/BF297fKz6qEvC1e+erSxuPhngDF7GKo5SUCyI4v+QHVftVmI
UwWM36Ytbpto17nhT+hcfSKLPr8jTv7VTPtMR/u5cDgnSSotHny+opi1fF4vTZXfyR6ouNSleDVi
lPQ6LXYPpnHABDc93ZLqFofozZiL3my5Pqhi5tOTPlR/AYQEXAIJrBQC7nSAsjaowmHGOA8Ue7tG
RW71PdH5W4BB8ETPXKn6PPW5InVPo2pYBrDBh2kTYRF/A02NR3Y5H6u95QxaXr3FXYJi1KnaIh5/
IPyE184Eer2BXVvExUzgw9ho9cD4ST3qzjw4KWRt0PfI8ww/oSO3cXZ8hg7MRHI52A+Aci+IQ2yp
5ezUIMZquLckAKXR/qnf3vV91Xo5O49M1raF6WMI9r5CLfuwbO6cJMfqkyAfuj4+4PCuvD2CWI1V
gKGw/wTGyxuP+Y2SKt3j5x4+MmuOGZpl/Za/kHEgmH717lQHVADPbjb+vIjJ46/uw/27OlXYm579
9tMOSIHRhpw0iJKrk72d2F0NQJHkaq53yy6Y8Q/2A8UHonwbOiVYY4ibn2txyVsrapwTyM8+5iCQ
ppqgvTvsKefSAZ6vCJNMDkx9Ae/oaiYgx79ajTKvCHvTE7Frc/OmQ055VMlPzn4QVSbEPJTfuJcT
DqW8Msh5cpW2LJkzUx33lPqjsohxK2SYEtF7cMnW6f21Myad7ocD9SgvgYWxML2BQ0YG74PdpnZ8
SCuBgb4DVFR1t9lm3b8JUaWVTA0N48iad0dRs4TI6pBNO/RgElfm51CyvozAIO52YU9LNkJ0Cdxy
Wwi5II7t6oHB4IwUgiwFugr8i0NLuWPuCIm7d6/N34RR0A4Y2TwoE2wCw6FyNzrDXb3Js95eBqGW
ZGWiuAhPo6QUGs7w90R3hJ2ajzlEFgIi08RHg6mnz/BNCukeifWi15ZnQ/67EWA1gcp6OQi3fJlA
wQ36p12nUchZGpHddPPZN4dKKcdTDb3nHptD7UrZi/6ksA2JG17ebQ7b56hW+m/AOskQffaUQybL
Ggd2yHqLj2rrHdnq8H9dF6Iuw3UwgY2qIgDRHB28plX611J+rBqacee+JZCD/p4fzCW1/WcWdC/7
vdVFd6MsJRg4mMHcRbOs4iSCbActxT3Xwtgyfb4oZeLDvrdjgck4gzrl/os9+2Fu8suKDEohi/JR
jAvWAOhrs7KNDuQbdoS4UVuUBFLdOgmw1WoN1Rfj/lUTwghoWpTbJyUWV+FDTgjOx0DvWIRRTC5S
Mqu2IYvxRxf1AqNDu9q0ssB7U3KoLPkgFovRM1Cxi7hUHEVTo3tOdgxek3gWtL8YGfNdLDraCdIt
7S9D/wS1ZG2UUlFP+QLlmA/F6O6wN6ZAA0c4Lbsv7OyhrH86FIHbhB28a6uafD2ReVsRHBMzg3VP
uWAFUEGccjpPVcsApybSiU4ygTb8AfBW5wI/5m3y1A+Sfo0TscBs1lC2HmD9M4+O0z6kOcYrstir
6D1vbAhK0waimiz03ziwLxeBkNH28jwqG7ToiCCjJ8+a6KpU40CL3Y5UiXhe7T+g+juFWnDmwZkQ
5avIg4tKBu9gF20du/A25D3tZtFJBOq+JwVRlRtZO1TSpQWmD4LNXW4TWJ1w1Xr4TLSzThvHXb3G
7BINiPSAz9WXCiCKEuDyXbIgleLYaGmhCBP09rMEkfE87aog2p9riLiO3fyaIywMK/T/j9Dt8UWC
vD63ncaRhAKltNKi9HrpNMJ49R1kvXJFo5ts7lD9ok73oKiVmLfxNBXG1xEvGFFXpNi2w8++aw/h
zHdM72ffvzGA3dDhEeOXXwkrY+EDYFskQzx/XTXnjB3vEL0X76iFAdnDA3/7GxiAXw1jTPTauAe3
/R6mnSPf5yzGQE80bJdbS2UFsWosIb3XlVs/fvSUYYqGNb31K8VlRkZ8ZjLSO2GXE/IqNq88iNCu
Vvx4Xm+ApLSH0OPGaTtWrq45XWwfn0PtPLoHjdBv/FCrclLOi0/IZvtXsJKQReRdUrIE/m6q2X3r
40sY2z0I3DvbbdIKDP1ha6hCAeHeAMZLOVkQ4AHCAey/8Les+a1la8QMYKHcyq2KXyeaHuCL3Saa
J0IMFT8zJQiLgsSPGAzyd4Vf2R5rCqm440RZIdrFO+1ySyUvmsBgVeg5becDD9tvuKQ/3Vjp+tqX
j1GiTtXPC/AAfay2mVcAokZ84NYExRA1VCMyQZ8UT5WXQ4sfAuU/9uyy4rEXtqI7mvxN/VBz8Fo6
aA2aYI8HhtPqf8UgH7y/8nE1asAJz3JQA3eRqW0mnULpfm/Eep78jUiuryceqFi5dIURGwSlZmj+
5PrAoH6aTjkkEy8SRV5go8UnnQnMwTU58YiDnTkbhpDks/BR6eWx4B7F4Vf/D4pg79m1frt7yiTo
vzv5a/8cAZMNvPwnwfx+J02skunFNw2lxgbGTwE7Z8QNFXeoO/5VmCwgHRfms3XerIbmIsDuV5UN
cVL0c8/eKVRY6OWcgpktYyOSXluqL+TtXN3mAWk6slmpABx51E0Sef3Af0bOZ0qGD+fpiWHDrfAK
mg2OpSJYJlmWPFZLxGUvrPn/xtwRARv5dfoBgCBgkdAJp4PT821qBA/QgmZLNNjldD4u1NdFNKCt
yNdiIok29AGAasQtdzKQAq7W0B7gLiWsdQHVc2nqVpP8hBwmz7O/y9BPlUtW0e+UM508sqJv1g5Q
FX93/+fKHZAGgM/Y2h8RQDwUzYriSR3TkE6fltSFWCJUJfJ3EAiLLoNaVrV1sg/sgALRlSjsgKeB
p1kOfjCCzZwvYyBhixGuEp7JSUuRRPah/zkbdlB86+cpfyECAL1ScIWQ4CPboyjRy/pxL8BdkZAP
WDjpLSal+u4Nr4KPSwhVSJaj5F7Moq5ixKiKibosIup82TmTc+AvpdXAlJvaR35gbNN3/QM0rTeZ
bEYGkP7Jajfzq7Zifa9RhbmVNfn/8UdU7DNeG+xeCFMIrw924vl8qHI75+7Lrq81YIyHDnCLq7Ee
y86x63trdQNnbbDL1S+boMGcQKlWtxPEDKc4hWKBazEtYosBIKICpOObm/3hdFV+q+AkNoGsiWKk
WIq0Dw/Bva2Xmuyg+58bUSAmJtniC/WyjYmTGKASR7H1mQQje2qfc9VNiHpUnD5H97YvZvK0ffeQ
t0DT3yl7+O9mZOLJopT4Hfh+anDVi61b2ipw/48/AXqHybHIKAk9aqsyAh5w3oxczKNiO4mN+i4j
pAbCUXfKLcDOMpheXmGR4GdDIvKKqscw8pZnFU/J7jpIgPyyvE4ponEqGsGK8ZRd6vozv2lZf3Xf
/ZUuWq12BAAjFJVGllwkxJVLA50paiJGx2e6u/Aoey1gmB/g2T+sB/pOHfnFFcfg3grT297nbnGK
Hk6yVq4xclltHPWz1MpXs50T1mT4kBt0AIp5ckpJM4GQYbph/NDnXYC9A2fjtwKIk2MoWpQCLrfQ
5gBToMDC8fT/7BvxqptN1vLgj0RIJxqdhkaCvlqIpdGfGT1D2rJkRVDgqQzpI9a8w8ea6HL9z7jz
cfj6eu+PSK7GDPRtJ/mmSaLXjwg1HszxXvfq4yP+AuuexunUFkXmU/EnK6gdebE2pecRSsCo2f3r
1ODAqA1j/L5RhKW02ydzjuW5tEC57WGN+uv/C6Fva5ovayGZjEH/Lme35gdvP+PwkQymyb9ymkZv
pMquzP0MmqUBCaSI4BCQU0ji6txk7RBUb6p3pX40T5lgYTmPxFEy59ZNV/AATKt4O9EZYfzEptkZ
L8v4xlhOx8Xw7q5TXdTZBHWZ041xCCtjxC2eNjyNw4Z92ha/jO6tgHDqytS5uU80qScU5mvNRfqq
8vurdp6zdVjbVwyJafoMfHzZHFBqC+qIGM6WZ96WvDX3akMJi7/8SNj48dBbh+PHrd+Qr2xPWoOA
qHlxVEdDCAKtoTVMMFtrDffLMTn4m5zlkJT7K11y/S4L6LpHWm+C2vP6hy5tqHuTIre2Ggx7e7mX
LmVDoR+Bo3FSJ2uscgZyI5HM6kVLuiCgojCjDor9vPVWTLCqyt0/ynwf02zAzriL9OHVb03uXYvi
rY2/C6j7ZB9080Fs8ORQcvSjoLo3m3/wT0WF7bZHZAyLgbEzMBTECBIQAWbxvFfvbyRm1PpjWgJu
E0IhLCBoDvxwHIT56hKxKnoNJ7wdDRuovbdEg6/Xhh6HBCniAk/+YBjHHo5abb01ORbTWQ/V9jHP
BABmAez026pCGoQc11j1x8GiSvLXeSO5K86vD12StEYIhHi0N9FeHUE1v4xNLVJryuoYuf7Pye7n
DgqxcvGXZEEFGHGFuTjwmvXpwweqt+mCTJD2avFi4Mo/57o4hRVQCm9CQgo4egUAu5+uYl3NEMdZ
6j/FXUhbRd/wFGr3PynLs497+hwQvC39Dm2fO05RzbdMHX3efNGvM7xq+akKB2inHSJSUgfR1nb3
WjL9M6nIK4UjtlDgtxBkMt3yq2xbwWyMMw/NcTdsQAiG9uSuKOfX56LnCgRB+gQmHEivO/QSqOtT
U6PAvAfrKw7MJ4uOP+o6c59sTqTlfxkSHhbGeocQaxXVIvGcpjFRjFbe77MOg+QJMd+fjuVEhE4h
1UOdrFegvQ4lVk/qoUpwtDUDvtrgefOPSwfWkU8vKmVQmkdQ8MqNQBffTHT9abGyBD771HKVwFHH
WaKZUel+dTIJ+Cgej2FZXZ7Pj6HM8AzL7nLJldv44YpFvqWI4uXuXZWtPwDAHwVJoW+1++a1Bgzb
f58GXeboaI9zKgGGAkj8RTT7hDfKeeRVapyg7/6cIXMGMnvn4HP7CTFUEBpKUSAFfblGLVQw/ZT4
yWNb1Z7siXq6cZtF8XKNwwXOI7uHFhAZcfPGqtRlicA2yDBSFrp4NtrE8I3pzX+kkCdEX/ryoZwt
eaIBWVsXloFJW160Kcp/PJMlFVUnsGkdE4TGDHT/k6E87T8YyBTbNQxvBNVIDd4qsXUfuRciaT76
4vaqCAgarm2BCVSC+w+/VSRWPH4HttWRijEVuHsiUI3xfHjJdA/CeUINyrPltd1xLOGtMg55uQBL
FkTViozFrOUg7/5+bU/LTtodceyTqUV1vbI84WTgjwq/d3rGpekG6i1Lp6jMppNNssjubBf1tItz
gN+L5cxkIWsebwHfKXMfVAdMx+wyNtFHev9nUwGaa0LZsd6kLtT+LBadC3Q4zgejVpqq8dlRkJC1
xU1U8Pb6UzdLO28vrVA/Y8h2M0uNjoaodYo11HNNkyjAdl+vx141wtlTvHJok4L7A9aELhZHmrSb
BII2gOu9l89JhhMzUtJWsL34F53Tv5GP5B4k/x06sr7obs+zMGslG/569FBOgL4Y+pHxNhOgSVeP
8HDFEAhupXGDoRwl0VZktDqEJnCb2TTGPlIYt7lbla3Ba93Nmx7NVaYFMQYCN9Zqjlp2K5TNkiSt
q8SypOhQ+QjvT/gVv+ljJjXTUNLYzgkvcnOsnlZudAGt3FUCR54Kz7KmkV9oIvtpElyQ5sdTpzZD
YPh6JWvhRwuHsIIWJtJa6IN1/QVOnRRLZqj4gM+gZpXiJkidMbF8qKSkUV3Dlxmbdau1ooGj1ZEt
KHGDyRwyP+CuwB9fFaiop3FxDr42kJl3FScmj1MtSFE2rGB+RAQKsCb6vYUdG+JT2bKN062aGO00
PdbxShB6RCVmbG7DPmLSQ6R3SMa8A7me4Au+QH7dyl3QlM8Mu7iNBuBNLbARpmB75sHhEfwEDDoX
I4uTLL5hJngfkxmTWJk9w22k/emaL784ULoZdM3JHgROVpYr93c8YomLWE0UJCmH4Xm8TljnPpa6
iaGKbtPteJp3xOGnJyjDQ+C1FvbikuKQtxO2FdFIb1KEYw9EChyE9njTig+VJjJ5Pcc6FsEPNNUM
XdnYnYFqJ3n3c/s0bCtL5PLOae+RFR7JDNhDoAGtBkeOom40pPu3DZXprT4oReSI6rykWadMPW03
mKHT2d8YeKjjQMnUDPcdah1qd51KL9bg+d0T+/b6IaXfZuEXEhSLI+nATuss6e/qbevgnlVHIB1H
Xc8xjdbUtYXfkkAgLVgJVfNOU6YFWxFZA4J7a4JyehNf9tAv3JIEEphdIhhqNVYnr/lh2tf992GG
PFHp4GhQOOs4Rs4rcVF1PCENoq5Z4Qs4y9Zz2QRvBJ0++WfcFPC7p/mOTRPYWd9Ib4eR5mE4xpfs
9uGF1Fe9B+CcYBinebF0RFFrLwWDcyrqkqDxJeWLc7YSPosdXgiLgAU+Ol/52+3bi60URv1sw3qY
6+BKwC2nUX8TSuz4cwvWmhsHxniTHxF91Kpojj1rJniRcfgc3ZjogDx+uUknXKxxgeuRxzFo5jcz
6tXo9PDagIYq4B0ViGED9/XRC1MHLyVI5qtYgbBSIuvIYcFGZUmOC6g2Ny2uK8Lyqr5ncoI9LbZS
v4+sizFI+tUrVEfFjIfemZH0FIWrNs3en5kLNLVF2ZdrWfN7+/oWqz+upgyDGO6dO9RauCG2S5rV
RgDVzXRHC7YfSYKk5nQDW7CzqeJih3wqJSA1i6x5c1MNbx1oBl4l6kwF42DQ1q6SSeb4Rg/sOeA7
Wt8n4p8m1rthLH7ik/sqQdybQGDf7wfwuen2uePnob+EEwozie5LmegF/lJGPO2E6IN50f/KjOfe
sWWEuazxbXVfGMz5hBKK+H6f1sO2z0Pb3bOvBpXVpI8QoNSeckqj4LoPH3lX5xf8z1QFK4rx4W2s
g/wgIzLJ6+WcdKowvuJhPa8UUyqVVnvrDNHvBkACi2rXIomfDfJNfZkM7Ng65wyYwRzuwyNfAS4Z
ovKI+XUYYSWjTokOostmKqbwld/eac3trA8YeyJdQdefcHdCvOQ2Asu7vj1CPzbQOWY631lu4hev
2VHdjqLOKW6HrguEqjSUW6oyFQ1w8d9gQOL3SOD9sibxiuHJjwITSVbBURd4CGQoZ1EWpRB0hOse
4z2FTmwMWWRlbvYktRFivddUfVZtK+ZtmzSritYOZOo29+fuOptZ8bryTM0Xm0nGwSXRsUrEgESD
ewU/tzyebQenYuIMQJ8hU9CDsifOFoXP0DUjKcyRfRCVldpPCYmm+e3TdQaSQzwk5vk3lr6nzuyo
R0JQrWgCkrLIsxiqOg1D/m0Kg+OAIJgd0gsYVviIPuZbU7ci7yLYlNcvxH7BsawRnl3NAXZyFd+P
gD6CMKfczLraKtPcJ416jwDjamupMrtsMIY0O3SD/ai7bnC3is+u4WC0hSx7WW4iIeNyd/hq5pYj
2QTk1hXpmmJGtV3jFM9gD2wDCXsBF2uh5Tgb5iXfOadupHG+mSkCa6rDsSCck0KlM5BbcGMAI8a4
nXa/S3LwYkRG+scA6dzr4S+As+rFVln2lEOlo3XnoXiBVt62s6mETvvfWX3+tZDcUSxyFlCNSahV
z+rwIN50FX+iwdaqjq1N+I8GACKnB68bClbJgHKczqycD0UGWTVF4/0fAfOCX6HYaNmcAlYBhY9u
iPBkgVbLtJHPZ/lnN+uT+NbhyAFDRCkqQc/vF4+zXzYM7zdDq1aJz8BuTCxXAikhKl5D6bOeKkQt
mnkxwjoZyGGgBlEdFxiggM0fi7bw5TKIV/33sKfxQcmxrx9JveB4SqX0VltKGz1Ptq00VARedkRa
9NkkT4+jBYWv7VgwZ5oq8whjLrMVabjev2AG/CsSVuszEdp/BKe504JoCTCDmtm1qsfNd5DHybkg
MUKgjnbww0kcSLeiRPnW58+CmLcskA9CUR2UAoDWkWl52Mg33a/Cn/v2ZFMtUKrzmFz4SHl4OG7d
ZZi0651X4nYhMhaX+EA3CKmCx54d8KLeLKrBo4zOr98pB+Xy8dXz9QnPvMw/rO9S2s29Maxvkd4I
V1QNv95c/cE2Q/+EWQPJuGOT1s1ss/oAE90pBXpI82hQccC4HEW2mDi5wUp1LVNm77Dr8q6BFMRb
dvFAELIqpmojNIIEiDo5AxNqrNWO6y4l7EXmotrgK4Bh1/F7GSkW3XQPv3JEDk6CjCIiACNFT3uv
Raf9NwTqJu/qCiCgBtZO8YLYYOVNbrlKs5hhQJfg0ujkFF0DACtMp3NLCSyOcTtwbYM0CzDO0muI
MkdrUqVUUAzXtmsNoyrFEXGKSwANQKTOP4mkPV5L2PN21miQ//X7rX+qzizq/Y/11sug+kAv2K2V
ZCzrA4UXFpJoV1me0iDZWbgW8dRsgjd+gBxsyC+Vbl4oiw46XGV7dXgjke59k1+v1q9dIbNHHYGC
Dy4rFARbGQcc6vFYl0596sVLPBkuVCLwKyZsAf82+WwPM943ABf3pmOTSQf9q3NnYxjwJfMwKblG
2NWqdKsozo82hChd1bAOFwpBBI00YMZrp0a4WQmERm4SfBICSEt/JamMjl05xLRq+FuTTA77g8Pf
gkChYmqjn5S4xYr9B514iBfbWiuH/LC+NVsaTjaMpvAzpw92wirVxKGAedCFNzqw7a1uLBnWC1XV
3nqtIStHb2h8XG1TmXNGXJ0Zbgnjw3JDDvenvdlXV6JY1a0YuUdk6sq5/wKyzZMEp39Yl5uwEiZn
3k3SxI3FfZiEGfmu7x0k6i4pOG5ALPcUxBse6t+VU2Q91uEkoGJe3KA0CfbrXcMF5JxeKJQLTQGe
bX61JiuSzWesThITsaUvDzlK+rO1V99M2ZCgEkfG5gxoCpnqX356yu40iOHGmqTMz16kyGH/w2z4
FC4rFDvuzRS/CnY1eDQAJJqxAmcZDnw8HUEQV5g2K8xOk352FhdTuA/dPdrfZV/tUmd/sWVYuVoN
1KbT3zV8YuMrWbdR79gSu02u6dEsZpzPZAwIGz40veH6y8cdRlmjDfPaz3P63NKftLvMoaO+wft/
Of501D8/1KzaqVvPBw6zLfgVDyN34Ma82vHgpKPlCJNOgjyeA41qy3b0AeOKq1TSOIGDx2EnMPC/
tIKDz9cl6ck2h08UAtWwL3on+/blRW5Q0TlaIz2KAwymOfWAOmfyp+GxH50dCiJIDlBYBUACB/TO
72pdSjXVctf1I4qBpdVxnlIVtZyYf6Vpmbqd40CvJWR1on+tKO5KztX6fhL5EOg8597CMxx24Frj
+X9U/Uw2UUlv78StYyfhhrxQcjeCHGbz+sZxvht0csugHbMH9ToCMQOFVpGsImHxaTwpa2VPpsWU
egagb74H4iqlSv8j8ZFV7zG9LhrtAJounLd/3qQYX2VODYpd7GdrR2ideJjYlyJ07v6bNJZXXMbb
ui5WiR/ltGvq853vngrn4tUp1l5dgow0k0XlKjl8jKUbKAmxv/6vEea4xYjEzKHO58jem4D8MHbU
Pqd+6SY4jogRPf2lryr01H1VBkcBsKG5xcdT9QjjYdTNa3cLVJ28Hwt2G0cIn0pdlYU2SDBv/+Vn
u+MGU+378Xympn7lhXMOsMWEzyuE22TluzBVh8UTjK8aTbMr86em/LSpjPc8phu3SAY08rgxhpPX
PPor5uWAqwOCGmOGJYs6nik7PWe7YXSA8l9HxSjXWf0wtPCchNhioQDfKnqjfkMAfrZCKl+f00tH
oMA1e2cmWHxUcwCy/ga6dItjPGNJ8TEawiNmlhfy3B5XovpEAQMiha/QFrVqWe+oh9w0RM7L0BQK
Y5CwGBifOip9A885/h5t2PL+ZrFyYKsXdqVM7GMmAJpjzLJfjhyvDVJLx5rDhRl1Gr5OdWn+B/g/
2yFIttRKQ8f9ZxW6XFUqL32dthkF7YsAuGXJ2TFT4a39X0qhHTYMsSdLZU+VfogphZGyzBnPt7hq
4oD5K3yi0bp1HPAknk01xevQh7Z+qjJYMYsghyVnY5AaJ1M96YieUy3FvhbVyL1LloYJIOpz/MzP
tUw0iPyfdkQB6HCguKRPZh9DGXxK7DgEBFImdNLwWm+Ql++lO4lEmmJUeP1VmMGfWepdHkVAhqX9
50y4YP4ELHTZnIVZiBB4Xvs5pi28RiqbdJZ1FX9nHPfRlRlbiwV2hsxnGq6a9o7SIpimjM7Rnhxi
UwRUIIMWHxI2T1M7Mc8bKAbeuxNxLeSVdQa0B+0UsjjCTnR9HNvCdxZSM8E88Jq29hWwavnPpStm
N7r39ldNCPRgSckfqwJKFh1BGhQ6kWIZWazGUIoiw+flhyfYXRWK7F7nbD3DCC/Hw0RMLeYd7yxG
GGPAmsukJ2PqeOIr+qadL9SoF1G+tbKTEdk/s2+aynaFttQUmikqWUVewS9HlcV1Ltw4Y7484gHj
+XgVDMXQ1nv2Buc5tHGRzs0/rB4PYmEu92OLOmOk6+8ljPIQ0FXXGmSybXqyiLLFdz69b3tnTGna
fUy/Atp6/uy5O9fN+z3fi3zY3zlXK66ModxzMCkOW+Nuz9rhfVElqEep/heU4NzpWwcCxgVm/Hlb
zm1alVUUTKB1JuL6eySH38rcw82ttnL0Z775btN8laPG5CAQRTONeO3Tv00bBucNEMVon27teBa9
LSw7frvJW1Qpf8/U+fthWhROssrVRf0VI9MI0DhG6N7xe93LF2eLaeBzEgMVyNRM5G2u4nZuM3Qf
nK6JmewYeaPso884L6pXndmEipirIXsvUKAV9xoloTTFNaRFU1Bv6jH78FhQWyO5QtrzBTEkP/Rj
r8hy9Xax1W0MztWzS15SVCkF2xgi6mKrV8GjvT1/njvxhgdYTait7v3E54vI7uWEe7kWNbtDzJAx
OL78K0xaXwDwrlURIAJJbzkDXOGW6OJzdDmobLm3t2QBoEkwxppTTUe0d7CR7VbN8egWcMBTmDd4
CwGG87QZ8bH0FBWjJf25y7ZmVm4F2zMogbxTQvrQpWs4zGjg78o0xSFxpphsNoXTHP906ASHx4vm
tmY5dcsQ5YUze6Ude+CEjE3tMqSJvdV/ZONwH49ddmTEwRzqbUi6nI1cbwIUv73E2ARQAD4XQIuX
t6uj8AzjwuMq8QpJYlK9PGRQRfOYqIyEqCm5Yz1/mHGJ/f3sCnUkU/DvyPNIg5XmaK8tb88v9X+y
YLQEV/oaUA5kJieh96+RyWAcjgzKviQAszD++YnUHWoO/+jFE804xe2Rdx2vX0Yq6u61DjtFFDkU
DPlravf5pEQYQAmFdsWSbpbFaQR9CaI2ziWLss7xZRgeeJITP4pK0VUf7XTy5Ef/XfnP0/5aLK0w
ms1DkGmrJ/A8teiADmTFJC+RQMczsWJhtTYJbPsa70efH0OAOtZQ6tQFgM5qBXbPndqQVtCY9djH
NLB4YRF5zR3WSZyPMxTVaFzbySMsnenodbVKv2ExBS3/Wyolw0NroRtiGo+xSzrTg/3cUHXg5zeK
ODzTB32DQLT0eUn3alFI89pAEOwSZGsvy2ZS3I7x8SP7VzZMK5SIHaHbRso3JIi+sX2Wa6DhOuOM
/NIS474/7qxzvQaZhkG7qIvRFdP+Bf1l22lW3asPMv6W4uXr6cg//KyFhQuDTY4rPz1re64vH84r
bjtGmoVvckTht2P0Cwf335Csm2M/LsUQ35qtl9u1HkobF0jpS7wk0SXgnipxDVbhNfxM9OvwC7+B
14bSUti7ky8yN1Bv2k7bU5oV4gtp52yiF+iHu9ujIwD4fEvUhEX3uTkL82ju6lTMJZzDp0vqfWFA
SaSG7JHnLEFlsuk9RzDcsFlJIUfBxwgSv1AuUFOzAm064x4eSF7PWUK+sKdyFnxUEypaTuI3tAP4
Dmrcl3Oy+yy6QzDKyCCJ5hDoTt/Gl5PwiFcDs4XjEnNZnbHf+ofaQa+0L2H+shctA2EBbwVU5Jfh
iFqPQZu+rOaorb/KYwKecWR+IxeGEdwcFxYx/qLHzurCf5G92DSpyC/u+0kA8oHJDHQGpCBaE/mC
2XtABzZFOH5IX5l26pVbqDj/2DfVtgEWNE+WE4GpOCf4L8sq06lCOtA1X6plPTlM4wJCmjHqi1xo
Y352kQRK89vY2Trg4RDiY6ZySm0Ttd8D0jRy/XQVRGLgVHvmyIiXqV11d5Mq+nrwRWw4fbdKHyNZ
ON1nH2Z9Jpv8WRaxpGA3eSvxoKy4Yk90eS6I7bV2pUF/fNyQynO0zIUDt7IcU8RUsU1lbBiwZbX3
LBEVS9nA9CU+TTUENKVD6k+vS0FyYPnjhczW7/U1eRIHgj4gLYzs5eXEYzFDv9imnJSvE5Ly4GXz
3CYsnsuRidiXqxIOuivijM5WqaNSBxSH1Hznlow0YAsL3W3iBXeet5ih+eI/M1plSH3dnGFEYTV/
QuIoqmdxTpzpBJpQD7ZBJo5Su56ixGaS2HQU8SlbVFe6b2ps/8EO5IUcRFNY/2y4XZ88hP/29phG
xAVUWxNBwei3n/ZlCo3V/YMwNKTRNGJ6O+jj6+P9u8I7z3TmEscw3UDP+6AQ3TvzLa1/kKwdMq+F
mH8352rdhzHkYRUTkBGSEmNUNpxh+skN1Udm4tcjX8aOnmoeMAIKYqJAdsJlNOxaESf6cXJpQNG0
G/CcX3W3FqQjXaTkb09d/IZNtdHVCgXZYWOs5/tmmlydyjlwYmgq+SDnyDksDG/QyfVuO3FUK2xF
16VJYDpmf8A+ItX+ErVcEt4Bn7urA71C+caceygllWP87oWuaakllRWLpVBiU7ayHQVuCNj8I4HE
iWUAnoxUTlb9Bi0ZSHzcbsCQyP4Gp0xrkJd7X6+oiaXZIVIP+ItHQ+6/TROJCZBJjZa428n+uNCD
TdRlqCagbeoFn1BYwM67aCy9LlXGo6kXsobaJ1N24156u6FTmTVE7MGPWdwnkfNf+yzGF0UtUzZ/
yoU/0WbIxho9xt0PGhcpuXRMCxIov60NKJcAvFBk1vSiuP42LspEB2Cp/6Vdax81ZiLS/5LMY74E
UK+SXrV9L0F57+I7N8qTqVkG7hHm928y02EcXKDD6vsCg9ya3z6eRUBOtUn2VnBwmILNx1D5w/Un
apANDJr5rGkydxIwsZzUuWM2yNeU5kyuvtfHD1puFUEeNrPLfiX711gIciDxCgpJBXxl4eeVH53a
mgBtaNqCE/KAfJdNHqZCezf2GTilNB4meC3G1xMybUQwo7Al+M/UuFSs6JRBksnddN1P4HiPxJmw
rqxcBP6HR2S+PK/pqHHghIU48s/0mkhpwAHTAOWs6zNwFzFyq5u6AFwx1fJR4cXzb9dw6F+VtEhu
yTqT+/rPX6o/eHrPFppEytYYDmZ7oLBL9/JSesEj02gRN2weE5XIigBrov9Hb16j6w3m9EHzpE4N
+x0+4Mn1nGxwDPRlR/02t0FiwMfRQXr3bfOniWSukyOyfi1yIGTd9be/9egq5rlFJj8bmRw1t7Ht
NBy0UrgzlKCw2E7x+WEjCEKPr1LmGBsT9aJUW0i3d6pMbeTmH+ZM9mUevbSNk8GIOGm+ID3o2LLG
wPk3urduloPqSgoP3uJDcTGc01v5gOpa0SuaRCnyavgmQGCkEGswtYFCRCCmb8mFjnQhxnCNH6st
xpeJm19SWdU9h49Oh9YMWKFbGzXq/Do0kgjhYqen1D1Ssly9iQ6tvNcyRIrffWHejpmJUu/eMt32
iu3IB3VjpyVNB+Rl6TNk0nAJaYOZ//P07f3FEhUMG6pPkWsh6TQEhiUWNBwOHBIbo8M0G+QAEiWB
357q7xaSiF7827CdId7dcxZ7+wOcXPKcMmFZAkLVZB47hYe0R/3nd5uy394wkHNpZANstR+ESnQs
jMRfIm15TBHtMDHQbyjVRKLs2Fvc56MojMo2LVW0rsF6+KpjLMN/9pZcfw/SVa+mXqhOG5xYbuZE
r3mYkMfPGwxA5WGsg9MG24yiKisCXUdwttVHOss516jeF5bDNOcQ/2i2nBpW1aCgZNhTC9nrqBBr
5ZlMLiHRV6GIcRME9A3hvGKkLtmH3VbbHyyMdZ+khIBKBHOl6oGjprU19ns6u8IK9AU7FRQrSxwv
RYOOavl1ZsVz5hyGt9AVygpdwfCakBtNhxX+Qc3KfX3JPuAV9moqCZ2GXl0tG4MXEQ+5T6LlQDAS
+ePTQOtVOny9NV1anZ67nDihOXrH0Y/DAbwA6Uyx/RovNIxXXK4rNSBv+0MDO/B0g+WVJL2Vlnsi
eQBo8p3Ekdp5JpZ83yVK64R8+cc1MWYVORIxixbRJ6+j+76ibX7C7AymwUnCkxQC4zH+e6mnng0i
23+XYIeW+xi8ykyb0yeEe8SsYcaEq8sjDBbQBkyqfJ4UA4YXp5jcHAcbJ0pD/kWhK8bCiZ8IxABm
RzcJQxhignpzdygB6tfwZcSLdpF1uhERrscHX591Q1jlyKQ8+yBT6WpwptRS03omMDWxEDsx/qoF
f5zXRV0uBF/+w9IaHI9HzJlWEqdti2HLcsEMBCDtOgXiNj1n8m/rWBERqUCSVsr86HHXrZRNiyxI
zB29Ghje6I88rXslhe9pKPjcLXAB+D8YMf6eFtvV2yRJNttOvj2Sw+z4z2p34NFpfT3cXq5Q2lyt
pidHySSQizZj9NB2e9/zwy2BYBp0UJEQCDr7BxwwCvOgpfKfl1VJDnKKIj4Q1Y2gB7vd2dYq0ndR
tCx8rjpHZak2SjUJIb09x17gL8KmGQROJIUGD57LqaNWOghfBY/hpWvXG/bxr6EDUAZiVp0Werr5
XCVE2jjjx1sp3U8g6kTidWcVI2qLEk+tqFgKXE/BRFX3EUxL/zIsYwqyo5wbrXZy9YwEbtgoQqje
lSR19l/X45OI1NFfaWvWmDAlHiDPnBXOahZ/bFns/yColddiQX1hvKOpV+pnAsix5o3mfQSB3y1H
oorN+U2qqIynvfWtADqvnWX843e6s2gny758efZGNsrFwpm2yAPrIz3KcShjpeixkdp4mpxMsXDU
j1nJhpq05FjiFu6ySQSJdSi9A6xJsZUIK4Xjd6jMIN0Oy9Iq3EY7OoAq9LwmqMZnBGiBUWdosjNc
LQujxetrPAyYO785QD5tt2D5M0qr8bN0Xy9kcYPCjMcmgx/xGcE4BkToIHDIqglZ5dYm1ZHd5IYq
DwcoaU7Wj3TRAtR691z8FOcvDXYs+u95EcMzj2Eh2YSSFd6JuxURJgPS/YTWVf2LEh8q/QCafLGE
BwiXWgHbVKFLbAs6XClC08+NqVBJeIEXQOJ28IEs3B9xP5yipGDiwW7EVv5Qu20mtOlDFc0iu1AR
12g0uQ6oB6d++BC1aGcT+r4I+bHak3EgoWG21eE8J8E9V2o0WVUfsCHIUBs796E3bkn4qiyXW1Nx
qPCsLwQ6VCWABOcbOSp4WFzK84ql5OyiM1TBehwGborKNL+/zEDoGwv0htazc6AthUavd32gxdtI
4ferWUdz1Z0Xw9Ewt7sMLm5QTrBgmAVr9k5BH5eCCq5ErxQQqbWVQBcsLYes5hLxCLwQOH3bH5j5
u8X070hZpZnOTptUYrYHCWiOiUtshODCnG64NGbuu4jGpGgXvL4BsHCRznnDKiNhkSaeP0Jvky+b
839RqFUf8J9bcCfZBDU1dLoRUNObzKT5Rx/pHdcsGtYMUPhCDCx5EcUKFIB3BSrlevyHUfUU/4eC
jdyzP2OwtNyut9KuvNRbGvKv8NvQRvrLtZL5fr3dKe5P4QNWCKYc/Ii72hmWZ8LTpXNmowgwwABW
yg4FNvvsjSkpGKqYT4f7Rn9T0Z5lukdqCGL9rLelArljUMz2zRATWKvAsqJEEISlWKEEvx9Ej9kc
A1Rhp4ovISbwvZj9swjXAxPJ8aR74AzbyDD8qeSomUljpsR+xoY9UK15zNJqlcsweSN4kowF3wQ3
e2zUYWAXK0YGcmhsXOBCusNTsDN5k8f05eoHkQjM5P0wvOpdGrCmuqEUuHn2sdz1CuhAL67ct0G0
St42XUMeeHyIyRLol/LYAQwW0Zb5EdgbQ6hBVWvPLvqlAdwqyfDbau/unTem2bfRwDVEiCVFIkYO
0iaTYuyI/kLC0UX2mGVVg5KRoTiCq1sN/lQ8pqashWBr87ya7VryjOvYmO2OCP0M5fvPO4g9hQAH
I6m6UVCN4xXdqDFctYvAoKVxuRuO7YNO1P69m5Qlh9lhxwHdMN8d8un/q5ULoz5OfZk7LAIIzFLF
RMuFUAh1JQil0yh/DODpE35wmpHtJ+dDPMQYfE0WX7XNlIgCmLGYZYRj4Ew6nhNkXfu/ooi+GlRf
bfJzD4MDQDkvnzT3I8xblVeBZpBgatJxGtuRq+cAGBmvBxklIHhqjtKV4m9EPpOjjthB8kkUCvrT
rfr6YtrGiqoruNh+bTj6xYzsfLt9zc/qzECiKIpW+dAvoaTC68qJJrmKisSI0eirqx9sEeKLcZsT
2YK57tAjd5u1Z7+fS1Ika0HbA0Uj1Ktef9INColPFfjcqacf1b6HBKjOaenO7fphizNmXmf7TPSx
Xr3hos9BF0lnxcAdcD9v7DGWUgw+C9wf2TA6dZEC3eEVNyUwXZjT5XAmQU/QzbslxDhMBls88Klc
Omv06PgHARyxIkcG2/2sYFi9IxbkxWP5epmKS2pPWAvFtBTqoyWWsZGP9AWCe5tBMTg84sOlCA1J
VZlamgnxtQtCx2OMgjDjbwn54QcXqnNLxWwDdXYXAFVU5GRFxh+15otqlCWXARckrfqLPqYEzZoL
qQluf+wrMxU8IPspYEboeJnlWi7nQ/XImqMEtIH+IGnSRxePfOhDifUzTy0nQzcX51jLrrYONNrc
nMUL1kq+NA6jfd6zm0PcoIur7UPwTNoh70p4OK09nvQK1QxdmykHzoRBKmi2YSgrI16KiyJOOuIZ
Rw4kNDAvE4L8z2mIMrxJgvFnl5Cj1uwlGp+HLAi/FG6FeS0FYSaKtd4Sa8/2VZcVqaAK2IDCoOE5
tWRs4TJqYmzYiq9jMPZLEw6BeJU8DOxQAJ/Aqj5VGAyCR5KXiMCKfT8KeowIcYEPIzHcgy/WT9Zy
9Iv6eg3XonhhPkttFKVmQYID+o8fFwngaHis+v7L2dTn5cjeX4Tu0I11EKonKDFjqCX0k8s99ysr
ews/1/0S3cQD9//NXcPm3CIb+jG9yxUziRcgCWn0oPR/L7E3ndBAjKqARUELhzC12myUGJ45923e
FXpb590uwmjEvKSWKiPEPu7pw6sY5CuH0UntrmFNejAMlwxgDrS/F+L9/4sfD+mXKNbgOrShuvk3
zC+92/I7jn54CG7DhQdUlHyNOqJo0HuCqJxFBBmRpfi6WkJHNbXfXI41yJRmkmK3vp2IcB3aOL+6
RPs5GE6LwcUEGfVIaFIoVZrkIhnWXSLuTTvzOa7CgIgOree7ZOLZCnTPvGFTogVN2wccBIi386Pa
5eW64keLszGyAhdc2dEY1BziXSz7qCaF3itnPvwu5ofSC0xDRPRHxm2oh1dhEW24GeqzvZEpy1g9
RjuLVCygeqTuASkhwCgu/ZCnvWeur+RDUGJkKiBwOg6FrdFfWKLTHYnbaaosICsJoP+Un3+sYL50
+0asVplUNq53hRvBRARZL7T9x0VZtUzZbMwrfOkclzt1IwazN7mkZKpnAjH1k/fb4Ik+fj3Jb6Xe
R2a/zeqd5YQN6ryHGFebsAgdY0U7D2xBoyDK54M/0VqoAkX1wYU5621T1jqpXqoHbzeUpHMXdzVd
tW/DSpDWkVyLuAGz0djfYGq07oW1AibBAdKCHtgoqcjwXzFIW02OFHx8LYVcP8tFBEvBYXUZiq6m
3zhQMineyTw7EMp1K7114XNa1pDlyMaTm88e6vy8YkCQg/gStVGFWhqQpk/XR+MkNyv061GjQuew
4a/T7VAKBzmH4TKuKChvhLl/1QYJcwah2Ptmw6DHFvVrQAGO0v7PZlS/zer5h+vcFR1afTeg2pR2
t1IDD3zWEv9RTVjJlKtcFZbLuO0/Xjh0D1SOosHY3IUbKbmvgJZabhmmCBE3qAOOcYBoE8rbh3PM
dbvQn7ovad//HrSHm7XfLCRiGwwJVdY2Yt3QKAnnNqJR1UJmZxLCIU7JrpZJN/MDvJ5V9hCpkB66
/vZsD8gGu1xuY6VpdPdS2XBj3CJL6sNCiiPXcWUrozEwIQJ7GH2FpTJDZ7/kL5tRW3AcDnfsQy9/
gCTZtCgAZHZd8IzOaB2ASOvbFThgLHc/0jzWCGG/7HCuvsvtJGW3yIG/Nj0Ex8qppTGQmeWTz7PS
gvStUr9KZnZKiXgQE7I1w7WbwL7daeE/RUH1qc2KenIfvxBW9Q13OuV1n/ymIyXVpUVNdLeJ+E5E
PbCYuHuY+Fr1aEQzGIQrYtu0Cg/xECQ5d6f+V2TxWQk3hzCZZdAjoGLDAIxDEGmm2kvp0pj+NUOE
9sjrEy7xstWJD0ivIfFG5l0uCeyCUtWv7tC1KOBMYT+BTUxiPrJ3/LLPdqodUlWYTB4lZCJXFJ26
6S4hku4qO5S/tOfZ6B3gikrVEMf4bpgd5OfndwJKHZI9XrI62Ua4LWSACEIW6LWIcLgNEODYkYyt
cevA2EaDPsu2jPMo1W/uKIG2cSTA33OGqGA4LjEuOmc8GBbV52PcyPeVDC1qvE8yQROfMWdAktyN
wCuqAe4OILr46Fc4J9TvDmSTMHUOPOI2q5xRriJYjZnOk1HYX13JQ1oZ12sPlNBRrkGvsY+iEL5A
tDU++FM7SHIMkh+p91NnEq0jvHoQk39s7uQ3scgA0bCstwF4IR+T1sVUHYUQMuYX+qx/8lcHDjQJ
4N2S/tKG2sl7gcSeNLnieUmZ/Mh7HYkoBPtN4+Efv54liu5utQCW+dVNugDtCV8CKxNWGk1y5W5U
FXXBxpXGfHycGHmBppDCpI96Pcgy6L31kwTzlsxtXMFJfWF1U79GgB7sPXrim23WH4fBzXnBwo1A
zEeRRWsr3hH2gnmMMofYFAgLbVJR2df6UYyywUSejgRjtqFLoY5mcUNP56mh3+CxpydCLz04OOTJ
oMQtifkXz9ssnHWRKVqMbFVsq2oD+ctJlKz8Y3fSnASNHe2JhNt7xZ0yLW1Yk4JWcTzRVV+A+5so
T9/mwaAa1hbKzV4kCeMzbhG7hccCh8zu4zoJrDduWxGpVXntQa/r5hhstPLDxowmpvFpm43p3etm
dgeAwPkiUtq2p9TXGiMsOeYktH/g/E+00ijvHu3PVMdSuHs2EUCq0iOTeiBYdMkoVCt+oNxrfPNJ
C9ms+GgJ/LCKCRa9q3OtPSZUaWG2ZSmqn9ddOWn+hGCWHUffj8lGcnkKpN0WVWKU4Bw2AnCEnNF8
il7/dxtk5sqB29aQFfuFaGMliOYRZhMlTDOruL38Q5sRc275hqRMsHhJIntI/cC09DruznQCMpH5
ItTm2YWm4ngjUnOuB/iuubvpQL7QzgCj74MmR2txFoDC9tmzxUz7Dpb+uqyl8SoFPqL21HhtB2dl
Z1Qn73JkisuhfLWQXIo/AyOUc85d9dkDOT+AW5sdCuBX2d4ZIhK95XjmeAjs5FlHkrf3WKYFo9u7
2nCYRCflKOQvjfJ1UZjBqeSM4kZICzV1gGt26VVogNabx9F5p/h9mln7PQJ4WMzuIOOtxmA9wArz
B1UZv2BnskJA1RKxyoVKJwMQEKo9OSDcchzHZeMn931t3TddLP24dlgQGuyNf+iMQwnBSNnnupT2
+oITSMrEQDlIwBghMzgt0d4qza6VzWxDby7SeEdljCuvUdxbnSDwWgcnaPst7KE73gYJUzdq2a40
5dHz7a9fNBXHm+Jse/4CnxJ5OXXxNMaFX3xMhgOIN/0kKWSUEb3gJiUhpjQwxPQmHAGDOsrmEdVA
wVn2H8FkLFYBzSNew02/sxbCX9pW+f6qxs2O1fW6fcV4L+U6vz9jmaPutL/XhB9ZaoAKUOX+Qz82
OaE55IqYScKx6itHMaUCXJLd+LfgiVW+607u/0ZxRDcD4+u4yEXPXLS6PwtiGxX0IOsUehM/RZ8W
MA1P6HDujmx/NFTezbqvAFTpBSCHVHlpX79jYG8SsmawIvvE1cpgpuuLqr6crOqW4Pr6MqHD7uvx
9ncD0B7xumL4xwiSQQDVg5RZPtwFyG7SDEqt4EilQFxMgy4G5Qojmu88y1BKu5HbemtgY4+eGiD+
MFnZmat/OMVE0YdV+JYSb76lAhwb/8CAw5CzTJAXmZk6dsoiUB63TZQAFZepDA95Hh23WPG2wND8
5FvkDyegUSV4JF0GYZP0LPdR9akaeN0m35EcizGcXlTReIjx7tzKlLyCK8qgY79L9con1xG2X/ae
MP4sgz+EX+t13bYjws0Ouxvkpnw16o4SYsN+Z16dkhnQT8fv173lPCiA7AjRXifLXKs6lpBvXVNX
GiyVsOeA+gDjQu7bdgmDgYI89ELWgJjzPe3kjW3XVhM4NR8XZ+Oo+J2vhEcYEwL4CFDE34HBFb7q
z8bq/GdcOGiRhtSE4RBe0CGthATmXW5Dco3aMIfolvovirkmQOT1fNL9h0IhjM4p12DX58Y2af/z
AnFlQHe1+xP//A1ZIdDm8WU5os6fWfm8nZnUXFN9DVImHJLkvRivkcfKzikTZuDxThO7xuBZQsmU
d0UPL2i0ibTOiPSJg/lvjKo1+5LaU5e6AUURn6Tpfd4HqSFLyUK8Hu1Jen15Or+MYY71Zhvin25u
g/hBDVfB5v+hY6lgcSfVwTk3Aw9U0vla/vTHRByJKzPL9JokbGZeOy/GUA/vWLC1NCx7k2rMDraO
SzFbOquLdDfHIFzPfb/+UTUkZCms62MyPN/VtY0lbjIQj0XPGHaZX2Bx+jjNYVgns+hXrt83a2aL
0MNTjwf940jpxLeee2bRp/A5jcrUwjzlHfQs0Dza1Ynhp6Nv1TxJcPCOPpxCTQQzGFb5wOIAfLn5
9m12hCwaV+JkaXB6AMqV1taunGAhrw/CqKqURDWSyhLAyE/jn5PLk4UyMTgE9ZAzaue0hr4FKYYV
5yS3mLLaB9XyEvogmIQ2CIcP6VgS25mM0iuB5YMWMAK4BUswKmm8B6Svps6yOZoUGaS85orMrGch
M4iD39Fl50D2AeKkWDU/uHfBmNnlBg44xN7z5yFlk1kG7X6YSs2Ty5o1B67nVnoXPy4I0/hFtqqy
DIMIaS1a8WihjuL1BvqQQTpgM3Zl1c7KNtfg9R19wUL7+XNFWxKcv8Qmuo484rnaLjSoVQeghYh7
UWx/I7rF/ekkUc/0PB/tL9KygI9aEbdrWBRtqITFAKoozBxHQlobdB27WvSvM/kNQrumRiPm83y3
qcaNNwFSwuMfpFGU/3DCuuJp15J8lD36mXEjVF6Mfq3hS2Hv0LlrkP5h4p09w3VG902l8b0VBQDb
9/3X7d41ltYHJhs1h1+FcqKYaJy0nmW0fV3Lwm2uoDdldEx9twaB3jSxxc4HUvTJs6sWB4d56fTW
k2p7VI9gDZmJ6g2AhPB3kPgl00DMxzA7+DPnGq+cnksaueVe1NFLjrHyDVjmIQlkiDcoj+slbaMu
co5YNRzJaTVxV81cc/nZGvoh+UFT7Ed55K9N8zWs7D288YmPYUrMqW9oeEH3p5X72sw2hsvb/JSH
SSs5sN4c3u9koiO6Iuhnd22nH6wb5zowhrTA0GnLnbz9GNA5HETeXInmY+UjVyBwKrsZSy7tf7TD
MiwFcmqEkHldnkUASzWxdS/AwoUAhNh67RXGeCjULjgbL/1YmEn85cpPMdujMjeAQ0qtKrnKNMWG
QNMwujzMNaiAJ4Gep0ipG5TEr8G70aMUBp7sX2A9VKLiDDs3hYqD7UB29KKu40tCKLyjoTgtYWw9
SOWJrJjkIbnQgzO0yT/zhsUiKb+n1a+TxaL/maMiUyj3Rug9jg7AXccTwi2kyjjXJdGZHJOWj2VH
bwiJ8x5IONHdcfe5kbXfyj6qeD6SbhQksVeZAkVTHpRtedeLjOBjKjHH+a/X/LAkJN/hfOvsqesQ
NPoCv3g4YCNrppgJQyGOKvfjhxK8XqmNmpq5FW7XBGAFDS9VVcBFe9E3NDY06dyY0D5ZeK0Co+YD
Q6C9eXV/CvfgE+5pM9Ntrzl7JlqrJkS8ziSgs7fb3XnFVqzXuq9lRMMlTFbAPMprg7eNUAB7iZys
Lf9s+ekkrJiKoK1Tq2kJB0th2bT8QKB9An5Vlh93ZbOK14UjZiLktDSoBRLTNqW8GbVEyo3G7Xad
YXrOa5IijvdDjpRRQ4aLA84YwwsL9pZ8LOLFhAVfuo6BhaIEQltRJkp0tzi/V70307NorJw/z80X
Bg8v4ptbuUb7QvWT/BABxMiNNkdvnLXYKp0aduyZ5UBegkm6nrQE38YhB/v2otiz6kMcfMJjALp7
xWXIGkeAqm7Hq1GzYccMQOfYh1jrXzCY8Fec1dfNcnzqZ4lUG/Vk56u59k+AGcCEizZtNIQ7BSE8
nfAoyNLJ1bPPPQF3yQ72hW0FKvfBr/EDgULTRcvwLegLsfy+Sh2Wz6pQwphfL4fNosv21tTsf4Wy
G+A0p4eE+8UB1AHlso3cj3hFjN2yUdInOKmrmOANweWOB9J43oEBrG10oMj7Yt/a45/rffxyrbTI
fV3Bb0AHmoVl5yJEXoqCVq7JJ3tUEKF9tz0BeZtCE6lcwsNL2tJrbDOy6uX15fy7sX65/GDwtNky
T5Wk9UApzbIH3vQqjt/UoDZXSAdvLAQMH/lysaMNU/qB0zVVeFjbLCj892LFP0SJyUHx0FtmAtms
Oe0Qz7jvDLbegrYNtp4cp7TJNo+zsJwCLiXjX4hq/41skkGqM+eoX+3FwfRelVla4jG0D1QMVQaE
q77iDnymzY0uvvJiluFI41sKb4IWIsmpwwHZYX+1fZvsbVNzk+9UNervnY0Z48TW8JhrC3v2/o++
u5oKU7hCHyylsanHAC9fgHR3eBo0VnvHEFSHmtg90/x478Qtf/u4+eD8iYAq66+KHPLML+Gm1vyh
Xf/oOCFcdHNnM6isRswKJIWPuZxglkIfxo9hFzWr0Rin2Zropvtzx2OI2nyvK2pFU1s9+AfX4sry
XP16oNCGNnEJqYWTYxYbfrR6KbRQlkAfsylqJHANo3TX6YkPMNNKeYIXLUULQjRHAs5mI40df6rS
GTf975JRK5DdZe00nVOIF8sHMezXHFS/gMcc9BpO0iu9PrgbyZLmrFPxvNfrZdwpMsRYspL/sHhM
rzrzvaJrSBTriIJTB9YdV5s2ZL2y5LIyidMYch8Tc+7U96OLX0dzYrFFMRnHG+grY/zWdH/xUGZ2
2aIt8ernj1WuyEENbmjLGaYD2zJ1FbgY8NGpqWiXBV3pUOvWVRalJEO4ONXxRpdUcsu72MkEDKvo
n7XwZelOT9IquTivCOX7osWaS5Y1RA9Bu2BRZweLoDpN6VbxentO1Dh2p5xfJ9GN65oAlDT92i2G
ZwL6/SY1TWOFIb6CiY+4AAGWdmTPVBZ0cOeMA8z6pOc9rTlOhMKJkZOP4dO/Ih/rmA5J3hHE6SOu
dJrEwTHi5GUV8oke+BE4/S76Q9Qdsn8UjyRI8FCY9l8bs1bVFZISjbJYcvkpFfwrJ9f7vWG/3ozu
AksQtz6pe9k8TBiCDkKkSv6U4po5vv1GZk+Qr4xxnABdhQMHa+EWI4nxK5QV+tk36/IwL+nt7ow3
MQVvo+b6DsZq9aW/J6KQ13zX2p6CKAfqYt2haxGtgiQrFRgaF0oAPuto1qTCXt29+mwV7CJcPOcF
KrRt1B2dmXC3fkOM4oPZJO4lcfLovJ9x7GiIwsNlWCHq0wm+i4Uo0AbGpH/mJOHa1BaVnPEi/JoP
Ba9dqIpX7zR1fn4q0StN+fKD6uoqr2ECcjOh0YMPrhV/jIA4/mebSTfbAJTGffleQBeyTOxgZA6s
rp6grSpAr7w3RWndeJxR1SK7Zs+L5CvpJKQk3Y1QCM1r1QarqrrYmvw/gs5r176emep11KQ64vCs
xmNj3QWrQSANc/UFLAKYpYr6otmWUBKE8RnTycNKdLZjWcB9AVKb+WTa3lLbRd5rHQ4QlKU0TGCm
ssnCglLfi4hrYQIFIZoKYp+e/j60IkI73bEzSWKcXf91LjtlI8kSK0h0a/mSROmtgRW58i9pVIUI
rfXQgW2ZjITF6aEDS6oKzpYbiusv8zi/dunQF4zTWkXqN7DUa0gmhsYcbD34ce2yOonEkhdsdGCs
3aCh0aEvmIC6vmMpQoXyBYyADxIE0r5wdQLlT/awb/afcgAqME3f7krb4zvJ/fV2ej5mV4gKIEH6
Gao0yUOrZXxJY1mrPEBRQn5Tze0V1q2+K2DktPEWHZdPh56FRvrSbLewXB6qpn5uVMHbXU6qc8IY
6AYu9jGTl0OOLlP5gZmIFVE6D6BDrYY2kXvcaA2EDhw9Z1b9VCKmNV3kMED+P1e4l8XzeNH23mNf
HXgQODLJI/44CFnlbYwQ1e+/5L//EWc7LbHpU1+WTDG987EgNCOxe/CfkLvogGdAQvd7zwW1KEwy
omT6b0o2gJDBGoavrfK7TwVKMCAhE46oP6BwoJhT+oKubQV9jJw9G0Y6k9vPEQ7gqYsC7k2XtO3k
LKdMjom44uYiX/gD5czGglUws7xhD5bw+29mlIt0Yi+kQeP/SIinza+KOIl5papPaB/ClxgPfOL6
LhQBcfI9wM5UjyM3iV33YOgPG+mYMO7A/Ky1wIG28yC9QlzqwytJXj5Tqivl8r4Yov1xo4n0aLRi
yL4BxV3jIl9EoNYGnu07QvEVoa7P9OH5TLRoqzxsDecjTqkvuN6p3HSKsqAnLCnyA232GyJkPMX3
lCpUVuDu07IicWq5W3cECRCD1wKfhE88wGeVnaYtBZZyJinvSjFMftRqUC+jcJkIaHKyWvUuGG4T
Czc8uI/ZLyYRf/YUBXvROoS+ps8sRlYBfkzCoLv1M8lsNS+MYqDJtnV24zGMoYzuLlxLQRnbCUlh
+7uh3oOzmoqOeyFm3jEpMi/nF6Pt6Ou/+sWdoBo0sq41KEzE2yvnv7LSgRI6qjbOZq3zO0FzPP5T
sEEPJfKw2/Rjr42w3xbVwfzf253t9PCas0sJSyoI5uptZUAGowntruqF8IJViRxGiDH1L3t157z7
x/rtHsfoY4ITm09cbCtxNKufiqinQZOmYWkkVjA9Mlc7wRbVU4PbFU2vQFOUFhs8KnBpTSs8sjz4
yOWpiNoxrWTN8WiQF4BdTDtTlpHkFwjb9YaV/puUET+sXIDjFCfX9/kTmGoyHv2PJcWFv44iFeqF
o7Ig9Gm5Foslig4xcpRigUhT+sSR9aySzh8ZgEgKK+iqaFeHUUURedIsvpHLnWEg12ol6+oR4R7q
SaoFN52kHg7HmHnB9SsBPMmGVByNFo4kf7lCGqOru+8eeR2rDFilR2NK/ArCuC+O7PVS+B4avlvJ
WmODkOA3oV61VwHHkcMJJIBKymGxW1deKVetY2dP52TjxL7G3XOP9ewzCdu61Ah33/1XByIiDR45
Hid1/L8A0CPCHfiTfJpYrFBMgtC138gEyfWAHzBtfMecxKy0enM6jOpPiI8ZO09IxSu0My5838xK
ePhEOsAOxMhu4KCL632HM7jwjDRTXhjCCUGqUbfqPQH8luNwV/3ePV5OzXbY614aWYfKCVmSFwJ/
ASvY6g9ff49FyRHxCFEFs4zJpH3Wb66/Myu9/R1L+UOiUwyQNdShkfcqq+fDiv+7BENBKJDA6PjV
sKnKObrawPY6ffty+D7hdBddayG63kZ0yMczcC4HW+Z/g1pfZJnEBUYzNSdGyZCiGINk5iJJrgTd
XuJ4YL68CJXAoZa5gUUaFVJl1G5OupLwO/JbwtSUF7+ETRW+TCPp6eenwcxLnLV0H4hLah1hpLA6
jKlJU5sebzFZNH/SB4BKGaAWVZzhQ+DOeNTa+LxRYah5Wzb2SwdQbyrqaAw8MIoB9a2kUKDTo9m4
0X858hrlRe2oxwphj5EZxrjb5HRqGaYn/VcFidS27c/kSFQKtkJqn+lk1SeFzqPTCTvCWwdLtD2k
xBZRLfbOZCDfbizd5uVgPVmd4SX/BOFG6C9APZtFzU7KaxPAVQvKYmEy5x2x0dzDR9/+KK5Iwm01
TdBIpzjetNN1dk3+asFlXnUsAfFUoG+K6lzMdw7h/rAgZKZImjfnpBJKFZ06YEwBGHd+bjP0nPPi
fcgnLswaw+86/wR6Y/+SyN+NWNVHOr72uzz6ORrIFBQr42BIimqPbLvAdbwyn/62LbmQS90WAgxT
GZPwntXp/s4S+gxt0CLoWV2Gdxu5/MsdtQDbL1eUBNUqbizZaRITnifyviEyIfFSFmnxSN4J+poO
eeMSEzbSiv8ZsP2ZRh/vj7oMaUUfhmjGkb49WjrqQ9YcrillcbQWZVGcRuDtfo5EgE8riAQDaS5a
puh/LOsetLnmNCqXbEgXRyH50n1ZDTh0hJMDOkBMhD9DSlzOjv2V8XJxcwJZcB2VcEUU+XFEbn7X
GIeuj9kvXraHQKuyDS0enP7DEcPfaY2/bjIOiqhAHJtr6dV6xZ/7oXLS6CeH4sS5YaiARmAU9NOv
IGgzxbouPhL91HdqpY6f3kIF08snNW5zX8D1VQtgD17uq12PicVgB8p7LoZ+CnAlzkoyN1MZIpLr
MmiPLj7Eow5HK5KE98oizwE9uaJNJudI1VkmWAqH/hTErnYm7tMOAZq2mOrirS5oi2Pqsqj9MQts
GXzW8PGqmN4gs7nHYTg4gYWx6YTlZ5BTsbrdx+vxg1w57aAzbPeNwgWomcW65iVfkIMipzcVcR2Y
HM3w894iMQLeaGAHi7arPWwIBvHngmpRFxuvEs1U06gP28nQ6nmuhICECoe0ttWqImGsjC7MXBwl
jaiCIf9jUZ+Op2+UUmom6ajtdYz2sy/2zRtl1Hb/pMUfb+Vy/11FLKdCbhGoO/Jhug4nDLJlbANq
AUXLNmlirpesvHMIZer8ZOTwqr4wA28J5Ipl1Y/BwBguCvluueY2m65FCFr1GkXXxe5adeiBcPET
AvWQZFdg8GwddeZUtANw5/43aeDCUr0DyX7ClkRg7JADWXB8nrcjlAK0IiZ/ketrHjh39+lpTR+O
uBdKsfkWzOcn7H036/e3XvP1WbuSQMv7ZsX5TcuALKB7xcezmsGEJHZKegLN4xOCptt7FT1tXxj9
IfeZh59/lK5maM30+9u9P+9z4VblV0bKdxcdmPkMPNgS+R1QQJH9jYCAGxlV16xEYEPeDHhuJait
duqCEn24pwhw5mQbvrRVhvDeXL5iWOCt87R07rRgWFqLvyNln6G83OPjEaGezBiGKWRyzZ+wBfQw
TisasA6Sdf9kKpUoWIpK9rpmEswW9Bfkhn2tsSlwM/bgjKc3iIxvxaQ0tARyPc5YeEK7l0+suZKM
hBlijT4YZ5P9IkbGYKuJp/8ffR9ej/VcyWN93LlrLzKjAWmvSFBSz7bDI0M7yQ3WGDrFf0GAnPaJ
aqG/rsmgCPByqzepAgVdFc2c58I3bxxBCcrqd4diSu805JuwuGBZdB1ponH4RYN+bOEpoLIzVxdB
CREB2ogItg1e2Jhw84YjIcM+GY7/4sNOo8qYIks2mVLJW2IaHaR971fPmskni8fvBWINNjUbdAFr
MsR0wJA1pBiJi5UjWDv97TCUDDtHciJD3x6H8cn7OOH4l0hANMw6DD5tedLqPtWG/YeGsXQSRpAc
8VV47HcAEWSd3Rf4He/4z6QIIhMSSOhSQC24K55WHsa0Ll5K3+9ECsWIbVyyXZ1FjvTbAK7atN8z
kdcSSckiDMFllbriLl0+z1K2vefhwzIDumS3jA+32ypndYCX6X7tkNxbrxsi0nTUR8l33k97HlWq
4/vPyfilagATvlTIZCqrjGFafvahEktHnskPZhdZrowynGs2UEWTxlULvmCMih5wOtlHPZ7oa2Xr
J8Q2LFDFX1ReQGin4nzHRQUOvhqFq5aAHrU+0L5vcDAMSPt+W+L7yooEDKLiK0J97J8+w96Ejfck
L/219cXVMLFXKy/Shp/O747ZBkzUSn7nXfP6BTDWlbHCaBTjwhEOT/fhfSpncqiNzUDNnT+clom7
QEdnvncWzv9r9zYyUkS3/7V36F+nhvOABakpknvGFQMeuERHk4MYolzklymw58JAGBf3eFAVdikT
LQ04gIsUpxkRMpIvv7r2eBbQkwuhIJF6DlYQltui8bG7KLVaZuuXx5ZedUMdN8VmZzOWfvLVZr2E
0HuxoFuMoOer67040SLxkRC7QIX+LManmOXaQJLd2g1HUt2yoOZ3wm9dHUxcWNvqSqj3A4zMI0Mm
BXF4sKH/VqVS21zbjFFEJ7VTPbe+VU9DUqeRMgMBgj7SESQs4rXfAWeGbuZ5bmHuj0GqaYAwOQbO
SMgC9ZKBjmBJFQ0hMQKGIybbBfP3G2It8EMGK5okFPbbbR1JmVXzBh8LT0fF1v4Hm3KncyBQT/g8
nwPmFkx7G6zczRMReTcZTcNMVbrvVeCLfxWXJmCAtm9zJq/mCSfojoRwZZ4KvInSYRTJoNoEJni7
JS8HP43HaEWhZ/60YohuxEUwsKOaUveMa44iWHjbfNMGO2C8NxjYuRxwZhIwk+eJ9rf27gnsdW8O
VicHkhXtWTACrc3xyH6gPdWC3bQfaFZaa1H5yKqJETHMAfWqjzPMsGJsBiSr76MkJkCWwSp7MOEE
tXiUUtiGmL7kb5degyoTF2h4lKbmVklDl+5rOUquHD3ltTn2/0ucC0RZhrp4NDRJU6OxKspCQoUD
tx4XBgv6K32nVSQbVB09OJuBtVOHscSMqun6genpUbq82kSH1O+dQ7FR7+PdgQ0N9ZQ4qGJYVAXq
lDDQfDt4/3kK5y4CyWDoVL82COdNx59+w7GTsHVCqkbrdUHM58VZfE3GpTDCooVtv5yqxjMZKCPR
8C+FJWEyNnUYDcNC0FlZkIZqmGVXaxkIxTqWOKWVtrAx7xA3M+aFkkczlH5478SHijdAzrpdYjtv
BBuCsB9pMjho7Lgj0ZBP3A7D4zna5BPmwKCYHt44oZtRVhK7flcVCdZju9Lww/Vyf1O9RjhIVgs6
Mwfrs7UpUJra2fegBVV784OaQ/G/ipokCWqybeE9qHvveZHmMp03HWgdmo4RYyuSc39aIeW2ae6X
yJYu0tbMqL4JX+hsr65HP0JVVhJ9vdK3fQlxKTXbTl9TrtCQdVYQ7PA1I3+ZadeMsphz5MamNJ3I
o7q2rfl6UcFajgAqvu/en0Hpgo2a6Ry5l/ySAzMfU4gN+UDBcBjMgtZ2EMNPKt+sal5P1P4qd1ll
9Yuyxx8dFQukdX6IQ7jnl8Dzc49XMKe0Iz/zv0o9MK5UOEoN3UnHywVG0Bvxsa7Q1WUjWNB3JTQF
1WYqRg1YWrpx//u764huidlCaQxfGO1oR0O+FOL9FKaIeB2CfpWUuxaLO6VU1aEy2H57oIsDTQH4
WLfVOxLlW5PNXcfYGjSbNSOH4z2E3AWN8xvZ5nMJSvtaN5cutg1t19KUQBoVR8nbF8w3Nzx1SrnL
WIOTJDDF4k6cg0IKBwSUPGzm+lkg8e2m6tXu2+KK4v27k2jNThBvK5yENoMHy5C23NcIZp9kh9rj
nyIzhE5IrtZ/IyL7M7GPF35rFpoEvebAkUYUhHC56OvNI9SHRysn+Laljo6TAFVNM08zRv6ijK0j
2e7W8Sx4e55jnK6U7wzfMjVk/Ppy4Q43dWa4vGKWFbuisGEtOtdG4I9MD/mjDVhOUH6cFtwLmRNR
iQjQiLNehKbRNfZb491k2ZBNBaFvC0wbXMEbM3CRL3F/t7nGiPHNVu36jgYPXWGZORGr0nGZh0Nz
B4vOCxudfsVmWMRXtZaQgZYFtJb1tEQPZmYtnn71O/pHZVepYaYX35J2N8a2vhEvSgx89grkM/W0
sHxKzgyM2f29AONqQdftu73VKES7EH1Mce6zHJAlITc7XyoJp9upRVZ9/sheX7cGmAu05oUkOvZs
DB+vMZx9KpT/PKSTygiipRFWoueFONSsux7hLaxHSlsfaDxQGlyfOQ+ex8iYYSO8zBCTG5eHhEia
Jf82nYwr7R+3g9iLVU/5us4cu6PPgj4Z/YFoYLf7ZqH1NNEAZ5Pm+OrPLX1ocNWo5gLIE5QA1AAy
MKNihulCK2EDBb4sP4XVLFkZVG9j19CbvGmaT60jpp/kKpukaV1Evfojf+D1ODdyDJbwBcmE+xuE
K+Aw5GoTAAWbf1HlX7804AzDQxyeTff8RHU9ovblXb/xoLci+c0pWPXg91aOudV2zpfY5SKl2Qkj
Td1LzV3mqCUESFjpCsqM2zj4wEAAz/rtazPdQ6NfSbM+bDBtxBqVJvfkTUJ3wi6gWNH0KgNu2iKb
oCt5A1GwoPfxpXDPM49Re2CRj+sZTCdVt954/b0Uzgnlpm7219KYpFODVY+ZoDSFqRp2vn2WiMeb
dGtAwz5n6bO3PzeNWw9pdwx+smIJrL5oykOi/rcJCfuNTCEm/6Fio/VFQO8xrqqX+ypbuJFaUA12
PW40b8BolHXDJyJi7Mr9UdIcBK4AWmJSGIN9GwJ7cin/T74BidJ2Xil4yW17QiPzEmDJL76hvIk5
wxw3NdmqMpB0KaYBm1yBY/mneOkUx2+IL9ESCwWguI56t/xbJVuXD5IQOuVAD2w3KPc8Sw4fMf2C
bRP3SDyuoKKECKXYwqTsFZYouyfuRfxaVTFvzR51hDXr8tbbrsvNDDBfeD/NEnzli3UWc5E+jfAt
U/lT4zVz68R0XVO2hJN3GP4nT7faus+vUF5TcoY9nbtH9hPgUonSxY1dqcGb0gf9DsCvSL35/FcX
KNEGTnZSOX7rJNWoq1tHpeb2iNGq93MWO2oFz0iJFgBRvfBxlnVVsTmnPWj11iqIAWkPYNUYPSCX
jl4T8DhT2+XKbNQD60xsjFMsbZx7JRbqYHPZAFhjY6WQNRXymfnByXWSzcNUKgWlnAVIoPKPE/hO
LTgbxUODBW8Bv9GntqIdzWkhkXitqD9tt9Ppr7LN7cDtX7xau5yf0CSj+faLrNqbvFTNZ6ChcI5Z
q1Fb7pPWbMi6dxMxJfZZFKx8kWhpI3FUVvsOR028PCuEZ5IY5U/hOEa784W+/DBev7zHuTMkR2I4
XRQiA1cnhYtQ3YvYIxSlWmFSv6ST+UNmG1OOY5OwqKUfdUD1RnIajXogTEOEvzqlnfCr7tGr4hP7
yBgO+WbwI0omF4d/OouEcQBqg3iS3lYL2ZOLXkpPYgl9HOtxz4RjFG5NSdFwYKKC46q++4KtxF93
e9f+FQr1bp2K2/f4XMLNKKKvfSQkucjJACawOG/SbB+rJGPrNYTkhJyb9fmEpCq6qOCD+Vf8tG2w
0hiIHeNwFQinXePWfYIKog4gT3SQ6LmDq9KlYcl+V0OWgjJ5QPwXfKlbyAqSyE5roELaBdhBaCiL
2dSblBAfikiJ7SDA7nerPfpEvvTqQXuKFxxn2cUAOznOul2QyuSHajvIrLHCFheebP4Ddjxo20tB
23TYsjuIwotHPGI/+XluxeKyB6oPSKC0yWNAB6lvo/cOmNs7CD90u+mq8UgIsBm9LDfm1dhv4OgY
idAB0Z1cmCRbSDwwe6Up+VlgeqiimgAjtDaYGu3gq3TtRmKoF7+WG9fa94kMA0KJJpT5YePKlvRK
eWI5Yq7eLCCdWh7TxXWiFBUnMuwXmLJt5NYipM6lVHdtvJPd6jjAFGE64yddCvqVtoCYj129g7eR
yVCzthpdyt7E7OQX4AkM+U/KZEis+HrbB82z8ab2FO0nqwRfXhzu4FwFGaKk82nSoJ5u+FXswU/6
BWDigJsmvawyj/eKJxZDH0MTBAXdr/vCZjidvEK7KKTOJP24XPVH68AFJ9/CmT1a1FxP1GDPA1sE
XLaRB75DB84HMuLMR4MnsXwvrncv/XBspnmbjc7VIg4pOAWWSou22gFyE22l7CLPdmgRZ2bdsQqN
OIMuctuhfdTEdBWxLU/9tj/KorJCAUCJBEeRl6GIwzqi2y0LVdQXiVBvXEQRSbChz0+8dP2JkQtd
OVKtQsB9Zs2hs4lGTs71mRgesmzXc+e//DUjS2trkPW5lO/w8dOBGk6aV+j6xAcyEu2XqK/JE7Ef
nplxdYFFyIPf+F18wzFmKOMYHjK7KycMNfflReNv1Jzg8K8PqfOvlQ5TMFtCr2Y15ZFycyt3JwBh
Aoq+K3B3DWW6vv/0O0lnu7+ocDH1WrNaO33aZYPyb0IXzVAmwfTT3NJNSZAhGA3k19SPRL8ST2Wq
kFJA4ouz+Kl4o73yJUKdTaqtLCb352u/RAbHfzrn67Z91+FpspM9Gdl/6QQYc1C6h2n+Xp7JUrQJ
eyueweECN/LijV6VSH+k6/1lpSM0DKpjRphrXhlqeuCpoGxSac1+oxtOMCiEbVtKn3fcM3ysBsCH
IvGKLBz8JCNoIa2y4Xx/cc7Y4WCbs0IdMhdt/Mrd1JieKxZQBCt1/aVihr02BAh4bdSKZ4ohljEm
7kcfEANnhv3EJXC4O7QXB6fuC7N8oPRCLErfmw+/3aQotK1lM8WOkDBDrzXrVfcAoi0GRBpZTeHP
47B2XrF5bynyibt3heQIZabPyZCnn2e87eu22TcnyrypyuzqM9EdvQcVitQZ5LC/AVrQpWY7tVtx
x3cgcyalzTlpPzAcD4Pq7jjPkMZY4HxvmUBMSdRQT/VMYLvtEK4vTsrPlFW4tUmR90ExuTCTYF/y
YD0T7cDI5IOBoHu6Nv0lWjcqt9Ym0JEsoSF1vGThwK9pmzrZh7oVtkm9pZ0NYMLoKxQAiBPNMnjR
hlwhA9XjcM13q+RLrNkQpNtC6iaA5m9ZR9oeQskkY8BN4kGVTBQ2CqtCVboXEFdr4sk+gghnX4iM
1RhZCHYIB170Royc4+J4vtIx16sBBYyt1bAcydiB59X/Esc7YUyhvuxB7hCYpcxVkgT9P9nOk4AC
mdLR6z/ucLx3JKjtlN0fhYZWFukIfOXfpEOcFsrCM8B1YyjmTDf7sU+UWRWIZ3Vu3t3885qb/Evp
kcpcHrBqiRFmR+5GKQN1nF162TB6o1xfc9o83R9SMcMW+Psyrrp2bRzdUTB4o2gCKLgmN4MapLad
TGBlLnA3oMfsWuSwq/erw7uX7+b/XtgPtMKmd+bJAS5Br8A9a6uxPtmVKHGfkXyrwK89D83D9GII
92/S1ojPs41Bpni9zz6/CuhUGSrzupU2PFJIbDyojh2gdgX0lE4/LSL8N/eUepjOS6989wx6/ubg
ZnpssezymPeo6CiWb7T8VG1mxc0U5fIZc5iPpVgrjroLpGSad3ivP1Zzt6hMwc82wjpr/8BWV3YA
RIr7PiJ8ZNG2+rPOWBjT9xgIOpUfeRaJ8llc1hvQ7KourBKGCOwzWigPo+LjV81zkXD5aJV7JN+V
UD24QOIXaC/TdjneXZ7EvFUn2RdZ9D5dDVz5/gc/33JNz1g9tQtn9jCyk2D66D9w9w1kmFlYNkBM
BEFObLaZPSIvxd0MTWHKwPSvwOj9t1N69t233S2eTxb9GUH36kor23LPwfDRbsm0jreWIZg4Mhtt
C9jIF5AZeGwnF8sW7Fz+q2Liqj4m8kquUlf8bRmI903gneq+fhs/XD/q/M7WpFey4YOvRY0EC9Ny
lNjiaBLQekgYEfjg4KM0re/sDLuhwBiTZnws6uHkcP7PcUo5RvCOCdbFC/t2nah0zt7UJwFefubr
i5hOvV2TyQ6FjdceiyuSEznyhjyKXse85TdGzx5WU96Y70g+ggNDK+k5mc/DBh82k0bzHnUM+I3+
vQLRGzUT8Vg5LBSTtou+d7FU6CXVE1JqDLP/iiX7i9w+s+jsXIAaR90S3bHBm7wVF+Oefun+msbu
rJMm071CrpBcK2JY1V6D6Kb2cXT4DflkCZ/T6lz99DGTC4Xj5cSp20ERmTXSkEYvZknJH+2jGel8
HRdQ5744CQLk+83EWeYsjhqIS+V18fbnKXVdj7YM/Xm3mUvpHR5e9PG5SZB55h48wqnyau8eE4Ec
T1qoolE4PGUCLgOtoxycFf8UhZLdYcrEZlkRRJC56CfnqsaQitBvRv+BUV0HnjtRUsMBCfHnrjJp
E0V42IkU7EelgOo+rZ8QcvZhCu0sGGUnAxAyAhNAlLkINdYvGLSH06QuIKenZpMsklzmCJUkCmEB
aLRUS3+uwNxTH+VzAH5rKj1UpRSafeO4Dzb4tQtXlT1snAtMDrCEDxotKJ8V/KUBLsXx5pQUqyu2
6VAp470RIJvC8o7paqMZoRrK+2tCp1g8UiKwVwUp7U0Mv7x9V7kS8b4rbgsSCHq3AQ9AMoWgtAhj
NLV+q9Ra6gnUDDCOuQ8eyu/yOcqk467vKgkJWeHdoiwH6gHWf/FhXSYKj7XtG3jxX/D4bppgXnYA
288AuyEOx9wnj/kKiiaKcZ5eXvBC65EkiUxwUVBuYioHGy1COofwUSvOdWsehfBQlnj9NhQcI4hn
k+pUzWy+tUFAm4wZ5xOG4GjsnxVL2dqkvx/5bDsvDOEj+pW8d4Ywo3SmHt06Pmmy/6HShqjLhojh
XD/9tah6VvuYw0gdIGSKYVBGzcWG7Noq2auAfkyAI7bHfqwS710N6mSEyOQUXiY9TngZK47ypL5z
CZlPX8W/dTXhRZmdUsMbrPmGhBql7b6bWU/6onvwqw0bjHgOMEqrG2v3eoNVszcP+waYsPnb0cah
8xJTjUsmcPLkxUTNgt1TFS1wQvZgiPKzmvOlnvOUUUUBIrsUOwZ9clWiu4B+HSR5w7lIXtIlK2U4
hI1QObWg9iECzOg7F3qLuHo1uBdJRe3IfXoLD6GmRd4Ie5fApUf6QTYTKX8OwiQrM2JiGyoyYW7X
O1ryumhZBJFmr7g8Ovf9OPdLw2/8xt90KMQ487jZHW43k7ITqTDjEYgsXHvRNdBBtk2DIFz0at1V
kfqwyiFyAKUjVLxNQdzXiohL1LlchlSOMwz1CCfZsBhJgJhmb+fVvEzFMsCsDgBR2K7LDz9E6N7r
XheWImTl5Mb+9uIyW4ReC6dQmk2imYxBZ5mSNtm/QSgERG7+IKc9o0ug4utC0u4Ozxs0gsbK6ny+
HLE8ZFhvRSlhvuYH0hDXAxhSinTJmX3H1EZuGKNiXL005BixESYNCii9bMor+qA/DdCKKu0Xgqse
EKz98V7pyJBXHQuo3cxdKHUxg1/QdE/MDZXXWC/Ra/sZZI1yviz1e/fl/tY/eJlNwDUCzeNULL32
GisGpZAN9t+fmtC0QbeY0+AggxJmbDSQaR+H83CQuq6uZdnuDRvo5Vzrsa9sGPTix4taBpW8zmsG
lzzzipK32akkbJfj8CctU4lidG+dRwawiOTLhEoIq6UYFiLWAxGqSOTKIWvPNUaqGKHWeQOEMN2e
CMW74/trd2CkZYc02YaeawD3nb83JajXGRe4zjNf2Ri/89DIDNEo0PQ4+SvXbzVjvF2AWn2urDEM
CKq7/mmzpBck9+MN2UEOpSHo6efiK0jao7SZxKjU+2bR1V8iiFwur4v7fA5qc2P5x4sC//RVxOWv
x18ws9soEI7NTfkQ+Q1Cwzsl+6njK8YVgGOm6ylZSsCvI/vrvh5o1QK1YZM8avbceFOsts+cYX7L
+MxDLkPEg3TvdFtzTj3RdfglwirxJxfiGKOF3Yoiu7YK0iO/ZFaugPm4jOe+bhov73RszDZs86QS
wJQIPR+2OTWoinnwwzCbwy8Kjslooej5RFRQbufXBHyyPx1i3yle1YnJif9GhW5oXFVKCG2znoEo
fhnt4uAuEaVo9WTF/JaWI1arR2oJKdV78nNV62zzJ7Rjz7wgyxyxOlY5q6snQn2UixEaOU2oRAiE
XTvMXZPSXywz+qido2peWJTrzdw9qz44cDnBdJsiTIRVY/R3e+m0vcOJWgrQiLxa4QzF14e/stzF
SMLq7kerGFKivOplWWtP1T0upZDRvB8hzbwV4GOVN9iop/zQsFnY3EcnR0D0fxwOKkAG6UBib2jP
pol1PhOYHxBd3MpDdyX1iDwWOteT0eqVsMnDXYTB8m41ZctjFu2FKJ35PMRBEqXNv/PdtHOMnA8O
XUYFEaygU0/iu0xDbqyDwlH0b86wiVzKgs/LTM4NJZpVQpVM3c+V10I9JXqazQsa53R+bC/IQDd9
+5NLtmUQ4IpEyb8bvNmv/AUDFTF9m+Q6Q6n61WgNoCe74FFSRanN/HIx5dcKRC5tmemSX7ulEpx/
ojzsLmmuTXqoR6cLSNr6D6S/U9Sf2r+2vLAv0oLPwB/OZykQ09xGDfuj6kuisPxbPNS9sy4ZT+Ux
uRgvjHwJ+q6/5kiAAEGmQt3E9xaezo6mIaECnnXHdma/SC5Fve/lB60MZa/rqmd/s8a13XU6kEip
3t9/JW2Jt9RBzRV6PJ32TxWKioDsmv2NbgQ95nhds+tV9l9GJfVsmDIicaonB44QWp1NRMfHmGm0
2KkAoCizJLDQuyrWb8tyde3Z4TJMWD6LTb0Cv4WeYmIKzgSAfIF9Er0XZAzJZaBYh7vCO40IR8oB
nHLnRNk7WyaolmGkp7VHyekPFGx2OXyTW5t4LvnF1zLg2tLkDgBM+mp2ltCxvNnrR58alu8w95lC
/My5r+w40sAd5R4GZRF+lJcFObf+u/oEHnzbCddwG63UgdKCe8Mwl+D/NjSEgyr1Q9BgA5xYYpVF
RKKpKK1ZnXonZMrvQNUgprz1yGjAy08s6JgdxGPUJtjnIJEktBQIbYm/Aw2eXQgbkZSl3V8epbMv
eG/j3SMDo6TVimbavxM751XDCBbObqZ9qYWHTTx7UHZN6ZFVdWwleWR/tYakFlcfsoLwnhHiNdkZ
cHZUdKH3ciNGNmasmY4q0WeAe6UhohFnnUwLRflFONOLN4sQ/J4igHTqGiR06Z7SxEqFlGw6aZha
Gw7fUrpl59YSis0MXEZ4n4DchdgQZ4WSJ7GI/76LUsW8gSrsbcvxMu8QAxDxsMM6hSaARkX25yVl
YC/piFhmT9JyNPjrTcf/0ygsWfPL33oNtQ6NjVZkGmGqWifQO2ZhRQ8BdeS2+uoIo02X9DRmdEHU
GC60XEKSGl3m5t1jpTz/fM7/R2TCDpWMCauX8yoWMAxR6SMEkqZqahEfhZQ1+v5pIAuvd1Pad6M0
hN8oOzpXpArASeM1L+c5sqwYRmDB5IjcGurM93RPtoxeFeCQzidbfdW07mbpuokyUTXOXlscYS7m
A1WnlYLSmW7jdaxist3HSTt4RaG1oGpp7MjolPDFgJOH6zR6RnGdSNPgDdpD4BTG8+5+ZEp2u0BH
2JZdg5nuIegUFy1oSi9vYcfyaS0tU4amd6BMyW0TtzW8h8cmmT4bczkfXsOm7vx7ma0Z3OC/8aOa
aPVe0ojv0TbOKdZySa6KcWuxcVKDQr9/9RXBjf9RHKgP9oWsrClmW/ugYIVnALevQ2Ip/MKSzogy
r2CHf2r9ikjyx3ETrbAMkQaaGgdFJQL61cw4Qx5h53RlIjDB6PTP0hkwro2tZxG3Feh8LXGGozW4
0bcAseECTuoUoUGxX1sryvXGIw1d5U9r+2tQgHYEmVcfMedH3EQ6nur2iymlQijYYmOIgApURy0q
1RrA3C8qaMCM4rSQSszzdJutQSk5c51ty12LF1qML4P/r+vJjQ0AdGi1Q6ie9lw3EE4CYalWnfmC
jYFI6yh+yiFWJP1ehgIy1yKPAnzRcf5tcJGL/UzZ+QLCoAwCtpeX8FljaU5zbK1UxFQqY3FssJsu
5T0GOAQEZiHD+xqO3CUtxo9CsbpGz7tMaj2bDZgnK30vdBjX41b99o8bgjbTkjmMpKyNkhMDOjiO
FQXC4Tj3tdUUpa3XXs14ROB8u59zCrBrY/FDKw0zoA+O0NvVw4j1ScY7PiDZclWXNwgFBhccEyeK
OtgPFCDeU5e7b73C8mvSS+1ZxAOHOIBl6M1cMsWuwLTjEZbCPPmCtfmvK1L72SI/KMY6wJL4cEIp
08+4mjNvPMr+gjsDb2kOxBrrSzr0gLVcBpp+VddXdXCaSr7mNf9HqQIC8+V6OpE2wknhtszUqNbR
uI6EKQdevnEPcijM8+M7oL7llE09wC6oqQYomjpjFycEvJG6CL/eM2iuakUM4luUx4cj+qUT6cKd
DoMeZYnQyuc/LvrqlK/XWsKiYEadlYIYGnm85dUpkCUFFempv4lcS/tNXJAzzIhZNinYQj3UP4TJ
/bO/PLUi+vbihInCDKx4Yoiwv05JlEwoHEmhKegrTxyn82R3wEY4DGyO3JFjHelXllmfwS/udd8h
9oy76yIvURYa6Wp2pf1QWoiw3FEkZcYWRNJPsadvdugEUEi7NkKrJrwY6xVt2qVVUAN5iDJEiVv0
CWV1+p3HznYi3xupIaOgYBE5zJqxe2cV/V0Tw0gAeMuPiyim/x2aMfnA8JD45xCX/kJUK8o3qnf5
tiSJSqmJkxdcnRMfqrx/7S0z0zg6qoYsgxzUSPzqa3KiT6iUr4De24P01ll95CA0YPL8cf7bDvLs
mIIE5GIowVbdLvTJM/Q2efglurEZnDahrh+aklGhenEoHuNzO/S9YvvI3llbR+C4gOPqodYyibBg
Hgah05UFrXk/kptt02j9HCL+5kM8p7VchDd5TBNndEyC/GA4uy9mW5MyPBjpTTIle0iskmctnlNI
uJHvxhlLmNKvIMCPrLjV60Hcm5zptYBNN+aV83mPcZlAmhWpznFEAHQqWLoda7JmMmMlWB4861SY
VBSnz9WgwKW/dObIJXUykAj9lrMH76TahUsriO5ojE469FWpBdhUZM1v8g73pvERJQxZiotUHnUK
7UR4cDpwmZHVqb83HZTS0zlIeIysd5JXdMUfYXUEFfcbFCCcTfnjbOyK/d0ZYsPc/QIk1l37fTg+
QIGWYR6E7EwXRVfHatj09IVR55tSCApRqYQ6eq7eY1OXLLEetzxsV2G0AfT68ErCkNmIKz9THKiy
dTlNVAtqWm5+uafyCKxAs8b7DfT4/5HPOPzoV+P3pfIPkqwJS3TIRToMWgYHbi87mMMSRV3zS1vj
V+mHDUnXUz3Ncz9UuM7/3Gojm22TgLPTKgSOTL/xjZE7jFe+Hh1noWnQAhDTYfEF4IxIlASQoEbY
zwWz8RwfC0A8u9ZsNt2U3lIF51bJFGa16NJVAPdcWwpGiZ/G2Lv/qSGlR3PVLW/sUGU4d0vInbF0
nsZxJv1tKxz/1lfxhN6+NzVr0rzQl6apbFBayJPQZZtH67UPcBSGH3DMCWS8IF8i8V0ZpBOv5HnD
SbfztFFOIdVbLd8r/OJ1AanpKyKH6jg/rWBfx9MKu5fP9az38lIZdVQXhf4t69j9Pr9AvmFwHQQC
6Owag/ajoudrsik9/9iO+PIcjKbD0CEKw8pasVm1qdjnYIrOYQGs7bY++hR1QWEyp8uG3+lA7+hQ
VYsuSpwEq/ttgcmzwtbPOPjGE0rhOB2Q8uuIbrBs9TGhDexiqKYNjFH6QQ1iMXgKlEr+J8e/rC1r
XwsE36axNsTlrV8zJhwuLYov1ORmHv4li+FqXDyD3z9ygi2DJQd9s+cCdEpIootdGWUR5bv53JBw
TQSca8Rs/DPaKG9gkhPcLzkd3ZM2hybpisfGFpB9Pqlahq8+UE2/EMwEKZEmvz6b6JD1R2PuwvEB
AA2ZvD7M3ICqvvNuRmf0aocIlrkNYvUvAdL44yhvETlT8fEJEAQJjkDPr+Y3G2KfCrfHOtOETNCt
ySkx6CCRxizSaaukMecIzNCkR/DTmDGdvIMh8iBXTJMtpc2EPuvX/3kJWiylhMaW02l0Nzjim+wD
lsHWsk4RkaPhWocqfVOVcJHGiNAeN2LHu3irfOU0X7M0yl7wU3vvb/C0Oqw18e93YMT7Y5nnD0vG
6uQvoMx25irtiYPLdzFmTytetgn9VA0d8PJz8kzfPqK3TDsCB26IqxfXKHpGTl79E2vpkx+x818I
kuoLq1cmB5dM4hY3yJBuFpccoiSCnEWMbXY4DrFxOFv9Q8QuDPUrX4BRw3BJoQhq6bToxyeqiY0q
lhF0+Mok5xuAJI9KzCglKrNj+C3jvxZHiUpN0zklus9ySaPmEoAQHnvAvN3a32bXRdP+bNCWF+c5
7npL7sIKvpse3biCZO1hG/ppBX9rH3bCXYfYBiIlbjq8azpNwlmWH99z7PIU90x+QHEGXkPUjy7c
Oy6C6X0/FeaFOVEReaN8ex4G88gZ1j6CxlfIy7BUxtxY5LopHyAstfwJBzLpFP4cu0QV99QCzDt1
yH1V3Rquuyn3NzMOA5y6fqcngcyGlvRjji4eYf2VZC4rZcAsAfzOppICbpq9nA09r8sG9naqG0hi
c1GGBvIp9EPi/wopRAZuINgnp8P1+h7umkjeXTWRplyEF1Cm6YjUpbRj9qBv11/4idt3LJwKC3tQ
LibVQ8RHYITRsA0LP0gtCC6KzwbqIX6g9FpikvsgD6s9Hfp1NQR2/aRExkrsQl2yXhUTCOgjPaVO
jerQaxnVCclB/UpxWHa1D3CBPokIPdEATQPghMbTMdV5wMsiwHQ5+r0vERA59FUIkGvL6Eb2ONE4
fSbSRrGkMOSv9LkijRdnAbUJBx2x4ogmEaYNzb4rpWwmwmltoYS4KuzsQnvDDJqco3MpgCkX63HF
604Nx9oiOK/fzE8aWtFACBS2o3WHrT4Rd0Gdse2E3JjrQH+O5qKCho1XVO5bDcgrnk7hNs1XTM1e
tfMp4Q7toIOXOMNPmwNVjRX3hTPSljO9XOginZYfr3ts8W81i09RESHBuddG3MJ60SWnRv8XCMwj
tL0jFVsaDi2uyRINj+0Nlxg3XmRqMpPALeWs0WUpPDXtxCq5VT4eyRDcAgi2BqyFumXOpyXCjFzf
oXmIjPdLIIcNAWYP/+O24apBTYswCzSy3c9T5dor2/BOwwsXIGznTheAnT/ACY99MedFL0nhpwGu
jSmyyko/7C70iXdpul19nu20buxKPMDosfDrozoqTMdr8P4OLH/s95f6pbLxs89tXqlmjqnoav1e
7SJqoIsyScih8r477RKzxIxlqc4GIWZmANOcFfvN8feXFnv0X/g7b6uqt9A4Shy57x1pa9x32aTL
gtzb7LyG7tAqNoOccbr0rO5d++AN7t9D6SJXZv+ecWAV8J9tbjTrWcDV+aiBe4/VU5ECokwyBiF8
cE9Jl6wW1AxYBJXf20v3qVLeolkP5ObO3+ERyhK2q1ewuc9RjO774K6Bm7e2FN6X15SL6fjsmBhd
Zkims2IwqLCUA4TVsx+hO3XjayW/A8iAS6mySMebdz/oN0uNwpGn5WbV7AHEH+N/GK0XZPkfSECe
lNGik+0ghoH9PuY71yjBEGut7XsIMV2OpFfcq3v7XzIhv+MMtmvLa/Kyc69HrkpFas8C6pmriCQR
yPxc593FxaCysijzYYerG49QPHZLiocwgkH/Lrir5/TJ3gun6rACIioHXUmusOct+sHWFoXt5zHn
VyLV063bKt1OIHhEy87XjDqAgVXP0SGyMgmZy2gxKFYzeGjC4ohqxyhp0h9ZzX63A9CsGQaHboOu
F7JKmIz92hi4/Zo+gDTzxpWW2twO1zsvDvMUATNwg8YpGhcnQjpFwNwwHOaoxuuA6GGqCEcmiO8B
ewvZ3p2KTG6q4hkfpkjmJMhixEeW55i2i78siPy0URmbu+p1swVh2DVmIe2BTDTjrihNlPZKbnSt
1otpIvjMGTCxnYoRk/lOb/GiviNMpyJzEBDJ1Pf+AG7TWbpgG4ODcva2REdxoTVZ/HlPR+fxyjbG
t0kEtmEdWtY17115xfNsjj/L833ISPZfM0quSJZeItTC3KF8ghLRi6Q+E4HXe42TzSHlF0h59im4
azQsBVIPbfPivxAnLEFYE8UEbsHvPLpHiv/r9kX2makT9PGPrIptSpMf9Gut5pZAZI1ZvQ+f+7tw
JBzsQwZdyST2HqjeDph99SoYq8q/nTkQ1Un9kBAGxStTI6LdHAUBpcz9s9HzULHe3b4TP0H7zebv
megUCpedXfDdiaZFG2orhzuKxvQNQCmJL0Qt6m0D3YnC4dh3V0qy3bmKxZ2qHzc5dZ/NXHD3kvEA
9X8iYBy9FPvxQTXLlFKuoI3QhWNRYYkQByfM3BZaVykTRmRH1zlubLAWnwvH1NW7bwRvmkU/2Lbg
losT2mH68OaS6SnDuTiBbjNtnHbufRynr7n/3DQ92irtYJEYqYTSFx+QB8F19uuuaNdZpzvC0Fm7
DhFJysP8bgQFZVFSXTVFnZESt68yL37BhZHA6wVGiBJx19oYnz21WYd3tv55ET+TolEYPPDUD0jN
iYy8vV5wN8DsuulM2UjOOe1cHxIDV1ZDkSZluHHv/SuK8Rdq2EI/flbWtBXLg/7LH2/cTdmaCT5A
goUjVoPyQxj89eMsnIMChdNLQ/8t5YzwZ81K6KhVycOcYifjBZNT4W21PRyXetIqGrWAPqUfkkH9
hZk+V5/zLNJHvRvbH5Xec7/ygPhsVwuP62/VvIOr+U9P86zIXZ/gTmyGcP0a0on9lmhnj4WBUrPe
pRkjqd1B/GZy17kwN5QMeCVi8MijwAETkwnzePQeg2GavcvPyJm0x628ArD32zSq01AasGumIvjP
r1BG9/rCFkdofcfqE364zUwe6po47JwDDrU/QO2CGDSyvDoMxqJPTYQmmImFWb53ghSLbH7151Tp
R/8Iu7Ya1r+TjPwPSBZjILkbzPaKI4VB76ta6D9m63hzUBiSHCwy6gomfbQsqcVM9P46K7QPWYBG
yiuJATzkDUJv39AqiVJD45LRzBubqsi1e1m9jbT9xjlVz74pyBQPZUfJtm7RV9oymYi+7halRBDh
9Os0+TddJWYTCvakC+jTqPGbgrjwaSZMbjmHoT1qBcQ05Sn9VfwKnWq/2NbP7i9j8ozuFW1T5SwY
migK67ZxrzH29Hs/7bkOL63IZUDUrizJlzVbgD/+ss6bwB2jmdUpn+1RE3beDH0TvmxbpPEe4W2w
Q69qvO2jdZclmC2Mk0mwsmwwWSmCL0puG6tU+ksmKfUJfZLHGMnRT1EV8ifA0E0W5R7Vgcpd9199
sMJpaaUTk0xSBwAr685aB5dzoxIHFvFq6qR1YyOGTwRu0fjKqIL+7gvJsGM0WvqDZ9JnYV+2kzW0
pw045jbxxRugUagOneBKO0dXyKkVSUff3MPzKA3xgeAzAlqYjxkrh9/euq4ijNoV+3aTLGHkQ/wB
OwW7HJyt0oQstejmVdI+JQEmvmuCy9vQicpKZ4FPmoFMy8MNi7WFtWITBc7SOHBJl3nu8YJPme56
9ydDCdPE+HxUABahq+oUP7Iu+c/c1K1LucNvr4D8Vf3U+G/B9ky95EFN4/9N34VLVCBe6dHmAzpD
dZwm/7UVz5X2bpo4jccyEfKXSTyUYuECMOKw5y8LYTrKPyN/58wJ160Ak/4UKmoeEmQvae+jLeL0
sh3I5VPhP3fRMIAhcC2DZkAtohuvJ1/ia5J/ejyv3mSuOE5jdRIvnrdkRN1x8vpGAJbpNJt8gcK6
FtwOTdx6yQLk8eKC021I+uF9mHXVmaEbqGCPd6dzxxxw1Tj9TMKT2ByDf0V+shjyHQFoCaqvyqz3
4rftLiBozSy3xQCz22/a8X1PRW9BY0d+W57fBqIZM05aBjB5b/ULPTdPu5RMbmE0LOVgsGr6i9Xb
VCPQZ1GG4WL0uJDg9eev+0hppYDcRiNl2QDVOyjizAjy1nbVHfOjRQeVNYuZHJNDVhK+prpRsTzQ
K+hZyqSGkem4M+bwhbCNeNlXRLGkGROMM2fZQ321ux9XrkPqcdXb++5CZvAtKdzfIfSEJWiXCzUg
m5wJU+Nh0HrTY2Sp98/zIns5AQYjcIPhpg9JJadwfh7H/NxfjDvOa5clAu/KJRuXbP1wnhG3I6mV
/QR31qiE28b+4CCHk3KWNvfHQT/NpB2wRywoQODWuutODzgl0Ut04ULkfMSGg2sRCRjw/BVta86w
5s9cHM9KUQomTcXZfX+zAUnJ4uEx9flATh418/mbEFgr+0FA5Mxx9D72XFHJ13ygQ7bk9u5Y3dNc
ZUmTlRWTfLgviyy3lx8KtBDJjuEDuGscBVxsHHp42PqqizuaOCecbB42cAoqJVI+jcuMJayJUjJn
SSRY3bb/UvkN7dnspRcyYYtSMND1H+TJvEUkmyOJvX/61mcAwN0Kr0ruqc8NvzWilr9y2w1PdHJs
NWvd+yxHTUABxNLvFOLV1RdhNJ+G3gLmJWBMpc0AV5vYxG62amn9oYgXm+L7aiUzAbJ7X3/UwaF0
S5VWBenctFw20TGZqGokazdr3amNNMVGP5XFZ73AqORT9jw2fQQIgSheCBCmo8kZAl3hquxpN9im
9Av89dj0gksNSbN4EuUAwOkg9v2bxB1I/krIO4B2volLIl3G3z5dKzCalgC5ThFcWx2fWvq3mYt6
1l69eW6IYTPgJLh1BrzwiZfxf4NSaTr2ULMOS+GqtlpjiCJFwwWNy1F640H0PYl/fqhHTKoWQvm6
jJpa/neB+Bw9FTrzUaSE6DIzC4ZLFp+UsY+Q6yetXv98KAbEvpeJg58WCxV1fHd3nRuX+4GH2Ia5
hsRKMy+W+TAjeTH90bicR+FHMP5xdYxBuLt8O4K3GbAfSstzof/ihqWoDPlKQ6tALgZA7bunoO5O
4cjNqtyCJHkjIdvq68ILCmh1P5TimaiEmvUUhftnxRE3jpPcrLKo0ooEDhMJuvPPg7LBqFtWPb+F
6WdlpKvADG/67THXWgx1tQCHL47uuJF8hdaKIw62H6xexslRPOWenhbXkQedQO6Fxz1JSceSHTJS
WEus7lEHvQsg5rSDdyk86/okFOZKnD7kqx94DlTmiaBWHxoJLxv449L58HwPwmGC1B5var5X+w6A
lKd+2kqkw9FZIzD7HH18361SNhlzS7vdbhIPqT78j2mKo4BRrc9BXTFo2Kl2nxeI9dPobHRgERTS
VBbGgw9JgaXnbFZElDntDZ0x6uicBjTAhAiaQjfbzIMZySS8GjDnJGiaiQTdbwJowigscdgijn7C
mzhMREVXvzMKAIfRsa9d9DGGcLQhyDM2NLLLpY4cdj5Ih0gQRZXknJ4VPu9SzT161Biay3V+YC72
92HHx4xnysm5lZYrEPDSRcd2yv8HW3LCgjDF4iaRnxOGKeDIrJz6rBWMADlTt2EU4rdrzvDab6h7
Sn+WPlP4YfQf3qmTSRE1wmSL5/cYM1fr+Yw5qVuPebl/10XV5jo771h6NcQlV5I4tPXCAN/GCOFE
ft7UAmak73XCxFNQ9Lc0lqlelwK9Tocxl/6Tv3dp6Z56FDphXhqt3Ssfn/YH4FuRbUhwJeL3ucFj
43sbk/59rZdxXlxAl84zUG7d2jrblslalrht5+u7hCGbYPfAT2WbZjh30hs+M+3R3hF670gSP+Iq
t5YLTwxLOoS1RtD/4cVddb8f+2ZDl2hV9qS3FoIKfUBijKlriwHovqsmlLGACLertuKyFoI7Wgxm
h7v11pmkMJWDD3rI2bRaZzSyZ3aJGRvUy2jEAiJYOve6vpNe+OI7K+pgXXKw1vA/EoOOs0SUR+Cd
C7h+SX5diNTLzxM0I47tfnhEHfGCTCk7xMeedgXT43G/Cbm2A8wwncEGGzfJeLctfp4QTDNqnhre
cMKCEXV2p65MJKQ7eH3njNfwu+41RJUQxglmG6H36uZzbksCxdCxBCW6ikp0YnWFGg1D8nRvJcwU
6ufIM1jKr9Uj/0BJRgydyr2fSU1p14RtpdChC7DxYrGDCVqLqtbweQSIRfwDOM/wrCuWg7qO/QMg
zX8cBWw0tkzihu3FqBQGaTIZ5lMyJgPgIIK+Muz3h+wALc/DJnhgZzEPNNBfydeTj9gfRu4rlDAQ
e3YzXy/acgvsL5BSB0BTMVkWMpY/DCfT2w4bTujSEuAKgSJieSSas33Y8TyePEYvfAIBK/EiO23h
tJ3Cnm4fl23w5PQ2ZqhRNIb2SCbYoo9vncIgPDNMZtb9QHjsQf5EhIUn5xEae7+QbKDD6WCD1lIo
ag+12kAoNiH0FrvIeZVAxyDC8waAj79PEC10LYekLjLg5BPP0CweewfVzmK4ONnEm26M+dAXHBRk
OQlKF4+tl8YU23V/FzwYEiEXfamY0+pUKL71JqJFJ8sE/XhFF0Q9viJaUms+mZpGldISQISFOcYL
SfWWWmSbX9p3GY+Vd3TrzPqSJhRCZjqIFuiQypRGGqMeeJYoKCWG97XqmAnfptT0BfkXxMNgxWY/
RCqWLJqMxHD7U1wrZOcynkESM+kCT1q5qX9lpt0OjoWBsQmmTq8taw6Pnfl8XJWRvcArXs7T8nbx
VUQ1n3j+9+/loTAoBzfQK4gOQ1fnrWm3jJ7VI/5oWiwAjxMewhjwDoD+67YIRhgNz1qZ6icQIFp7
cxGdqF682oU9NqEPEWykR7eU2Mg+KAA35Y6Sq7OUpK3rA5UfwRz1KSgmZaLdSUp7QbGdJjAB/3Sf
PY3TCqUI0F5KmGGFvctbqMn2M20uaGxmR4/f8/3lhBhsgyTxWtERFAsjBUKj8oqSBUMmO7QZ13f0
Bgwf6QgOZ7nXYKqc7A64Me6eF3qrH27iE6EGynl6k5XJ/TGXrmA8cy2PElmaSyoMQW+baWHPBC81
CTASENNtHyT2GJ2HJ+/eicfNh3IAxqEJevRVO97EQjBZA+/E4U3YXkrBNI7DuVJWeS5oEpYJdq8r
TB/oObwj0qAZ5gXWrjs58ddYtXu60dV0f9bAFFctKZm3+GuZmnRDZqjH7ohSMY1X/2vW28kykoxw
kmpS5Hcb4kjXAmi4ImqnSO053rn8sER+8l7YJykqFgeTXo1B0lOhByHOXpZTT2xVniUoh3bvxWw6
k9jDmaiGx/3rT930wF47bdqC3cK6be+A6n8afFqe6yaYwO4uK+nYdNVi+VO0nPnE7ZAUbYVQIS+3
YD4XbyQtl5ve13ivY2iUwLoX7Bru4Uu5hiAytyhQ/MQKBgJxeaaYq0JUOlCzW5KXXgzqV44TkUCO
f9046xkaXDW9igm1cWxIteD1SbqXyQU61fsh72QDLHolc0tYE4XuBonpXxaMQFnhhltgOTclcwam
LxMjtU1h7Qoga9dWbiPBX22qadQLqGeU8s5icbbG5iS10wZ60FO0rFQjnyu9G4yNbUgiuc1+tBEd
neRn7a3NGDQOvcf8RUoNFAZMFfem+1ON1Ex/X1EkqmaMJeklsXeJt0iMQhFgWwnyz61IRzSTYulN
Glm/sTS3jebL8nwQNAUc7ZGN5SIr3Jwm7Le2uWJAEJOtIFqFDM3jThCOy4lhn71AWCnS3pXEBF+d
6VJ/15ij9lR+B3ULiD2skRQpW7cuJAGiOz5TYOLvzI0/S2TeSEambF4/iiMm0k1pQ7IIAa/w4EMj
YxRKCyXodYdI8+H0LOZ3whWKOAnM2Ufz51IYB+wBdoyoKBClYkSU2FyiMn50RX6sX93A1iwKO9Ur
hVdYZE+/fi/ZvT8lmHi9ZE/NsxcikGuDX4NH0SPa/DACS2f+f/alInsk1g+OCmcNH8zEvkTCilEu
k/o34ogBDea95TIDg8O1o3+u/NmcKgqKEed9aluBLWIS3Ljll32dozpRVwVb7+MKDP/ICx+lC+1n
FLp+TQkyjkGrazhYewe6n7RuWpksPTFenfjeUPO3gqgmtgeKO5pmRw4t3upiRvLznv9A8thFmHm4
e1eMPj8U1XPCqlh9vb2RH+Hokhj8VDHQqNgivl+U0jypl1iD0wINSJCg/QuGkFBjj+LUGZSqnh2G
w7O9Vnw+5qcKI28BoPiHk0fbdIQgT4uWex3x2SY+SfCp115IB5+lbgIuJuxrQ7S3Uw8jRSkaR1b2
k21MgUYqeIcncf8rYdsGpob4HH3aUQQH+vM0IvFywMbIO0jNcVTRV22kFo50tp4xefVwm7JOU49i
OSm4y35ufPvVTiJNGGTUc/DgXgeTZqRiO+c4edEPGGyFchy42Rg3ISCd+QRtgHVNo1S7eurpy5n3
P2cuJIN2DqdUT5OT/WcvjLe4ue95MZMlJr2ASR0AcE80GUrmHO4Vd1LIfx3JmuchbgyM+uMVFt/V
dqeYh4h/dXxPt/4+xFCuDHCgrg7tHeyMvWE1D1n+uv1DPv/zPfyPMbZfh/dQcwuc1vCqRQzKMPa2
a1IHagf6+c0ZCDSDVAoO7XUnu/geDnvF/HfkFgdD3CjOcDWf+K30uNrm6YRvTsnmkygryTj5BVUh
2gX860CgHBg9ZlF+kp2HQS8caQcQ5vZ+Hj2/y96qzJ6x6bDbEw1FFCx5nfwZo5BbdyoHFZjLN9AW
PTul4wnq5X7tZUcORqNqZsWyNFfFMeaWjr8/GWez91pf2QspxHdwFWjWVOFn1z0z5bUxy7xZ7/kl
iW+Js4adtnMhwF98j0NzRmo+faLsMUQruuBOfsuuLMUTSv4/YK9OcWCtG2tUoYdwjPVz6Qw5eKl1
LUcg7T4ecLq1FRCFHL3gN4AbQgyWwR1yyo0/0G8e6nKYAZa+TRPK+aVBSyJZm5hST+y1UHBt0IIi
kf5SZOTacaldLGQbpcuFSNJp5kTYEVyqUx7qUDy32CPKTjs7adrmwH7YpLQEeJ5mZ6NKNHzznqx5
UCEAGzBvnboTjXWgtOzJjdX2hqHWdd+3XrRGIrSQ+LssupMXZQOMAt23uvXS4eO6RFuaM34dnyya
djo2uzqt/MHxebqqPp8hiIHEEpCT4BNk2EAa9k5+29KbPmBCXfFW6jbZl64qoAgTHabTg3cgV7Ke
QCriNnzGMVb+ovpMUCnsAjD2FV0trwMS+6a1dTHYVZNdqX8Cx/yw+U9yp5fGDZ5poWJdEwRSqqup
fB+hkdlbp7bQY6mGsI1n9R+BNrcoxjXj+sWTdWsV2M/qCJSSvc76nZMN+RGfCNzRvQVzJz5hOf7L
g8Y5Te19B+a8zVYY3K7o/Gab+sT4xU/jU8K+Kk6f8f99d13wuY4BGd3EdsVhAZx/yGoSw4IJQny6
fmWl9PS57eGftXop2hNKCZhxBenDKzVsXHjFxpEuUP4l4f6Bn3qNvg8xnVPoOdeeFMaVZnOettLz
TlzZOG2iuHV+OnC262vtRPDfQMp+0lCM37icLWISgrJSWYHDAgr1TVbrrLfuh8R+Ht3v0u/FnO9N
VfBq7xT14cQOgVX2/ZfRn+H/buKE6LoHiBvCKBsCUzdRPdpWvuCzbfnR9f7dR5KAUYh7P3/UoYeY
NEt0tZ4nEfNHd+2p93PNE9v9reXxn12B0HbSFbZN5g6Tu8k1cnZ63c0p1WQxdwqj6jtlFsObrsmD
/qalbO2ruoE+dLNxBDdQmJPgbuG7XDIGUqiOAdmkoecqdZzp9y77OdZIXploFQLj0PLJNR0V3m+D
16EiA4vA6h6QB+I/oU33igMaDSMm7zTx8iJIp7bIe2ov9RqG0Y42qsoUzAw8oupdbIIg+ujP1B7Z
JpuglD7yEoxlDM12/xRejXQSmdLvefU1JESKOnwGqMDqEJB4i9xrJnFr7ihyOluELLWipAQQLS89
jBXu/+ImPREksGeEVsnPX0JdMTjKWUn+LyNjztx7VaLA4jgNkUTxzbb2Ptsxqdau0Cl/gWF40Xzd
d+7PilyD+Iy/EkkajkoG+Y9r7MK0yQpAoyUYquWY0wfllt+fdYgE++pVz8xSitHt3gIH2C1EGCHw
S1yRsSIWd9ekOOwk2NZpYEIKaPVcpB25kOk/MX4dH917q4lfF5hMp7RyCptzzCshHP24zPm3tcQN
yuI2gUM1pzwMqHoWzQuOuOXul5NBrlwzRNI6uYjReTtGN/IipZssMBO+QwohQX+gkP1ggmTgf6Dk
YbAnpRh06LwjTmAlTuFPiTBwiDjKSiOsx8O9ehNnECA8KPHOXmXMKqbt8Vn6ke7loIfpxRrDF4aJ
6R1J6n/mKbJ+5TOcEEdqIqDIc/hLUFojaOiA53nBRJmG0HD39haXQz0ZxFpDY1yrU+I7ohrqaUCw
akaD0uS9Bnh8fGJnlkqgi2Kzyw3zI5xra4beIHx7VRzNWNwxBlDrzGCytwSEq+FRzNuuierLmLpF
br4aUm2AFCK/4adxagT6H8YysGE7Mo5VM4bpm1/hKQOrdDrCcn9LpTvNHNYOmaviBSTOiyvKB3cQ
Og4t4atkaIlZvQgsRr6UoKVEM7Aqb59laqAVW3Oe+V2tOKkgnvAEi70nBUH1k5008Laeh/vi+AbR
LOCSe/8bMDAJdj2O7QPi6yf6PC+ZJp22gOWpfaasNfilV7V4knxxkCWRx1LvQdpwMD3XpgA32qJZ
R0iS+sQDglbw1gosFtpkKI5RA6WzSgGatAkRNglX44eSwff4+SdJSvLGwXStp17kT5lYSQ521Nzv
u47YaoYEoJnTVVvAcVZJOIbpm5f7mkGGDqE72qBlkh70JRjhh3ADuiq/SqaZoN7XYIVfntEAanv+
HY3L3MNQVo9hP1aucWPgCl7rZalazjYKVwyKVMGsq4HiLGZSGG2VRflJXugFJATh1SwjNn/CYzL+
FY0c7aKCYsaVE7WCKUByalY2Vkmb1dcvpdnyz25aJtwdfBSF5zviFc0xYX8IQYtxfiJ5LljPYFlI
4mmiWNr6JKv3El7//x/p/zRJtz1LD4T0DUpIeBWi6s3cCM1CjnnUdt+WZLfOUdU3po/o5UgL3no9
nhvE7JZM2m9oqLDinJVd7UgoCbbp9YNfY3G+BottBAN3LEUtoeUn2E+64WBLVR+clY66ApQa0qmx
DiXIUHNDy2f+HyTI/X1a0Il+iIfL3oQu8fLcMWSlKDbV1kk+RlyCsOM1X8ZSt8dWGg7Erwa7hvIy
2XhBIga2QYuowEHV17/QvPYyTgFFUNGdXbfjkbIPMiChFUqYBfShYr7FW/KheOJixLBlAraRtYKG
Q5EoY2VdYb5BWlbRV3AE6s56MM+7p4nn1nEvGxiQ5V6KHA36ncvom7TMg7CwCOh1trtDINWlXNBA
TdTFZ4kByaZvR5SBAwZ3B4xTygxVoNGHyY/VVxzxyMQ93l9zJPLjRHZ+E+qR7JObjgE1V0JehjTC
dyN0093nNlqU/T0RX9T1YlJAM9mgeAQbMP/XfsEtd+pUqvAhm8bRRm9tqSAHNZJ6Q0s4q5Ja46l9
x2ylXNp8EbIt6lkMbT/QBpBZvYTEyzY9MwPEUX5/ToLzXx0ivNhNT15Dw0JeAO4sn1jANzNjgP19
qP75tkwnEZJYvrxfNR4EsLr/18XZOXEw4/tItfkBId7s4qO9NVdOKrIcaxzYBuxoJHC4Tbfjg0rd
W4qR4ITOwzI+IMFPHucsOcpudruJJB8CntTWsZ73UyEXiXDe/sRB9LChv/kr3Bh9XikbogPpVLG+
wrTjv+7gOUIP8bYEWJ+884cg5W/NtzsAjUe+v/ZTUrkkeU2e8RKDpVSmzk7c1tWx5U5qK67sE/QJ
pBxGAb/Vs1L3gdsL/k2QhQ/+nkyrP6JqnjQqpJoYVHZnirETm5H+m40KYyzxq7H0nTQ7SQG9zHiV
VXQLVeNJQbAfOGWaIshR6yAzfpGNUmtocpS36/LnJ2I+RCVV8iT+D5b/5naLZoFmC2qx2G2ys96N
YLkZj4+w7G+MuwbzddxddNtOtWCicXJ7sk1ItAijRJBZsgQp7bxSwcDdOBPKJZfYkdB0rjcrTBQd
cV+AHrGmOM1KuBmk1ipaodmZs3k/YKAeYX2eK/+ZhZSZClA7FbOJLLNTrlY7lxg9po2/dWWwtSC2
hrE9lvZMYt9nlUGUD5mFjL7vCy4P1vKyyisBBVq/2Fxp52No3LCCGNk+ZYDD8RiOV4IFJjYlMB5p
N6m2wZaWJWBFfxUBjD8iejRUZtbDDpK3QIz4Eu51KT2JIz1oI9mAYzn3vwQ9w46D1Y/2N11n5+Fn
i9oyMd/2oW2QyUVNCory/qbrpNXjdFGFb2dr1VYnLU4DHHVW9LWOAmQ42CZi5BKDWBRsBpZMbZiz
0UJjEOIYdylM7w0sHtPRdV2n3wtPlYrSxCPI5+90L1BUEqd93o5wwrMKSxZ5xDdaut28nJji+zD1
Ff45Jz/6RXdjExzl3wcYe74Rjp0IOJyZ+2SOxjWtIbYprRVcJjTYVCrHJ3M1WKXgOsGx9fXuG/sd
WXHhAS4VZIf3K6viRMJHSJuLwN8wpnOi/oz6q4aRO4yv+HhLR5TC0qEJYF87HWjLvE6amBkGXQ90
OHpVic2DkW6hwY6aIWNuN/r6Qdkb3QAQaSIIY+F2mtCt1BM5vxvUDCI1OuFWHOGtXOX7JtuDndVg
O6N5JrMdMjboVK1DG0SIoR2wIc7WelekmWQrLWF/3ALfHLw+iWH++cA9oToj4afytNcDoQyvooUM
8XKuDfBuMzDdtvjy0me6XOaETFxZEsthMwJRHzWzU61ql0ecmSppbfZJCt6CElSXTzQCiPSUhRBs
1OuwNMbauiNmbGaxa2ACokPaNok2NlAd3fpLCugjopVi2qJ4yXVumABSC3MN7CFOXFb6QK1vVlNE
oxbQHiApTlEbVWMaiQO2fuS3jr2KEF//y5IZYxtDdPS+3fw7iamDTptoqrdTUB0QCf/sRRFC+3nB
TxZGYAB674LhydkMqBToRRkaPSZU+erxUmxXwuKaUH85aDmaDhECufc0Ij3OZFx5N4yfZ0tfDWd4
MCITuVHhVIId3EWNyM9OxUtnBkEBY4loNPWrBLFrX6L8yrdqtbHkHsLEKudZJf+welmiqVxMD3E2
9HrpPINUNy9cmZFlQsUtNeiFXQV3uSClEoGvO+Tzu0bqAckINajdW76P+HAF/rzZNIbX4VJbufWQ
ljDBRYVB2jlgbyYzxmyfgljoPTAGIHHWBb2pi0hOzQdX3ltSETHWSXVnpx4dwDu/0OPq8BIDB2R6
9VB3vwAZ703a5j5ARrV9caM3jbEl4mvZgUoQ+fo+tAB5PH3Reksn1V9A4jD2SdzqT/zf6NZlwh1c
v/RQX+nlLA+2nXE0uL03nnCBEVCy5ZrFQz4YRJcWbSPTikIKbdmSzfMYcH2LYKh3oxViawIQLotm
/zHzsBQhrooLI2V8RpqFSS1nskjhgQgc/8UmDVG38pHSayBAe66yCcbolceUrb6ZECMey/4IRZJI
liZQl/7JgumuMFjcVfRyrCha/CyhQvBay7gQB480AdFvOeZlllT1PSbxxOEKu7lAUz33bNcQU9L6
ZcXbfezKRMwRIuHWbhh4zS85MCowVVgZT840nP4zlHZC7NMLcOKtLFH1t5jy5TK49MgYlT/OEPkB
xBNv5NlSMmZomGc8mR1h9bgpIXzpfSFqHPVOkQGo8qwsqgWV4/2JROZ/vF8qwt/eglzYsTZhrM8G
3gX4t4nwr2oLylM6AgljiRh35cFYRTJmpc1QbbtCOyuYdU9xyxwkvdgcpRLQdKbKF9bZUdf1o4KS
f21FKZCAXdPbWL3VFaUq62uLZIy0Og3HOs+JDns2ZBfGxiZEwk4eEvVrvRKu5BYZkC7imtPEppnT
cTPkMWcToimX1ySIEUPrLjKTYN6w42HmInUthStPT0MbPZkI8nZXY/e8W5zgPF8yZ0gM4Glsa8XC
llEq6hS9UtVxdpW0PiKGbQdIy8Kmq9UdSPMljSbI5aw2MMoRAObeRUwGoK9ykG7OxLPZ8nuhmgtX
95wnYb9aR/d5UbX1D2lqUrn1VTJKbBDyRiGXK/ao0QPL5ly2ijMIfZgdiJf75FyYW9AiiVEt+TwR
M5ockihUIDfyJxyAFUGnFT4pjjhYSyihrDWo4MvY8IWLaVaQOpngIW4Cs60/2f7H66VtfLfBNLWa
wJ1Gp4ssGYPgNuGr8JVhF4y67ujYBqFmXNOXGLaaK/JilHkp6onp9fBZj2XqAT68WDLus3h+yy6y
Xtkfmp5c8cOSL+JzIaO//Z33z/gHk+gvvKad2CkNxqjFTpyImvPUOzQDJqUpTk/WPMYZBDKzfBAr
AGtAU8+hUQGH1GT5e5lhoZUjZ3lZ4QXUDGt9/Ugpyz/3gEz7XjNd9CYlkQLqnT5N3Uxxn7xfsa5s
+93eJxGPOkBDcbjqOrec5Rcqk4Nmg6duTvcKu/vO8f80L+AutyBSSjppBwEPUxhAaYodfxLEVi/4
EnrejymZ6TtJxGLsxAWim8HBxkAAoiEKkix9rU+EgdyRv0WC5h+f801D3macmPqyVeI9FmzNCCJp
QrA6gYmh7QM8DD+9Ewik7p+ShWASQ1BfYq1+qurqCW4vGwD2aQNo1n7sBB7j7m6vqLM+r74e/6tb
1IWjC7EYzWLRhsTQveMg4eDwZq/dmbXTeRISEzJVzakMg6ZJdl85gVTt7z6eTauqHazEZGjUWvPN
x90WxwLm24yMa6AsH5DfRb1NZYOGt4IKpDYlbiTQps9sOuOGG1Hu5eWo3I5wGGYOmrovNwkZc9Sj
tLS1UPl6FcvvR/iUyBNW94D86RvCctNBw+kFNfUK55IWChIN4FMnpghKiWIffxUNOjInFhipDU+N
sR89Hoq4eHfliaE+00h+kIlCbpDMePbgoyFuGo6pJ3HDIVd03URslSQAiNyWVyGR+Iu4U04DnhNp
/X0DKBlTY0tW2q02azX8BPfGM9PF/MsmTZiJgZ6IiYGfJVkGvIoI5A1YWFIMsOxyP9IOEFkKAlwP
71Gvb7BAm1GZ5Okb0mbLRcBu6uVrWwkZABHduHKvFW9g7t4FpG9mjMtKJj+y2tcv2fTE2BzDv5E9
EV49XXc21iLoPFdJ9dS9QCqgUq/cIM3Lru6gaWRmEuHiRQnlJIlCQp1P0jtJIlERZ+h5x++Y1aeQ
ShBVi3Ze82b/29ASQMvDennW2u4HAMD8v+HGVZzz7xhj5SiUQdXYOBwPGwJNz2ca1CCoVhFoshfm
nbW5M3KKYPJch74VeL2chunZv7SLAKTA0djWdVlA5VjBnOtY7ncf+fxLVVOzt1PikYfFzb1hdXL7
DqxT2eHXgf8v6Fe3yMab8Q2D5zuVJYCdMxYq9TZ7WZ0UC7zfLlQZQQaTEzjyutAlMUzic2YX2rAm
XNV3Vp3vNvMjgchi/agI7RJBffpBFTgokQqWjI2gc8s+K0Djzdt5+9hi4/ljEPBfeKXf+e+c981+
yBYvXL0oZ6KTwXPbdJPv1rOtLAP6MlXjJSCWD71rekBUEj9eFiCBH7LEIyZ59YaLnnBnp6OhAbc4
DkhS8Dvu3IGDLR6rp3jgr9sqi9zIgjsfZcYAivEgmmpNzDwB14ycmfO6BhpPgXi58cpi7sjLSGhB
VwZfF/FcDkqkrCLUgW0st+N3K9dKXRcsAKmy4My5HQ1Sx9sdXZQmu8DLS7HeFZh3IhpI8wMG6i5Q
YDn2yHQ7L7BTv7+43sCDQnzeo2rHayK9LBruNeo60uYn2xNrALWZ7jI6QcF9tMkSgly79TKnjNev
4+GMs14e2YVys+dUPHctUqFdJfQ1mKjNfRRPq/CsWfdCX7mqqRTDctyv5WO7oni2hfmjHnO3L7I6
nMzhMUv3HJW+/hHhUZmRFBrZg3mtAwu2BtCkzM8L0K0Qp2OFQpZ8rXSw0BY73Yy7q4w/HqQHsg0t
4oiHM3XBbc3l0a0Ckkuz4rx+U7y4idHAPqb0oJfAGXgKqb4AAlXB0dtY5QrEpzHaJ3GqiSA7Mu5m
Gecxh8BJ/P1g0ovcAmw+N8TUKapCg48VUo7k5tr+J9LBRskR1bXqUXlXLiKo8SICru7H2B258/zf
MayInscG/Z4xmea//X0cEWAwVTJalaJKt9yNZ6nkYkSQbFpn31t3qmdjBYFLsP8Pa5VmDOn44HkN
z/9ppFDqUV26dwIfKrbaI0vFLx7qkwIzIj/BMDyDPxJMEYsibB+onOajgS5n6sAyzOpkw3H/rWfy
S0HKI527HVAdIDh3cbrCh2jBAMOgrsOmD6YFZgElKl+JRVteRTmRdwTF6tfn0Zwh1c2wDfE6+I1I
+0Ld9lTC3LDijvUvAXGMgugUJLOITRo08EBunbvm7VwVzwZTBfe6cYqTMCiTG2+zJhr9H4Hc5ytM
etyn02b0+QJAyyQ1oa9x01SDIa7cjf6t8OUHf7lTFxhfStNczpj2Lrr4Y1ulQPasfssnunRzBvbr
KeDbYBNxD8nbHfabqwGJCDsrtU+CKT7c5nL1I/SxuHeIO5/TpOU40lQHbTSsWsiaBueSBNTTu9bl
WLH706D+oe1e49SV7bPytqa+1y5ogWR6YWPwHO7NS9pbGDBJZ/u9peV7lE5SY3EdQT7VeFOvpwUI
1TnPKU4WWlmH6Boyzs3pRpZC2LtOsyojVRZw0QOYx1PU7ZazB4AAhsonr3+GQo52P41J7R6CLqLX
FjJ1Z0P2Gzdfyj/C1r8LMnDFt+vWvNgGXIxFmAgQNhP8bR5rNV8HhXsV1PoLgauoIdHpjAadq1Hx
K4fR0W0gHBDP1Lz3KMdhl++7L2md+XcQopXMPl/2Z+gQi9m4EjzSheGpjNOdn5K/LrzOfN4e+8/2
Hb6J/M82PaGWKaJo0gekkLMbMOiNw0tgeRmLOz9wIMhuhpdpgiEe18UolKYK4Mkf7Tpf7yoZBAN4
M9bujOSYWJ9GPvmcE9ofemZrB7NlI2UfTHQBahaeYBDUZR4BJ32LiT6awkUMmr35Fbhf4QT+JD19
eZVFETlRyPciswz+xWBZy5nIrW35GjdUjeR9RKMQWgRvSjx9Fw+IMhLXqBJseiwUWxPVwCYB0DOs
VvezRSk7/XN0oHK6u7RMWJIb3H6yqj9Bd9Nfa6LmI4jaqWbitWxbpAkRzuY7l9WbSGtcr6pNWJH6
cRlf+lv2TCa0GCHlE7Sm0xDNvkEHGYfNy+938ySBL/D7AkE0w+fG2rerIJlGEvH+ksvGWOeAwxsm
nYjzg4GkSEp55cIvJ4q8ajcPkCr8QoDE0OYpfgponACvuVdLzl3KIPmfc34NGC8z/bzEYIZFXd3n
HSFYyiSFvw+CxEkUXbeMriqkhnBKP4NrUsK8Y6f0ln2TG+JqG1YppQLx77BoeCQWWObMRXXFCUZS
9IcmAEPlcV7l3GC6z4Qo1tEi7F3RP6wwzfZh7vp9x49TYNyjh45NUgMmPuyl36wycTN6mdMdkpsH
tT1kmho2yRMvMR0xoB/fqSfrGjfjDs6/CloOYnPY+PXEwxfU1pPbrN8TYSrjrdEzuQI6A2TTwonc
QODl9qJ1AUo9XRkdCLfpCT+BVbr9YnRE51Ky5R/CfysYBAIE7I3ZEFbeHX9AtgUdUXSrm2g5wkbl
NSnVaXwuTtwJVoeThauhHGMrBKrPd6I4xPcE9WA9UTQSZVaq+vZ422xNqsygoM3gMziFtGVgf+yq
W+pcbqJQ84fgwducUgyNMgXnLb8AQIzj87+N7yK6/Hrbn5MfkraqwGrPNZi2QB2UZZeLFu/WU39Z
xdgNQwBa2tQCERcY/033S1Lp2iP5l9KPOzo+iG37rq4EZss+cIzon0LYrxVsnnXOtRcomOstkf/W
u95EaycA0jjJ5qBjnKiXnOMQh4JBXOlb4R+rVbnztZPtyqlfhW7+fIn7y0dpUsJxjRAXRTteOtv/
eBpbWf1lDxCfhfylHQjY+j8/qyveil2ae82Tsnvoe2KRJja4/npY0f4GrVgSeJqc7he1WoKIvCsT
BfS5Rk2Bwn4p81/VV6BObv0Zc0RBB3DqWPFoAeunNCszmt57WxQGDb/vLpc5VDiVLfvac9RR+4vE
Xt+AiePAoVc5aSNO3WcC8/w5WQlIjntyh/XQSpzqALIuZ9JujHn+8X/tV2a1XAeqcPOIWqNcYEQ5
1DbSfge2owL/jTIHzxTndOaQZ/oXxn0U1YYoFxdwDhVZPvlfIVdA2x8PtLi+Jd5odO0OahLpNcb7
ZMS+Sfq80kHWJbJjJo5GPd+aqgK5mtb0WCdRXEwoK5Gl9yumEarE0y6Plky8KeYNQm08AiQfCMRB
zvg9MAni7g8SSAQeBnj1JP7NMvpoigQWouhjb0m3geVct2HW8CJMUuRtA//ohFQvrRKoywSk7upI
Rk2LUevbK6Vc2SQnYfWKgxfMWovLZyzKV3OQH19wgIOTxSqbu9K37RhsgiX5h2xN0YeXZQN7c12j
vKQt3N7cuyx845pEm6Iars6FlXPco0TfCYjwI8Q4PSlP0J25g+zuBBRm6S8sX0CF2q/GIiqbgQGa
9CewhO/Q02fCmrTjE+nJDXwuosmWV3yF7l0r1VdRjatoRif0tj3mnVEMZhTdZlGBrGtTw8hnDYCi
TOKZgfyMXtEhuiQqcHvuIJByxDhPXnMWsILDztdzLtI8GRNT05Gd0VTsnJzW99ONzZPy6r6NedVD
NPWvh/rK77BWnBDEwcOAoP/cSKyPIGpTo9a14LysydXMDoiUHJDa0Xm7hvc02xBg+1O6ZkeilxCJ
y7uEnjh3reGowoAolroTSWQ4QELhXefCZJK7uC5k+rXqbPInCRC6hMc2jnckET8xfkVFuK29Z0sl
GzVG+E1XVsaMhbKAk8bbPo4bcxx3/vd15HXCW5Mkg5I6t6iYZ0rAk+edOCW18mXtOMfTi3jI6k/b
t4g5obB1UgIdp+z9CV6h6WSs7S0O2QwlZR7DopQmBRfQeQnrhYdT78Ddd00d6uf6YQEd5s33+ZlL
IZF+x2aAEH1skxa+pAwdZSOqViPy4zecqtUT92bCEfE991GF+2ZElfm8WDExAUJ7ZzLkcpwtxguZ
zFiw9VXEBXANrOGMS2rVZAAZ24YvcXsDR02NqZrv8JZgPDzHDxsVqNS3b9sxiiMGomXXSrt98Mnt
XiXvIQR8ti45XDFZe2B4UgPdPly7CZTaI6oBkU+aKKUpiYnVqKTGX2Cc2DO0/2ZZQn4q8kFh50XX
vpIF7IVW4LdsuGOIGX6qTW+Jib7ERq4IAmb9qNFE9zds5D0A8ZEYBRw0KbITqkyyl+qj1OeMKmzt
BYVv5LwDRQcvgaf762Eij/KpXE5+HJ/SHzBBwAghVKBNWhN3N4sDUX7JoJhnx2Phn8V2QWp34XDj
xWi6oEOiGxhN23Vn8KY2JKw/+PAFUAE+rKKY/xF+IJ4tByDTvWw1WV98zqmsEnSRbI9lTSRKiNPx
AriMzobqBEs6Sedz3UfVFJ5C+ask2GwhCMWTnS2s7hA3B3sK62eRP3lc0QIo0jfqSmC4SDApffho
J6RTRqssizsVAdAId4bVd0S8u0wZPGwr+muF0jL2qInGcIjzko3pf34V/ODTkHHW2JxmLiAtjfBc
zr11TMdFiXtOgJ7zmiMgehtKQTFpPMWqUQtENCZtBe++xDBsXf6p9WatRMrAQyiGAfK0MEnj2H4p
CvFj6k5un8w2Iv99EMtPhcr56XR1yTFnRrncxkj0GKxC6Bf/CxMYK+bzEOg/RTSoM/JXRTHNDjPE
X7cPBax0ofaOq8WBsF6lc+MXn7coEDr1cPjkLc8219j7zxHlkncYVQnSzZ0Jj30ADdzwJJPElmLR
uHIzD5RtqcoaOhZhRYWNUAtm9ZduK3Ww2tcCKm8J9Iy3wafyu//Pp+VEdVQjGHgRuYQRQYEztDAm
heJrNBltPXnvXveZJtxmXuWRDg1Iwd7uZmTli8/HKsHQZvfnLUxqtJIvwJQpVpIuU7/Vfph7zRTI
hkz54MRq1+2Af13dn6ZQKkCqNZ1B/O7FnO0brLbzgzrQrIF9AlRWW+xYjplGb6ef4LXMU5tE4lTh
aq8cM+k9aC5txVjivaQy+XH035xBT13M9kWpEPKJFCyR1cUaG5kI82/0roNjzrU/ndoKeAIQWrny
hoMdcv2+RO0MnLxrgyVsdWEjtZbjvvPevNPugmA9CLN9pZBcEsrNj/UD+iSHyYp3fNV7hnWgSxsi
DlQBkwGliWfdXqUjrriz0btwIM2lGsdE0mzdXNwbQsSpjWUMzDD3roLnlHaiwgFFUze/EZHZbi6K
R43XNLkYpKI4du/GCjKyOAu/qvUZEOIpEgmwV/duc6HOkzk8NcCZkcpB7cWARTmqb3jcKNucfvVB
Ngl0knfqH8297Z7wep2oCrKuj683VE6VnDfowTPGLLlpCZrUhZoq2mm+U/kFRS83Sye7N/TBGKow
Mc9i0xusb1b2JNL2MEhpFCYekA2iWLtQvspaIMW3ENLSoeRc3sCBAo4CI//dgRtIAEtUsSnVRHfb
4lGeQp+U2spRTj63ZClCM3r29lUIYGVwdJwLOGoFRurECvYcENtf2YaeWUbvakrGb6loRhEg+Rof
G0g13wdlANJk9ON5+jk8w3iEzIYcjN0/3uS2M6j/mskoa9bGM8VOTov5sib+gWH9L8PrPapaiZLY
SZRrX9DhmYzs/QFhumJbLuk3QCJN5WRXp8Y0pFMD3fsbBx/hKoHGyzkFkLt6jhJHDjndJGO1HN9w
DK2xJV14W2pmCXa78v4b1hHrL72paHAnG/jpw8F8r1WSASbCd5C0tDq7wUTOWMn/LTM52ZPQ/r2Z
84Hn1lp7N6Dkuz8TCpn2IN2Do0vYNJ0GdeuGExjk1yJWzZlS/2VdFRr3AiHLmoXZHNSTFbUej5Ah
jwFPMRQWe5ap36/jvxvH9wBokoEId6enziMnnba8zyaoduEexR1fbEuxfi2Up+bf9xO6Agr8suy+
7n6Qd4pToe8ETV8GrAg9d+JW+cGxau06aQgPySBpTpaKL7Y06N7+50B7kZHDjvjaHRhhmmhJ1mQR
O96Q16eaWdL/i32fzVSPHIm/V4+WuV6ZW27+evcbt6ALtrgiV84xyJjfPXz2lxwWSIpB6xrPIxdV
i0maV7Y8FxS4kCSfIiVp18qvB5i5GjncT+SOg08mW4w0C2b4BreR7coj+TwF+0b+dSKkk/ZQeaEr
6yD6Zw/K35XStjCrGG17hzGujfnuZofklGaT0ATm4XeCF1toAkeCaGbMMbHy4tCk/RGv3nmzgg3f
EyzYzlJjpqXxowW+5/kbZazqlEInuWk1ZKx7UBvbjJaygpuH09YDRfYvAuaF+cX9UbjEZpDyE7MQ
wqyefM0R2C1RFs3ImxxEHaQYO9KUBSTAX5ximKjUo5hqCeSpFb7/ca+eVmMLZu3HV6xODv9y1Ruw
DEg8j45CfA/28ynZDkBUrT140VfQIM3C1oyS0XQHlM6ehwImNVAO0V2UWoEGscu+jQyySXeAR8vq
PSPC+CDWuCNLbTBfr0pucE9ZpEzu1fZXLyOHpciCXHx8oJd6BWINxKp90FMdWuAV3iMJzvpadnAz
E17u4hIBXVWxZQOaI1zq01g6UJW3TEGNu36CSYAOeWUxJcHZ1EMwbxel+4u8pfgcmP20LmlLnLtI
NaB+sUlmyHtOozWgQlGqDDxRn2azUjyTPjT18EqamYeQSjbTxpStblU8FtGKxH9VDABG3MjCFgBt
5HC5JEZA8d8zI0lxrMmpV8/v6+zS1YWX6AA+4tLourfhPtKGuzdSxtDNxOeDbzHcu63nPODaUaqQ
BB3Ntr6gBaL5zD8ZE9BzXRkLuUi0GTkc45wf0FVWhuT+KfwHpkjaEGY5rQGj27IZT6hWCxFnOIG6
GpkrmKHLfFaoJbkR47GvnwjHNHoYhB4nheYKmmYXI9EoU8wGKgAVtuhBb0r2I/Fol9qkg4EZ56GC
ceC7kXRJeqclj0v2zOUMfen/z4Uy0DcuxV7wn8/89uBvD9UY6AeMTtrh5yptcz3buY5UCVdEPZu3
46DwmrkgoLbAzTQAmYPaPup21ckztZpGRuuGAZ+hypAPbHj5m88TeArP806ZblyNmi9GlsjNAsVg
zOabpTdQWsxPuaej8L4okezk+jdHd5x0/MmsmJ0w8+tztRkN6DIvybgaSn7Jh28bQVsRM0JyO0Dq
PcFfISQB0G3do3Vl79T3f4JNLho9HzeAQwvx8YHUQr+K2k/h0hIcTopB2mcHBTGVXqStUWQpw+68
ZxcE/Jr6lMlCXFDwlafnjx3xzeuNXABFF0DhLrhaay6v76WnCbhBrOVjANv6rtwEHlOqzMyEHAp0
DYVP4LLJp05XULcbPqWAzH3U2Vzhc9ER9tHVk9xmUYjgRrlb+I7IDfWUc0mTNN9hR/SelqToPIwz
TrYwzR9c7cCZ4Ga5lqRkRFsj7UfRlsE63Jv89Ln2l6U27QmUGatGl9ybG0lzu64K9XKkISs7d0ra
TuVNUqxiAb4aLjtKMvng/s4YgNVreNWIkm4fa8/3ywCBzDze+E6CixrCBxeX9pkjwCxyMM6yrL8/
uZXesHeqqs1UK17cq3p51bqTl71hYa1P+cEH/YyoxXccjzTBfWbTBuO2vzziYNUUJjdwLRxyNH6p
p3gPDdFqXaaE2uZ5SCXmUkfFHQGXlqz9ErW3ohXsOcBI5Uy+riN3N7ADkH7vyqJb9ZWCpn0ZY3Rm
A8Uo7Byi+hozl7zmkyrRn4CKDvI/Yjg90LmtTZv/u6ZwsVdnrkdRFO40Ykb4uXOBArmjfJl8RefT
v+K1V0NEPmJU7pSob/6JqKZS8v0cTqhRsAOtO92y7cTbJVbxUNrc3I95UxATKSSMDbl7YXChGGRP
Muipb3PXOXclX8kOKMpBIFefDEmj6VLIpQ8pOluj9CwhJWN/iu/p0b9pUZwfmcLFJYVomp1+1LS3
2a8w7BGOKYEtrpzRLwu00D1elb9WULE5fwHdiltqDqNaZC25UFjtBdaBxClOGDnbO3mI4ymiMM23
SabX3qfpekERWGVCXivF7P3e3bYNX7/Cr/2G0g+BgckkhTCV/udgp3ULw53dXaFEm5dKZWS+rS7q
oO92D9eYFhw9N/8aH/MvPYoa+VBm7DlxJ7KQHuo0bobwLA2OmYnBZIiCAP8OS/aOqcEYnCtbNe+h
Xu81SU7dTdCKDaZyFhQqnKCO4O6T2aSzcZ8Ec3BHh8Rt3kCT11C0RCSR43uz6fMafh1X31ujuPkW
jpolB3iKNfL+gcmFfjkPotERytGRcxR7LvioHMOs/tyaOCC14Am2UDOuBbArCmEMa5uhEAleL/fI
Be7C3Nlmb6JnIkmAvf74BOwhbljg3wooo6xhajpBJ0y/msHvGNkyqxOQBX2MrjjiXc/lWQfo84JE
CMRpBF32ph5Py62sN3ksG2Jcxompd0+6+41BTofMMTj9OYi87qoq0p4p65Ie9z8/6AISo1/iXjz5
avcDQj2gxJQ7spLZaIMO8oLCvXp1Wc7k/MJpnJqPsSH6IkSCPLdh74sdMUo3dfV69ZsMP0bMDsG1
JnjTxvpcd3g5u5ftj0IGoNdime23ITn3/X2j9o1Pcoj2RaCnkJyzK4MinVAgfYczuo95/cqGMdRY
8onkCZMUOyX1ax9NDYhQXlcx22GLZcOmViXrHSzCuzxpJ3GS9IEdZks/Hv+69iOGY0MEDuL437os
MT3RsPEBQK+GOxuPIFSCPLm3gN39ak1bGeAO165uPy/I7XWjb70gS8+ZwjAghkVpu3Q91EzHu6yT
nysDqioXHu470DEXaBiJLCR8SDN9QaxMLnZkUzCUW/fJ2K5oZtrAIdyG8GxAbFSfbSY7DAiAfBSH
y9asNIo8K9hFFT5+zV4a8ch2fHfvwI9JVmYo0fwuw4BacVdnaH9W6jbzhqE6boPiH1HLNuwyo2iD
+qSBPnVxJJZzva7P1hCVWeZGLI1Is0xxxLuDP2RDZ0C9f76NRdqWEtt9zInTaBMSOeEiXC2Tjg7H
jluFDipx0/1OCQoO3vhf2rruowDm49qMkWEiH3vXktwzU9Eh3ilHBmwXAloEjAmwwt4IhFUuW7Bn
fdqxyvWqp8a4WO2z1Rs8ub5odXwByGeE27+WysoEV1G0L6nzPkFkaJgFaLB35xylKvd5AQhwPVBT
NkcX3P6UH9cEN91LGWiDW7SdB0kF0V3c0/JJYeigPPlpFZE4+mNYdJQpepnJNW4NC6ql8m446CI+
sfKkGSiSgpCC4Sehw99GSfNHCRXLJLptSvgLq/4NJZ3g9J4MrximVfqPB04AD0IY+89CMdM6T7Ex
XMgGTjDxFgw4RjMs2npnPEBw0YJ1mnRHpz+hD0sv0aCN0XbiTXH3pFSN8cqi7jafPZ2JavbqzPSw
fj7r9cDq0luuXfpWHqTTvOWPs+yccu19jy8oFrDIVdTXec7xexzmajXuBjTKG7fED8f7/q0iGBH6
Or+ngXHENhhC82I3rcy9d/pTMjMQIwktiAbiPAP14XxHqwpeWoD+P0qjMjxw241offHQblqiaHnN
F0mRtwRWKoUTw7P50rssuDGFbCjiFNGrXPOUHoWMv+ihc32UB2xMD6Lpc9QF1r4k9i33gQeLxwJk
ltGb/bh/5mvwNooPm5Iwyc0KpFKSgq2NnuXM6OSNakiIQXucXyJGcHjUlP4mEJ6YIzPXNPO+3r2A
qXpfESRBoVW82OR77pcw8yiso8u2pS2yRCqIZC3Pz6HDigxSDKlv5VxYm+aF6Dz9qa4ZnErUuhJZ
rCo2iTsGQh/2ZVCLpBVq0W9gLq8kcmwztXm9jDdguI6J48btgsNj08//nsNJFM2sBMmXBILuKnyW
QLl9rzacC/ETugamW5NoLQOOHR7uaKRM2OiQmRvfJnOnRJByqjluWAsca+PpndZuwcBN5h4tz5rH
ABtn7RSwtGZcivo0Kv7riIeKZYZJFY884F4qWJ2h1/rvo2tw9pdbR8WVV1jSftOJonVM6hmrkQ/u
+L3ABmxr8Kc9x6tOUg9E0GHcY8ZNj2A1HY/wD0BQwLrYeW8Ar9xHWlTgw7aDcPV3lDcEzonVATWc
x+N+3laWABDO29O/pe5fdMZvKugZgewumyDiRmkQTZuc8MeJNkTYwIV66sY0QwlNncfFBRLkgfJx
XG/YqSFVIelyXbf3LDjCsF7+JZe/Mnim+bdWTeXx/aHfuzEvBUsqNv+aD5owbkjocG+Qt9feDPh/
D/tvUVqJByK6EyW72+nBf+zOrLu91kHC9cPcu25IfuxFezYOqWmY1XLUEwFhAsF5HZGHnRaA3wy/
jvfvsuzdGXNIOUsyCwm1SSw7oMlEIDNJmH9XVvPPDMRz51IQEHliNpTZPRRIDSm0gQtVNpsBS20y
7ATrHA6TBGOGuO3PYaYq+bqlM7KX8CIkYwJUjBxdhvG9I5C/waJAv3M1qcfeIS/ZOkawkELmxdbj
dFmz5vSIHmxNZC9CDi1hcBJMls7YRv/1K4o121zeYl7o7LW2JgKPeYUdxmKj3xHD22J0zzl8bi1X
oWSCfONRRT5tAasTi156HInPppnwj/dHkXobACrK/BOwmVgT7VcsXiOKGmSCxPLmwmrM1bbXRIBQ
tF8IvY4z8tM9GsJ6fQ5cSrFArin6IIhpkQCvYNhlmCJoy8IsjQReVvozyPPpLv63R2lpU30pcKkE
puYQds/MavMTWe0C2VLb7BiuB3HN6xOYBGJR0UdtJxy0sHPA/dWw+Kk3pW8KrFNs4HLMs75nLYBA
hy25vrDVeYZK1bljueFK+p7SfNyhnSiQRC05KqfhDuiBchKEJ+0aV9Li+l8omRCs/tANUaYTF2NA
6mHFHv3MdR/k8uPYxbl5eNsl0PZv7x3EeMAufL4w85m67E46ZFKVxBqjZInhGkwdhiRVO6JBdwd2
Czqk8gCgjl/UJu8RIj0it3TG/3Oy4RiUi3K5EZ3XkJ3DlwhyRD1pHZMWrStbviV77lx+OMhhmX3t
y2/RLfg4YSNuhqpQBdFvlRwypn7mIOm+V4jVZhMFD8q9Rfbr8wKBB0uQJbcf3Vj3iCVCLHxuDxEQ
hMq+iG0ELvkkr0TXIhm2V3haSdeifD9MnE8EagsfxUKrXQ5Ma/ZTgLl8XU4Ke/5Bzq0x/D7M2QI3
0fOwHr0ZlskCzWepgSFN/fgkLXxs4LWtY/54UnsaczBCUTkcddUTXmmsocrlN3xNiBaA1unJ64vE
LAUbDssxfU5ilR+e+BjVG5IYppqCUt5eQnP3F7K/3/YzjvChBT7Y8hqtD4ZMa0Ftdi6BdfKkmnIO
kuUI3mh1FYOxp+p8zXDrxN6Z4nuuDB4tmh/ZIkYhrSqW2mVGxV+nIAav/n9Fwaf/0X9n+t+SCteT
wZzh0qqudEllVKZM5WtiuiJ7qhY8XkijpjF8kSznn1dP4/+TmhkGfstOBkBsHbkWN2L8g9zBWGT2
ixh/27+o91ClPodrqkxyT0xek6DSAxQ+xe2VLi7OAV9BHEkU6uryjnWLaS6faWbkuI/kiaIR2TMX
rBdxb4CPfoISTObNDqaQ1Q7+aBdZDEV9QPF5AudJZ6uyW3WWF/1TyJtEaUo07PpaWUUewv+EPwHo
gq1FHm2m7eigYYF2STpzEqxIKmfmX6DCFp8ARFIpetEBtc1p5AKWOD/Mus2rIngRjLyPWe2EeR9x
/8wltM3KfUwMQN6vTa52fBaEja+dvM+IkVjEGnRhdZ8MLxbOUYcZf3dyvl6PDYparcITXR5+CVkG
JHM9216TZqwbhw7kn7FJO9kO3Xp8yjVjIDl+v++lbiYjel6PdeapfZyE+tF5v8NDIiBrNs0iQkUj
REXmQy9s/hV/DpdFKV16QuHu1BT1No208tjvmalilXPrxpulugOKD+0XEKEwdxLM/yd7Kehta9s7
B0qhXMAFCeE7uFkxbF/iG1JFTFWjfhbcus1Lf7SSY3JslXGd9LPF9Z4a7a7J5AEP1nq76hGRISXd
d05xdEKKYr5OimqfZjuilRMy2QL8IkOhV2gTbNdHwF9amschw4pIxF0TKWWUc4DylO76oMoqDU4h
XaM9Wkky72MVaxWy0rla93nHkbmriHjTMIiyY7kzoszKn36X5mVWwtd7kA0CjA0Tjl8T2x6XwnE5
+zetvvvTYL+/roK8Qy0zSkju8wj/majdSZaEfZSBL5ZU7YgEb/3usJjW+dTLA1DQfTryaLkUSCaS
rGkn8EzALk1slObtjJWa00XD15X+7RtARx0oHS5Ay2My/sZu+XbXJOJjE/NGcDfuN93R8Zv3ctxA
JM8aC3amUWkFLyDs7YaRGEL8B0plDIfJEo2Jr8Yx9aF8+aUCv4ixoRQNRV6tdmPGD531641y2Idr
oWyI/gjd/GK65VWWhCmiF5vroMiCuXY50jjXtPvbqWmyT/NDSIX559pIeAIyFM89z1uPmpu3ZYHh
QsN2B/hZtxxRsOO213kBjsVIGNkHZUZooXTCUkyWA7ujtEs/EcurdrWLfa3JsthduJehq5ERtmpS
GjGOTJNyLBtBtEuteYNK87UqGhR3C+1P9IZOWMYCGRk1CK79Dpn63oL0eI4E7Iuvt65ge7BJAH3T
UgcHOfhkKrEpMNOAR7whotz7+qAFckfRx2WSLHcy/syW2psYMWoPoMFzoU7pINjwM4sYV0+7lQqR
x5ZxeeyicgChl+u5XheFmtMMDPlEJvdjxtHEKTVlcfJ6agi4n1h40i0BDHdYg2Uqbn18a1oQmZsH
AkZKvv6dynaZK+E6thwInoeNDYwkJD2vVGoh2wpeIU1W6Lmpa8VKZl8eIFIHqhKXFRJ1eMrY+PM/
UAyXlmU47f9Q7uSgGvj81SfzUFbxOTMiSH9xno7hNZLN0i2x/B+ORXZehAijUe2qFIm8nAlyI1wy
OIP9nQd6dcYuXeG4+QgVsRezTNfsZtQ+nnE9DKwdtLdUqNE4gDk7AV6WP5bWnPvlJG4SWAAE2B2d
gmZgLNpNLje35Uf2ZdtsGVcu5tK5wyb/BQRv6/NiWzXGuT/X0R0CDtESwI/1inXJyUBeflw8uHzz
Ly/Jwey9MZV+PuBVquIM9ocsd/BmkBuVbY2eomNXjpHj014gBAtzok2F/iAmUfC7AfiB4gUVrw83
2cj4Kd+6Fif8WsnZ01nKB62s5UPSl7lZvg8XzuXCKsxuOHb8Pn5K2bcYUfvFhVThWxl9hkb8ndOJ
DurVcHeKlOMSkNosTAqPL3err7uGexQWhadZzwbrqGrITgswit7FfZV+rOtqceKNFkPZsugRpovy
FO2JVz0hBqB3PddQYXPv5ac9Ka5oU29YN5GAk7HADmWMA5+YJJsU4yQGnzCcdPJTuzrAWl8dBcQy
zIfRD3mmiw464UxThaK7TTh2DkXLmm4eRcfakVTjGFy+x5ZgvIf+JGvrQWSaVpG3dxPF3iOpU8d/
2JuXCV9P9h3h8BwwDkH8K0W7HPlI4UJZC6x0j9F6RSMGdVZf1ei8O9hQ26Z2u6o2cRyTecHTciyj
x+Wfdw8DgazFukUvXkFlTpkWDIPS0aSuK0oZArzbLx7FNKXxpGSOkSDARBhSWH5WCr0NPNsAvzjg
ftXNSadf+iPJmy7zz6Xp+aLpVsRJqAD5JQzsOCA0xTZa0J3a+ysgBtPq2biHm/YmB9bwOkwwTlpU
ptSB4Ktt18Qjk+e+3dnRYZK6TIF+6yXtarq8ijK5SW82ZJYCWU78IWIcOYJL13PlwuZrGZcDCi9x
yQVmLNY32lQmahRPJYNSze8NIw/9muqpr87uOWUl4qj26pI4JiiKhHW9nhLbcFYce2e1tUevgBPL
zEJoHhCF2xjljwOr4guSMZ7mkiBficmziCy+qXK36z3tNCaEiWrPtzSzA8cJqNEX6nEKwtyLQbjC
jiFlOLDVf+NinuXFpL++6IBo+A1QXw2FKhbpQyCM2QyI186BLAWbNn0LkxfB+qdq5SHfGiyHVLK6
QgsObPD75RXbTOjFCTMscRUvFBy55aE4ymH3GzTlTF0KNX0iDeD7RWo/IQdziM9pB7nQLrdXI8/I
pyUpY6vu9zJ6r58ukdO3GdB7enYscJ3DRiKqUIrMtV+Tm4sZ8l18RnWCrhpkm39rLpqMOSnwizEd
fgCkXAeQ+CW/giba8JJ5q9W28dnEhSUGDDn0GmNcoY+FaVfacAtulZkTUF2nlc0opyDPZgqED+7+
SgH8sMkoANQ3L7YuANa633Z3Pa6NZbnawMbpUGDlrH/YMmYOHhyP1D/GUVVaLkdKRb9SlKsc8WwM
HDet4VOk3LZH45kQDU/eYKp46vlSuyrAZb6bqCsFjIYJ5WfvLYlVznm7cDdzYx69RBBA8G0YPlrv
GBwWAESoSUXRjmh4XyWj+K9mfUVSKjpW0W3q8xAkotAX0ameum7fhYVwl691hfM3hc6SHIBfi7nJ
LeTx86XkoppMTw6p8I7/7sziK2mzP3VHufGCgdoA8pcEwMKPCrm9LxiWUw1PEz6NAaYFJ0EBnTOJ
5SA71+0of69HHghDPxJpdLWcHbF5LLWDkKfVsFc4jqjqM6aW+QCLvCRFtkEdVNUFl+DcWOPOvRsP
CQySa+08Aw/4HVObXrU5W+wfikaC2yAgZ2DUDHLC3K2BtV9nvoDhyekX7G1x0izYhujeLBTNOQq/
1wZWCV829D+K7lTuNObGnRdEV4/hJ1FLuqX3z1UnOOYaunanKc48fSPWy0bzvrYrBj/XSZ0rw+lb
GmeO4O6cs8N+E2gQS2ZJyAkSiAqdRxSmtG2Z7nWRsqKDMndnVCNpi7VzcaZGstesr09ioEpQVnfF
Jn6Zcaqb2GVFtbxH/VLKjexfzM7nkwAnwq1ETdoYaMbjEFt94WjgVmyAd/+hr5iTRULeBjnLOWKt
wSmaYHI/P4gYinYfTOxygVTItE0ZvZIvcGz/lkDkezWLwdZaMMJ9qLUah65WqPD84i5SumraOjLU
mCV1qAtWQdQorq1uafvPtLB53EguWqEbbE8zYcJh5cHETaceRd36IYGwCYrMhuMWeUpUw7KLKxBp
rILF8cvkL+txVyFoijHJMh7+GKCc2BiTlOwFGZdO4VQ3RkDWaoSFjbZe4Dn8R6T4rhNZN2XWWdX5
nu2oRP6Yv9bWnLRpub9UUDnw3TSdoptuLr33PQENhfVKRRQZBOc4dBAsBtM3cvkEt0Ag0K/VLfJo
nhSDVhMxFaRlszxc+a4/7RwtlOAor9qV4VzRnVt9auzL9EaLdygE2qhO+R7YpzkY/CwQ8ifdbOaJ
62Lda9YEsL3h9Cw6Ir52Eip7LJvoJaDDpjrgqEs8eHIZM3/UEXVkMyJQ8CXgC1YpXYx4CyLfIKZG
B9cap3bVNYR4V3CGgGmPkbT3fZI0u1atoXHz+Fl+c53zEnePRvQyu1z8Rra+ToBxiiWZMJzJ1Cuf
tUCuuDmhHX3SLpZyianwc7Xr4cK0KrErv1Jki/JfyFKpJuanXFme7i36bI9MSh+KlCisQuBz9yib
18nVp/8/E+io00Jsa/N3ANr0L6M8u4k65kQIPOhqtoRWPj5O6tzn7mIGAanznpA4ZJnXE4+t/Psc
70kq45IuJjO8dYgothejsYWKF/C+7CetMzYPoHGIR69P2Szk5yw0LZRm6yNEqA4SNkgKDIKZPn2g
jCYuMRb4stLZrYLOi9aIKVjDhMkSIsgXzUfl7iiBw6Wo8KIQGfnyCeibfu03l1cEY/L3I9BH2/o3
60iuFKG6tQQFk+rho76ncPrkic3BqmEW4pWI9jwG/kevfrudAtP5GNYuXpZyycHJ6tsdXan5XjI7
drR6HESGL6ejCktfFAFW+TCaPP3D9k9xJopUzwYkwYi7uG9OyfFfaMFTxSud1mDdEtspoed4PnnO
IRgRZ/NfDdf37BVchc999b8sK7fclJ016CQkiVMEuyzt739saHrkrJt5I8AmOXE89c3ZjE4ozbgy
ouMIHN+ajsYB02Eu6DSe06bY3x8Knc3Z/EhPl5elkqmdTZpUhbOKndHGh+aqRxsjczNijB1pQk7s
fnlt9H4SoTox7Q/D0Y5D2yXVQKmzZvlI1SEoNn8AFICIk3k5nOX50geschbVBoSK4e5zFo0NDH4h
jdxlT6qBzWcW+Zs0QS7jDvQxmIRJ2JEjlY7pN/GyA6/CuilxQnRjxsQ3IC5rwFeVr8uYGJd9w5wl
UtsaUtsQfexs4gctg4SAkN93pkADF8xesF4x2MCzCexZbJOtGWT91p1SBMpUUIaTN9hGDDH12svF
jkDr3iJR9NQiVXwe10DC71whBf1KpAgrjCEInUuk/941uyEdHUo0TL2s4r6IbY+qQRlS4bCu8J9W
j07LvZtNvFrvQTvyXz6pwZ+CJN372GFeehFQecC4t3h6nKYwfZmGBLUmCCeyAa1dxC3t+3OTXWko
Y28Lhu2Ci/7EGHHGMemocCNlP4u/KA6qFFB2G+X1YRIZv7Pw4bWAFvnQ6xvoYBisCb5sUs/UtHqN
K1p9haUslV7dAbN6s6iC1d4cbjTd0+3aFHqrLryK9sf1ZLzaIQcA38Mu5F0m3ztyKOs5pGd97/aO
HLGs373DDeWcChbKpwNd4f/mtXv5SP803nyJGZueYcxMyrNV+kOn7NrOTValu7zT10aXToCKClPI
nfm8PkDwYoULpHElTmpKKDMAbiRs6JSfMFOWXudza0xt9d5AbRNugQ9LmG82mTTxLy4erbZfABgb
UdMKCYdHw0kGfgL2DzDo2qvoSo/4Q41PUDaZj0vdIHpLAu/Y/rXSqOED5jy+/iuaXaUWNbkr9JsU
Yj1rufihFwoBpkbDXtBlQfpqHkkJYs6eQCcyz3h3lDprUnaWpbtUrSQZFKA948fNKw8a+uHrOu4e
zOm2vuIamxegSwpfynHaWTeOTrpA1EbP79w+Uy/8y+SFbqSt94LArOTckrIabpsDXnKwu4jbPmE1
O1AqYY/wE9C/p22+AlNEkYPN7nlJr1it4BaP9dVZXFe0+uy5TfgTQuK7HzToAuiBx4F9zxFr0VYt
ccR03ns82wpbBkbZrQaH9uaQK9Xp5+pbxOE4+ocgeGmHmb+zFDp6t+a1G7E9NrbtfngjP0pDNlJ+
64apK5I6Cu4/dkZbLDxp2MoD3v2NrX3UHGqj9kRD/Ek/hRtfUjhzq7bgnns/Dw2SW0tIBdF6KCe0
RA0ljXm3tIiMSG8TRtQ6X8YkZF27V/gOMStCo+uPmbS6epMk+tNl9Y/czAjXuhp+tKtpHz28Qwav
NvAffnKagU3RwdzvMA6HrIWyJ3kl+r1djHNeHoPMXcZ7ZL2Z6X6fOXWwyXMv0pk2tZjfLBRVlXUO
C2/34Dq22MDZf1maOOOO6hxrcbU3qX4cV/MArKmbqoDQJqtwFYSaKoKgeQHc2pRTXpimWtUMeKe/
ZPXlVyhIR8komuDKPpcmpHWJnnjFS7SHW1k+d1BuBbCyGa12mJV4pfnlZVPXnoOznm659uiT/Blu
d0R70naEYzmXkO9SmWUKeWJLGyb/4LUEH8ColNsNzbrIi8cHmDhNuD/DOgf2wSJXyAvFEsn72xhW
YGq6GNr0gGqm3eyLr8WCqTJ/Mbd58mpZReROSj4IX673ybFlmjBu9K8jMIrAEos2c2neMOt6FQRk
nH/Nl7OzSr6cYmLK3Xyp98Trze2NACiMt9kVoIjYejj1h8dm5XCfsMvEiEc+XK5tUVNvUU9SxQr1
G2vKCEiQKdmHgUAY3w4Z3D/8CCSGvdt4Zx7/ZVAhL8PQKxdSdUoJWh3iOHOsU8XeIZARjSpVvRPS
EQtO7gsy6OIF0BdPXyzwM8BDNuGgvvqRrnY8Ux6H9Gd4L5JSjBgjhU4fb4khegVwGDTQYtEL3P6x
eF/RiyTB0Iz1yjGVBlGQh0U+vPYTXQQwhnKslo5EZeZHE2aQwDICqCZ+oHOk/sPPHmDxKcOHUXPh
dLjN2d1i8HNNfK/2jRPyQ4b5UCg1RlFEszzsVCL5wbdYRZsQTH9feifm3yY2MW3CL0Rq+BqPPVPy
zF0V96VAfro3fcOHYu2lJ6E5aarJaSuAErd3crhoksfuocXspbN5m1uA7UX2iOWrB0G62dNJCo8y
GsH9ZpLVnXZ5XQQ/1/BJyB9Fy0EBRXISg91/hH4m12R3PKfEfEsLMOgWBT7Sz8kd5KACQaygeSrU
1khDTp8URKE252yDJaJa5Z8pvOCKcGM49rDruvlc4ZWaWf/P2XPCGy89kc5wWuaD7O+YWGyQbXoM
kunuqKK1ihPpQEcFaq7i9YPNMW38yLc2iIAMpiiwNxrQ3jlGJMRg5g7+vUle5I95j9tHaOKa5bqo
h5J1CW4DBhCmginLfmeww5QMRSc7iGmREvJPCqBW0cRjdFA+2p7EFMTunGHb+U16zuvpfpIfaEqj
y+f7iiWrBB8mHn/QvDYJHwnMhzMs0j2BqBDo+NxdALx1WzF3n2gPJVuIC/ZunR8TqpUHjLReuQ/k
7+eepsVjBk3arPMOtmd5sT02ItsHcY11JPZW5tq6X2Bjbt/ECfNbee99t+C5KGe2pjuXavOe7Z8S
P/KuK0WfaclffKtJDU5hgmPPlZl1bHqvvmnmSYE81xgdZONv8YBzN5jv9v0z757p5Sal363cZ+fU
b0hePWb994jN9YJl8afbmy871MqWy1WocwkSrEdsRBpgtkyPT8TDlUbchFf/HheoCi3K/WG9+tZX
YTcGKA0UxdknJeVf9lzI6m+rwgq9ypY1jurhSoYLm8tyfBgHQT5ZGLmWGUsEGE0oArCAfmOHDErM
CKhBFmcEoPjL+jkozBiqFAS+j+FM1ffH2Mty2XAKdjZ2HD6YgsMrHbnd4GEBzlR17Lvo3uFkJzOh
+sZuRZZZzLUCHoH4m+02PmLcsCJIx1MfkvSQ155+7PwXCKXo1vTZLy7YM0xMYC4YYzTgsPknP3pr
busBUU6URz2aHOvAWYcMLpfEOC5YNBk6rLt4kthQ1Ovsu63vBRlnbrfpnoNZrjBmE6ktsWWk/z/d
y7Ga1E2tH8EUQqUNoqfbj5jEk6mqAuNuJtUWCsl76/v3ZxpyxGiUcL3Q/IqgGTltiQlPuLX+J32C
kTg+GYh7v37fjv8gmqdjvK7ySx5LO5Bp68bNNejqr8bDXyGVz80dAHt/jxGft1yJyTH5mtu79edp
+mCKNhYZnKzZwkSUYkQILoOykCaNwxiqrjgL27mfdhq4gWCPN7tpbcUA7J1e302BFpuspcwL9jd9
eZcQgw/6kPNR7uVr2TnMoRVUhE2wZ4xV15+q8RQRBg3vfERu6FNLvXIs3/YzEjXcb5RF4nISTeE2
JnFyHjm4GVl6uw9M7MweBZnxSVFkiKIvl0bLC5IA/KGU88paAf7EQjN29pJrvo0bmghmgktYhWkb
eDWdVHI//EmlqFYH7acmVsyTrZlxIgxwkr4Q8sweNnLMD6nvNoSAyFO3oLR+z0n5qgZTpqMHX2gf
0lQo+Su6u+TPqKckMDXa0n0ZP1z3oWxD+40AqSP+CMr7nccrKeoneoNXVRddYS9cRLvAorvAosLa
Jw0EBZmmGRQPDRZu45jbRyZuNX/8aDl0bNUP8QcklS5M1HjwwE7tkzUZbdBxXSriwkTwuFFSBeOK
93IVc0Zd+FbiUqcKrKkuXME36xJNgGbhIgLA1/YWeDXjTMfRfZLWw1+W+AF/J2lBqiBEaFCCAuAb
CRr5z2u8pha37/Bjewb1z2bj0rMY7NG4dDuJI75Evc9vUZQ4RMkAx3HNV/+7MTKOxVFhNww1K2MR
3VeiytS0VosozbskkuvJ+9nGYGXSJDQyBJHa6htqD9nHVVGmqOHcF3vb1V9ElXgNwQ0aQgVVBjcD
IYBxlzX9Oi1MBaekpUiVQtKXuHPdhr2bqJpXvUOUHfLW+tO4mOppZb2Xtj/v2UaA6xDenwbcNUZS
Pjl4ce+T3Aw2eJIBQlY+UUBvtQqY0BU7+En+i+faK8sYFtYlOqdeYdxoml6OVT+UIdOkEir1j/+s
u3eJPDCmUIixr87S2LFg4z5hFjdF26AkJ8cEJyveotgX9T83qUYMKuyFV+xtZVCFvcEKYntYYF21
MCgQOOssXts3cxCN2B5M6prgpg3ne8WmelNm3ajYhFlMAhunuQf8S2EwMSMnXg7y1RIgeizcgbjf
WrCxOy76DLu/mRbuaXN8ucFE0yUwYyXKxDozK56rrbYE0h4Qc6r8NRJjk8dQYAlUAO0G1+7Q6x+B
Pl5nzu4GofDHUk08aAnomAHZ077wmuFeUzRIn3b45S3BCck5pLjWAVoR2YpWckDb3e68VHKnjNRT
JazL8+KZ1nSP5y5hV8QA0CmxSHCNiVKM0Ks6HcCaBZSfIgcMni6KgSXQIbRSzL/HsgFKZXh4laU3
8WeesRVejzi7+jW1KcehhmFkVwiC/eni5ww+Iah8CTLVpK+EnixfT5qiBUt5huIfmQXuLdVy/r39
Tou6WBVsCjK9XKHODjl7/Z7z1j4znKcIZ3dbinstQtVdZ0PFdCmUX2DmjsU2vYFLlPk5v+U1mhK9
68GJeNKmA+aJ5QygbODC70jHyXJnb+C/BWCD+sJ9I2I+S0qRy8GWEWkxalGPV+v+v3P4bGSMFEOI
zE0KyIB3LfK9RfHOTRzOmXGL+S0C61mGKcuhHE0TvBesONZwE+Z92AjnqfNHgJCyJrb8mhhw4/EM
XMt1LKJFPKq//iDl52247Q87an9H2strOPLkT0NP9xhJ3U9e0iaXU2/9Jbevf2ysK/K8g5yreoKB
PBg6u/MZ/1Cd0uPwb5D09fNjDhUvv4If9LPXrMElGJStka8uu7fCP04xqz3QqbIYBf+qWM75Y8L7
PtRc+RdR60L8oskUpUTH3Ehl8trCF1vaK9Ot9KkeXFRa1WTYh4EOxXOqqJxuU4o3e/WVL6uglpxa
GQ9yYbnqswaaxuKtb1aUCfrMEMXAm8JfeFajEYpb9yDVw1TYcytbf9nUfpvTrkQrgfh/CFQISgtF
VeBWiHe3a9RRQpVLxq83qiqhMmwAwYXVKBdQ5tjChBtUkZKwb/yMbvCDdTmTkdyxpge1tKtmCFtM
cDITPDi5z26ireHDXFNMrPEKswVyZPp/ll7x9wrS4tIHieWHTFLCNTyPrI1Bx6lE+459WBIbMOMf
qI2/ugOrEhle9zHglwWVVsHHVZLQjN/xx+QLR8bBd2/arEVYZtjUBwz45p51s0LB9FAd4n9WDXkM
gRpuxDXfpTkrAyxTnev9HwL+4D2ujEn9ipUpvgjdVFc5ynOPZy2N5cH30eWh19L5KYfoV1AOAoJP
DBHk9SQn/RaLw5OIa9Q8B//zcNy6/C3ko2iAgAvw8Jmgn7azP1UqIqfutp0qkF+Y1qpqHVJQGzBL
V35MQSaTDHui3O1fWG8BUcLG5wycv0Dioz37zvghFw20bwhF1wx/ybL7a4fj7SLRKOmd3MgCbpBi
lGxYBnYXSczED8fg++06X15rNwg2z7sG43s3bIsKORPLbz9m/JQtqjTIK6+kVoGLkZ2bH7+udQmJ
7l03F5yOPRjfkO9q3+xR9CvOKfR84iY6ahSGHoIhkCtvQrXfefzaqGmck/bDqm+nt9g3dPUxlALm
tXbT3cjj/rv8jJdf9J0j8Waa22D6VOuMOTlic2Z/G9sKRyUPoHn7Yrx5+K6v3A8NzTV4ks75rUUj
2QlchiH70RSKBopETUWXdh1LrvF3TQsJSkqTh93poIIkpUjinY67Jwyb1tiI0AuJRH9jPD02KXNR
Dq2ig/we5dvlXnlsRhRrXldpFh5VlcZvkft2xWs4Vhh08vJHlcCfZm0FIy/FqlLr81PMN6yxw/F6
DX7MtagV7ZD0O33hkjqWgtzr7gbCLoXR+2wq74j2L/K0IxSb8J/tcvSGL09zpLtf/gdm2EGbQyc4
oBSohGQj9qpPRJU0m7LpIzZPbptQOuTVIfeoUD7N9U314Y6G0cmXL4S2LT6Pvbh7/l0UCvOGrRWg
nMgdAdpkqNzNdWjsHaw/4vcQzZ71dVIOd7mlVAypiAZxSNAOdpB1eyb4PQLZJpmltoK6JGQnWGpo
KooChehEByLs33tz88E42GcHnxdRY+kCalhPCf8PPjllWOaaPyGdWhj7vbJZ9HmHxEdfWaK45CnO
/SCRD2lE8drDpBctQqSfStaaUon3uXn22bOwX2LUtHSbXpptLnscre0ziPAu4QOzbGcdNL+oDX3Q
zq5GeIasoSkgKMRAhwNDORwdkLgM9F9MFoJ5q+kDaTX00ppRlIf6WE7Xlh2c8xeG/TF5kvUWezPq
WSZnEmr7Q0GQIpbLq5D6HCAHn8Kmqas57cr8MujW5KF5FSndlf2EKdIdUtnvzcI1UDGNUO0nVVDZ
RiaRjWUbR0vq4jkGFjehPmfgiUpjv5gwpXvqX7rcHC7j9J7Cb/inorpIAWMXRLnWLvY2RO3BcFjF
/TsXsdYDmmbRhDJpwdmIrT9s1opPCi/cHeiPyxUIw8o2IHyfZ1pkSc1SQVx3do9k0uIDhZJvR0JP
kLBg2lFOFrov4T97IWhRSkx+Ev2IHTFyXdKhcZzD+IOze6PuQxZ2Smjs1iikll64aFH8bfq2abd+
w6Z9Xr3Z83fh9OMm6h11LhJTmJeYKYxS7USOnlbqHZmW2AKtGWgcszLEiFuDzgTmVbW1FoQgTBqP
SKDKdvSl3GkTVVwuwPaVz05bd+aQEco37X7lXalVM0s+boGVNGbBaqG26nwnPeYfin0QjamPUq0O
rJsfGj1P5X80aweRBE+zjaro86MOapTMuPpXDSGLXZaGHqyiIS+a8Ylan49WMuApOv0tkmvS4EGI
QVZW1WbuQ/YorcDbKMslC45kZsvHsFZ31seQQjcHidZxzj/vnNebca4smpm32jdZHvvGNQyUxw2J
KKTs5wXUVY2ZCNOjz6FirlXJ+27n5UUwxUtv/eo2IgAJ+OWt4LKE9d/NcKK6Edi+za04y40GbbD9
AcOsN0OAtVKEBKoE/Q0q+wff6gCbP8UMIv6pZEWh2/f7g2+x+JsiibFmF8SoCDbShmUplDzPph6J
TDm+tHgHrAVSsfG2RwJbreOCTjYeUuUSmvhZP9MTXDFrZepX3SAFDn3arLdH0frRg2ngDqJCUM5/
veQnmLt3towHsIJJIY2d/jZJmkb8YJHeicbRHNNYm8nzkAhoixj3sAOMhXjf5ccOIiwdPkq/fQcr
zfZC9G5LIQ82ATSPkZQrwqrpWbRX6var5fMy7wr0WN5vGij5K95Y0rN2Xo40vVUeMVybDxH+FCqS
xm+O504KhZCGc1MswJx5JB2Dt058RX5SWY+ZCoIgBjIco+gI6wFNG/rBiV7Wr3oyRSyAZ8cxP7S3
Eov3Zqh6WIE/d4FRCPgzkJfoFwoTSPPIP4x6/7bXSPp8cnVBnQg8yA4GenjlnVYjHqjUmbZlPgAh
iYTnazBhwmi2TQyWsgbwSWnVgDqk8dFS676WJNJxUKgGYN1GVB+z5J7Jr+D5diwUQDPmiThkgUIU
oPkQRmaJ+AB1vfLCh+yo3tnFVStq+gX0+omrW09MAm4E+QGKKf3RpvUAyJ1uQj+Nu0z8T1NEef/u
Ko5HIf32W0o1+IkCVXJAFoZN2iWy9ZX2Wz4wVUCoiNP1N9oseZK8S6iBFz/5Bc6v7nRq5XjE7zxT
04whxi4M+3VmRYXXesADKHk/wbS5Nf3O5FR5lAE6euO1PYJ34l4oHDwrG4rLQaO7k0vbbTw4R0fx
pupumcbpxbdWPjLqcbVbKjmJkk+rALu5DtcjSTzv4o/3+rnH9MD69xpZAk5eVyhauvRS1/d4bQuR
m3t+fvZMnltGICEfGW+VoJTyt67afJMVf9pilST9b9rd5R6cj0LXDEoesF8aCrOJQGxwu3DoT8Lm
3DYbSpeHRFz1QUp9LB1XNC4ETFup1mnQ0M0w11xob6r63J/4DhL/i3hW81RuH/fHeq/G1tW3/qSf
zAzPgyxfTHLMWS2V8fO+XcKUbGbMveFBoPUM3gQUzbXvDfQpnhoMA9OCHTm/qVwM/ha3A65l7Yy0
d3RRKBN/N9TU8jYbE4tNsSZhFrf2h97bM8UOzHwSsSPifaKbNka6+yNH4p7ub+dEH8dJCRxXAx8e
rftAAChV2BTmigegZBEyAVwvEcKWGfme4q82eqgWMtyPi7Chhm0QKkBhBc8Xt4x17YR4lqCytJnT
Q4HK7pFv+wi1TARfgq/iLP454HiHZKSjUYxAJokRfieHF87SDPsLikoeKXMdQEEGjDUJOOIURZhC
E+L50mjmjV6SdUwlPUWerLHGTpY/9IM1EIY/Xpf+VjfKmC0dKJ2A1j+cpWIEYjtVCJyEswLWuteN
w3mvJ8CjfMyyRtxkkxSm0YXZTNHM1C4qSyml8k1uc7+z9RXo+8ChGD4DJ016zRPkltr3XPmRJDBh
lLP9il++olVhVQrRi7jkCkod4LbOOp906nPjjiBd2T5P2O64R53QgxUdon1rUfXjmTV26u0oAbO4
FhRwx8gwM6WVn6VVlC5K69PGAgGtIcW3NZ5YNjOO2zto1OlCqE6RId1bWCAAXP74NG+AR1XLPZmm
vz5KS4WnjI55AtHhyW7RHROf0NtKRFCwge7HwT9H+hDobPsFDcNbC0tweR1REqfC+jqwmZZtQWiZ
6UghKU3C+IAmc2jjCzKY+EfbZAz456yL5I2kG0j0fdxKVVVf9i+vK2JjUY3ZKYGtcwIbL9yEREY4
usMG2nKlINFMSFls9tb/MuFzsPltHIdhM/mhFVryMdJe9LB1miHrtsWggsx/sLcwsjD5d+s6QyRm
jjZTDlWwBOFH1fETXOQ05FBU6gLoozh0TOF/93S+e54YNYvWocPUx0XS2O5XT9iHA5M8mGobGwva
mze3OcjnRtvEIkXqh7fbasP8AKReU7lWmj62ZtDpfyp8F16ltGAmAJnv9smNUJN/bXjHkLkj/GuI
dCA1ae+y+LGBnvNr7jHoKDgBDtva1BOpB5v3KCr+Kd8ONwdsSQ10WqrLXkCFbVBj44KWZFP49/qT
RBS7zOVv907Yi25Twwfq4D/fkqMVbZRtA+O02IoROVlz4Gu5MfEmfIcrodt5qJqTthr6TW6qliLs
y3VF4CgyzHcVgNl9WDqN0toJ6msk6SDFZkkfvut5aEOBXZD8o1B5HyCr6tVf2YnBZjIp3wCMbQTz
XkQV0M0G8QqVqAs8KDPfhngjemMlwUA7xFR4C07BdKOgbV1NJqcmN7ZKf5ae3a8T/LshHCH1HKRG
ZrzOaGl45SUfe7bZLwdi9BTeJHcX//CcwiW532XQZvnBn+4MAl3V7DmneI4YrHzu7BQp3E/8exiv
T7hKxTQjl6ufe2GdHsEvRgl8Gjgy8v5gyMt8KO4KqPZ1LDXNyaZyp08/DEpTJPndGQjaMGntZV7Q
7xXnO+VWA+YEwP0OvErhLXvLGFeV4ES15Jmv8zYMv9MPNejLl2m/El8iVfutECxwrxhBbHGVVsxY
2SANJ2fYoYlEQwslRADLlkbdfGs8ZZb+H8nxTt20BMQvsjXNrV2Zc+nalblPAqqTbCEwFGZsbx7M
9wIe5cdNKjfPeL59BM7kKeVPcMjjD9IZNrK9v3+B+mwpXtHT3SUOXHe+vEHz1dqIQ3b+4AqT6Na3
UxZ4wcc/wEAHQ7/5E2xH2LMuWP9qbaFQNXhWMhay7V12146a2pOUNjEqVZN8BqT3HPkdaR8kNh3h
XonOE4kuGPKeeSL0wDMBIc4xcDwR0ntykohhDpANeDY0jbX1L5cLsNthv0r/gXzrJX3Rf0sIyN5t
wLUHQNbW7l422S5nYYkzQiBkTBO4u2oNhg0z8uYA+azehFXRnHi7orqWtB7fS5l5gvGG0YT53VJW
E/er2oKInRs3wgw3Y7gteE6NG2Gc0q54G+qvaqS4AGKMpmgoDLp212GjfprttSHvA7gtS1M9sRDx
SbHR8EeXLl4lqqe8oKQnPnLqzWVYmivg8ejsGGb+zgoYJ5dV2NdLRGgoXm/0CJ5cw8HiTTbLmNYA
FNYDzMKqCPnXkjtRxGwoqobtpbaf0hU6SfMDJCS3+MGUH6SWE6z/VpLoYq4QqyUT747xHL0peDpG
kyOEuQ7tyMu0j2jyZqThpEBWEs+/3M/x+/A59OU3G6OzdIb7hvsKeiSm+eJA4VNN8rkXOmWaBYVm
uZPBy29BZ14J+S1YAzFGmk3WAST+8xwKjJh/PPLHMh2vtrsGLYqeiJ0Axn966OE3lTJz70XoyjB2
qedOdnOILbS1zpR3LlrkDDYM7mOY8fGq90sQWflqMVDKf7WLbl/7tHk4oPqPZ4/FUxO5NZQyA1mt
01C36eM5CMrQimGKNGDn6LUQuqV4y5v+NwnrSiwmfzk4QnDv57nP/gVrpYqzIUlrrY9vWlehTAOk
ga/KE+p1WxR5L8+ldPENS0eQLJm37o0Sn6PAvt8++x3/sdgQ3Hf6lKLrz4QUPx1HXuA6Rx9mY2co
izAl4jJvTV87JTW2swYNIZ44PNA+hWQyPuGIuD4ppiM54aVP9m1SMin4acY3AJW7vecaILQ33+Re
LJKMvGUkD17MrOPHGLtIGwj4IZbMebEAGngz25WDtr6Lc1bwWSAAqZGZ4HLlGQ20f3eltU2e1u5j
g2qdFQb/EaDZDEKZ8M1YJihQuqXsIiDPQR3XpS5xZrlCRkiFEPZRj1DukJIUlD/jf3nUTUE0dtQ4
R4RHxxj/wlm8s6ToWST0mBedgBSCfwbVmUg0SmwwuoqFB2REQkn+IUO8MmjCbYIzPjgecogj7DSg
f9mE2XLQcYZmlz83tW39KS+2oAPH6bVavey4F35ZBJs5GR/1ZnZoMmek5NmSYYAi3d3ko6cYSdJO
TDr3Cmg6qa9q4v2ucOBQ8Wdufjp7rfW0KMnulrwd/Ry5LVliAwh/S5dXc6VcmNR3pUyPxzEeKUrA
c0dxe1UvCxYQNqtwG9P6zp0m1Dncs9LmAbOQm2yVSWSDFPg27wBDYh/Esu9i4JPcNPI45HQOVJ0D
vXXq2H0JqJtnxlXQvMH8DcVQDyvtuyMnJALDeMBhyaJWPhlNbRslC27iknqjGzVjlEvodcvgalGs
39SWZxQU91MeNF/Jn75LVGGG38NZoKJIYdSAuIyOHvYltPQHkr3zDy3mx8mcrlcxaLgfSO5uJLxv
hgcmYLtKskcrBk04M4dRdJVbkt6GMmVobBwgQ7cc4i9+4sj+OiICFwqdleP+EhifKVDpfTXdjSPv
Iu2ybX9Qb8RtQmpacWEnDcgwYNl4oPuh+nLsZiq+OhFrsj9A3RzC8uwHeCMAwVf9SbzxHg2o3P2r
hl2XLZdgJk62LffW2dYSNwoZfYTIGfw0oRKJlfcO23zSv6gc/DyH6XwC4pKM+lSqN6FUahbt+6U0
DuIoEKpaWrPR5+rUO2XLgP6/uvMeHVWZDJQpS7rHzmFWASvUHCLDZ/EXPKQ4lKckHXwP8dnFI32D
HK1A9kxSvx/vbbPZnAatda5CCOqDyB8CXvo7oUK9tu9LhiUyEg/4LT8mvqwn/NdaBp+nkE9ZdgsV
leGjAXSVDNcE0C8lRV4AHY6ANcll8+yWFWiyyHlrEszqn/razbSyQeeP3ulMcsQVjofiDk/mOtcB
1iUoRr69moZMHHhOfoBXHPPOJj3oZQDuO/z289nxA1fN69BC5NFNYg9tppdy/JC2v1C5681YOPFA
0hCMe3LipGpv5P/83Ys6cLxGiAOrkyoes9770x/QI5yZYsHE2jLan4zJ0hn0noxwJMIKtQrHCU+u
8bR2r3LyYlOVSeIlBLI08oEYjqWfrJ//v1hwMiFFG0itFwmhjJVRHvKjb9aQvofQTNZOPgDKwyEd
LMc0evJZyX65ZS0oijRRWCvnOFjimwiCwNs6y/OEBWl9DlucGNIhMmLo1KvjJfpvlOl+Vzia9F1s
qSICKdnNuwfm2nODji0Y/kXBkXUaIQRE5vuB5cQmJoIL4yL4Hc7knQdZvv76LIFvf5QsbFFABFgS
jEr7pFADEG4/AGANgGsCaSDDUqZT1m7q1wEVwgGD5qLMBoZauvZdpb5ggtAwvpx3gCj7aMtrtvz7
A9xF4saADVmbxclEITroaaM0e8RCDW1niC2hh1EL5TOoQ98Xa1CqNKQnfQjASxF3Ysfzbf61knu2
z336LspgkZpTZ5r8+6Hpu4XFNnfi6PSMFG9HOAfROQrLmfeADmffPmG0j9OZscHz5ykMFAhdiyes
+qx0VQmIrSVOGCc7y0PnE57Tl+Nuu2XrurSfRc4fEFQXtbjQ3lk9y9EZTsuVVrZJNrqPMHo2W/mS
ekEIdCHcYagWdOcv1vWZB5LfGKr+06z3Im4N6NQoBXqx9HPxEpm1diQdadWCED+XmaWrXRR/+Wv5
Tu/NcLj1zGq6ATF8SDffzRYBIHow3A6n1fPIHl7Va3NRuumVK6TP/ESnTh0Lloe3M9d69DQR8HDB
BcanMKHwK8AXAFOoykEUCD7RLODwYX8utuE07Del2QILmNcg60V+OUUMeNMUldeQ7As1pZNpqtqu
Fn76IxKkQZjHafcQBc6pJoyvzYHyRCDHHOqAduuYtx+elv1+BMTjyhR4uwu5tSQi7DBWYYyVRJfp
B+rlD7uYxvX38aO6q46p45N8p1dlKauZ8q2zjEaCQ8LFnDzj13AfUK3wmZeD3lsrq8LaXk5BThh1
NBKFdwnCW43rOxJM9rqro7qIXlHRnWbZvxRI/QFjmXyuZb6CV4TmUWjuQTW4BsdahtDTY35vwYRj
xoF/fAapPpbT95Q/Uj0hnWorX6iU+p+D4ZH+QjVmRIOrmti9lfeMvYkiY2Xlhf4xsFJbfT95IX24
3tGBtrzlFwhEP9ZMRL204Hp4bdRsqfSBLvISQo8xCo6rt4GvEbcX4p4+0wEHK/JcwEHKEs8aO0Ml
TFT+D8nZacu1yaj/qph4v6h4tx4XiLvnWWU587x9iNz2uy7wSHVGqBVEk0oziS5LDAthA3iCIY3U
jUR2qErtxmUT1pt5tHO1BLrTT8wOeftlqUOkPChYDuSmNplrk4JAZzjsiVvp8iLng+X4RNcM8TbK
NFB+RbWXlNeOaGxgXa7VFdHDP/7IMm7AD9tRR6zWNqt7Wkxui/r2HDANrDcCvJ1OP4j8mQKl46+X
p20NL2CX6v3s9XA6r0Anl7ahgJrcaX4niIsm7uNpkr/+VZzu4e7qXeSmvACNd5EV0EW7hGBO+KVQ
7EDmN7llQs2/5ZHV8+7j+so4IaCla3Q58XlfvITh1/fLQ8Y9ynJltdQP7Lpe0PVuP7RKOS4NwaIH
PAyRoqquIxZQ2wYd3PwKOGjZGWzDpJAexfs4AAfX/LebTKVOBwu+/QEur4DMq2NW1dYyqqBKRCmP
UROz/qfo9jH5d3hRQxVDTdo1HhSLhElFJz11lN+EBgY8FRzOm0ygATWGVd+JgCLcVQfTbSLzvXih
RRWqK4AoDA3LOzDu5lMl2+/RUdOVoTYC71OWya4XE8uMAuHv7jjWm8GeKZALBr+Ged8NbnwsUlxm
YrEWcKRGd9crF9+zEx0b4qUOuEliLDzjngKqQtoFKBCzK8pQJHkC9CszZxIPSByW+OoWxKEP+YvU
I99LXfcoDHJzvMLU+oWZONQP7bMqv2ZKYAzaItHSMHKnIAPaWc4S4KO5P0KBANLkItzCEH8PGI/6
DpcUZuL7u3EXBecREb0fmMIDTZqTMhd87tOVAmMXOwaZI1U6499+8yXEEh9HXaQePM1eg9mZxr9S
3yKWf23ZO+5fHUaKnhOhYGK4FrvnJMgzRFmmZlJuiiTGCSUSQcNRG8U7Un4y5Tc3HRtdrCBSheGC
6RPBYHmLKTuQHTGX3DnylXQKBBjTAhKNJRrN/sthNruC8rDwfLVWWB+M3jbARPPYWmyl/uUE6LZK
iIrTuTjtLAGAnAzOwmYO0klbrwf3zhSwSTA1jyhrwwV7fPYvbApIUtVXdYZk0Rjffzdn4sSVOHZr
R7CgOqR9E04aEAbbdfOX+N6sXnfrOtCFKTm9YV9GJRCg9/GDiWfU55P9alH+du46xpJjU6IfKD9u
sCB8+jASiogZk5hIDGYLGpuZsYzViTQose7vrn1qAsyPxWrkPKCwvQJ5jZSgU0UNB05Zc2chwarw
oD1v0+tblcTxWzlPEDk0Y8JBv6ddpKCLsFsHQD7eC81HjFn1WnKOaY3X0TuC/m4B304H8TCU1v5W
rAW1GOppD40qe12FSiK7TPpOiCqoDTEqNy7Dg2i+DC8/u2/W4rUDEGNubTIuTdlJON7gW1wf1wwU
XUhrdmPdthFFCiSg6JGV2eoY3N3W19OePaRXZ43DW77hSJmwZ/91aPkwNiNQoEHR1K/rdNDE6rc9
n72oGwr9b15wfJh5jec2fWdh9OrpRlj1vDGnz4LHT8QcYbgcC4iZ+ADlFUi91SdEENJ9yZ82/oJg
/pgACbb4sXS0GHjYsLEz8oRAU5Fv2BbSkAY3w+6yVNwFcafjFh/yESuSRAMlBX8d9WPh9+pY68bg
MeTaL+RIpPl2kOGjkS95sDyR94pZmAnSxtdjOvmcChPakf00z+u0pfgel4OmA3NIMs6f1qVCmN4q
90OLuwN0mpx57aFjsCBzwno/ZhuaIBvJySjxu42Vo8Mf68dYoKW5T5SB1OgeoZdVA0rkhcvmEYpC
hrxdxqjF7J4gA+Guzy9q8tQOsG1BTu5ZyGDnDd6upqz5TPv4quFYrO6JcT2GbfSM7zINXdyrsboC
VBw7fYKyzxG9tN245yqt+OlNW88wnqspkI54EiHK4c2DNlIAyinvOHNa8AghGqqqaDu71izZzUO3
mUi9gSo+2DHd19V4gGkKbwwv55qUB7q9ecm/FL4J7G1WlNCV/9zmL+Uzu8kyFqSgBbrWJHMrTxTN
io0MjKXDf93mYX7FIBwXFgNoRQq09F46Auz49VtRw67cHXS3Y4qc7qgz9nVvJCAse5iDXSkfgvJB
gOA8oKspKEgDq5+ksQqVBEdx9gOwvakoV/J6R2aC7I7UsFOZFfzQLkvPzO7jjqpOXf6K3Fn3Ws9K
f7tHGHLkIKOWZJA4HjmXbuNdAO8RLoGhq2Ux2NpVXl0c2NsjUEPTvyJak5pEp3+UZhHu7M1QcboY
EdTmgn5fO18hvdNDZ+0ghVjVXFfvjhM3X4jRSufvRJo9MlbcWUtZeveiiLFbWmzQqtQhYiXJ6voV
zAn8VLoeh+/vv9iAVIEpDSgayu8APrZwrfzoAyXAnINKxD1s1RGaFpPRHPe5UyX7fc2CVa8896Bg
XmTgDACoOiMP64rgixrurJEqWZ7V/PQFf+ghyDjo2bxKeYRvZ3qy3YGvnUAudF6EiDvWkZhBWM30
QI5Dc5aPOLeP4LftQKYd6ZWYXopQgGYeED5sg8m0TRQzJNqnmL42nc6cu221EEFaBDgY8WXfY2hy
8QWGYMIQJJiv7HyiFOuTzzDsBlg8gOJzY3fvMP8cMKKvwncEjZ07IY2Mc98XNQ0Xof8R4bwBTA8D
HecyNcmEmokU1UspZmHAyebUIgpXG9E78NF0Pjwcu2qGiEd+EmfWKhG1gUubHd+LOs79VC93M9fi
nDsr9UCGe72fv90fK0yJd7TUVGeYzaOCBBDkVy1kdAsERGm9HdzbOrTo2aUZJSlSZym8Ti3qwNTL
nIvv9xmkjAxP3Lq5NAAtVWKMkgkO+XkegWVZcegqzUpITyz53dnxPyQhF7vKkIlDKDIQNgWb5Zgo
ntqi69yG5hB1DJhP27ka9QoGHdzWZBefRcrs4KIkdlmvNQfS2JQN6K3RtYl+kGMEDoZLMSbjNegk
YgXENXYsED2XzhpCwsHT6BS/ZdCkA1aWpGl8aUj1A625Qg54YVDVLaTuy2Yd/UvIfY7XSvTiqmoL
wxFb89dFW3JcyzMW6twEuaYIxA63goC7oCCu59PljaPo6xnOCyN7RX/DCXhsA4DdZmCqjmsJ2UJv
npX+l4SgxJYyx4qpMpOH0h7zlGfTwkCJ9O+tu08gxG+YF2jyUOIQbDCpm74KYXy+Xg+bv3WGwH0x
Za1LS2bxr4tsZgMNXO2RK1U6M17tcr33F3GKv1LxeQQ7AQPmZlRmaqx0aL+QBu8DkzPd5687LlYa
Juo34IiyYhp7pfFyFcdOCtBTvYsXp8NziafE8O7wEdwCEqvwDtTE3dh/w9wXJzUIA96y37HP/tmE
NMWvwb12tdF92g8CuAiylEvSwioyKkd2K5aUhlcvwasyjXuvQAn43n5OUKBDPoJ/FwuLl+8dIKSN
3/xITgwm+JOq42jVfaojzeal+D8iAQS0lkwB7UjlA+GmBNrqlPHS5dNHsJ60192g2V6oJYBJ714p
2P9yMIY3sWsllPD4DucPIlgcBMpndn2DLAgArn5VODG44imU+l197H7jnEmCP/Bz1PxtpBo7H+fc
DGplwALOn9YGxQH4V6e9PTiFc43XaqtE4lVAYRIU3kMjPV0BjB9MY/xWGLZ0kqmGxVczb5SI5Nzy
FA1MZYoLsbOlbeR5L+wMnXVDoOAcFwoClNSuMFuTDVXNMksXlINu+sSwIfsjRMywvHniq59xUWxj
HdhN14KCe9BpvGgh45Hx8oMvczL7dpkkUV+LSSCbac3hw8enmfm+pd9QlRySIOootLdsNzNy9DaP
4LLyj9RbMILUmpFdS83zZ9jS+zzkXAeCTi1J4yFpiGfIyJxzwAj7/Yd3uVj1ttehXO0/9X1Dss03
Ui3YtFtHSiExtlGU7W4xs89Sq0rKc4cZ0mTwFj2kpJ2LVoRJwuJDrCUxChUfz/Ny+gUf6XAtjn4o
FFZ7JGre6ndxvSaZlGv2LRElTt7bliVqs/anWcITRtR1iOR+4rnbEnxXc38xMBea5AzyZYTMSs35
vOZQxL/3J5dLWg8N1yhK2h293uAbHHDeFMZgZffK7/DTJn4y8zug9kMUUa4yMSOSU+mmxcZgTDqL
wglKDLawW5ztSoiDgHWxWj9Rc1USMaLIno4YQtnjz3gCFh9qzsPkwf/lq02OIUmGZqwFtGpstyN2
tU6JlgUJBNlUVwjMgk6v18WDoJcX3zK9tVNpGmZh/r52SqAXmaP5Gw2VGyIvYlRlsZ5tHyHbOczy
0ogRoTSs4acvvHdFE3gm7PggCUwOPhyN6XT6iEm5KUznkQVf8YCZh/XOS3mHUoW/UTnZO5IgfN4P
YPGqQzvP5jxxy6MIoIr+9Svr76K/G/rphtPArCV6dp/CiVlESPCZUQLid2Z16tvaAHOUkHeo9WVu
L4FaZj/iwJhimXLgU3R3WFsnIHx7PZW/ngCCJ8K4tFvw/VO5XhBVp4hI8QpZA/UY5VOwEffzdFMk
PZcpk1kudQZ2GoEtQi6cDZD+L1OMv7xKqmdrX0WLWLUIS7nmqG5R7LKRpxOlDv11bKErU1iIA6lj
6czcWKUvHKX52Gj1X81G/amFhdz9gyfao0V9kXTzLBoVvRXFRCxgeay2s22Tnz3/xr3Z/gtSPCG1
gwdhi7NAj85bPqkP24da+A0Wc2PRJ8/OBhzaQStq8WpVlQpEmrVbmTwWsMM8Q+hb/rZ6GjwmLtv/
YTPMR4f/TQwhs//PUpyjq+4qS12l093qS/9eiNn4+wsmBuuMl9yTvgsmCjnBqesQVS1LBVLoCbRA
ZxEB6gnD5mvEzp7qVoEbYzIUvmjoqZXb3/bHZWH3TQY3T0vJtiHogZVWIZIDUcZink1+C4wn9NVf
jBPiaaFCTxVE6YTUo2bNjmFGyPJWh5EdrZPUXyxVdLKKIKYASH09c3usss0BHigqXxWCalZqtgGG
8avJcMJVPgPUv0oqOCtJYhXVvUjij7/yQu6lFBkeWm+NmEedDWB7C9UCuzznOcp4ms7tKmnQFDpI
UjwGYikjusbUaMytLSSskMswZBfeIaXS8gZ0NTgaFAIejnPvRHqc9pRcsFMHzgTiU5o1V81LDp0s
tueSkZp1xJ0GsY3ci+y5TCvkrjwqDmuYPlQo2Ky+9DusgupzohIbJZR9XFfPTagC2ck/wd8f0Rup
0M2OFP2aRuI8lcFXFCqrUGDBLBUF/et5vkP01D8GzOqeH3K5stIy0/xSkTaUEaxDMFV3IVPY492p
7IFptU7CRdbKLVIgiYTNEpd2owj3BwV95wjXpCn0HJk1iDIgzDR1cQNbwQQM16Cq1hMkxQ3k5EDH
tyf7vPeIAwNRfN03jWyBx1sjTMUDZ2K4vNT6QVKYEu6VbV6oyYORiDzscvKZtBs4jbOT2QkUptZq
pFSugG1ouVhZuZamNTeTFNn6Hn/VpoSa7c3jIz3kzRlzuwqWIan7wdcVn+h/C5tpudYuKUy0SJW8
LAaPXGiyPYR4PV2Orn3ER7l1AKj6CykaN9mzeQQAQTZmH3DXLjK1eXWxiOGSifTG/bkL7Te9BlHR
+a/zkNpe0c/3yiTccEaFHcvtuGt2aZaehqyr1hwAhYGmGZZ/LtAxlEcwBeeH8yUSwd0YIZR1I/KL
7TWiAMWgC1iu3CLBlurlM203/lbOC/lSXRfJNHeb8OcmKF7hK/xmjjnyf/ekJKEIMLEVi8qgDy3R
vpPNVzkdQSpequqaeCCT8W0bPss+2+CFnxdEsGFlEVqI3e4icWFYv0M6m/9Cq9XLjQ1Jlmny71Fj
ZeKMuu+zBfCFcJbs0fZZNXsTEi5omwYUw0oGKu7y7qaDyF6C6VNa0gGaedrU5xvxyfckOT+et9Xm
+NPSvdHg2lIv/TpU/y8ZB7Wf/DgRorXwEE38cJaB+GP6sPFN+7u55aI87Zp+q7Xes90sTUf5RQcz
e7lP9V6PtupGszd+q5pNm6Wb7sLT6llfof7A1xW5z5s8Gf/KhKRYTb/eVy5JIz6fhjHoqy2XJK2H
9I33qAK2CAkgNkLyLPu65YrLCaPj9S5kv2iJWQPdiTNnZOfvw6EqznK0LD26vdGP3a3dO3IVqPI6
xnQrCMjMAnrrnc2ItZqRgfi5zMAM3feD0280n1PFWGTXEoy+RerDX6hdirsrhSc3Soyk5PQUz61b
5q3gy3AtozNJjO/GM42goFrmi0DRTO8UZA8a8XsOfPjy8cYvDrTzIHc9Dnza/nIpq9MK+uhS+UiG
q6YlvCcgU9ZyoTLE8l176I/PM2a0dzsiI0x46jq8kvhMPGW/PcnHITwOCGZBnw0cZ5YqUkfcZjbk
9Q72SYGmdnVMRTibTOZuNz0EjEp/Md9wFuMtJurA97eRT0znmVhwd82TbM+9N+LRGTZgte9RE04r
+ZBSCOjcXmGVD6lnJ8p/HkbCIddiz4pJGJ6jUE++wg/8TJWhPeG/oQUvO8gIifcRChDvBSHk4FOx
SRkdqaM06CqYsJfyd3eDuJ+mFUN16wVmmFa/bEpK4DDuC/0UJx+dsBrMm20ADZupL1KxDLwG2+kI
xkUGtl/JJGPOwod1YmHAzAJdRyVUYomvbB9mXqItDBBaK7tEBWf61FPZu/wkRLD7h9Uakr/2Dw+Q
cwNrZGKKIWRlXkGWelIN7L6HW1AIXMjDc6A53iOqnZQYdpwj6LQGqN+HKciDJGIJatJi+xcrjA7i
XBp7ZZ7OXid31Hyi+u7VLL6Hc0g7MeKSxytNzkiXdG33Oyf9XHM99ziTGmWYfinQ0m9T4bUjJ/WG
wrEbuABEOqr9Fc5dMxwolqgc8b4iM9aFadxFMiPIamSrYLMaLBbqHJplqIwdyaWvB4T2hqPzclrZ
XDLZjQjPL2oOmjkz7r/tJxy2b2qVSQ3p3bVLoOF7cL/0XcWI2WW4w7OSkD61E49CJqbzpYb9hBsC
pTecWFTkKom1fBUK+DyKKZi4Bg084CRROsWMk3pQA/a8gmQDjl1EPoznfPA/gMN6ia9LKDKTeHMA
M2pJlf9QS9LKLNq5zPIlAXj1GVu9ZsTXyIXFfOGlcq6bu9IKn9UKbvxMzaV9FqL9pp4tLvXBHTWJ
Yw0tghIDNrpppFEmXmYOssDf/POS272IoBWLdZPemHbAFfgp6KklWMhHh8fmEcXCDQwHTYP6E5fy
CAVlBpb3Q+2xNGtiJYU0zn8MZZQlFsx9ZDy8ZHJouUJoPXNdeRhEYKn3dLnRgMylN8uOtR+DHLwh
bNdNIndBC4s1mbrg0vOevDNZZHCXBMx7VLY3XM2YlgRF2IB1Y4osQhbVH0qG2qZtySLjgo5D/8az
ShpB+YPwM+fiCF5VQNdEfSuMYf+Qg8feZ007/a/y9O0JVB27vzh9//gQfTO5zFY2YxFMMa1/0smP
ee8cgwV0oI89kBp2wg8vq6xfDILKY6VrrBgvRi0V35LuZAjfT1hM/Ug0odh+x0Wo2qdJSRZz3nD3
LrWU5au23ilb6+F3TfBAhZSlqVV8voDAFIQ1i25Rfs67lsU+bvqmqmy5gozl473vKS80XL2zNmfu
bSH+Jr0kKzQ5b9+4BPIOHKQW3k5CApXxzHb404GtTCQcfSpFxQXapc+NJ/fA78G0TgnKPZkCTbgC
MRBOqIAm+EfgCFxMei9NBW2n/4gNa45fYPpZXGdnUxYA9mJvXJ0sl+Azfw80VfGjIzFS701v5iLs
++VTLkKtR4NyDNfoP8Erosd8zj155V8YhgNY8RuMPV/vCsSqUmcwmIn59pAxxVKCrkjv1v0Jx6A6
PEXrVAkpBbPKZ25doNkeuwm5FX6OZYgIYlnGVgLnDHwe6howw6vSWIXWpUjlmWEKO4FkDu3UAAF0
XCrU8l0qSTrmhzJ9pUew6MGNYtzDrks42tCQbFBVCtYe48a55RQxzsE5CvM+t+eYUT7m/UZy8w1x
GzHXRjono9vNzG5BdCpMrZxSHMmJfFEMQLFsTKxxIN50H7mE2Yumq/idt8ckhJbvTYYPHYAQ9jCI
2u4RzMSd66mYXm9A8V5FaiwU10IaNu69BRZ9zvnTQBtQ6ykoaIyAt9kCSl88SknKKxoLiotkChJq
aIbm4+AHZ00YotUir+u192H2VL867iIfcCTb6D1HxB7ZJV2pOiejLHNQvEshr8/byEN/XCPxSKT7
0NV1zr5UVVT6z+Q4++/BRDrXdN+mHywyl2BJRo+5Mpv5cGcglqqgzhirGI7UzXmHlxIZ2zw4zkgc
fVbfX/7veSa7wFT07gnRVTy+8dxcK6qM7O9T/A7IdVHWDfOVhKouXUcx889E450zgnMSVyqQeatD
O+GxsiBLTciDTp+2zmsdri0tdvRGF6KXyLWPG5gx6uezKzZ7TG1gbEN5YOICwarZ0XkNzPfAQYfK
oVpjPFI68uN4yjg6pW5JBKYgpBvahRgVH7q+dqQD3lAFc0HqecmmznME/mNThR/GN5S4+saexHjo
CCMQRyy7WCTcV2NsQcmyuDwe7WZK2SPNgyPMHLXjwQxQtFfnF0ijlBZXk+BoQmaKH9Sr1DlOBT/t
sgGdOim7Z/Zm3zvHRxpxrKCYD5qOP/0j9859UaT9FtwByEldTjUUSp5l+Kk3QOv44THSmMsoemJo
D8uooT7aEgMfLMeVFnRnSxz/6dsfPJPN5MyUTLKpkAO8SaW4KR1VqP9CujocZYf/SvjcdtHi1xNX
F7LI6xhPuQYFtQm2I3wdfBXvoI0A+DySzdr84SeuckN96frM4FiU/CcDOtqjnoXOf7+EySVfJD6P
jNEeS9RfA8P2V8oV9psyKR1LRho7Cs6QW/6LPANvCX5vGiDdH/uJHy8xJTMPBdcZKGWBaqu5sKTv
bSsvx55U6Y2WwgS/ttpRrCTMIVMHMaHoehA9TUX4vBPUrXq8dHEkmMxFNH2usI5JIqoIN2909mLI
paZkoWPNNZD/jLdc1VfCF0NXBcTp8vB0OIxLwFDQl90cQRkN+O9/T6f6PO0Ta1s/PsFrSPE2dC2Z
5QdcK5q7OWXoxYb1LXvijTkn837+xPNSe4Q/zvi3sjeruTdITgOO+ET1fqSfw4VzFcm20Evw/wzV
4uMCGiUh9R8D8eit2X3U9E2unW8J4Fajm2H0HKpUG6ddpvT41QJZhptfEXOAYIfzKxrARUCDkSiT
a70zDYWxtuUTKLnyYXArqlxLG+uFcKXgQkrZ41JtrYyB7x9pejvCY1lepxfYfP6sON1TuFKnj8ID
5TX0MZ1TRwc3LiV3GMIJ2qvc0TSooenflT4oFlphffkEKsGXOYMdROdeNOfNVYEc4rzgNOpYrNqK
49VEcSijp6l9tCwMDRXax7Z1xWPISWNCa3mNkr3zT/zfD9T3FTi5Nc573kASHi/3DY/Phtm+bsIf
1uitH0RBFbEcFVNxXvF+I4Z+d6l+qRZPuPDRXg+/qP29abp+VioKWURrvr1KZ1/nNfrT6x34MoeK
rUgTv0A9zeOdUcJmuzx2gF22dBwvL/6ddzJjJsY6iYiMcpx/qIgbO102u8lpsMt6W4go0nYve7V/
UQA6F6x4SFkAZEDvZeVoHHhInG6Wz3zrBgoribKAGxHfCVYJhQYPFDQs9nUN7gBR4Q0KYbjMiQAM
A+75fOgCYKb92FoT6IR1vHcUyTsux4dYZHayQbM7VYJzbf/BrhrEoh6jjiiwsvMzB96YHvt++XQR
fEksZRcGhwXCPBwAMM7fJ7s90hfOwj8t1H5JBJ9GnzQxJahiQGLNZfSDqhoasq3x9vEgmo2Css+K
1CU6bI7ZSGGnAsm0zx5QUBo5AUg+N8YTanNb6H/ENIMOUz15vOZulnokHuuMeg35y4SgQONaBzHU
F+0+YrSBDSK1eOzlDWoGwovNe6S1cF8q4e/pqWigXo41Vf7mtb1hBAjFPIn6zcVG6zBBsLvxZVR/
O6Tx43XKuQUqscJQP2NocCOHclBjfIGsjepi6MGM+nd6W3ksojZAGtXXzkLntM2HNPBhUPg79DuX
vDMIIEXzOeXR82mfQPOzDq4gKmauxFBQUZoF2zFvflTxNvHwfIJVjfFG4PwzdYVWwGf8L8cex95T
ZMX7wXj/p9qg2In5xw6oUD0G4thcXvDZ+68+e9qSw09Hpjg+F8nEYm5RzL/VuxeIF5+6m8O3sG/n
+0m4dpsbsiPju7bMKkGHZ/sGZTrojDka+sF8l1DHB6/I4OQvfhz+vK9W6TySuXChMXhZEv+m5LTk
KifaymkG0QXLHg2WtSGIv3tA7vAu11qKoYpbbCCHQ1e3ppxkieis3znKMf8SjDY6bve615bCRwyX
G+JWY6XG+pg2ig+spEaslMdgR1XQyrAQcSwCWiS4P0zV+cciWffIWo6vbbWZLnzUNzfdWwGTA/BB
uUQnJUpL5jc8gkNBsEsoidgAh338VozgkDY4s7Y127EGP3fZNMUSvEUEbYIuQeFN2tlUgPtLFkil
kwqLOTCIksyZr2iLFyU6zrpseoCbX5lbaypa1E4BLo0ArBfOz8gAin2A2MLx70rnhwvTpoRS0sKg
nLRiC655bqTrG+HcrwOcdJpR3/3XsUiNgTbdKOzbd+HIRt39dNpZRUsRNYE9DWtA6mEd6InbpcaQ
W0JEEykfYjAOK7lkf5ggvOSsTwU5dDezjkJyMgx7CvGqPTRR7E6veykTzeeKU0/eAzOpo5eaB3QC
yT1Xvw6FsZxtFt6hZuC2CAf8b14hDXxYcscmoLr/P+oQLjS+ImODkOL/3dVnCp4Pd/MOd9OFslVq
aOsOLoTbAIr/hvHoV0eqLODTO9qkZbFX6PqrSdytPRbekfxypbHpgARByrO3pp9FxyBJpqkn263R
stDhPep2XHUBObJa0e5BzmPxaNtHvXmBKZrKIax5/N3r5Q6dMElEDhSD/m30rQjuTjk10L4ON8WW
VjjqiY0IvGEFAj/Fp5iLSFV6b9ecfufefMnJJCYCEUCDz/BU8VQdKnD0KjM3ySKCdxTFtUzm4WCj
cvjL1TR+ACnmzMzl3LPCqdlajxfrqAv/ReF0l2UZfjDyR2inFB39N1TAdsfUygPCmsfnUuMjs+FO
C1e5NRQZnUKU5uBFeZemFYMrQXHQOnoNgUYrAfklWmNm2Pje+Hbnqy5KTTm5aOj/Rc57KkDUiJgM
vB0WR6eRNYcwwAHBOvJoVVc0/GJOucQVEe11IfDG8lY0Iw++6pZvx/M1oJ4OmHYqnQPN06KcEVW/
P8+nM0iQBSacGbZYm7t7bnRjYay05QgV/XanoIXrWWsVbyNSYocnw7/8CuBAGgWSR3YiO1AUYFIP
G+PB7B+RBjz6tQTzjgKSCfbzl9jRz2Gtita2hpK4fjmdsDXp5/j3f9e/CUZrlcDUYRfxSOPpl1F7
+4HfA+qzj1Tk89d7JlyKVHddSu/qOPz6LRUwcUltvXYLHcFuvZJFKbNnFb107L97ia9RzhE6+dvY
M53YpS5XOnjfdmzlqb209LyxVRE9bPcM1PJJ9rwK4od8AepEG5VE6pbSnGV1wTZ90VVDBTO5Yn5j
MFldIqkoW+OoYKIroJjAsTBgbf2B9KY4tmHLln8xYr+4cMssGV6ABF0Tkrxm1/v3VvFvbp4BxDiT
KYcazbmzTFLeb9P7s/rxBopyCeybXTByvwNn7zmEytijrvxX7AdTMi2fHt8xK6JNRit0asWxqdQM
wCvVFl4q27aA0gaXcJjvl1RS4XT+DBzongDbjeP+yuf6gYUltV+/Xv3QMf2MFmF6zeb60neWMimG
9LwyZr3jbCMuI67IwD32hmurol1/JMeufOnSEHEjqKbJzudocThSTWpTnRw1ed27jSsRFR5O40yy
zfZWKpTJqL0ehSutzvn163RlTba/yOYG5RNPyBwqpa1FhRhLNHc1jsl4Vfxn3jNc7CoBm1kSvzfi
dok1E5iikOiUyyGMHsJpsDHtHhqg3iDO88MoiNa6miaqH3idNW2PDPLy0TW0fztA7vohUBLP9/Cz
Tql3EBzBmDwXUzj/A27F0UyI7LNxzMFp5Wz9b01vCaMiSx7BkZanmKM2bi54UYtg5P9/hf6gFoe4
zKawOGRXrRIG7Kf4qqaMP5A9JzCCf02ALknmqmlzFjde4cVhl7BM5hDMH2fMaQsFrU+e6c/d1KqN
ZQUf7IvP+2VzX50pfd6mPhjNNFKCtxb4GkON3aZZrY72pxPD/LwaTA2K9zXDs+VGAODdKHF+33m9
AqqL2dxfIZjSTN3TdnI158Vece2dfqzy5Wg9WSbxO4FhJN5tDe8IhcYHi9Zp09yrYaF02PnI07e2
3gIn/5JT4JuOGsi1AKpmhD17zbMeanKRpWWYcJ6NIXwcwPY736XF7TasuIdLGYuouEG4aJsq9Ouu
V/8ye00LjV+V5GxntHDEhsLrqV6/222qyKvp0A94vo9EbaIVAZnRew3GBVKzKkF33Fiks5Grky/r
3JDP8rxwRVH3l/ekK14mgNH8U4e5RNMxl/MezYRy901BQaXSp2WobJWQXK7dsxO2Xukty3sou1js
WOTMNKswqk7EkC0SlE7VvhUIGCV9FvDQDr+cOYF8XZ/fDR05ww+bDNNeZaOfNkoWqZcjWk5SDitB
WLGIv+I+HCLxfLQnlJQImgMANT2FnMDFapoW1TBN9Qepe/4sQC+KjDMBA1/1k0BOTnH6SJ4qZ2Av
M+8g35swDanC6h7BrhgayfFbafkgMEpJV7mqMAe8D4zmDMiUiqvVb5UMEgPjlWrSXSYjXm5L9qGN
sUi2uxPzzg/em+0Il1U0UC6ATOwoR3RRFHdhYgLfDHPSj9fx+5s82BLrX9T5ptW5ms7gfR5NoEGE
fK2ETnq/nTeJVx7GMVIm6Li6O65gp2Hy/oNtZndGPRa93wzMuovnSXgPOQv1MiwHAfw9dkku/r6K
pfmziNdKuc5sZNjeLveL242XetfWux/Id6wA9i7VZ4MhUo5hd3PR42hCNpFB/kWsyOQAUemTIK9I
RlcrHtSBwLPB8Z5RSANopJ0t+15fJMHl8f1RG4mIEQekinrwOze2UDzJ/09g0uAfXP5wNueAfZjq
dkQbPhGRsgi6hONr7+KjDWdNpwg6W+hJRpRP6hsTxYDfGCCVaurbBsL1clNnDaw3cj3GH/sV67ZD
iu8U3x99+VA6uSs5FmXbdMxlHBFOCgp0pTDIknnvN9Je2A+Uv1xa4k20yfrOs5q/bxwmxQSWQRTG
jJikstIzRTLIlOEPeevTKT3EE1bfZHYSP9orSWd76RXvblrQdaKCRFZMtTXj1poYsqltbvS6gSAc
TFBFBIG5fhT+DH/f0CV14P2gaGYb7ozuNLHGhYJ/k3t9f3IDHWKc00FzoYFqJG1ObWKyropKQ5M/
2xLcPkQlEgYzMWrvSbke9I0SEQDOaj/QV0efn4gOw7BBzgrtWZpNhI9s6gyqNoll5mjuIsCmdCQD
FQbBfd5sCNKT58maED1G3CRAKGBnCjk5BW3JSsyxWxJ1OlI4UIdUIIz/GVAtGVP6MorYZ589sEBO
tUJVJfLYJCg5ktRBZ8MEnXyYlSIlGszzeI4JBXNrXVN5dtnHXabzW/vJ6srkiVv1bxGlqVncxM5y
o+FoO796we3NalJY2ur008jzAXePTB98euE3XecCFd3bR7HgGidFk3Gij+OMute1v9aDEZL5TF+E
z3K0ahlNsWeDDMXzaA7aGChGWE7Yngp0QfY0VM99R2lNI9ORV2LQ7W9HwGYTI/7r47TT5XIQgaxC
TuM9t8bojbTIVmx1WdT8Q4uuq6o8PxgB55hvDCRAeSUB2Xxe0WTg3rNwkhyhlIfOvhNJeEi65pu5
VK8jdbr94T/gbqyRgYi+OW43GycH8OEQbez4HChyGnZvOr4aCyOVs8rrkC23DS5EKCokJZD0/1lp
0XpQE+m1cLO/hPBwQJ5YzW8x4M8WnDm83S/q4b7ZnTfNEaBgnv+ytLUNYKvdmj2yUSNTFOduD2Mv
WokgGFJnxiyaS63d3EC+e4I1gz5/TpVJPl6FJjDtYz5lEWmFIimx1tvLUE76JOYqKM6hqOPS/cio
eT97a5oygcevsB/lk+VdAhRTmgf6y64ITDGQljckApCsDhzdDlyj2b3XDqXl/VWlKjjfG0GHYFoa
T5In5AaEnDoC5vtNzMBBCICwpGAil1mG0E87+ZPFAQDbxTcEsiKJ6n/0RO4LNCU3xXpMkvDxFE3D
VIrkMD+OSmogseSlpHqb2daHxI3yW4XkeexIM3L7PZs56T9rMntf1tf8voEc/+1J15isX2Lu1g72
FNR353fpRIM7Llfegz2cn6mWmppQ/vELYejcnOt60ilBWY3bsL+AuVD5kGROA+hPtw9cqsMycneT
AtcyQ7iFSBAg2WbOHkDZO5Fj6hw7H/eI2mvtJRW/z56JhcnV+TRYvML9c/T4UTG/oT22KNXpVx+a
8xVpVs+iGed9P69MeEpdX5+CmB0eFPqTfK2escscXCKD+ATic68NtO+nEbxnCForkxkcAY64yCmH
rIKnI3De1Hm4i2a+3/8fCciQ8Nz0WQqEGL7XL0nPDjSASnQaTzxQ6a5GuamM37V7ncZrFeniUQlD
H3LkyMrsoVtYPCsA9oBDhhiIUoSwvncjVeZ2QzOjZJlDaxvzlFXEtxi/MNKsbnrMuEFw+jMXP4BO
eiflBgioJKVl0hC9nc/xD+BKleEsuhDXQolxAiL1aPLjZnZO3lLz5UJ/xXK62O5H0lKxTGcY/a4d
WkgsyM8Dm9l8+gKG4yR2meqlOCKGeagsXLO20ZcX4xGyaKsGbvphKEwA18mgJ7IjveeSXwUUfigA
olWfa8lSLnuMkbxHQlaTW+wh2fLhj0kl+gKY9KmTsVjcxw166oLQnTfZZMHzvKPxaURBvPJe75ks
c1xaKmjrF0cNHoyN6Yrpnirp64nPmVdHxpPJ9iUw8XoSujtJUf0VZtoPtv/RrBj0iF6Q/YBG2NBR
bAX7pz6ihQSd2JANQE3njRYNdzF/n+4G9Id+mdBCFpLzk+CDAWQMK/49aIk0GuoomVGahY2/51Jg
p5cW2hEnzsjmxx7X5zT/FNwBbBWZ0NfiWp3BfAsf4EAalnWTIjd5wSD3Hdtrf0ot2sg663SAyEYr
opf2IFG0Yhm+vgqPssRnSmxhoyF297gDz44jgGBkKndpO3827EHv9P1XzEiJPjvcRG6fofpU6x50
T5OrvFBRIku3xF80mJ1jTV9w1loHSisGdPQSiq3oyCq7QNBK4bqkp9bPJsQr51ySgjlSPk0zd0Ep
PpHiCC5RU/ZpS+NIw0GTdRY49CufgDV0dJTx52YXB6DbET8fwky94S4c2OjnEr4rb2cYU9HUpbWS
0DZHZMVSNVy811b3cY9WTGuvudnlgGa/Xhc85XB7HXusNa4f+SsFHBcAu4H/TdRpFCVVLIJCY3cg
No3M4aXTOVoStBwtwcxZRAf1fAkMDkj30JwD2c8oLHYD85xR1/Dq7I0PYxKTj87rgJlG+onXAAaf
yDRy9NeZm8PL27IWDaipLDKbL78+ThylTG2Q6fwJMSwEPtg+JYKL6rkEaaLzQyiZ3M1MVL+8ChF4
G1Ce5Yh16h5Ojhr6uJrsbrz2vMNpMOhk5LYAwlaf2KPd4xEWZdpoe3h0UuPFYbtrHvsu5NpQdEuH
REa920qRe+8h8xBFeNNkl4YYTLfiXQxc2+ILFOfk0EI0FgcOAZ7RtdIZG8cuMwGFXiFszj934wly
tSIDRF+jiqb+KSD/l/X90yZd/8/OF/rOLwiNmteGyHB9hZBU/eyjHNF29gXsk+Tkrw//2mPdLA21
FdaZCBfYKY33jBEWoWnJwROMBTg8FXjo3/3d9ueJvN+UUtubxXKBja8FGQ0xtVeOHWiphDr1BoLj
2bbY7TVMr5SW4W1MOOCXCwU9L+DAHURHxbajgu86LkikEmKMrDb4GINZdJ9j/ePNcNmRyAdI+H7z
6xdSe/+at2g1cMSfx3AklatpAPS01D6GoTwIYgnLi+Z43saMDMXwxl4J2xuWt6I0MHd7oQdxml5M
fXMgT/RTgMxNSgE/3y2A1yvufhmsewUfwb6soiCcK157LzNCjRJhU7WAKudCuBR+4WWI016qz/9J
b+d1mJjTdcjShyG/725h6/LreQ8tTCDpPbBQP1BihIE45ba4xDMksq4TvCKgsonFg2KvTN1NOr09
23DOEhV6cdSR72NdxRZ3rinGmqKLK8V5ijRlK+7ktLTMnoRoKwtyx5rBDgYupdg8NLLrcgZ3gv1C
56TZRFBliB8YdpqqDMuwL5dAOY6a8XtOi/SQVSSuSucSBi5bWi4v5mR3ZONXdNuk/il25Ouzwxrt
2Ni2FQFMCdiLPhx5amEXUCVVXEudssD+b0SHSE+UrRHb4eQFj1Y3hGI8b5QRcIV9qWkzLzbwvMp1
d6/TRcOapbklJsR0H9aYVIGAwBXGm5wj25FqphfWWoHKfvBfKMbotMSi+29Z7P+NqFxwxa+62OWJ
FNHmrHsAEtrHJajZJ7eSEo65CFQ8aDN7N0pAeECkytlyoEWTl49nJ6KoNK13JsTtXWEDW7Z2RW5I
4x3M7PEbaw2p/hGYTVch4ZPlFcGoOEM58sS97p1h6Hm7gEUleeGgfMo1lnPXopQVu9/il6l5SvIe
rPN+44ym+B+KrLTY1Ztzgv/YDWlE8zczyNXUnt9uHsihE57aUQo9nJWd22C3Cf73+8eXWlWqJWln
55EzsJNnWzo7oBKibsMihR9F96lYRV4EFvcuuv3nO8Xl6twJrXeOTDdiPMAoYDbHhmK7dx22iPHW
xftvKcatT4A1SO4qs1sr+VejZNUa0KCoLvkrY9haB0SaJ3M5KxIyKFsdfYEMtLCH0juXB/pYCPMi
cCPevdDOHoPN01320TbSt8gFWxALd3upu6nV9atHXij7g7Q/kzhlOUBams6Wsnol8r6WgI60AmkS
EmPcBkV/xPKCcTBmEgpJsvUiHWvhUFJ3rpZ0lGX/nPxLYUD6K+iRRdqiGZpoV0zigeBYsHnunCss
ig9jpF+6PY18HmorABT03+BuQcImkWY4SojdxSappp/UZdY2s2OhLF0cXe8st4DpqCLifuByRaQ9
2bdf4KGvvN/OrYXwnsoSUF+w+CvzWpaZw/WGclV+WInOfKoVNwweC83tZJC2oJzdeMHPlJsjmzsX
OZpWEBoadJPOJGv41KitpVCLbpTf8j4Kcp40brm1yHHyBp0vgrXGYV2MtSwxL2RKC170F/jeylLY
4doT44aY0ZGubsyzBTfmygU3tKXsmdmskG8uzAv3lshwEhU+bI0oQvZPdaiQKGToXuFISKBPZ7eT
aydQ5RdhiWcQzUicZmIuGfPrwMxEgniGzt1THwdOLuV0m1Tux/FDq9sx/NZrQ4TbCA6w9bfqFJ1E
NwfQt0rH2yGzIh7BfBC8oTleqbdlhBV/TczaMDB4HzcRyPTol8Iot1MgJIRQFHNA4nGXrecJTVjx
aIixe2PLHd9W0wBnH2mBIuNUgKh0MH6fXfD4/WsSyDFIZeGn0JfU0VMWKsKZeRjQMfIUZwIe73Sv
u8leJfLawlvcm4dqVz4oaod/a3T73XeRpkWuCmTF1fh13wSFgD8zVddveZk64dESMAKmxSan6wHc
k1MSSaTCp6DBVPWzW14qNrqanR/bs93EjkFj80TH9znigUqjsYRC1fsg6PRMsExBFx7Tc/LnVl0y
nBjEAHikRYyXltQi2EtIEjWFfS/2pYm07i6mAtVOrLke8PlKYFsTRpWa2rDV9pKy0rv9XIPVCACV
44YhyADB2Rd/Ik9EFLL8r8S+DM7W37ZPDF9AjbcJsLgie+lILOfqGz89qCWDONHZ4ffSQqxknJUM
DA4cox9WkRmgA2JE85HD/HFtmKGoK9cUsvKVPOHf+Hc7cofC60KpAPsp/zLiqKgzZJHwkC4nCPCA
uvRUKO3nqnsFKISrERb8nyPNYdnhSEFP7LzF4JTnB23wPZUayMaZt5qKv5apJCyvqFwn3NnDh2/P
zhBPddt1dYFtHGk/dGsLafL1KYTD5fqB0zwcJ69jCL7HxuWjSXFz2kUGzQUjbgyzsuWuBIeLUN8m
UnoZa/HgJYbQpOhYG+jl3mgS6TYsz3Htnh93ew7uvISGNIBCZPDV8gY2AhPxHLVJ+nPN5C5XXM6e
hYZkH/9CLQTb5T5wdl2SNTXUFaNzdypKNsY4KPI/b1XEut1k87vKhHgLZGDBLKeTCOpiHBI6bvif
C+gqs0AIDLt0dj0rMac+EMJAbB79RR/2Ote/Xso8Y9kRPHJQ2tIPi33kkeGoTvIXPg/waJcPzn4a
1JIF6ziqi4BBIDe8gnyTfc1F6Dexfdk7WDkN/N06RDgpxb5cf9mEyCx74tfyHJgsvDq1ZrvHzSId
xgTL7jy8mbbbjWRvdOAstW4NjntcSCYAOGOi467K16VveiptBYRPonj+30cYmr2NNYdOyuRrF1ei
nH+620V+N2qODMCqV3YysRW40wVKj2+aLX9JzKOeiY1xCrYazrG8Xiob4140Q0JzP/EHkqACVB1N
tG01nuy/q/uxVX9jBNfI3rAWGtAEFr/5LMUlTDRmlyECxq17dmohLHaqj4gooRRPpOqxYSqaiz4K
L7YZFpdpQ/ixDL8qm/XnjjN/l5desSy91tYD3WyNOsqz0hXkohy7uV9x4y+Xh2DY8eqDTOt9viEI
cjROv/yYtLu42vTeKsdPtgV//V2NAxDKA0hd/4mwI4XPo4wUZ9wOaE50RKeYp1MIGCH2pmW4QjM5
zkB+hFMiNBw1VmSl0OnIXI/mCq6kW/lRlvbhD+u9IwHSocWC+16naPZdGvm2ZYQ0xWhG9fLpXqL7
/82iJnf9AcLMYyu6ixz4qYOnC9isnKxh/h3NoXW7C0wR/EmWOfaulRSPB5j+y8n14irG4JnksscP
Qe1phbNmKnSsJb1rhZhZ9VWkzL8kd1uV+s+FW1RUTa+77CFKKK78S4uzETYh/24OTmp2f9yw0+xk
Hr+FlIIPPhOjeojamy4DszW/eS0xw4tpepFJj59UmjSlw6keVwh2SO1jRWjkWR501QcfuDC4agQ9
/vgpkBmGocHFEuGDPFXeZeLWD4iY8n+cMjNoDAnsu3YrS5twpDXmUW/mNBa8/eZvdpBJoe2FaPO+
AFlRZt1sB5u9a1cLXLGcE63myvsspwR5ho+wuMUPfy5oqIZf4Nvm580/RYSIxkznTG8wGoSFycuo
MFApHmLlenqGv2Gn4tP6t+ZEAyAJ8GjHYuATqI9mf96Sf50yLt3e+s2fj5XD2vgUvQwhF0E2FLbQ
f35SJ/OuD9ADvvHiscsu0z8MIlbsFdpqYVOlRYMRdgpAVfyT0RtIhAsL6w8bke7hltZRbq9qE5M3
K1bUlYjTzROvtXSBvDzXhj92Kvl+KsJYXsjtYf4y3HS9w3u3pZ15S9XiRlUR2GrLIo/TOEA7PZCS
P7ClKyb133fZ6WXaQs0NnOggXI87+3GurnIHXJtAY+kHQDULMCIeDx04FOdaHyVJUen0RD9OUo8D
bvFrY6H0tHzyCB0PYcJhDxstiY6fm3tEAmdmVGW8+YwrKOY68WN5fwxfAoYszcI1nUialqr5Pl6Q
EwAE00Y/YnlHA1o3hiuE49+B1Kc04GnC1ZHEr8/S9Ud2RVPO+X6DaVPlfvnAblREDhb0dRPm9/Zs
NZ7n0DVkBg4YqVonH5KtSuY+NYat/YgYH00i09AnFVePwDgC7uZBsbKqqnjAmgo+ufadDwDykv2x
JLBuzge+5CZGkgpWShJDkLuJMnu3zP6jHHPLuRULOeYku+7ZsZh8QKoV8dCtZoDgkoAZnX5b8A8O
SOAtMsfcM+gu5SElR3pVyp6loOJmnzL2yJ+BOhipigKH281Kn1BcqEAmrIPENoA0gg89dzLeNRsU
Z+v8Evujwp/36MrH+3/wySnxw+vQ6WTslsV9aDVyq1e3xsRcVo+ALiAfvop0H/zeRsT/R2/m5b6j
EHGo4P5z3wehnkW2QVJzQzhok4EZIEt0p946sv8QAGWH5GhEiJddfvav3uWeeshPStDsEaf0qxSL
IgvprCwqaR2y7BKTwuPliOE58iOkthx7sLyBUQVdQcdpoRgqlv1jUC/ROvSoQdOu9RRyqSRSyyX9
qVG6aZ6Va3Z+vvhaClhB/VqqJ+h3W3MTK4AgOO/FWHx9HpGOgyt9u1gqt0Nq+NPPzOO62sSh/cds
2x+kyOU1wkc3QF0lzEl2fR3YACt38y2ODUBWTt8OnlFoMqlmCgr0zzXzwtsPVaXohV/by3v0nGdD
aolChfbffr9p4hew3oWQt1PBOnZ6XWKatEerhY6KkNIEI/9PWHSCsmyN7EE7JccmtkCono0/WtnS
15tNkx8t6cauDPFNjM18NwJ9QEGS1eIGP4DC0HXFSy6beUHvZtwji+4fRGDbGk6CUMhOwNE3Fxj6
YnOK3/l7UhBewuO47zlw/eQDUsqkHoldcQvGVADBe+zYBk+bLPvAu20mQd0rOdUEQZQQcrX6itmn
DuF97J7l8/4p3vfB2HNMU0ELG5X13WdAR8PhMBr08maLnuUx6VABTOEdN5oCioEueDxRw3J8tGOw
Bo3ltxXAWBK2hMDtZu7vygp5LdtMbJkoGdOg3GBah7mPiqnxfGj7PkcUCseieN/n5CN/dgkPEvg6
zCxTYZVxIJ9HMezryEUiYI8mYdJJmXqekXTuRaA0EOYzwmS2AN2Tl4BLqDgSbmzX/S2a5lD6+pvB
Z//197fGaGgL0blw2jvbOtZCynkbTLL/Ok0EVe6etvXj98kt6UGj6Kjic/5UGhBfktURwPQssQ13
F6nkRzPxphInc9n/Tsf8a6UtQSC3E/79vJhBJjbGajfomCBv91Iwh3qyS5gZ2L/z/D4prtAqdPA1
awlFijaimMkyUhS4CmYFKVw69Rl01UXwCOrVJLxJVjl2o3Ao/DKbHl5Qc4ibaQ3MsNWu2KNUBios
OrxB9D7w+ww4iDZQCJgnyEhByzYvGO6/95+2QYlv9S81XOpsQm6yy2zxTQmq1ryG+CAoUno56a9J
Nipb6+kVtdy+sf5fsWpYyA8oaHq/UyYXGctt6AAajwSsuJCx9Wt4jIjuGpIhRqJZvsgn1bJrehYx
xvKt41rVT75IFg7ePX1V6jeTWtIaXe2Ufy1gGcn5RwuQK8xOOu2AiLNqPZs2VA3RO4jim4JDfInz
FjKMnzeCYVaCwP2m5QBq9Zke/WWM2BRh5wCtauMBhC7pEPd2DAaneN3oUn+Ht1pmajIvg8wuCwbv
VaVxAGCPoxu9lXRk2OTXtK8RTTdXkbaX7KkQdDazn4BY53RZVJ/O2g7JwOtwCCwq5wac83z9D+lc
jzBwQ/6pCxkU2RI/hMENybutR5H7p8r5Uo06UiRQJMVkCq5fjQg/OC2ZAMH3zgsi0S8KXRmQzMCD
DwvCIVLSPOfB7i5N0hsWHnSmgtZHQDsSMK9O+QEeaPqmS3rKn4j0VPbAAB0h7b4JpWsGnHQjJPgy
AlQrl0GdezdxfMPdQW+VpVpt535r+/Mr10UQB7oERQZ++UFTpVo1U1GMaztO9eGlJPmw6Sdy25jI
6L5w+mfuuIJHCgsxwDhwCVVXvi+45mFB6PZ8MtBo+/jpFkCwdBzxdYYajsZd60HhmPe38FNAIfOh
FFuNHQZFNoZ4h2/KQEKH5xS4QPefZEwUVDt6jHZDagDk4krX4NiLNDJbrpE6H9KdVXNLVwCeAYhN
9zjYq3axo4eO8Yq8quBRQW79ug7I/sgdBiZYQmLqEGWL0/fAhCOuJLD6pCMLQ02UOcxkLT9l99sW
+pPaixXKvBHs58mGtO8CPDGsm13Y5OVppB2eFC6V+r2RXcsmVyKhTgWdVMd4A7zuyOSzDEa/rPZY
uibJ6U//2jxE61VFxpqcpbuChztNHABFTXesOgOO9DqRF4+sEcWgEEMmGlg8iW6ztw9POl6pKUca
FoeJRsoJWVIxb38mrBQLiZY+RRc41K5JJKGAa4WruA/esgsgtq64VdPR8AFn7ubo4Dcf+2BLAc9I
m7UG5sMcZyt/NNf62QIVjyiYkfGFL0UMet8sYpIOkD6St+mZ/iWNb3k1p/wvrL2v+SQSY23Y3LCB
jRRsTkCVdFAfAGBJbAHaFSjpibBdJT+hdAbIjEG/oitqnLyNVAiTzGTxxthNcxmOPjLhkjQMrsAI
XLusoq2x46nWkr6HD+nmJOUUkitviSLYdHq0/18IsZFXRuewCvF/Av+CsqsPMaRwvSC+aFsTEvUz
0fYjqKIzhPGS2tDJN+fx1wu2c9GuIbrqTiOg+Awb6loKLKTgKjHrhth8bO2HFNQ/8aJdlf2J+ubc
ZxMGk/hEZhP8hg3W0lICU9obzCD40jtK1dM79st43/4jyyKrX5pYKl+A1RJ1MyMrmDm/ZjOlIVN9
4nACGCuF8tmcNz736R2xCaJrJ0Kjd2DHfT59GeMkzEK0QZ2+4QayUKh8qVvCOlvZXfde71IgWDae
NdaMe+7uVQ67ifeO1lIJKJjV/Ihsp0K22Kdab1E1N1aXVQteua9G2fjHah4PCvhTB2TLxXuAcjFE
UU2rY6oh4L6gLZsEzdybiAUv4GEEcKglN4z/VZoTkcUJnh/RjkD7rVbqwS25uFSx4Hd/aiIibcpQ
ViwuMusHCyU1wuEZaRSTW0gvX6+GLE/BkhE8KzS9Tn3y3Br7qKmzxrAQogghtOfgAwyPAdxS6bXJ
SpHGG2oAoFdVpbhx5BJOa7TCrMYv/clhnlhE5iSuEbyyp195bP2vBH1HnISbF8iVcGEk9pq0P/sG
OZK6pkpTtv4PgjDI8D9fjVhHx/ZDH6SkQ5O+5yrdkD0dPXGRoIO4qwwN+I9xtt5rEWQyrLrLyk0y
4OV74mqjvS/24dgeSWEqEJaGO2PNQtG+5aOVkFtp0L2h6b6h0PsGA3DDsKibuPPYPufLmEAOSTz0
KVP8Vi2NYuf1eKrmAxdSKs8Mnkxw51+B7gqkkgl+uOjFWWPcWroPMJPg+W+qtUDcHGcGfuzsWBqE
tUhiRBA1YccaCZfWvsgEwZWVBgL6E6ng5Ry8ziq+sLtxzIhL4kM+Qga4xMRjecGB3ObOTprwG/S5
qtvyXoBma30SwOINOHcYV3gbnErMaiLjz3VyEBukNQr3Df5QYPzWhEurU2AaGMkiUI+Yc+iM93u7
OEfvIbaN6hbJd4U7n2IccEZCi/hsUVfKKn5I2KxkdI9qlrNviFI/HHLW3RIUrOGYwCzovEQm062O
aHNBCzKddwLARcJ9udx0dQsH3W1bDsXosC7vURoBL9oOoaEPbquUuzoe57Pw0FfqdLK2F8GTmfZc
DKX/oneqr1HYku0ZfypNvWrOhcWRft4ATavhlfaT7rNw80lM7oX9F6HPEaJEe+V4EDr56I96KG65
LeXuP1vEMIHIxq7S0PL+u9mE5UjzR4u9Al8PPCz4qBnnYUS8ouuny0/1D6RDxTp15IHWqPwJZ4cu
e4vuhwEcW2wTU84gcJPCkFWIg6v67NVZJUlvj/cgYr7iEB3FdncwUDYkcYHsXDPXPvTX5vilkq0S
fqUZX4U9SwTUFD7n3NiKFkAoLZI9VdJGVhcEFtgg7Q6UTund6wVn8vF9YFkDZ6l5jMEZegstnYoq
rTcCjZ+7J/WRifM6K1zOHdkcWjV08jiTTmOD/w5JJ8dd23Gf648vTAHMpQTEecwls4owb7fF8dDA
UikWhJoto1j0/q4TA+8XE3e15tFIfJYMEt7wPOezTAEphdXFxshI7eHBIq54UdCGngQRj8ejjoB7
13ez7veWl2pA9H560r7RcJUIBp0eY69BiyhqyYkgtCm47cY3DwpdoweS83PZHSN/tv03fjMa/gwc
aHhhkpXUf0PgDtZu3zFbEL/H54ueVtxXk0YuMB6CaOO3TSf/FixE8KdsUzrKxzM2BRPEcwkH3L1j
oJavBaCRVFaTwAyCiS9959zasyoKEdqUHRts26wGlNgOyqZ7Oev8ebence9WYQRS8tx+FW+ywMPk
bXAJ0CFz/PbnjbpshQBtBdpqBj+z3qJdCBiGKfOB+po5WlD4mXL1hFCglZXnZFt92eQwfpxqbNr8
goKGEllf4UNCeLAMNxDbJe0UsU3KgjffEkmrEXgkPmbKBxL5PROQXRTA+1agmS9NtCq0KgZ0C4OW
wmBNYhgG5IzN+v4LlxEVAFl0X9LZpaS7qIMROkc2LVTENm1uf5xiWcRtl6voVZrP2gYT5dE9VtY4
NlB9lHxqVh5E4RJBgk0a43O5g3Vt9OZ12rNJudbFdYoxCb1WFe89sKJuJlEsUCJ7/+iy0szrSqci
ADugWros5dt7sQVK9K+9r+uetnniBwCabrk29D6tnpup9bk4mY8JTagwc0WercIvCtGH5UdXyy0d
84eaRqEBxajesUHb7Bz+IohuTOJUJPpdoJ1h73EZio0JRuFAwk2B2eAYS3e68SsMAOp8hWsOPLh/
FrFbzGmaJ/zKvx5A3PztNJmUhTRDZPagDssaydZAkWWJIDFzlEYfmcBCGZLcBY1WaU3O8EC5RhJR
sXKxulQbxOHMXT3IR1RBzkvUtaQbHW3vaYcT+UJFXieaJQEC/ZWliMcrSkKC1l18H2V6yzAor6x4
BaM1j2hjyAai70H3HMu/fhKszt+PLhJr5qW0CCwgS9iMeqQ+bb+t0uheoxzOTpUXvIuVCQpScmvr
3yjCaVtDHBwTKpGIpF4/YG8TmuNsMzAmTFw/imdcPV+xEoREh6B4+thoPREISAVrOSMt/wOnsCA1
xJAcmDYxEKXsa3vOyUuptLD3JHaC7FmQyMrs7dLB5ZdszZCqVbDP1VpiTeaCRUYarXTV3mpA1W0F
uuqYN0reLlfixees0Tu1/jRGDE0iiL06Vl0XGm/mqO99XNNAJOTbrLcd09mcPP5x4Rk3uCpWmmOx
2Hgs54DWZH3t8DPZE7aOlOX77SALT/655F3pPfLZt5+Wuc15EX545QUGofI6/lvxHMhzSBRlrk9l
N//mP7xSgzPjTd2Vfe+RjtcYOeffL+YY+vDjJtQE3FtbPhU7UN0ihAIkLnwAOkiS1iG5R1wsU7dE
1KR6ONfYJ9LBHI+ewba4zRdysiqGZdpPMdosEdThH/my2h9mYEV9fWw78KhEhxsekfrsX1UKbDKV
Grn9bbnnYF+o4dQY2zFOWbk7EaGMl/9M5fr384cUo+j4UXc3epOatB34ovOfgAuq2Nft1ejN/K/c
bAs8RZWWWRKrNYyTXGwPu6aiLRgnMWLd89r/aqXTiPJ2lJXSPLAZW01i+QB+aOLqAy3cAyDHoXeW
5hoF8ljOdQD1vPNDv7isGqENPxlEWTHxGdSs0y2rdIgUWu1y4ryzvj9EUVaDqsNAsIVLhrxk0F7s
p3CAbzF3ljGb3wwIpn/yMnOR4lvyCReiGdu6nfWTgS0GBBUd6c8ym9dMgKoBUo1pk6Iv1IyCHMzu
h6jrdLVvmwaDadXyp5XwWrCJ1fJyiGlEw0N6zp6q3D5LIqT8TfhVz4dLv46ATzlXg9t185xLkyLD
J6ZSpK06y9+NT7g+xtetCHGwwWUFcvBaWNETYIlh9i1AKE5HYBGi3FMC9L/FiPx+W4KTkYqyuB8A
QkG6Rp5OPoDH3h7S7g28RYRTW93rnJexNvdmQkjefoL2DEPRWFhK2UPhR3bSENBuLi/SJJuGPryU
EG7wsh2rJ1V5MywLOki+t4QP/9hq6LyECWx3aqHHcccS/U7dnRc3CMbF7XlBXiVeGtFUCbflEWZp
rJIGdPZF9uTiR3U0TaFg/5/hXF9oBvCLeLiNLXCWsBzQZGubcvg/5hyZVSv67gm/CE8VsnNZETzh
vu1I0d3h6QScC7amauhKDWgXdbIFbzlcWRe3N3NL9nDjeVgsZtA7EfIu8V1+zZymW5HGW+gwjK4u
qOmrSAzusX+0u7Oj8GxCupiQnHvaVKVj5S5Stzd+4KfVXXdVlQbizIOrYTX6ShG7uWi9Vyw29CYk
OjkDyFJxIBHO5/fbfxte/jQilXgMKuM6DKqvQcsw+/CwIYR921A83PygWKju3SrYpYlHoskHd2oJ
pngHHMKLuOxM+7nv0PT9rndwi233tIvYV2eIhgfcBbb5gWqUaBCiKCfPceKHqt19TEE5YV8vj7yE
qS98y7pLKHc1mVaU66BPhh2QIEHxi0raR0IXYEIt/16Hb7W2fbprMCvnEbeLB1YmuuFvbCDsD4j6
tI3+hoUkDpsof+B1sUsG3tytUi80oWm1tJ3DPo06mIFqSMaxpikMOrywbL57ASt2lEb9E7Xp+z2U
iVXTGyREV83goimvVxgVEc1MWGwHgwjjl890ePrzzc70mvWVQ9FOqK/sixB+UUAyPT7JU0Z4K4iK
gJ7KbgI17hniXDAqwn43sS2rlz1xk+EBHcml+/0qEAVppxcv3ehW0X/NYieLh+O8MW06UXVre6Yb
07jTshCJx33CR0kmIew2JILMQY01nh1l8dj3z4diYpTECxKqr/h+h+uyKXZSO3sFFldDOgPCAbBK
LQua229kET4q8Y48tT8iCfevYh2vYANqSYc60cje3Gr8fj7BXR2bBfMfetaBjFkouJNVFwkZ3XBN
iHTT5t69hQl79AlALmnEg6hO99uGXuCjRa+DvoVpTvc8FhuQ6vslpVkxWvpcd9KaRwQz3YNjyp6M
wgVjZn/KvbDK2Sx8cs8l2fl7p1HaaOWEssHfMSEGH5yV4nhQ7aK3uSmguLi/3hXv++y6ajxoTJZE
eHNmBJF6ECFO/b6ESStUH26D99IB7TgvlDIaaMApODETUaHuyPk2Xm2+6a4OHayv0vvc46WWnXX4
c7XYFZfBylwcM2bvXPQTN8GUO4hLCGHa85AQAfKR6Id+kZp5DcV7TzXLsfQIuH1JTLFxOLrLWPtl
9bwyVp23wBw84jY9ozML/G50JFR06s18N9YV2kekcQEbo6S9CXF8NBcTrWMEyT7DGCytz+hDerpg
UeNtxl4GxUqM7fth5eoVDK4ubZ0WGhgY55B66RGmkPxrxzYGv6qaDUnUzO0heSpQLQLFSP8w7jYd
7KToO6XO7YUA5Z4KSJUXIIi6O08pX6OrPhHq3GLcY8XvZxC2iPhJ7f1llHgy4j4Ht+zWC4Ck/uqr
pYi7cH8jcIf6C+eUuSiVTHNko/MnyFh7kNRJ4RwEpACk/7rBz4yGJnttnMP6zXcDgxMsm4nlSSoO
d5el+IC8YxuSMVytlCP/99XLKOT6+9DLPQTnNv1YebhtEnM0JNqnRTj+p5UXCKl4KolVKeF8DD3q
vIQBjZ3HDnrVaIzh/7zLgakSim8YBS5TFnm2AutK/k4/Uya8bZQ+p8KTWJnBwYKtX1CKYQWgzq+s
mkplfwaBM0cJMbmRCt7sIaIAXTqmGKqzYOvwoMJ7q3scv20W/875pLm8SpnTsRyu1Ziu2WTB1lPl
qHZFLFXcNosXG4Mv7SNbKsuuEOyTNP1l7R67vYTEmMxe3iFnh/B3vWXcJfByBHNG2fXk0q6ZiBrf
0/MWHIHE4HnBLI5g21liINBPbuqYVEH5xtqhl9svW001ErQxCkkSITqoZWrxvVqzplvICJQqt/Sq
52Noz4Dt5z7iH551FxA9Ip/NLPvELsJAFqq0nvDgFjkjDqH0Y9dKLgpSBtbjKZZfMdBQ8YEj3IIj
+esnYgzzfyP6mT4mVD+gU9kKN8gVJSGRdKpnOLH/ifFCD+eRPO3XEehpiaeCDiZSm3fyoobkjl2B
G8P0AOuBq7eCzp33NhfFuoBtBuoD6Z7i6Xt72dZWVEyPr1GyZ5hvttdwD+GsYZ5Pf3Wmhjp51p/6
7bGJMeHzbQv1n+Ukv6uj6QvX7nEjAA2FLlhO6533qZZrijBoVgtI3n2WVsul9HMLwWBkBlCzfehh
uwejh6Cj/VmqW4yBEof6caInhE9KS4vcOYJ9xgAIVs1WOJX/nJQRyNunQEWaXWPrVpblJjEZOqOG
SHCoCKLC6Bs3+yTR9yEKPrB5rGfEXbYLFjj5v8k5AjHEasETtCIaIxq8vBTnErFor6UU3noT/892
JGgit1W9R/RnGP0BXL25O299EyRO9Ffc35KtBsbO3I88H5h1oiLpHtOYWk/BR2iQ+ujY1Yt4i+Mt
waK/+2Lzdec/JUN++ea4XCLOOzxehTqgD140GMF5GUGYa6u5h1VeYEUYaLu/NkAQPMvuCAm4Nhzq
1gzFpX6DUuQMGGFEmg2lKsi/pJCjJ4m2jkasq1CtVEAyAulHgGUp8Zk6Q6LzqIyBBTgvvoF8cIT3
+2mYtJBmRt81fUaZ9XL9vdP96fMwJwxQEpvb14wnIraxnEo6pHLZ/0t0s6GqjxY/3cmy0AGmY/ox
UegwQM0PUV7PBPCjPDYBTmfELio3oxH9uKfJbmz37uoNTlw9GP8KYTJvbZOFtBKN5MbL43dCvVBI
La85wTJIW0w3K6OKFbbh9TjhHLVD7BjSTBqaDsA91Gcsisdtf9F/5ej6pTTZFr2DZw6DtA4bfm8J
XRkWABVB+UOKdOmyUCPryG7Pc7RVF5oawOC1JfSCcB9xWc6mFtX7Lw1YZoMOF3TxsVbd8DTPKTCQ
JjrXlByLC8ndp0G8wAsbXtz+bfXxykffCX1wpIrSi2NCDmFyMffQuZQOJyLmYQnGadb4n8/tmy5R
2KvDNPL35NCWx0KT7Z/wIZG0J59+kgDwCrpTrUyYXvInvAUs+5/kN1nfhEhVuUjxCLEHhlkNUaAL
5qwRMW4Us4lGkBT/z5ywhdA9W76YsCBIO2pByXY5c396WW+mn2CVEzcuj/VUtqDThd1g68MmqWzk
FnVkbQG2mKpfBFsVkDUeG7UFDYyZYC7y3kZAl+BempbxCyN3LN4tRC1c+DFXP9Abpgqt9+i+Ici6
zYbsoF1ldJUGEIgYBkBkYc0pYEHfLH33t3G4g8gpXc8CPed91LEHqRABwhal8j2i6KHtd/e7rE5w
qYn/lMxhZ+JF13WO2EeQTXOTh3yJsTi52OrNyhapFNNZNZFXZZu8fdCWIxBD0C4AwRCMIg8l9bKc
E3C3gWBAlFqdTQIVx0rGER+LoO5e/JQGHnnqdIqlpKzWJT59fmLocs6ILbm1O7QH3M0KDceJCIWi
ofNzqVMc73MRPVlcNK7JANojoEABasxP6bZajCzkhkaK1iKrDkKdL4CcN5rYmBvBH/9XVVcy4rLQ
1AJ6ITssGghrGdpGulhiM4qVh1YkyN7HyAItg4QqhCDLrJSktGaLDXZlXm0MeAZeNpdYRzaQh+bF
uPdbv4Y9LNNPZHemPKr+Wt/r/1DzEmUDis/HHiGgnI2Z/oMllmPISlWzR/F9RrAIW4FigX8vRkrO
597z/aH0DTxg9UtG+F3IThZwpud6DpSKsACnMURX43qNuMPqf/mpxrDVwlYloGl/PtY/6dHJ4w4x
m1D7cW1RCfVxvOkizjp1XGeD24fWS5wp43IqgwwWm4g4JCYhsvKCY7ArggufbnbIAZu9tb0aCLe3
vSCc62h7nIvsv7w+Ue3f5Psu/ItBkzmKxV+0KN1JNkbQ8I8l5/c/HR5nFF6YH3YeSYZ4oHrpVi1i
xhz0J+vWfbBiEjPUlP62ltEnqa2BetaMSMfjDR+buoe+ZnO7KB8RjbuRlh8ioRgpjAzyoAj8Va8W
SVaUyoJDMm6/Lvpy3Hm2kKEQSo8o7/PF6jPEZLabyZNQgQn2gL+USJcOcet1f5yWI7bd81MFRePw
eAQGkLTwaCkEcC864rxH5CZNIc1EOhBHiIR/SFjEgPY/2iwmg8Q4AFOV/7KHD9C/9YxHqOFe78fM
rJXwviEXCfOUCZawTmPmHvGUgEIKZjNJwqqjWgWls+4CsVipG7u/sjHAQe9tl46SNypvp0nXHL4q
vK3XXv7d5tix/6qSheyOcGyJid5yrRxgzgMYdef/whwStp63iwyumYgy1NF0QpjNjPtxAAf8olyq
QX0zQEiXswWOPdkUzzHqFlTzgR+38PwcPfWrYxYKnaPCNXie6vCo1NDQDWF5LjjEgvZ2NHNm4WAS
YM/Bc2trczgMW6wrXb1tY2OUAKF9jw3fLC9cXplFXoElV00Ub1DF5Nu7DUACoVl+YXLeVbCbWVoK
EH0Mnua+AhjagYbbkG2rGnz9GcBI88ucRsuPYkbwtOQ8No79Yg8ywaEzUYTj50uVptN+Wduxn184
84UjU1/8KIhYVqSW8aBaSLiGkkYWbwzdWLAi5RNdTh1Q89CnLmlV0Rx8HgeFXtbP8bGqBmC/N2Me
VsUbww4JuYTchEn/LPBgdfqEd2IOXsnr3oo6DOiJI0zr62bJ8/Wa4rE8JmRq43Ive2G/xWd4YR1/
YOvl7Fm/fbj2CytmqSeAT4i8W3wkt5qAU42KPSk+wc0t3O/tjpQ2cU0h/g0v+dMx3Ny3d1LNr43e
TyWQ/j3kMTJiw7pR7urXWXKcNvHBETYHS2IdEsOAo69TpDWe6aqUPldnqAoq1JqMqyoRh6f0A1kL
CpYMq5dsBt2vSVoltHhidLkVQAdzByeRh8Qkp+PJ9i37L6HsTJfwAg7RVWw3b5+639tqfUurQWRf
Mp5ZmP1WOrps8QP9HR5lKp0sCbOq71d2a14eZoJyxmX25ASS0y7TvYR1iDpjaMYyQZSFqcFcSGjX
hySHike22EuQdF4yaLZGE4oOP9iSPQcM/PGzo3U8Aaz+pFHuziSSOmUykufDf/1HJ7MsSHwONi8k
riW1ZazbxKXh6ejAK5cnokqrrqPV3anFToVm1CWkkoW6J6yqWnWemIQYx+UTvTOAkidRr1D+RZ2V
cVcSGOmRiwG+raRiXq07/wC+jkTNnLav1kUrm3M9a5Yq2LEykdkB0CjkCTn74Wy2SBD3ulRVQ/6C
zGnwoHXPYRoCWE73rsvpD4h7W5s+Xrk8pXl141YHBXIkndlWziZGr8qhJCs4p7Vf56zB6YXn6NGw
yOXsFADo40WLQbiOnINXZgkAZlezMfZdR9hUdBDLJhW8cbBpQKgLb2gQ4iWgTFVudOVZbKVIjvGp
4Jch17ksoS5o3lzQf6rHSS1hUSw01q/qe4DS+eZnAuGuGuHdSsePlX4cPrwu/6HGz2/DncjaxU6P
HEXj9t4+dyQ19jKdZfp1Gq2WjtzMrCdLjkqujG6ehxVI2uYQfpIx5EC7L0qt4aURg/5/Ju1AE/FN
UcHoIaZ3Jwpra3KLBe/QnWwmpq5NJjyqkAEs5wBnh2CKgu044EHksa3EvM8c59Hykyg7c28yFj9m
Siaiz1IKY+3HKzRFXQVCEKxHPPqW3lQ4Hsb0WLxkv5IH7z91WIyVk9xZxOFBh+5gAyaIEiwQj7o1
YCOjihkyBEai8fTzsbtLWkk/HMKVjX3SgvwjHy+oRKGuEx56jvsR/aLcX6sHXsvbMdI7IqmK0Fw1
+OxaP+OJsUReclr87nZ0e6MWnDJDOuGOH3Xns7h6V1Ng6WSXAZBDWxsWEIV0cu8tUyT39KbG8C8l
M+GDdI5ZKMaHp0kYlrFnjt2qlwZJIQzEXPcTHunNwMgW2oYeQXHpNnqIfPSmyp+vNg1c5+QOGtH7
SNhs3rS15hfcuq7LL0wu7dE6/xcWPgxoN67Cde7h8BEBO8PDgQI37PA1T7b7MBAVrlzZSvps8t/A
mLWo+AfxQRDHbbqeUgvT9SSCvNqZzbgTEh7wpJXoiCbO67q4gM2LhuD9qu6JFYzmDOQb9fU9hDoA
6Utx3taWQLAQh9A2fcn+Tq4UBHrfTtkbkK0cPwpi3bZCsP6nuF7sKeaOsq76szWM1fFskctPgHgW
hNaVPUQQojeGMFf/OuBtxZtchAmimbLTYXTNbwvz0MYTIDF0OY+eSakedpu0OLYQgENTHtYPJ03I
wPWB0Gmb7+sS26JfIJU6xX3UIfolRm8NUAIfApGW8wD9k4LjUZ2kUnOtZsjl875LBRiv8XvJbZys
9aluW2avgjJP/yZ3Yl1BypTUL9bps4+/6FC7YFd3EqufM1OWRDbWEodJmpjZ+my7/DoYPskTLwGL
K4o7ziks1Jg/A/3CQK6gSI8AmeEeUXC8rhcOqrVzo7aaGOkr0ZW2AJAGhzO52HdNcBuyXN8P3B93
S+2ATRR5H01LEmAne1P6AF/e6TOrTEQyFTG7AMf2l4PjD2BnacLzKLvxHfz8fN5HiR8Q+mbHVNQr
HnAvpyihlCxlCY3gq9c9TMB/RXe+I2I+FmQQ53w033zEPVUWYXm3E1iwyJe6PHI4DZjxEocuoGeE
Qimr++Mhsy5MiJnM16FtTD2Gx9o1E3WVASO0F0g7jOLgjy7ZqQSFKn1oCjuO1ooE7+d74Dab6oqb
Ig9ufy+IdO8pHDJZjy6fnNjtAUcu7F4nvbbx7AqIVIef89GP3ExIIbB5hhFQ6jm+D4z/yxaP5B0V
1rLY87FOxMjNZ1LNqBETx6LZNJSuJUvkOY4fk8rDsWizxV8LyfBrlyivB9SQHPnaJ5l/GvvDuoZP
8xWkLvfry7gZ+rCIiyhFwRhRQsQJspsKLWsZh1m9+6qQXisdptLymUDPKc/vl/Nxbtdcm++z5A+b
cfX4kIb6m10/9TcHvJWwicT+WowUmT044JqCQ/lohoUSeEQ68lb91yf2eX4b0mSmPHNSo8ajxbjn
rf0nYQluspogPZ69BKeMYQS57ej8LMAvQJ5S+UIjToeCBL/xd+HdtAo/KSRlKNZYbAyp+8fHr6Kp
Iu0Pnr4TxI4AkyanA2/FGIM1Sgx8oa8oIpG461txFoMKj/voXAZP42GI9fsFfWc2jRbdFOmT9j+y
J7lFEe21PVEVxS5HWcAjxsqWnaK4dkjqdqH8dpeMe2pMHhfsaUaU4Zo1235R+tSYY2BHmd4HB5Bu
QJXBXD4tZHrv/zwgQw2budkENuCet+17mNzxKu0vjyf9+fEVwGBHZUO5Ru+wBM3RxMPwuA/QMO+Q
QWtnHrOC1yv3IEZ3eI5k55xXOKYWAtbT6FQcAH3xK9b1WZIjqziHjAs3HpxfI0NFKAxfacbADMS5
Yv7gxh4VkB4gRRBk+AzwkTi/MV1BeFuOpvsJmtk4/i9IyaYWys/OE4rFnCd+1NOkI6cat93coovk
9/SElgkAkYPMNWK5+iJZI1FRSand22IWRDM/hyZuliHJDhrmX/8yF+fSw5LhqzU2NYG2wnOhVG7+
i7maXVq3bZeh6lkvOzU3weUY7HGbt3fn+NmbligeaNKKPUHU8zhbYguNY+51udp0rHsTnsSHFU24
vKQH1ld8a/FYYQ3+7ciOgzokxc1IiMEJokdxl44KNv+wKuWez+EXvcPQJb7inHLclPghOQU26PMW
f/2OzpxS+KnE6XUXrrZ3RECFJsDfRQh9KpNdn2try0p8AjxhuM0yh4jr8ojIaXKfxeapuIQ+67Zr
Y5U+aJrb1Y/h5TjADpJErhhMmidCOUahWdl8BMqXN+0fx2TWgvq74FGG1k5gb76xfNBUWp0RC0Vc
6MFDhYJjZCNzT9AaPMy6LtHoERpXQsZduhCVLTw4kGNl3k+IhygReDqFwsphZEflGi8DQxZrKdlN
2qKBN/H6L+30Z+FqVx/YLLk6c1odbn911B5YyEpCdf8VxIa8SaDtpRVuMTZ8lyr/8kwCp1O7ft8D
uTk0DRfRv7BaGuvXPAnL7d6eLqpWNvDGwxsQdf/XZk4wRNUsrYrY2+EHm9zlGB4UYJ1FWKJKk6kp
UAMuY2eVklICTURa+8geIr81wrsr9HziWTvhUsDs2fkX4Ej+uNqxE3iaZOSmywGiitm/Jsihas4/
BF5WdltoaYQcVOCDgOAk17bP8pgvYc2wNCyO5s7Unw5ogo6XuOnlvDExyYQaOKOt1dDZXOif1lxD
5hxHkF/ZgtnSkzgSU/Oci/q3crlpskkf1F5Hd0bYLbRRNaLS4BX8Gl2E+z82LrGlaMKjjn9A839e
9YkvwFlx4BmjH1e5IAk97P8LbUVeFLb6cHr6SlqrG8J3HQYaloRO6hAaiUkuoSfHlcW2OCYr77kS
4CaGzmadS6j8TY6doUREA8EvvJulLdWqg+5B1JnQn187BoFbzaiyIf4z0S0sebzsd4DOM4oFL4Ie
1xWScf+0YFgC1YFoJKaq8yWfQJ9NgEIcahqlDQgv82kHXFAQJ2ha4Euf5PCE7GVs3giiW1zAsi98
x9bvbef6DjJzqLhs5XQxIGB0KuHzrwhlkI34VRvdBU/ozX7btLNkIMjfHmw9/4JnnwTXO/BC0wzK
oi6iVfdNYMKotJyhmcvaC3dpgZkhUafRMaFe3ch3FCrORrCEDwRKc9EeFdmYqjiao8oClk8cOIMO
4/6LX0W4gyqp7kBsWipWvIMZVYLkGLJsCgvjI/wNvOBm+EjCLgnWEIM16hX18uRj5Z2alTyj7r2S
nFAM1Pt04XUa86J9J7U2L14bVjpOr6FiqA/oKey4T1VwMeYWTamB5PuKLM1+j7DboBbxkKYnBc2a
KXKGY8xl5o8mtOHVh2NnvSSYa329CcVZXaB8b6ng/jAQ7WwGm5cp2Q7ZumZHTz8iBA+LH1zJulgU
dvMufoP45Rx8PCqje+IqB00kMwmEp3u272OzIrEtdokDG/oF2bWooTHol9HZkPsjOZegsoryw2Ul
hm3bcD37QZc4hSXmgAXKxKIKlFkog4LpZxL2OUGB0A6fdXKWW0T4SRa1aW5ZinCLpqpIEXIqQqfg
H9sWLmPCM+bxr3rhtX8p7ILJhBo8UHjB+pVM/LH+hkYEz8k7hyETGICOP+HwXWRZcBb4901JpX7Z
GsE9njKuknCC1dM8vDuanB6f9ImISt3TwuB60rLW2JgQIofC3+Y6uUn2cngyM5NR/Z0gGIIBQ4tQ
CDly9k0A7fZ+Ae1YcUvFt+NoEE7OqpiG4oXKBgeNfasC028iJhP7FYiFe+6ts+MSY7awPeCyEtTW
MHAM+IfVAm2HkQvjA7l5Q4T7OL/1eDiQ2JpGXYYKSqbedUgTF4/4Pmr1eDD6YuCs2piuNfJCGVQN
8Aik/+PlhUok9y1y+gdTe7kOoB3ZNWvIvpdvFHt785t0VjC+laiiq3+piE4UErPkTl0LQ7CJWNWB
T8sJ7NKeuL/aFpMtldcZYLSo1MpQGO1G8lSECbizBChe9VnZwK+UgAXrJ8zIMF7HpPqlZJunNKeB
k83aDJDaPdH4Ob/r+nbdvOdVeOK67fO5PC4FexC7X234q/FrXTQcY9GAkVxiZdh9ZcyAr6ER66Nd
b+jEgBcy5c50wldr2yXtJISrKj+muDnWRuOj94fKozRJwlpM3AAuH6V/UkrHdRSx8yloNd0+pnhN
DVo7o/xts1Dwz6+pibSWiZL2FN5QrWfhyI0l3SqfdElCVoSt6GmAngaE14dyjJnTBIzpHOnFXCqE
Ohyc9gk/EItW2W/dw18AsysE6lQlN7ZCm1Hg//SnUNKBhQQpqHrzwCJsflLiLHVKUGx+UasVoJcy
XAKy5FliiNTLyA8NakiLtH6JAdG2FO2sjHnzl8Hz2CBbhuzZZy3ZrDtWGIJ39Tm+B8doNN6Q1Clp
RGPiJmMwymXA0l/VMlGRBi2a62D9pcr8+/zKrekBovEdDMofo48WTExUtXEVO/cdeO09LDhuDxzL
EpF8vMbEaCnTk36hO1TzKUYmtTruitg+7pSAGyNVE2tFiRVIpHqWeGNAqMcxIhwupVQSW24sD4HY
csuG1gw21kF4WNOwehLJzdPPeSYNmxvAZ/yuWHfkjfdbAF+6LT5z3PEDFp3+bTrRCi21JituKJNr
+YmTIOag0ty2bN4aoE9jv5UCekSb8vyuZt6KCclbj56qOYXJsy4R91VhFLUi7YzaFyWneGy4gviX
LL52/5G/5H3c86FAdjyIkoXBVkC41wdV7FIARbz5ssBXsutkZBcE/GMw2a3a8tmfWk4OGT0c3sot
byGTfytuxloa0EW9sI0NFKHeNRQtMH1Ag3jmKfLd+cNDcc5xg5vVdKsmCt496wqFerLOL3177jCR
AmSiDfOgjbRQxvCwmRAVYn73iKOToUIl6Gh2Gxc09lthtgan738P5ZDxcNV/hqlH+uKQ2zXRBjcs
IkWSfUJdeLJOXHxAi7xJFdvbfeMDP6ALdylC5UvrGpRP+j1z5iARq6RDccNDrgyL/qoEI8lTtiYv
Kepd5mSFyQ9Zz2UKNxVnidj4LWFPUYpTi080EVTHoec5ZQ4nEM6LjUpQ1+z07utIkMRJFIESJ5a2
F9UgejQointQ/Qq+E/kyjo5ifWpup/CEdUTpne4tkpgE2qZENyiyWU/Lq3/HtUun15YD42Ola+fa
JT7vXe+EOjv/3nMSV0wHruV3UUNtq9fyuuKr0DZvHVIn6bpSfW8Vh3BFujYM7UBt+m1/Bt1JAFCd
oPmbf8KINzTC/nb7iC8+2A8Wh+yMQM6o1NlnmVXP+DQ6ffxM4u/X+iOu4vOFeU6IyoSS02ZJBVMb
IBEcOx9vdq+Vnh9QLv7IkD31OTtbGMfmww0GfYpPB0yWDxH12g0R76cXQY34FNyq0WvbkCrpj0N6
SmvSB6C56SbgtzYXFoOT4gmrxiT6XfflE4lMz4NI9SXsyxzYmSiaVqwTZgQAV+Varr+wxnq5KSkk
r0LvNsybTtXv4PKP4lbLm3cWgTt0d2dxFK+vf8Kj4UkDlM5kro/SMvFrTw8/FUWVuBBAtyG19uhq
/osdTqohaKmJweqid4Vmn8bybHSpYx3V5JOggLoQqgenTbCzt2dANB5C7lk1RsevjaL44Emk1JPm
AleWwZbBb6u6dxhcxbSvo/ofJ6a3FUUm9dBVA3TcfjiMoceU6uIr4IYQcQeYUsca4a6aCQzvVojn
bZXzxO1A/fM9Ru3ElWjBafuWgFIuYCPxhmJNC0FpmB8+GeHgdF9KtfjogT4LnfNKK9npWid2FVwt
l045f6BVY7U9l0cEAU5csKmUVDTZuGa4iD9WDXbJT7mUlckfisxgvF4r9kgcRhhjT6RbeHKhll5N
rizdNZKIK8W2wYAd7LanjRL0+CKjJ6YX0qzepCQjHF+lqjMQHEl2xdHeZMjyei039x4hmMMJa2ry
4qXiDoP5CuHkEgFYbFJeovHhQzRRTguM1qae77jh16z/MqteERzzH/b0Cn/a6C6lmiv2SX3pxbTU
rwTK8BH5YVWKwvfViGzA70TQfuFdt4vR5qbOsM35T5E3uVUGOxf/VB0cuU9N2I1r0bNeVH4GCLZx
Q7xu19UWLtuOYocQiDZ20k9VGpV17h7DmDkAnEkgn36yM3VY2UnVgZbj0WQ+Fn5Fk4iLuASjN9NR
liNQ7T0NjFrs7LUUMyvBAr+NVSe1iB0CDiH5JkHCs+y4MSgP9BKr5U79kEnwozVPDBobV4wO6JLN
ufbl1mft/tEaKczreE6Gl3UlL2na4aPCpmwVfw8nvLv5fKApABuYbERRYo/z3pvmRMvsajbdW9+P
dxfV4cp6L1PIYBLxyH9Stpv1CtS+vZdbRrPCYRED3KTn6try0ifOiXg9cZd2EajdCgQPfbKV+CoB
NAZ3eAmr6Lf/Y4c9GHSh7D+gV5ErT5YgjfJeSqKKitwUba5XLplCPQtXH2U/gmxTX/Mx82rio6W/
bPSRVXvsWjMoVSjrZm9b4IlIrI7n+2vAgCIXVebPImDrzqKYAYpYZQatvZnPlSCwWoafTAvUBEf4
ue7YNLgmPPGEoAp8iLU7L+ce8l34usIXspvrv0b+l5BN9kTokjSQFx1cFxU0hPoNTkiMBOFBjXIc
DfA7ozXo7EWm0/CnKiMmNgfytQujNbcU0b6TQA6S4PxfCwoy184ZD3yk8DGGKgWnd8hRUcB1gwgX
Ma2pGI7O0+DLGqnBUsc3p2ldTeiio3ox5GUQTRjbxqeCYhAfq6Bd3T0h9Kda30bV1PpEF0Tfzslz
XmqovMVhqt5DXHKUpCxwR+iX2NF7Y3BPt5nh0Y8twyfaVcJH5YloP6nQdXf0OLkTS/RMV+oir4v+
ifYvaBNzfKa2yBRpz1msnixErq+7wWnB6i/ThJznt0Sm5oRj1BKQFJnD/Qhs3w+nIFw23l6PKnlc
wyvCf2usv5TZ1RI80xpg1Bco0qxRcoOOjoF4SK8W1/LiRSUMP615NTVAEIiuxtRQ02Mz/2ghFscD
sIEAyXrpthB+erkJz0uTI3aoFO18jmd1JRiB/IZuVbqXr5ZpnB07dsd/a6UTxS0eYrQgtuPlK9ej
qAjVp4X46XmmFiVaW7oQ4MFtruNiKk2l/vIryL0heGagONdwFac4gpJZl00A0+h08PF/8e6T4gNe
EfVR6MMPseRMbksKCrGIHNF77dWXYght8hzmtpu3v8wWxNLSaAVyCKcYVRH1KcjrR56oDcjBAnfI
l1dCburXUcexOn+8T1h1pBkXrJ4FOrS8v/Z5B4n7p7ytbrsTBnar7LcAC5VgFHVk4OXilW+18OCb
t67cIwSBOsR1pQwl2gYfPvhkNDmfCnYUqi7tCZGY13u9DdwndiM/jYI9MbbC4wcUgeVBB7yC2J3D
HQb8wVK8r/KqkVuNhqGJgY3a5RiBaH8R5K66q6bxsVmfnpjDIkHT6A7YDPYtna8rwo1gx/2pty3F
R5QELtJaAkKNMv4lywat1oaQcfvoPUwm+Gk4jtPU3IjASOCBBzuKd8dTOZ7pz9LKAyI0PD8ZJ/Vb
9ZZEBCm3R3zw9NDtCdoPjNuGoABJ4osCl9sIIjM+MhICE2o58XKfeq+veHGD33E8tW4Ps7BN3n2C
u3LC+WV+K92nxs23ZqlmTWM9tu/aI12tAm+tn6/EPBrjdR5nT/n50KX5NA7EZjOS/7Qjv/kWfOZD
OIZwzE85+4jSQZ/ccgeJdCDyVx0sZAEQUbeffcA+/3SjhNQbYzkMFbLt12IkI22OrE5KIvt9pf00
BrnAf/AO6mMpWyge+c9hTQWrefYkXq4yZPkEsx4jUrL3hG7906+/JoCabOvb1IyzX1ruvqpn6zuv
XSZqRzbRyr0quBiQVX4q1tfTDhSRADzT9qttIs/KEzGZbPW6gSb5lnAVE9bPC0rug4Drzk+cZAQu
az/Ef0y8qGJ0GwH4FFNytCD3Gs1WFLDIUGo4TVxa4rXnZTqselH+usUAcjvWs40kLJBdeNNmJ8u6
J1VBWQCrqqnl0GXZQdyqu5HCIDXel6xlQMkzPIsRn5NijYu0ghwOAwbemRCXw0c2T9Mz4A4vm3BS
vigb3qhWkQyv6LpsM9C6kv195sPTFTOIVBJlYGtZhi5aEgPkeyBv7em18xoEyXLwbzIUQ4hhu4ls
JOzTP0fAc4QpbmQms/6zdc/SiCOga38reoeY8zDv4ZoZXMa3o3U4kzOKReRJ09x4/WSuZ39C55KK
+w/XVlblK2feTKSgLO45iNt1jnnw652gqPUMhOOFDEGLe6QJNdLsaY4pZWRYP8CJeBZOjGNjXNIz
yN1+ySI+U6Oz0jjFzxQ/kclkKkqxeq5HXZC8R1cBDPoM8JUZfeUBQyCzWue9BWTbQ7jHoJtPkY5X
FptFBFrywMyqv9VrlV/9P2rdaPoiHRoKDHXE45pUdG9o5AQKPn6sONWf7ZDbzBK6BehGH7wcb5v8
QjlvBk1SSNPT2gh3RTSun0ySk3ZnQm6Q47wOvV14ElvzzoBUA6N+vjcm2UKokQj6GOP3me6Ocn8Q
7B+8mqUUwbVALfPSSe8BBgghS39HbsIeF/wDrPdySXpBGlA+dIJ3BAS86imRnnmsD4dft2azkSUg
WuVuHK2Oct/1PfjclDwzFTBZmNb5SVJmN0s580nPPENdZoNz79UgMheaOvbrMb9Q5ROf1+8dN4o2
7bJBAdOfPOmnQ7RtVqxmTj/Pa3+hbuXR+zX7kDkJqiYnuebITajPPi8CXabGScxChnhMxmYP7iHE
9H/JvFA7ibhiXjdn9UQoQ3ePoGpHmPONoRlticjNQTnSjS/2cZB1hSVqYcfdYBWLZQ3IAtatTi4f
/ZKZkmRkOXVHGhQtxHwEjS7/YYEp6sLTrpIMqBd7/loTMqQX7iPfqn1NLn8825zxPCRUscW+/1fx
RmNpiA9A7Qa+cErN43msXxJsPjXaQ6FiF1IAXEct0QXPfal43K5GvD9xjKVzvtoY66GfHdiHVKgA
aWVjTKXZt/UqqepqLwZONasSfoXBMtINEp61jpupD/GvrCsvjCl5vpgg/pBOEaf2oqMNhkMAa+eP
8UPcBu9/EF6AremDyXZEsr9g73Eu6RJoX0kI3FwuFBAs+7fII/uoevp+eu5pUg5ibkskM/LU0yCd
6TD53lV/wd6wNlzDcwOxoScP17DmGR7rUznZT5d0L5Wr2XY++yMyhvUjNb77AgWG9gaNMX3aBJUL
eI//faagOg7kGbD/sJN1qZB7ppSNcfeC7FcJnsj240Y6vZerLYQ6hQPnA05vc3BCv6BhOpIvJLK4
ne7tt6wUKx49H65P3ta8oZDD4csKsc6sZyePiTkjWO/W+O+Tgv1jQtMfNQdo1lZ9wG4xszr7YGtx
6elrcu5LQDoYGNf3zH+Da3qAO+QilIBRqlGKj9vK4FN4hHqYGg9hNNEq6pxcG8kbMa39fKODRoRp
y/a9oa5f6IKE+m0w8rTktImmHWVuDgmdi/J6HvJTrMpcsJuUG2FRlPAtraOk+Blt+LrvkTmaQ49P
r2mDnsnNCSlHEus7cknHG9O98RA8Ujmf5XWTz9AdPPZUnhI9emb6qjz6TSf5FoMyCZ9kF1RhLeeZ
aMTZ2dLGvNEAfss2GPqVySWpfMsTc2eQWlcFNFgBZf9xsjTHY89U8ghF7AfrRM02LmdjJ9Yf63gJ
jf8I1iEObQkzueBjSJfYwK5oLm/MJj0bVh9m5o7GRSNr0tKl3QeAiuSoYETnLxiMmQk47KrkUwP1
6boPafScciHuguRyfPiJsRM+ysQgux+M0O3LuowLUTSTHc93rnvYGyzQ5zt6oIOCuVNmvFT6ZUrB
Sw0iclZ75WsDrbMZNFBmLWdp2/rezvZ6RYIIYRMEZ9WZKXjLhTzqDD36Nwql6N92aM3gPyPhGhFJ
qNdbZshfpCHjUX290eFwwFT3gsXShKxpqUH/fmd3Y8ByvGzQqone5IvBskup6UFIoUqfu0IGFygH
gXb1bw3aTgKo/VD4uPe8jAjeoqYkrzhsnUC+uGQNXiInjPxx6odYilHW43a+qRjNpk9Al5ZPo2jT
5CPXcvMYY3zS0CzfmpIrlBXpx16m6XXRiWRqUOVLGFhUmjKttwn5s0YEQrpDsSk+d0y+0J1mA8UZ
hpYT67boDx4VFxCPRRKMxbfcZNBC6i5OwuLYSx1bULJuSTP4GWhVOLzeTS7vv/GBR+WccMHxFdnY
7x08I9qk1q1Fd0MWbl7+j6vUAUvrq7WhbxoEoOgrWCvNi1wTpIKeZrSOQ4UDcmTUdBm9UCLKJsK0
0VYzL4fPOrrGD3yrK4uOEDPAxieOxsqH8aEzz/FaRawK4/EvldnYaxaIcVenmD7qK1eEmMuqg88p
VEZ4mswgrDdWDDo08biMrppFAfDr9s+lPKbE0DdwiXekaXo3kAXK/IUy05jSXwHsns0/o4wDvPt1
29wOrAasG+4vPQ7TuN58ujmkjBdcbk9tF/IKqPuDZl8c74ku+RVvtYYKyRAVBDoyj57UnWxShmbk
uC0Mq40gYkqDx9wrisMwxfGcpO9Ft5wVOB4SdgQgOPAgCsseO64q3hssuBvWaBRRGLtbWPS1NKzE
2zJ1iO8XDAmL3zbup4xW+FyB+tcnfJ26xY/Ud/7l1w4KqwS9NLNM15ikNTIuuko3/Uam+jawCtqR
06bRAUWiFRRYi/LEgtnFisGFuOL74I09MmzwISerqQQISoAWybKYDI3J8IJlInkbuk5jnK6koub4
CIK5ih+XpNKsZzP2lbl/sLgko4RQZQLjG93B7oQjEZNl8isTkrWDhVuXmKwN/VUmbaSCx4FLx1Q9
FOm3NA4gzDnT8jRtcB3dFdLqteNwBXU4ZQrlddJvqli54SA2Ws1es7Nj6dT/BJA1qFLzFpka+fBw
HateaF94e8LodvsJYMft/swjiti3DmlY2uSjoF6zoN6eQmWzYq9gxuJwR/MA88AJF/Skd9d5XZ9f
aJeW0Ob9Qn0sEF1ntOnY5bjPG0WOiKZSYiupEkTHDpZfVWu2qxxMQmgYSrLIicQFPvnZBHkjggYc
ifYzYGmt/h/8sDakqJxj1N30PzscSSeug+D/GHmw39aHsxqT9M7Dy96eoWTYFYmYnaCFQhfT2J/S
rKz1HwlokC3iWGkFG1/1US4zYlpV7WN0/Z6a73Q7fMll2Gx5g2WrqSMUG20aecVhP5DExYqCb06U
R7RazfRmvH/EEBJ/gsR+qAzNZM1l1XWajpRTb92fJ7ooSTymsXHO//7yHpzthmJ1SXLdIHgxN0JE
11f/hKosEWOg4HShy/GZ+0JEen5wqTHjmXsP9i4XT/VRM/j5I6I/HYZ2TJFAMoYYx0r1dkWnoQue
Z2dHDYlcGaXdMceA2dLjpUZ5KhNfulbV6btui2ysKdhF/JVgExpZB0sTxXCgHz2a7JJxngoasWpE
1bfRymuJC5iDAAfHxquVokn0YSXuOxl2pga/k4rYt+Hz3n/odBaO0gF3LFF5Xas+m2bBCLevGuQt
cSAorlM6GHug/7YTl6F+jC4ZI1pLOx31sPGAv0fiVVexByBL94TLbIcLG9fwy0/yzitO+8GCL3JL
ThgXfjC4boThIMJ/kL/R9veP6zmGJM/TDxtMccfHwlueHOrX1+XXUR9JeCmriv2zaPglV/FzyYre
gHsSBlLKnS2wsYnVNg+VP/DV49RKa+1tEtPN5VVhJgOkvECMA8otWhn0wPRlGS7tN55U0HTKh+vv
nGZ0/yTNIJxb5W4WMIDfZy1TMVmsNNjAgBWvA7i4Z1Wxiq+RB3S7K1quQ1LsnkU9X7+HXspnvLMu
qHyfHNgYqyQ3KOfNpS4YUr5wdVLl6/VvEop55FpmgmVz42UW7YleTZ+ttsLyHXwOeLEGB3GwU2G0
HHV9LNdTct2X3m1lM4BRBGpSn9/xHk2kmIFnjx+slT8zZvg4aPCTOUvQTBEMjHrLIqM1Zro8Mgpu
CbIEniJw9LKm5zswT+EdKSAyGHa02OnqugKlBN0ALJdTgPaiewsGmesM/ctZTfQDy72suTJ390b5
ITVqtWk5YK+nr/wPTl4sKnpGnFBHP/kQDrhtJM5STrpNWwp/9RJIqHZ4N/QOheM2r8+yhS0Q21bt
EsRsPsdaL/79eicyOrvNzcHipycYYbR255J2MDSpr/bIprA8OIRGlQ6bYBe6bNStahXSpEPu1eyF
W65Ho2EtcD//8HVcKoX3en+I2A+R7Qm18YoKTtEi6d814gPj01pRntarngF0pY8S8E+WMJK2c+w/
uTUk5WjV6DCCmw94rGVVCM4q50i4rV43HS7Rr6IiUhDkYwO22tfj21Be0lcFj+57WKTQj6iqs1UP
ECVGNbj6uaYR4fh4gsMwmdPYWs4Zt+gWTr2ZU77qwch6+yisC+UWHbI6KGod09vU9qdL84f5B3EC
8WF5GD95wE3m72jHOumIpNCakO0QvAW/TOG5LYBLgaBTbiTwQ55qCanEpoHuIo/5pPiojx/60W1b
c0enZCjUF7nTzq3hkrenlXh3FvaxCZ0/Br5TFp6/J5r7FDNNMWMGOtdnV/Aaeqot5GQ1W3Nq1mV1
ZnKDAhc9B7bT49ifDiFUMNf4Xv2vIoEpOEhBMAi+vsxROTMSi/DejnUsfn7FAa/wBbfAN7nWm2g+
nc5/15TwkGlk8jj9FLhNpNdfmpenmYfPqcM+TtkNYr+BQgGukRnF1IPZi1FQ/Pe5RmwCmjOg33t3
s951Q+66ikLiyR36wHTlu4Tixm67TfgAXg/vO8UI5HMFkSy2O6vBQsCnEktPuCwmdKne1JUSm1s7
7/R8A4RCUCcPKJgg/YSQqTPmm2RuW7zi/WQ4zLNOWJO5BHLQIzwGGijs9xDNsG4OUarAX/OVH1DH
9CTrHVaP6hyUeZS6kpWJyfDJ2NnS9Z7IIl2ffrou8ssxOCVbGeuYLaioxQfoc8OR64Bj9jsiUPVa
/ONJ3e9yB8GwK5KF9qB9JFfAzcwm4o2ku0yCg9+yNFhbw1PhPSgaWmx2fXfymeMETzJDgAh3pF6Z
8XWXKASo0Y298nqhFnEBcrx25dLNPv1rpO0YXdSAWJm8ZbGy97uKHoc7ez53n4wc5+gKnmu8SHcG
pWyyopHCOdit8lfuWi8GSMeuC8MTvdcaT0I7gdzvtGD1gmh46xQ3Y924GiJEu0E4CudtTc04e4zS
mv9jAOELCPkx/Yj058GKZMYqUl1Bu6zSLwQ1rV9n4PeTbhGL7LQEr2qlITg/znUv/ORGnKIyqqIC
q/nrx1jGVgJUkCZHb4J+u8n6VyfuK0bZ5Ya5FbojB5cwzIP9E5gmUc7GFm2rp9mysJ5ect8BVw36
nVjXP0sR/Bbt22j4SR0mBGUH9JyIYqKO1E7OiCFVxGcJXXVQIuwvYLytr/XP4t2XEJ6TIPZrYi7A
+bMErmDnxCSVUPEngeWyziBnaTw3F0htZGppU+dZxM9yd62bBqalYZ6dZhAqASf5UVjxpCn+bCwj
MieOP8YqYNll89mVJVqFZKF1mlZWsvzqxTKPbsgKgJHRtgsm2/QxlB9HpzCl79KtoZ7Tk8B8po8j
FuByf/j1vlyaBky5wPeWTLFqHhJh/KAi3cgZg8Fou4mt+Ikgavo3ntNiX0YEVhWU9ckeyCzqXcJN
3owXUdpDHzLzp6VfK4Jg7/xN3a/jQIIUqRMX81QWs2gxT/jatcLqUICeunlMcHSlZ3HbqFO/vZSY
2s+liQHNWDNTShYfpllDYU8mLjYTU0oeN208QBUdwWWJmDCiY3WY3qamsA5ayZBdvGYVx22j71Y5
6FEU+V3n8YvCcdwvCJY5Ih9OxDdgORyNMOfqRRjVT6SB8f752r1fh43KDqM67i6s+PbA29ZohmFr
ACw55y8LYpCXm5C0N3lm9InHj5F0tbVvZnrMwh/32ey1nxhUDBWDfxJCnhwhofHYm+QirzWur7u7
OPUmNfytEAQb3zMM3urAsokuWiJf2WMKabsSMnaeMzNBb3SDDDwy/4SKa/yX21e21or9E8ANZV4h
jjNDWCKBIx4xcv315NuE7Eg+ZY5CQQ96MfUgCqxfeou/UZAr5wtLBlpITP0OaxypQtWcGZzhZ+04
2PK5oBzJkGEydi4ng8f99XC0+2rFlcylt5pcjZrCca12oKHtnXKLnTl/KcSzSs5TmTLoibDi05Tt
hWu10tZTgZclv945DWQqYpldMYYr/AFq1BeJ0B7iatYgsRy2FSZaahLJQ8sIZ42MFEVmHrkS53hl
xJoesL5pIVMfNyjcEXnMsM+hnXFjZHcgieIM+coSXAoCRDvUmDj9oL2SQuoS6iir89fXiHgbRAys
aiHwpeLlFfIAgyPcd/g5pwjddkCYHXByAhd5J7F79Z7VDF9m3l1Ezq+LaiApxH9Ql7zVNpBGNMRK
nEG6/c+r7j24OMs3BCDdYsoB7AIIRx+oId/Rcq6IK775cMrNpvLkgiCFKh9WCiLeHm5HQXH2kPDK
xZsgYZtobY2GKVzHyqNEhNohe3J7zw6OoL+zoxPwngzx0SN3jrfoP4aPQJZMlnKrMrA6OsSms/ey
+IqHvsn/vWjYClj5jH5q3AbXrj53XaFK9Jv+dI8LEpqwF/zt2pxC3YMKiypXEe0OuomYByQlhzei
jglOrms+DJbZSJMX/4y18WLtNisA9/o9G5MRhViHeQn7Z7zBhT9ck8nXvctJsswj77aW5+xdN/0s
gYMi5X1zMzBIUPxoGVF2wxaqC8zoSB/8Qiz17R1VwYqmYE7sdrF84KiVscs6X3Kmque2xWB5Yh78
4fz9dVcdpow5bwdRLk4AQbtmdD6qs9ne0yIiKH5jfdf2eU0mM/DnEcMmWyVBchHLClL5nmymQb2L
SQh5beSQBnIY+6ahr79Es57TeYmqhZ2eZRgn3FuaZkyFfKyTo01ah4ViAkJDu8YxO4bqpfMf2SSH
ZyJ7I6Ta0CPgRzwXxBtgqyaLfsCS3wF5nvOOdgWyW62+f+BBuYDDppaztOIG0CRpSoEZiaJMTx9H
JusvtSYCfxNDqlE0Q0ZhYvpIY6/dSrNFOdNsQgaRzUOXCOC0Z3w9n5j61zChJS/GneL5PtOeiEm9
rhCgcOABvbTk/Zh8aU2+7i9zp7iozmxqdag36mpg1Sj9sSS+BK5EpfvxJHX35iE+qL3ZOz9lU/nr
txCyx7G+gtkqePuOt2gP6Aa34PViNrrhA3zcBiPPpyJ/aAmBUMdd2wKwPQB3SeTBvlQYfuKQfLjg
0NwRuHDdp7SvDFToj5Qa+ERnBico12BG7jVSlHHBtUjNg5eRYPfDjC+IQ+dLDJiCPFTyFq7MoCxC
sbeJwSomnG847u7LTKuDTTVXjZffbiznDkEqYTpBJPXRMT04zsXP32spH35MHnyNPxeXOxoFSB0v
i0FIzQOC1sePNmmWO4QKuv/SQL4wFtiVugA3t3sunmq83HdrZUhgbrmzNMEQy1Pa7M9YBqLUFx6O
y2NX2i+3+QksvJqDAaMu8vPQ5nTBv4IW7zq7NFNx1oLpGXQPIYbVgtjLv28SyRsszu6OtFg1zcrN
KpvA7VSntaNt+4GcYTp4EPaBXesdYMoQZupK9bIjn7Sp6m2oh29hohQyqUKe+n940V3vqL3ESO7j
FMthdUSxeqtCfQIyrxbnNZFtGTBMZG+0pQZJFOhzA1I/n55uihXOGUR71O0/Chl8qP6MhlUZd/jJ
HjoqM6l2BdgmB6UC6i4UrblA9K7i/hP57arqU2RkiTabyrsXcCkuXujV0cMCErhBdfacxsr66GeO
UOQLfFuG/irMlvL3uVmKawln7bcli1tREmxJbK5jX4GYChjzwmUnpdQclRQxCfcaarOcs169Y3CC
IA/oTFe5n0GfvBEP5TjoRbgkTbvYR1PXrhY6ugHLGiQ8yI8vHhmiftYqWK9mBWXRlFUbS1VM5FeM
FuFb0SKcAjXKnkuaeXNX2MrMaloHT7IOsD2RIj3CoCf3KE/fZA9sEAyzJkDNDJBqO3FyZ8nHf0wV
4+xEIL3fRUrdv4GhALE/8sJECHSYFoLDNpsmBX3arTDkwNFpnDfKsN6cobJm7KK1aJnYyhmAa5DK
wQX48wQPMlAWHZ2/DhZvSMDF6mIAzFKVzbmCK3TId7J7iP9aGrZuOBIaA6hLeBCQx9t0X+LkAdY0
1hosihkcn9VZ/ADf7sm0HaSCos5IoEIpMJUGJ/gqqbIMM+SCblreKVG0dVFNuqH0Zul2/2AqVlX3
ZRQGWgy4tdKFRLheV0A83GTNh615PR5stlLcxzJJJg3RdPRL6FA0W0omdkSGsbYyFWT646RbEN5h
Ogg6PfA+d8fByaPHxbwi3jMeC/Hk3BDrW3YdNWfc3vnMyUpAhTUkCFnUtNvj0r4QH9sWQUpuw+oL
bxIrzunKZnu26DBQuNkXK4PH4c4IfM6fTJ5tmiRxk7/u/w98JhU49pLoewxpiJuw9hrUnhCs9p5k
Xi7OtJ+zyY2G5WI3onYoUYtAe2Oi1z+T1tfFlcv0sfioI0E6sFcoAZ51fUZzQulP4ESMwUZArjqN
PIrtaF/V/HG8+wTuyaC5P+qRGkIL2QP5mi0/UwW9sQ5M3PC8Gh446gViO/+wSYfVOXnBLBO3MOdz
hkrAGcjHjq0l5R5CR15xwHU0tokSrRt5xgUgILONclvl8xzlM7lPe+7lmogWutFmuFzMiL4jrVw+
fFh/ez/WSGt0TK4lJ6uPn0+cO1Zt6EuNI60H+EZtu7yCf1CjTtU5e5TRHtkuDgFboju8okEgFV/v
OU6B/t5ZKiI5reF6Hyj3OqJagsC2JfvZ4YjnUmVH1N6Fq/c5lkpoy/PFJ7XLzcms1azqJ10i/O5O
D1hoKAzIQOMzFLEzNwfdIeXThI7tXUqrj3X4dYo2QmRBQfkppwm4FG9PBSquoCMqiDGVn2skJbzX
wjq9lRhvSxLSnx+p9kKfhlGUWN3IVyy5XAaFMOFJJsKlwTZXkdC39NcxYQtBxm8Lc7v8Bl+BuXKD
zOnUXSitQYSisa1WO0WkLmwCT+SHs1CAb7pXuQR2u3hHC+Y+38vSS77jgd4JmkHUeLxa/1nuR0Rq
hTKQUnv1iwWq9CxqG4zOE/mhbhrLDfYw/Qs4wDakf+oLC8CqDQMoLPN8dwLYlskBZsMfrPdyjoke
lQTEyfd9ZRZJZCUo1Ufoz5iMOuOfG/RkTPcW4IhNM50QQH6XuOVdxnof3FHgHfPGqpCbdtreJLvX
WcNuIf4A9/HGzP5Mod+FAqRc5fktj+cANUW6SXbaLOUqj4qh+MzX/5Mhu8D8bWeCd7A6XWZN+/X1
BZw7Szr/lz7WXy7zUgKqpm4Ypt1bNwEXjqWvnzGkrmb/qZqtAIZzsmnasdE59DJzSMAb9oa+Rw9d
7sDoZWVF4Fewf+FYLk661uUOu68VpGYIUcW9hgFrMfb8MdP/lB1KGmL9yHGZ1JO4pWx958WKxqow
3zLJZYpiKj8YPvtXQp3TWbk1AqKxLy2/hIBPeS1lKdwWL81sSnDGSZU2znqMNL2gqTJFTwwB0Feu
wqUdfvA5a49QZMX9S1IQMnEqSE0+ZE9+ORt42PmpwlTFSCWcaQr39clpJUPkerLzh4HKT7gG7kKc
SAUQkRB4DB3EJYgZ4SiI6YfuxUqf/WwPGzjx/Pe35vV/c46PloKEXQLQFfsUX2gbx3+q/PUwsNTR
wgOAl8AK4nYQHz/MfmMAi7bIdqzKtyPyGhY1tiyk+LEOduUtdgBWCz1QBILRUU6+h75sy4y2wOuF
EnnZkb6yuBxHC8K+S98mxG2zqx0cMqn2MCl7UUGv4d+skTd3QeCZtp2fTs38Vp7kVUOYUrhVgIq+
Hh1sv6jCCdSKQQMaHmMiEXr83OHr4PE+YHUv8TBL5Zl1jHR2OoPhlGA19bppk6u6gDTrQAvjXEZR
BvR0l1v51cAqRf5/+CO7wxS5xRSYh/MFsaAVdkjSmJ6pUzXVJsyOhQlDiu1Y4r5tXYBtH/lEzR/Z
g8nZoKPa04Ja1MLXOTLACmvmH1W81FVRbHzu4OrpF4LqTv1+grDGp8yl14pVh0ZWOOCIVvHy2kkg
hOxmUlO42U3JFMsDZNpq/JGiWQZEzgHmtHBu2qvMZEYPn9xPdvL8AcLHHn4ozynK2gak4SQl8s8N
4qrFldAhaC4pA5Gn53xpA8ZRA31Er6J7XRlaAOUuuUrPh2a5p6+nv/coYWEnCS9dR5t2M1u4airS
pGTIB+7w+nZamcJLLgaQqFSBYP8VGV75b1NUz997L/cb0PJYMwwjZCPDixHV48tKVN2JceWyGe28
5fsi8jTSRX0XNxFq4ux26vxbp+WVPdpgJ6h1duQUh4hscuCfGwqjUgn53H1LqChDB9wQmTkOqL2j
yl4lHJQtA7alcfsNptKkBg8cnnpYaVXNjYVxGlmxuJhMI3JWvNvksLi2QbBg3oTdWZSpuxpZbDlp
L+eAgjnEQS9rnKG2wvBfwKlcKOeRTDxc0EBUtsvbjtIIL+8I8e8QHgR4HHmqAKBqnFVujG+39ulY
7pjG2wGbt0IdDnLFHOgjy7BomTIGSPmhVlt1yL9fTCADeDrX2T+3Yo9hOBTFvJP+p6NOV7+0OPps
eVf8/ZQllZL+23Ko4UUDfs2+3Jda4MXR/L1Oq5dpOLPqykVE3EASCWRoZVu0mKaZigiZqBVc2mhK
i7HaT6Sj7CqlCsinLVye6jfjKokfqKxAf9pCdrj857bBRt4JkTn1HjK9ctruH/O+hzDZfc6e0glY
GxEX2TsOqG+PSnNpKqSDQ+a+jlw1Uf8cFBVKlxTjigxLX/xXXHIaqgQboNd/ho3oAl/zwPyeBhIP
CrNql+4VBxciZXs7l+tbEQvZ8WbJoekUAdIJHBvtC3AwUUVDfY1GBkiWOyDIU44u+N1KwcYv4Dim
pr9dqzT3YFhMGGp1ExUEkLYvcrOLNpcZuXUhjDJs7m2iAwGjO3Bs641Pm/lcXUXkAJiwPD0DOvNJ
3ISO4+ZOYJADgcnyTDCrA4R3AaSlFe5WuISZAGmBeFJQw0LDgD3YMPFS3wcXfi346ybs5CQn/IAn
bIzA+QcrvXnjhmlezYbN8m3rZBc/LxjLvNEC70Rwy2TtkGHc+WMWkipFAZmdjzzdrTtKXL6vurg1
UolYeYKdbHK+DN3LM9iSocQzA6KUdLtYxNpjFpA9WU3VrmpFdZrG7XyJltVMXnyAtmBEuhMJUkKF
ZIqCqhAwRD1s2Pk84wpm/3UDcAu5T4yQ8dqXyblE/71dBTiCVGth35AlTD/8rpIzRnUYc6bIolKz
hcE2QuVsQhDxAQRX/BdkOyfkGrF+ZJIjL7cVxHJuszlis0PNr9CiPQL+ghM0lBjGV6uj/a6d6mG4
9PW+rje1wFrKcC8WsKWNHb17nCw5M0OtcHul/Qy1TdkTBMINlnjPE5im5G8JnCElKFGpuyhjPOQn
dA3PmJwCQgJg6jqfFOc6J67SyPX1nYvDp94LB5ZPso5XPBzyYl2cgC/phPfwsNBy79gs9Lqb5rev
LVsdpjCmZJlsEfm2p6V73glEUdWniaJ5GNpw/c7FO4mm25DOD+kQwSgUFEGYPcmGh2HHd64TBtzw
TYLKx154yYsb+ys3xBGPz5XmWJckNADYNuN91DaccoEcXmevhGA4B/2xkyABXmBSakwalME878do
8sLv+cqC96IL/nw25S9XWQ7ndhJsumgW5c6mYfPEITt7MFQfDV6Y54797XDr98C53wMqpmRp2wBO
k+1LZOUQmPbl20eoU89FVwErPrYGzwTSo9vMOXzHW70OWVnaRw2o/26SRyHZr1bae9dKxyxmmLUa
el/nn4Sl2d/TMqelzuTYxOfeglje6h7XNOfsnF2k/+mxr/heKbCuKZWUaCYS+AE6i0UE+xcClx1s
r5IVMPAC2HW5dYJHV79OX/uqkRY4z72+ZtyWVlYCRajAW6SmUoIvw0wne1KN4zLhaoKckyKCqdxj
1gcWQrogmdcrGlS1SrTnNU329pilA4I5EtUKrKKBenWtTmOPUqUWQ/Bjm09wnb027b7nRtWDR7YH
L12h347yRPeWd/A1Qkcw/AQSABFRbPSC4ljUQAPY+L08UU+cGjUXs7AMMsEenluHQuMaGmEmu7LB
lhdskQZ2bFf8VrITHIxG4ArGBz3D5nca0pSnnXKMNHSdKV/6Lvpfa17Bc1E5OAHX6J7w8mHCVTjg
pI9hkidhaWXw1cmFctOMwsO9dZ0S7Cl1CS17IZzyGLjm15DwsHbhbxtoqZ+EA9m9gya78KQOXa6c
2+Ed8RV28HlOKhFIuxA+Vi9sCRZY1c9Cje5D6NI09i3VZFFjeCuydo0vMYWtSNTFuaWWqn5ujgfE
Dg2WcM4tyM5OFoWxAVfuuI2ELBt/dpyG/vCdYscW2ejQlifbSS11IcUgfYlylVot5IJ8K/1011Gs
fjbCapahOh0mJ8Wa/PuQgcCtw346MyKgRCzI3MmeB4fjoDercgKF6rhe7d/RcdHqUWuyryMQKHoj
jLAr6agoqCnvFufKkUaX6MFeqOoGI673gvmrXaCT3TbX8SuFSyhm1f/NXHE7IpK01aQGRqodoDp3
KyHRxSaUe1ltbNwLZwWcI13xK8aTe8T6s7dDYBuwyD/sHE4dkjsbLvmIEOBhkUX+N/1Mo5z0RhWw
qp0YzOWvirUVhcssuWILOiZq9xj4PqHU+6npbJi06z1WOno7hW7nW4mAsWuLYJr/Z0OeCSxpbt4D
LL1m+Fqe3Wpk25XOSh6Wk9n0vrWUzqeuH6er+o5vfCfEQwnqFmPDWBgDN1iE5jKnx1dkiW/BLAhh
FjoNJkTox+oBcZ9rSGdGrbfqZowjD81HA7E9lBiLK5AV2oruY/sAnemuirI/tfbtfz0/jWve2P7I
ZGqZz6nopRZh6e+XwtX8VmYkJrGlk56ichYcUwLkjLyJT/T2ggUw80UY2OJFhBZ5q4eNYTCE5VJ8
tKTtAEKJmD4HAQYBt4WqwkqcY1n9eY/sSTvHyOQ5QOHIj/dZEuilIF+d+3VGfZnHzqvnt+CLdelk
i9VfU/2v4+F3B46iq9Q3QWM30Ve8Siqh20H7TcUqF0lWMLXq3iGdyPO8V3GoA5p59N5spLahA8FT
LTqpXPM4hACNO9lwfqpETcBdXK5xLN6yXwD0CWAdQR+tqZdhU4/+W6J2SCpffrOwUiSSKsYV922f
bsVQfAuY8ZaPRELKIIUdpKKT67FcdMSYz124esc2li424Z7UFUGma86UQahmPD/VjPnNUPIOmdAT
2uBHg3WliJsDACOgFOQwn+LvRFJPGS1Tvy8kMculVAUUHAiGBEknktDlYkDdbkkR3gQKhXykmDR8
4jsCmCt25h+2u1rT16ujsZwc6uB1w7OmY62bPUC2oXiKtQK5dVi0asRGcsxgwGTLLod1HmtUMjYp
ldUpA1Kv9QXCXPzfogpdob7ni/XTaRBOkojC7ymXkma+1qtrdGA+jh0z0y3JEmjO3vGLeEusfrjo
wIkRYoDfynx5v29cJ/sI2HOQoc6CEUFYwk9hoxUR8LpkgigJ7GzEBcKaT2J1WGp3Ag6UCzCMZnz0
ooR6RNuwUTbGtYXBCSizoHeAWXYR5vtdCa5VG1/56UTomWWE+6E0D1TWdXtF96T2/S0welop57Rc
IaE6Jc4WIeCO6nb2AdRuQ0hLSPpanfAyF8rGG7Sh2RGmwGiRJ79oAjLQKC0QGpIKgcvbKA0Afd10
Cp4xWlXab359fJpthSBwOFsPpfzf6R0nx8hx8nFaH1bvoa1gTpC7P2d5oSd5oSGm4m5kbaVa26me
29RpzYC+9V5rdU/yH7glnqlhS2/OeE3hJMHYnwuNjp3KZVQIwOchgUXukaYrLK1EMiN9EAoavbz6
Xph5t/nuOckuEsbMD5+pxTIxwtAcrUypTN3OXcdr+h7CF7fa7pPcGCpjkSepDSasiDCPdXb9XZQM
YxdQQXVDE0KK8T1i9YRY20kSsFyL8KTwaLuJ798P4m/PcEoLYHUmfoCZzXu1Bwu1Qbrl9BYeinra
9/WIuKE+K+HJWIxPsbG3+2c5glHbXsBBdf79iCvO9Vq89ezJbwuBGcB2A30jJbwTP7hwJ/IEZ9k9
7jkF9SkNyY8ksYlD2fBguoopJ2vtpBZl53IyLIDWt77jH/PtxTYuH4sHboGhvAa9/1kcEPlgeofy
69qCWf2V4qWfMOttXdsH1vn3XOmgnWyUT2tOIsyKM0Av6QCtTBWi3oUJlnQbkJO1+YtkwOB5p+Yu
KpIXd40hLPwz9ss9p2L3Kurgi0vBhTmTTuzWzBqc/WVnD5yuH3dWcmrVyM9JAtmbxsiS1hVHcwu3
yAaZC/dXaqSN1+TosgjhgGwWfyXjYNOxjby7isK6ABymaY+hxpAI1l2ZWrtLKOl6GpFXeq5P3JjI
sGZ6JM8fwTXo5o1wJLmU548kfT6avIYyTKrKf8+RwUZK7VDW3qm5dr/wz1ZAn63PZRiTa5mwmXA2
BmJyN2MP9Wdr1GHjprOkxy4wk7k01cdPA1yPMlvpp+svdvInIBiWh6fPiMOL/MZdHrOQ4lah8hg/
eBwFTIgQDxzYQE0rKwbTRLWwn+qS+kOaTHtmd4/Qjf7DnxrELY4mLGF8xS7BQ25cFQd+Gc3cEQB+
Wf/Ci2sHpwK4T58NLmRjuyBhuKtRICf2RO0ETh4eZFbTYtLoI+iz94PRZNTVX1dnNyVfBfuKt9fQ
d7quehN/fAOgjFZI8bFKLx5Vm7A/lmG3bUWoj1YJsuaL4AadKF8NZiqfflKdJlg4mjGlzzOYKFgd
LVk0hl3MnuNVCzsYySVFdEC5NFKjzLxynGBpfPH6VQyQ9f/dpZlEiR5V8d5DnHCQMOfH8AsQP7ra
WpPCZYhgoJx7FYjijhXymcIiU84RoSqk5vk4H+sEaUiLdQdJNprYKxYZD0PQELLlMrUYLmeweOoa
99gbHMFriVKl8/797oeKZsXmAZ25XQexECZqLAt3ofw9rnzl9mQMxCnmm8lUOoMOqtnYi/jgb5XV
z1jgIzhmdUIrdivJwewKTX9wgstw88IPGQMGwK74tH9RXxzhbJjXMxUMk9IAjTYg7ESa2ttluZJ/
K1lVfLPaY2B+NTnGBopn7E9VrqAgjKfn/RNif0OlKGAjKZ/5KtbwTEsGN3SqN3mNIhpiWGSaJB1J
E9jvpWhbOy6wgNqdJV8Q9ppaxrx+HD5Jglj7ZzjOkCAIhWjQYaDSIMvKFaCDMluyiVCPu+OgIg4E
mAUcgdO2n2SQLh4Sg9eaVj6m940ZsseHf5ueBD4J0geabdiMzgQi66VTDBVaZUCtN2uwYFS0fBdA
ENCjtDSy7vOCDV1IT72Jw0G/Kw7TnCwER/Abe8+ApKQuRS9Ycrr1QHK0shId1n8oZFWMuL9TOPbE
JGsihgQ+LzqV+lHS/omYpfcaokZQN16ehF1d8+YfOp+R6cne1fvGR2At6JOlE4Vwf6EvocYPop0l
brky+8sUbxZg6TWMJ3eNDHOCIaZE7mGv5EoKafn5jEh3MHdnmUqMo+kkxeOvPxLASla3teA3b205
poQY7w339COJXFMp63iOG8HgrLaNr1nS70ppZ9cmkzLgcIT4DAOqLiTaBwR4UJeuCkOuLcbTMo0U
ZUuSt2howsthMct/lZvPraps33v4HxEHqCy5wOfAOHoZzFHeyMRRQ1z3bgSlYayr5kp/rYmrPiUF
800P09tjvUL/2m3aJBC7FmNqkr7guernIwkdb/Fg0tDRjmUSuPckNsE8g5adlZucd6ZG/cYFr9XO
18FXAidX2q0fOr/EIsl9Lb/wFNnD+GWHh8RX48Wd2umoR7sOJ3U8b3FWNMXkxxZlgz7+d41TszEe
TwSovah5Daq8S/dvsSK13vSDcngE8Oh5d/99L3xCmrx6yf6Pip0U8fPYi3fmqm3SkZmK5XKF5KE4
CYn55/9uzwNAnV8yaem9oz6WojPM1SlmS9JHLADNK0e/iSAzGEbqBBfnF20MPlf8F2fKPmMbVTQI
zKR5RLi9kfXEt9K0ht8AB+U42OoNBrZtnVSB0icHjS04E6ZxxBI57W0lLvqf4Ft1K9ZC25HnoSJA
92TiQRAS1B6aTWfpzkuqONGimGhT8CD7rVH6OPdKKOxZmhPh7mX+m8CWKPkjXC5ZBKCRXk3dai27
8mDHWXlmBn7BpkiaxmW4OXlMDbJW+C3QRtEBaNJjDMbVPCXaLkij6IiujDDN9FtKx+PMbvl/bu61
JK6OuU2k7vR7nBx/vWG/zSvIDvxQIzcgc0olVQN6djtCVbZtRunNo211cRMjmaaPZ9QPwDMQQEBv
qqQaMwNMJhOzHORyfWeVnijlaiCHY7XPaaG6vTb0CUynAovKD0Lg81BL6oNHNVYOqn8Dw4KywL0d
fx7Xo58n498SERRfqQUPl3KGNUyQABZyqCiBLoslnRIpwCoyV2nKCInw7qv1NonKujgVg5DycxU3
v+uVa+E/q/axSdDbY2+4caLuD3vZ4LJUJioCrbfty11CtJ2UBmD+b5fddf8PlbiRc+fsnmMFcvHY
z9yxC2RBHPCIQeEWd6hhZEmS8QjbF+tFjFYhaEflsP+/uv8vpIMIPvNNfLilSRMI6gaLIj0N7jdX
MzUkLX6Rg8JikDdfj4K1Nzl65lPFYl8qyds2K/w6zj3GzsJr00i4WgLJx6VeafHjAe1cwwcJRHtb
CpUsB8FDaOu3MfthmzkoSFMkKAzf7amIKLX1l2Sa8VCsn7U7ktyiqjFmG7PnJgi7HA9XgY2af/N6
8ljgMuzu1vTl55PVcd/OTtAJSA8UC/viIwejzVtNpBFsNap2tQllhh8RgsHfZr2SEdJN16MROlGN
KXO9Ld/V0cxdWP0JLVAHWE2Dymn/4dj9P3ezUp6+c7F8o7i6TYEhEyH7fzU0ydQu3p6JiLQwoUO2
o05FCPYp/0GnVhFZ8EMs8oHDMwdJZKtGTcs3eLSBqWCUJqQmqwLzvc5hrMPweO3CNG5uHbSS1J3v
Dp+GhBsk+faaoc6i5RwWvoVnOWVy1PzLBiLRQYKs4ATXfelF4uR7jA8NBpsk5lAQREiT+87lu99p
c7pzCedCn2YPkr7ycbrPeYvgXrANfX7CV3J5ZYZlwsAYXo9TNtzoy2ekTF+cmgoQ+5Gh4j899Tkh
36gLibC5afizTDQh/91WDsMY4eVCwrKrw92jx69GafpEaHPNmmK440NsfkW8ivuyIIn0sOtLkMiD
viT1VmVv2V8j2DUINwF1/AXqIcdVGISrBZSc65Ds89fXCwldkqUfCQYLc/VgKJ7NabgrWtfRSsah
FRexC7Sgv63gnwF9BVHl47cTXYU1H/NGMb7ufwStCFb0YfrqJ4yyrvbh2AGTYJu0kNiIiOyZOrit
xaqrT6xxrfB53DYgGKE5gkjbi7gYgIVRpAXQR4jaDmnhYbt0poDnjksDNolABHeNE4L74urt5vfS
dUL4zWcEUZaZfZPXONgENAXlg5APafHb6jpthi+1pT8A+wMIFnz6fCoqWCg5QNx16chSXgeXsBkQ
BbpG/GeR3ZLVAnj/DdsuHhVF9/feCGqKUxwret52VNMpLLbnB5Wz85gd8HX0NJAPxRaWFdrqwKa5
u5R63auyiUOx3HL7OKbc0e10kH366ZnJflrJ6hqbtYzCkIDWEyYeQpv8jMjDSc+6dlZYom5iNKmV
G++y7JXg6WOFmV1uSHWs55iY9lRHMcuKLWDZtzcP0jwrY+3oMRCyEQsY7uk0zYGK9dcYA6yPuzED
TH0xqm81h2HPTwWs0yRaOpdckyrsHyf0Z45nR0p62h7cinvbull5Q2dot8x+3tYQZ8S2S0JQ01b0
b9LO/jqRBMw3XrUHdFukL3T5mazz8+TkPYqXr+kQNBtaqFSVnGT55Zfw9D16BzqKXdD/+0z7aRR0
aJA6UcgyWvjCqGjcihtRPHNkoeJ3XV6DNOE7F8g8PMFV9NMfq6A7mIMcFvTTS4/pQ2Q1Mrb8Go40
+zgvggSrouSTQlA40eoBmT0w9MJE99aUKrp4tkQtBnYgWZSPL67SPcGN3bw94BMSaEHWvXDnOevv
Tye/HOPulwxoQUTwupbS/RLWCMa8xOAWPPvjn3QgIBd6YukRvOPWOnt5BByAqUQN8BTW3fZSiFIb
m7WQOE1hAL8GkaMKQGNLRjzAJsyxTjomEkrgsOtQIWaXVXQVYczmBs5T6w90PFnltP0KqwzCUc2A
TuS4aLt+cVXaLGaXiXbhfxygu6lKFlHbiKoB87m8q9dpvXF/GQPn7CsFH0fu+jE5384vHmmHLXj0
NVduIOPuGRu2+B0lZbkUDzdw1c87jxUClzP3ZHg8yOUTn6eY0Zuuj/rRzGamXNf0txokNNQnSB+K
//OzncgPrGbX3inlcJVffwYO2HT7m6yhd+7O1qO59mFvF8jH0iooZKqASlpTNVoAjA3zm8qEmi+2
lmWXcQj34Fkjpyem+cNpiQXKmXyodOSNrGvbvWdtBpfgvoJLHztQ8SbuqlrBK8RSPe4D1n1F4A9W
ZVZXUyRBrP/2mcuskpBYkJSw6bQNsqQ1K7mhEcJmcmhybuW08arj4co5X+EV/fWt/eGa2OK0HYT8
++PpPOqlQ9JYSa88q2LclCJf4+rrOpOCwiVPCUoPH0DosCQVr9zkslYp9V5IY6PUG5nPK2V8+usP
e3tiIA8yUfKG54CZyi8fNGYuVRQnQjQJnuN9e/Ee7l1Guu58gSRqoTDeKMhXWTQldKzumdmD9GeY
7BsK6lfIj/JnjKPyvwinEt5NDIw82Tw5hfVu3TISVMJjLepOlwuHVZSZrEYfJVkp9UMjO+NFTbn+
msQx2E0rhDuOspKfxnOCjtNc9blnvCcO1Mzbq+H+HFL/V7EOyFNXjJlr80G1hT4OxQqNntB+ea3y
g4U3IAv9hb8vYglpMJtJSOsF7ECpXgUNIpCf/fnOnQpuPVz3aRsOthXS6rQNFvOpvfyoPh8jLCFn
XaAlE/WpWkcymvw5OIPfuRuwhbIGYEI9OMJmDQEETsaSWDLWAnR9RikeZzRC/a3+ugQ5BtQbFGQk
PeEh5OZ42EX2sL5OUCH+VIdA8VH0vBGO+M4UMp7MPGyE6b84xDUP7as+yU1UPdLD7EFWSYGRCjYk
pzI4AYsl1YTyPggge2ihFPCdxeNTVO58YWcow8LTWcfMH/k6QE1veWh3gG/OYLzHX5wDb4EqBo/L
GM0BYybMS40EZP4i73NEFj8eD2kOSIX/9H1kF8xe2Mydy9+M/YHEtLnubjQf+xpHlE737z4dXZ18
EhcO0eN4laKSx1DhWc+ZJovu007yWXL/od7pE7yT7R09ygyJLgvndvCCBQjrYLhGKX12d5J1s4f1
KB5kElKjaM2U6kSKPCRlhExG+Al2pSHSaGvg/pkp1ZnTLzyW7jnxp0t2QyKETqZK0mgcsWt+fAko
PgWzk1/HAMoB9//Ih2g7wmLOCF67w9XQ7CjH80XkgCds0jWy8rEAQNv9Y9uOZAwKftq7Q2NDNEB5
JvgcWuq29FUc1UH7FDiqjuqFVhGLIFShbV30HdTCtBP978LvN7Am6LVUegTRL67CJYK3EZD+nrce
pDsndqvp2GilOaJKLh1iU+d9WagvuvO2UFd2Laus2D7Kkc0wMECCRaXAm/dVXDosdwrfB14qCasD
1zeYCdtC7BtEi6FLhueFdjVh3t5ESgsLA6jLw6LuaZtA3AM9y84XvtULlvjJJiIV3NiGdeqkAkF8
Dp+KrFO3jKZK+BzqWSpoPZLAliw2SzuYYXDrWzieKy5JHvQG6x9qfd+zgthNVQntLcQYuXpH3kvt
tssqqO2TOG9Lmj71AhWcxDC9Z3OJEqRPdL/0PKaKCSHNVCDXuWNKX9MKIOgJdb6GpIvaaLWarcLX
kZareS9mOyy2x6Pfj4/FQsAbNb9ozOq1ATIyv4R9LliWS0ojSCO+Xs/Nz6KkOzxkOJdIuOIxWgrR
FAC1HfW3govYIiBb1QGkg3NkWyhzlubaMxj+ofb/qihc6Tyew5mF//sD6ZjpJuyPnuoasUDsPfAF
EsfQTPyLDlT3MzetKgmIeduzRiGdJTGjuGnNU6IxxHf2pkoBqMRuo+jZRTsUy9TaaK4F9vSN+NvE
BDdkquGCLs8TxFG0vgC18Cjh6jxxQp8g/HkM10aH+f8OQOvNqRKgopffZq1F1dMj7X9D7bhLA2/O
U/8zAreMTsxKiQu94otvnMsh5zYa8sW+kHqmoataHSkCVmpPEFQlMRBKK5/hGIBh0vrI9yRsFPdV
E3FQzfGieh6gciIvCgPL7pEuLY7zSf5yM/cu60d6WB4j+NCTePmN7t6K8JGpHnqtx8H9z0Aye6DK
icynZAFCk0IUAT4wAdvTZ4Qda2gVYvr5eOeZs22SvIvA0pkaE8XLZYhdQSKZP5MTsMTeUkLZCCoK
byEHaglbjy68SmxOUf8o8GASX3rJTP4m3VY2opJ/04REJwqIMQn6TePmcsHEg3qQrY04bigf5/J1
oaZXJuH3H2JJOq/HiWBGVZKrtopFO6x3yC1W9POJG4azDMnMcmAH0Z9R8ZX/NViYEDBBuMUR1LQV
i+wg9t2BjqIfRgQuyNS/x16FVwzY292Nz+qJaY2cO+Mfcg4ujeuXQhlZdzXVCaK51CO3pdiRwBVv
eD8HApQ8s98RMVO+vat7oxb/LXAmzzJiPhnXsKyo3xTYkUIJwnxAt66K7dhAlCEV5DmC5z3Z1LVT
0zipMhoKHU0mnb/RlIeNBAzteSVArUQqXTDREya5FIe/jPkzINq6YBb93uINSWA3zRCZhjAWGusr
r5CwoB7NXiQ4iojM2ld6B9yF5KyZHnwAJ044pBHaSg3BTGnC5J8QC4Mq+1jU/MoY1rUIBH2b7Xso
JisgQWpvW5E6mBxUqcSsGhslBQ7aJ3QhroQ6R25XjZM0tQJRXQe6ZyycY9KT36ox5qvoTsxt6QeV
sTX7qMuaDvWcfleBmWIEJFdaTZRKctsJFlKQbVQFMojB6ABdB6cDjHwGa9WGJzRU+j0mFWp/DFp2
1iOMiU6/g+zRfO2i3lEuDQEo1Nfbro9sjWbeqavKH3Mz9TIV9Fl9GzMqmHq//vb7AsiH0sJ97hBg
2iAsWclWY8dgHDvmNt2Z6FJKaY1zSyuUBmaZVHtFErvwAt9DrnKIlrZcpLWpW1+GoDR/nM2n45P3
b29RD5QtljnAJbCNrsFqPLuhu8XRRYyGdCl2oWR/b9mtyxxYLd7luIDhyJsVSE9hviD/WHzYxp3a
xq7E9fA/sp+rHAXi4P5z31G7+Tk9bjCPtqzZlUTiA7FLdkIpeXFGoM9566MwFsan7IWfzc98jGpu
mpDq/cFJJLsciajxWNXv9titbjRyIAddxzAytHbFq8kzOWuCK2Cp/qBCnNdcO60xsifCtsTMOcZz
fLUrA0yuTRYPL3GW0jJxyozgofr2mjnLDUF5QCP4DFWOYhIkUDTTve6yhw+CYJ3xhn4ikJuoI2gg
Sr2mqnlxlcq57nl7MP3jjR/rG934/CQQ28IYAA0HmTnJ0twhMu+5ATvoSI6/a4tlmzdaLX/Rmt7k
ULB8kuc2PkJdP3ySbFu5dIExP7fyy+tBhlj03OQ6jzZuj/jE59nIX0KA7YVqVefpJYJmJG8EEoqW
H9tyrTsKQe56tfFIW6RXIsNPCmQRmQSecn7IfVBaGXLox7+Tu/Tmz5z8kShcA3XtVp/N1Kp2IXbS
0hGDERA8EuhpZA6GjrihWexi0nHyLhlkaDlR47HQsLonFElcBtAnqOBocnjGFLX5LA87VLzinO/q
5C3kbfMySSWJ5uMvfyFn0pM6M2c2hJO7a8X2uYWzhtfJPz2A9KXtkfonFUJEAgtATTXlz8z7bNjR
RN+ilHMh6cJKMhN4OTyH9PKfOTl/2DIPKIjwVqKEqYHJEj6FF1fjBhKElyM5MZskPhYbXcV5dein
OT7hYLe4JxXuvNeNjNFwa5N+nBkRsC3ZoncgoWjkLN4TZR5TBdkmUZgRWuQsN0abmkGL1cES+LW6
okQNyxQkJ0jll7xB0mkWjQS0e8aJdvxdEArq86sep/VnyI/YDci2CneH1a7Me+JMuEHDGVhaB0Bc
LP2O9kA4bMRAeSd/cy5Lsb0sLjDW/wZSou++HOKZaFdoz3+alsFTWI1HTMeH1AJcr8mo1NI0+vOX
vXTFoHKOmSVJLNtUat8mroUYwBVudPwCRvHZduG1DDBN03p1JFPasSnlQev8F9vU/3My/7fzxBQN
mLIaHnXAGZVilM9IQN2FcL7g8xN8oAVZnifnLnlIXNL7cZ0YNslsJqawrRZMCS0PIbVCy2HmIOTQ
cUtsb46cs3fcRpQ7ApVutMpmX5eG2ep8YHSNwwqfAHNUQu3Rj5kg74LsWwKaFSnY5rcEM6ryAdDT
xrTBgah5CKIq5mgAJob7eCEpW4miodMCsoRER0kpVjKohxgfmoQxFdQQ6SfkJlnduWtfQ84g5xEF
xXuHhhZyZrwYpen3nQq5tRXOYQfb0chkMM/b1eYKs6fU8db35U8xZ5K01Bu5RxzXLiw8t7084IjO
lFqDG+29XtCGWSeAsh8ejWgCaWGEacUnlyU4ajeTm/RJzmqKbmBwQKfjD8Pf1v1oChUhQ06JwMhN
nnUH20ZqBaUrCqhcjZezer/RQoul63OLhZwKuGcw+OPqtL5EOOKJR5Pv5YJF/9T7NJ+Hdc0YrsKc
pCdKgw3gyr52IHmiVTyQ3LoSuWcZiOWY1U0BJZBkN0NG93iSsCumECQkeChVxaeyiLGKyS5vAjtA
3gSR7p2U/Du4LiWC00VWvD9FSY1ogJMAk3Jol56+Wf5/4rbcyAzpO5MGUyCsw7EfYyQ6iKxOo9Rt
ckUR6U5TYRre3Hvddw6dUyI0STgFftVIlFkR660fYO5tkjjI3CBo2EcuKoDm6bFAIW8SD6bCdGvK
eujBzC1ruoDYDeAF6o1rGn2pSVGr7yMzxg4LaHi/ceGoX8ZCUlmv7vfl5IUDyKaAdc2/MKXTn/b3
ANj1DFcynJyeQFSoF0SxdqkB/qNeYtzhLuZD/AXPyGpIMfeX0TW+KnXNznM/XoPeRK6bRgpPnmYz
6B4B1SGYE/6TT8cP2KJG9GYJqYWITx6W8nTu+5wXMT4SJbN1z9usizn1+quXLMfJE43inl8Am3Y1
pfVsKM+T/uJODyK6anaWzlEqs10GlpAtktoZj217BUuz4pt+LcsLKDj4LFCdPJCZq6Eh9sVlj2LL
/HjpORWRf0j4INBhdT5wX1qI/QAok2MqLkH3A/hjBPPwIb0pjRUBJ8fVXkXG4b824hDXCNjZm9po
xWfFDZe6+zPpbFPjhF5gF6kdVCZy1PEjyDn8ta7m1Ops8HIaEyZHNb0kD0Umi25nWhnt6JX0pg6H
+C2dFxw9eYyHnpMOQF4Ob8FjMoeugC5i2vxi+RoeArcQIqtkYc6zIMdyNfybuqSKa37A2GIVucX9
P0jHSKLb403FsZ1ll6pQQJDyV0JTFKLRaGiWh9vQAigmYAIoCcaf8mlYg54VKpdL8pqkziiw256u
mr+48sgX5PrV81pAn8i7Y6xzyL0oZs5ZhosPdGZ9olnLPoT/+y5EGCSZzAEi10wR/W2piU9+Bkrd
9wQApxWebKH1A8gbXh3m0nEnDd1xDosI6YiAY5oEXOqltEcE1yGuN1HV3ug4qjz/2Prj53A6dAFG
Kxn1RNOIf5QaJ92R00/rq1Fez7Qr/BkmTXJq66tWx0na0r79V0izOawLlWZ85TVRAqAuhCgum8Fy
pJoeNbM2arBTALRQkfrRaBTIhGsVFaf+GjeO7pRanvBFzVmPTcCb3uutMNH+uJenwMqE/wNOBKek
M5alEFbdcUyzLQbjFtVEipWBWaC9cxLZvQquMzoXYcPSilaFpT1rQ65snz0eN7hZXUqYUERI4kWW
tycngFqByhRUXiLHXn0r94sIUnKFrKViAnlqLTyscDDZPfUNYE6WfOI83sRx024KEmSkjUKkIAej
vLiCulrwrkuC8lxpSUbFC97YHot/L4gFlzNDkWJJ1cisa9Ti9ujbXfM2mUrEBd+MMqyenZCQ9Rab
+Nhn1x5Xkhsgvp239vCaq3FltnMAL3qgQMGKMz856fvsmmgBrwAHdrP1ZLrUWjBFW5LubrbvNlVX
4x/LUiQZ49R6aO2q1wHQpe+QsZuRuU4qDBSOmK75ozOwauhSi2IheTMQ2gChvJ9Frdf7SOtevNjg
xz2BIrdd7y2tRe+088FkD86WfaCmOFnSe8N9leBr9/u7t3oRTYQMkm+TkRa+dmAM3JYmovw5XPhU
EgoZNGLbYPzI7xW/botM4SqcbHneVbqMOZNW+h0AQKzzqeULqhCjEE6sKgbK2fG8phMjI7tFwxKZ
gPqlfeo+Kc35HHYySXjxNvMUZvmHGpCwks3NX3gLuYmxPUjQw9llEodV3rT76O3KWw/FX46Pp0l0
BJYSWjmExL4xFbLVMLop5RBwO6PU/S7oLcMzqFJCSwibtDyfmZ0kKiYKhI9ZrOkh1xm/B1z0UBBY
mrur8R1YS7R5b71ayJAvu2fMdTcsEfsTnblBkCNiNv+CHXRezZk36q1WM5Ykb+KJUaGr7y8uvGeD
jBJiFSomCB/4ukKKSu05m1Ez/z+WNHkwGpVOBpE7pUUtIesKzvz7gVITwVtz43UbADWiFfuDdjns
+jl0EyiW+v6OGI57kJOWjTLnrm/GXu/mnYE90fHgMBmeNe6wjBX5Q7DDOnfU4TUmapdZ1japx93f
yFKogmPkfw/RlnZKtKl6sqA7mvG+mLkYyhCPuiuhhk9UT6m82rF4JqVqoYjKNbjUxhLpjy9SbA9+
NzqIS9le9FIYvFlePrd+njePI9mels0xgTZ5atdZY7sk7ykxuNypCW259WYiJ4uC6JnxjFs8+5rm
aVJ2RRkWuu6sHbfgKoVpAd6lW8HEK/3dt/s4kBvclX4MjbTt4SjLbrBR30j6nwym8Dh9RNxKNyFu
bDusjwsCDCulzc0tqiPqfBnaYBCTGuYYcH6pOzcUWOTf7BlcVg7bm3Pz7wfN55nQ4On8kpuqh1a4
26lhe2fWBPthttJ3/+n0BI5XTNvDmnEd2QFrUvVt9Qyn0jxwIGF+oqp4cFaThNLP0/yMFR9JXARD
pYw+1EIxSbo7Lwy++uojhdwCKafNL+XI60aezzIqrGSNkrz+qg5j4Xy5jy5qa/tpVAcM8ORAoLQR
TRw7UDhIlc9WPYCON1pdE1q8aoxEaqxZttABKlQlFszVRIs2gy35ZXavzSdg5rwKVoeVzIEj9reU
jhBifsfPsmULxQBxEOuQ4EZ8IrxN+1fZ4PGnq61/06hnDmrZQMxX/OzowE4iDZ0SYJ32OJRLfDgL
15x0Wj38vV1rueUS0cIuYvnIZdUee4lTMXkIK+uBDeVmV1/tDhF6LdoojxTfYUYZym/Qwmk66QX4
h9z56QA3U+QBDpvA3Iuh9C9p8oUwO8UYnilYtO9zkq9fbuxzjKHhWiHtqbd1U1TZB/jZZKdCE6Md
nnr/8d/wpq+J2cK+c/OSWHyRH2gg1H8QUei4xyzoD3zgp6i7lDxEgyy3f04ePZVh0MRodrrY19ho
6TR2SQCWxj9Axgk7en1TpEGW8RpTf6YFw6NYPu8DMxqVKTl+vx3rFdEcWqwQ6le/vrF/w8ft4Qfk
pnnFW36COXKHOK2kQUexeqzwTyls+Uw6nqrtRD/vJjXgnv2pL/SHepmQsxxjhtSoLujmLkjbwRlr
ytDdutzRNTtEu6/xTeyrhH32JG7Zx35MJHPBGelT5Gsxc8NXqlggQAcOrQSM1xfUlqsQtNCeM2Ak
UpWRqJpLIXEp5gk5xGXgX76ZqHz1D0S/r2GwU0ll/li9hze6BPu9Woi+1OwZx7Zfw2cFRGgsAY1e
ru47awXjptUBa4PePCnmZuQuhj6wcaXxCi9v+bs6U4OjhBsDCV2DLVFbZ3UfYHy2NPR6lWNjWIwv
CvzHjlN4/pztalKtBzztjYj04R3KSF72FiYcWzp9yDAfv11HyAZEhDmU7t0Jguu9yULOiCdYw45a
ZJ4py7OuVWaJbP5VQpBMfTeKVJpwhDg/SOQLmDxT/YoP5sh5GouNlP3UfXhmibRQNBsQFGIYUZSE
PVxcjySlrcU2RYNYLbamBOSPrG9Riruk8v1UFXx8JfkbXq1JjWmyIWFMMQ7sQANIbTeR2+dkiCvZ
RFASclsLxIvCL+905zwBkNFvLK5goY040gnYi9lfJQNE31yPma+dPYPECvwECT1bZEYdM5zTzB0z
4g2ShsIA2h70TM6u/rLkka9wuSwJqCFHP1mf7lRElpHHmOzCNtW3UdWNfrRNtR2NEtJRQa+M8Sk7
8SfLmBe1eJFjCnl0zdvtjrd6oc1a8o2v9vTQUkRrVJ4mXJtieUstZtCyq0eFfADc/9eqbdHHuAeS
gwZafkA8IqJrBfYmYuWV51I3LUMk2LF089B5BMGDDdByuzinRtBNkTmBrUds5soQsTTm8cT/Sf+N
+DNESsqGsVgq3+lq+Xy6ghj3/9XoBMDIo0jQU+bGsAmFf7gQaL/TlnVM42GqlS31Sw+bPusLxB8I
BepX6hgfZOU1AhieBVyk1T07kLSbkFZBx33RyaoITSLzzm5tSCobPAqWwsh7w1ABI6j+ez6CIdEs
d3UlJs9KaaliWzP6ICanqwC42glfOJD9jp7WSw2EwqURkgBB6QQbgHdWOVCDJFfLVwgBHWh1gqtq
9KbUTGxOoQOGaEj60REkgoFa04Ntx026dq6uFBOcKNq+ICFFHaUc+TAnydyOEPJ2NhZoM+Uy9R81
PzIqYh53fDhVHsBsXNYCG1Qc4sySusX8GQNMcl43dyHI91tpWiR5deSrBP/NFP9jNBMAgP+uGTy8
n1dLlPfUcJqdNrd1feAxLchJ6BcmxKiBGg5nPxoxAteSv/9KngRK0C+enNE3myFCOb657EbVsus+
UJMvULKKu9RzrialCU746FEFKvX+7GmDFwzEcbyd1nqXO1XXgAKQXR7eD6QvheVQU8Hq53AuZ9f6
Yz9TxG3vNfx2F2qRrY+XR9RUhW6qFZRJOeGUzFN+aE/sbvsiaEHe/fAqCs6XkbPDtRLpJzA2DTfg
s+2Gsbc7a9lEsCxrSu9R4BVB+6uzYGop8WCs+sEfQIKb6GOJ/oRHwbXodv7qUJlGAS59cFjaR/OR
z3grDRSYwLAd+B9JOXqKyzmWM7k3+NqHDB5p6mdNdcJSf2EfXxLPSzUWyEXq8HvKdnIY62IqXU6h
0F+JfawHJ26oAIl/VydIiO5ky+9a+tK1Q7FT/Tdd+npAuMvI1egw4KuTfxJd6AJHQoOOea5MEaLK
P7l6eLef5dihCtuPhHNioXOVkuGvJHloyXVttK7k1EbH8Gxl4x0rnUwSpyKbABdKiS42RJY1rtAE
YXiOAQk4Eph9mK//RKzwOm2Ymy7vhOsSLmvgGZxl2yMIUan3gdHfsmYIMnKD/+XfRSO3f0MtQNqK
BD5+6m8n2591E4BPinF92ELytNhrHB+Ykoev6U/AiAL0MYUIiJKI8fNFTTS2TXlfr6C/D+xOhNLZ
cqjTPMTttvfz0jy6+iTOuuBFil26Jd0aVz6VvaTouRCqBSZwcrqeacRYSsJgi08Czfi48goCYEYo
UdNHJBbRQBxdsX9zHSwRIu2MFhYtKpR9WZmndG6XOdz+5bAZKT/iv33IYxqS4mqXRz/LP50Q22Vp
bnZ6yZoO37GU4dD1a4hr655xVJl+SEGuXrbqs5PCg0VWCa123z+tzqeJ0EkUNItg4YMguiAyH2Dh
LJp38Jnf4i/q4BCwi8Jv/7ZSChf/GkVF6sCftjSEY4t4aH/TOhgnmMvAn3a5NZTO7CKVJfvPKqIA
Sp22gaSxM50l2vrqFC4nK94vz1JBaF+BOzr3AgVczZgOgGwwTchFZF8G1HOZYri5UOzj+JiQRgUZ
EDZSpezbYooq36TuA+qGas+6fSdmomXK2R/5AyCKsz+30sRsyARJ9VcW8lloK+wDEp2gndr9thCc
HGPs7dNIEi6qwFg0vZiTJPQpW334hlHN0ik6XFNdZM1iUEI7j7P2K1dvo6bas7h1+QTa98lPVibW
f0w+gMEWppZpLfoEpQpQORnmQXd2s5OHakUxYgagyQp1wQcPCFhM3pcVjPsvbnW44urienLH0o2R
tXYzyS4n2g6xcMLyhPvQjxi9UMCF1+XQAQdYCOKxFlRevAgwUinffUWV9KZGQS5+J+ieUGeWIqUW
3bGlF9JWi01BjYAzb4b0TADhwbXCMr7DgXHO2ws44BJEQFev7t690rTJeSA02d8lAwrqkFmTYkgu
PjcE1z+1oTMh3jdNDm5ajKLx3Pt8OBYIlTLRGq1iznV4H5GuKQn5rpoPQ4roUAxkn9UVa1j2K3I9
v0nVMet4fX66NFBX6eJpw3Xw99SqLGI/mFnSF1T9z0J/f8j/2fP6udVOq3ECL6X7fmtEXgR3vPn7
JQ4pjBbhrihdPq2c/PbFNmvUftzmC8Kr+wkL2d57FJI+i1o3M1Mree/rOitzfx7w+Oa+z4bF5UbV
yIERZOxEMU/Yn67VZCgUZcUgVQzhGOXv0At66O76iT21pto032Nv/ieo/bOPEl4+rAb0LPbqBaoM
UKHF9kUBPCLPE8+YNs413wlMq8GbCTGsvEXiec3FW0k8r7yyivUJmuPq5OPBsxosRjOmBOTL/2fs
Fv3G1SFwPKqRoO62QmyqEeNRfEFyqaeZxQ4FkZCob06NBpX1hLeZCsOucprR33xfRtwObn38tQzX
9q5lc5AF9lHgMEyHOYMA6svrvchAF5QBruRQi34e6Eo4xednYafGDIORXL3pjyLHCbT3Jq3Rkz5o
WoBawJaODstIZlzqBHgQSuKbx/Fq3j4baI91/EsQcSGECA09I5gCaHmDclC9RaCotJt7GsbSpybQ
KUwKVzPUZENm86auoH4SKm3ppB3PhRrbUz5MEcAKqwfziOfWR4JMN1F6rVMILqoeUUC2UKunOPYK
0zwNeR4ImyuKdevMMhqSdvvyivxMClVAG95J846LCU2PXjtEy0sFIodSIdZeCv8wb4ssG7f3cIIh
M4jttP9et+rDETNPoS4ll9vEFtOOZX9kFh/RKICnh6kAUdRRmr8p3dCgp/G7jpJfYsCLLL9cBsyk
dbDm5LuLkaqzmp+I6zVdme+MDG/yufzf+3+uY7qPN5IIj1yGkyGkyFsIt612x15JvjQbh2gaD/wy
lgTMIenXoZMVOzCdWuw51RtIyvtloi8YpsTt7b99gmuXoGiOMnJ8Xj2nZZo1PY/7RsvtohjR6HKT
Z0Vp/qrhq9X7ez47BbWnW+KP6lv3r6WOVqsZbM49GR4rIlaTRaURlVHzvzeW8Tn2xIse4XRuZH7c
Wm63Vai1pz17uoWG7+HpdblgUWDFk1SWujzgJykGOMOTXuNitu+4gkThFMYHo6sRt+53O2Luyg75
dXyTZEj5kq+t0Qk50YF5RzqBF8BQ+zKRmCxM6Ri928dPV8mJlMPrd2EW2Qzj3BBQChJXFWzrKp/3
Pq/vqhtonE85risGTGoy9RyVkkZKWiq96S7XqR8p4wVBvSwYXHQYDO15JJBKM+tIyrMBYwB8Bmav
4fq/RttHsfQYImg2CopZuZbCivDOtZWSTTcyHqAVSRIXqJnr1dsIY91QbLhkpOLeWVEKgoNV0c0D
96RT+hYDLq6HoSbsiwUyETWpN0BFq2KL0d2R1CnWCKJJKvTeQRvUHeIWQww75onr8MgL0wakJR2G
NFjYyDNoMZloU0D7+Xl8J0r6I4oDasDHL3iFlsSVnDBg6A5RreYbrOuy7WiAxj3ytG7Sfu61a92D
dFIPT8FN/kte6RUGKfk37zTeedqbTr7ZsuVuX2aNxxKg0K37z/Xrckim+UzohvPQUGOV3ZyicUhU
6loViMNSj+55ZjnrBCka5JAjJ6WAqDPaxoa2LXUX+bs7plHRLEsmU37BIyGc7IX15+8fuQIrFVxM
FQ3Xv4F+3vab0mnUjd4O3F3WjPL8cC/qnJC6LzlNvnY5A0riwqchIHFwmw1YqNCQde+mCpKS3gd4
RJ+L9L0OCHP2syeGId8kN1l0J1tBi+kQxHknJU8Wovcc5VbZZvcTInRY8inMsUwF9T48mabNj774
undGHLl8L38+nb33KLxNN7LetmH11H5koi2oYt9Re5ytC6lMlaMVewXK4un0XZHfxjfZZY+TIIqF
WynhrSheklTEKYVVTDuYqEY1FVjxsjTQbFmnTqXXiU/Ta/qpXgFq8kbT3YtbpcroAVjNn4Fe9Joh
OMJrpuTUt7LAl9+eGnxH9VcIKI76yD1E31T2kbWTSUPvgixvxRXe1+8XjGV0Mo/cWWPSlysaptak
k8jXloH7sRhgwid2VkCI6AIzISGkbklxWDQ+rcXHGDXPy3SS5il/EIX88WqqttdVtRRyrSkResN+
PZZ34uxjh/UzXSWAaHKjvi0TAHQGAgc1I2YekGVbZUDQ31qz/WkVoBtEfPHPI79bYg7KBgzurtga
TX8XAvNWVhJlB5md9Jz2kcWV/sEo+8/rPR9HkEviPAlKsCRFHqzXOi3ZZKM8dnGpR0F1UDd+KI79
+9rdUVp4Z4l4BYBhjFuJVrwNT5+ox2fRo/uQ3ffo/Cbv6guSuYCoCPio1pClshDh+6c/P9Jo90LC
TvYVMhKlREoAGVU7QDjyJJVgvjVXj8l6GlAY/d31p7L97Q8EeaQHF1q2z4DGUoTUmHaY5mH8Aibi
0pACEGy0DJWa67EL4o4L0LL8RwFfHizbhwh4qfBzXjrD+ObGJI1ZxlQaUjEqc8XMeud+kDL06+lT
n5mwvPIxOhAMUvTO7VeA5cEUt8anv0n6EZTOSWp09MCSka4+x66wjABqJZr6LSgtNwZ0WlLYHfzt
r5LmXlADLrllFjw5znxBEU+LTbyIffHOFFbcjTst7yHqme9HafmgviMwrLzq5DBKRRFy691O7u9E
UaeiPBAHywxSHuL8LgcKkrzlqtCG281K5lNSH0sqv8hky6ZiiTsm2wMTFbxJoMEhJtufoHY0A+cG
V40mNaN2nwAT0Wey/2UuDGnbpc6m/SHsIcbj7GVTYjAyzZ2KacJC6shQGWQHvwpmjTmjKBTDSE2S
25a3Oduq41b/ZA4Wcpp12DFr4R07vZI99EwDvHKJEua7WkEY5A7ID+0J6lQNqdetVOt2yfpkHHPE
skfJKVVve0r0Px+g/MO2Z2qKyLx2IGa5JR4XwPVkt3E14omfi4EgIdOxqSA29LFzgO8I/cIFueLQ
YR4Qo6ISRv0QduZ6fzm4aFjSGN/RBIFyZYEM/WKfwfLOv0vdYZINOPcDlw9jO1WZeZ1IduF9o4Hq
HfG+ufR5Kiy+MhajmUO38ztOJrJC/79uR1GSAwFC/Hu2/tFMelb6vO/6n6l3NC+2XfFNphgMrYhI
ArQBQ4OB2ape6yMtHQ/c1A5arULQSFu75o7Il2EAhxqNpsyoiwwaVqZFXurMKhGgb9u1Fi/Rvo+1
bZthYFu/+nuHQ80RZDDzln/NsIb9T3mKGxXJHCg8AY9JdPbUEFyUAUEuzyM4FbjLOFIeSik4DAj8
iZZ0Cdd8Rt8QwZgGODZxuUzoVXvJgzKaUL3lmDRfoh2aJoEE7TWC4ODzMj87mEGE44NFelnfvsda
B+5/WsqjDTL0cfgZah+jbk0noRs+rFl6/2u7Uv4VVG2Wx8i5BIRAQpyMt5cYUqsQHEM2S1sCqQO8
R+5qv1HcKI31uKEtU6dKkLnaLizXBcId8y6zJYb6HOjHPYPzAQvDVGuNgUGjqREmPb7dxUyY3O1N
1CmlF83RsdB38ceKPmc5a9HAVoPxFecmOG1TGy3byS8YBdBjPBDH0kAB6u5rarvwilLys9ShrPLu
PkZUkhFf4w00MZS79Qe8bZqa1wxXcrsNk6AsfJIdPsR71qphGgbSbFzNF7fj5FD6BkCj0fExGID8
vrn8f0nFxiKq8LKsJUZar/6tO7+Q/R9GVxMgzRZhY8vOlDxw2K/RE9Hg15l1e4eoQxE5A4Co7mtb
POdMxALLSu2mm8KU7l14Fg3Sc8Ut57CKyCrDO/V1rbQjY7Eg4leyn59nTFtG/wPNS08XOiVho00d
Lh8ES3CETmSU7Fz+6DFxXFXUq5H1mNCR9/7qyRbV2vqP4HHDcGwljHDI2c2fbfZBQ48lqXMojFcT
kclZXzAgsKW9AHa6CPPDjnFcxY3olx3JXDEF/PoxjEYtEQsIfBVDcG9tFTkamFuFn2+m0yzcI01e
VTjYSM8TfxZFJUZG9WmrwiQzORrPd4mde0D7ZhnQuv/5KjObn7AffVLGQLKOjUPLokdkkMBm13pI
pe+JeqqluqXVQgneTUURHfdoOjs1WKDOoT66yV4Qf7TASTaU2O3WUSNYZ3cwDoozzfw/QF8+kpUr
xPIdnjFGRYtonxtz2ryUO0Pi1dguxuuGF+ZaXi/6wtdbfEvQQQYVX8hgEhKl3hvkaNeVc9nLBIIb
McFRk+rHuN2XbESnd9Va3a/NDWSKtTY9I3TRqguKwGaAoMoykiMe8J1jDoRht0MohyYJ/sdIdxKQ
fx6kUxwyKov1fl8QEob/lfl4GOdGCYnfj38dL8L0ZZ6fOorA7uu+I+vEoPyPkI/vnPtCAlhKjnzD
GJPi4siSKR6uzVJp32SfC0pNuxEHOr+tnyHNv/p62JTh7ZKD4/nnZUoCZXGeN4Q6FODmCazzhIiW
gVubdQLPNIHEhqqg/VwS+zGHtiDlkP/cinDcbMP7+H2CPvnSJ+biTRpRfzU0ADzmczQ5jQK5dFvF
gtUEkO3szqEB/U9jUwcx/64ZlmyKUjSFYgDUSzO2VI7CJBQNTUEHWT6w0Vustash+qRS48s0uXIg
g5f4TmBDHME4sd/NUNJfDrUFWcUuacttPEcSxuMb6v4Va+dt3wnuxoL5aKOYn6KVtmGx2ndp1SV+
cIiYvgxqHPwtdpflbqNDaMLwLdcrYNFUVgELt9fNpk+oF269xa+YrCiS1vH/CGQG9VXDJNKYHeJW
rOEBOS6rh1HNN7N/HOEl7wWuDfs1I6l76KSU4PvVtiptW7feKC36yRtb3jLPSe+sTdz0TLqb1S8M
/9OdZYs5oisL3Tdvg3r+ztyfE+NibMArAIBCNbh6skbKSXgVN9lqz7X5k8kAaTDME0sFKQ2MKCcU
PDvX4z0KTqx8JSVQCTknWrt/zoknPAfKCop/+NEKZLNMiTGU135D2htJyh4FnS/b/i5N+XPjXaYg
qJhRYJhL51PRgCA47upz1wIF76YlSnLwW/cF8UrTG81FVxuNNrwcSFToSELBvm5WfA+K8htCy3Vy
5SZkp17fP1N3BGqH39iq/seXraIAXP8t8T0MNUyklftTbdRFWND8TW0Fzsys8MQm3rD6k0pLwDC/
NQPqTnyvek+fQ8+9bxKBnF2PzoijbCMs5YFBrazsd6UcNyvlCSshF7Dgaig1xTakjmMuJrVdfJN7
HdJStayDPHAE6KZ8C3IQxcGuP/yjnIZfVmOcWsZGchDW88xm5VYUr2gdz+IQtZ/ooDdGwYpTy7NW
easYpgo+xlLzsWLb3VJdm0LXut7j+w3WKFnSN9+sy1bN5XrbXOD1BazULl7pMh7VmKU0XUu0L/cC
tMP4/SvDffgbazYK3u3MOsKvDoft+9S2Vr/gka+xG//SrERuSM2WRENpvJ7dNaB74vzOCTkXX6qZ
OEZzqpPTNvpXGCt2R27ri/wt3ud9aMipglxFhcnPbFkBLYkBIBpcxwc/ywF7s2semKXQQcKlaXJW
RLxBMIh94XqGS+jTJVbacrUIWD7pKfh9nla+VG/UGnj3Nnk733dWqGUzj/5Fr+6oxGJLLOZSYqfH
T+hrn0AbLgJx7TETyESJ676vSEtnj3VD0KemIrGm92dltKC7QC/lGTKEJdwf+Sl5FArgDKiYzNzS
+kT0qvPNNEk2KqKPg1ReDyKdpM7qPiCy4urxz3g2RdrPYOLUDMym1UMxKfL6+Nr4qZRL1P9dvCbw
XV1tPQq9V9SWfhjg+N3iBGuru/BjRhDjwrwFZA4IvoUyAEBp/NuJlAU5xM0CvtO7/Ocso+JDUwe0
e/+N2DJeRrlKFvVKV3m+SDB37E67eyXFVID09VgYlWiS1wsZOalBzkFDSurQQindAuOYjp3PvUfM
K6D4cqrrAvFiXDUNV9BPSYJSmZzwc1S1a5mAaGbUQtJkbrs1x3/A3LuPyGJ6JvSdMLlYRDGSRUWU
w0hCC2kvPKXmNAyitTRD1TDOMja5bK0cq8MYOb8w9KzZGW8Fu8tfn85+TGR/cfwgs/HDxaCQC5+R
hsTRppWZbklVUhHKVD9xGnWzQYRJXgDUO4wEJrLedWrNTH2LkwjGqYDA/GoLVMWTncRLPeoe0iPm
MlS6vpiozkJo8Jwmh+mueeNGk3q4cwsAXqQcHV/9fOEcCDJhqkpD65QVqZS+90JbYfava3fthoHa
Zwghgtwl5A98KLxl76DG2z78dfwKIOaFu982eI7ayPmuAvoYeSmpca5v7Uv0Nls+mt9UZTCrgtA8
kXB+FbOEGMjr5iyBiEN4ikt1Z5v2rsslZNKVnrUc697DT9ZSm/8/+qmd48b31zWnmW1uKW1RA81e
ss/xhhC2uw5BJvtcWv5VDjRfclwHpcWd6SUYaj5P1PB/tAagm8BG2i+96Q0l8vuZD1A/Ef+ejBjv
aZflsRN169ma3TttJ2JRMgKdSZRhzCo/oURWAsyuIg3q83xn8dRLf1u+fB8MRiroxqTBePQidGvO
bIMI4bc/Nu6acuqe2cOAVI2jG0lpS26ydQhumCvmnPz7dCwuo9AeHp0kBjG/B1FiGJF/BSyt7aob
HNlFUZqgQ2O7eTooFu5RjGoD8V5cqqndpWUO8OsOGtrTYWfDwV8fnpzds4tOiFLgMGmBjxnSUZP9
N167U072k6akn7+ODkdv6G/0yjtSGiG5pm2DLJRmylIHUN9+Pkm1OB6PcSSvFhagxpffG8YQDY9O
GDC+YKR3Jgs9kSG4vczUeGt67d2UUJYN83SuzgsH1FoMnF/Y/vDFMWlSrBOihfzKjYcPk0XBTG0+
ZPHZO5z4xZ2wwW1/ogpHkcuYxwxUMIoUv+j9rc7zEj04dRhvIftfV6+U92N+F8Oo/BhoVnMWEisb
LU1HToPGF+iW7Y5/GyUmHOuOV8YTswZ+U/tulRYuWv6wrtOOc61Pdmg10f9uHL2qKVEyt9N0nsCL
QYe+DmBTYnwbHQoBC8axpk4EAR5oBRFIcUMgbumAj6xuEXpsI30WiW8QviAZzts1/gwrUYoAZHhW
KcHV6BiskMtQYev327lXoqSXfFZyHJ3SdVugj387dktdzYl1MfltdjqbJy6z+t677Ko1y3zE6SqM
bk/cUm540CIKbK0X7PEykEa7CT0JVFsuEl/xfKUI1oHuqDOLzEnuvcNLa9hp4Bn29ROKzWo2tqJK
wJUJJrV7Z1Vetkc/GlbffdCefcxNP8SB/rPr2sGedfOydDRgNlhZQxXkS+fmYuMKxZDyepxm2XOD
j7eVdJM2idx1hYaFQfiL1QtiZRxVpqUKRl3X8ioQ5+EbZ++xZ0g9FCFboUf43qRQaDK+9w3Mmfu1
NIX8EmROgwJhDmqmbIdQGbI31lijvCFEZJMCxJGwr8BJMRr7SyxGlGzm8Dc/wYDvesHdg1kGT6SB
0UY4gnzt711YqI0qqZgSpZu3PxsYIiPR1R555OI6hrGNMUC4EAqMsf2V1l+yfP/XtQfBF1VgEH2D
WgeN5B4e9sT1aDMjqcforqtlqBh+IcGChIdfUsw8Q9sEpp52jyVHaDbe82ncI1cGJYZvL7+/qdMn
z3BsMST3SWTlMGDN4gr5AYSWakSvLuVjgYmQJ4lzWkyZ0P695yqA0bKzk6nRyKJXg7p4naJ4SQhZ
KMJ/6E0QI+YcpMhxNpvmbNwGcx0BK+52BkWqZZdH1vzWqMMNR7w44n7KtWjKXOX53VIJPDp3jenE
y9EKXksllujltUkJOdUPlAeys2IK8nEi6Gik1OfAj/MBaes1t7i3FF/YCcD6ScDMmZF6ByIovr8q
skBL9jPaKsRE3Mry0Ku3tqzWeWVgYoSD8Z3nA9lmNosNB7YKtm+Uz7d1GhKczffvGBKvlOtoJjKq
ulfE+LQmC57oHWf0G6L7XwZqnKrTd8vNlqYRJvXroF7gWKGIHu8JWPamnqX+R4xrGYi5u25ngXTd
bS7qBXEkKy8x21G3gY6bHIxQUlETPT9TfSqua2/DwUOMoJ+Jpek2rgukL3QLjF7Z+Dv//V9ddBVC
SEHHdG7K31rsP6U2OXMYprnlglWqprNpHLOv9Cphw2QE9xCBhK6ZOrFnSQvUUWa1S6A5yliohC1d
CLNaT89s37VsU1kzuumYjGjZKbjvd5wBxxpB+hdQ9pQNZV2xp3Ge7zZxTrUGztOWNJpLhb+PM+Bl
4RvAo5A4xwH0sNeznPFyV+6/RAlUlHpuvzMyUhk1Ii94BzNE2KGTw4qgNaENYLmJJO+5U5K2xe0N
CF01ucYkAaaMQr1G90d7CmjlD2Q5n01eX1KrF+QzA6////o78tNpkEPpC8OTK95zYn8BfDmACeS4
6ULEYsSs9+SI/UxWG/RuXBrxYA4ZZEZomtXSID/K3mdHhKZVenMyJIMKhNgzNvZ4HAhDhuJ5yilO
s+wpVugAlOEbvcP/QEAnr1VMFTrV9+AK7paGvA41NCTvtK9VpqlAJl6GpRVVI1TOgXCkeVxkznJJ
9orFXWkG/umbFJCE0T9wX5H0DHVmbwPg74yOdbXqw0iN+aBpONfXVscVegOQxt/7C71EtibjoMUi
FPLKCdPjyuq4cS/kyGigYwk4cY1Wp+2r+fYueoVdCpzyQiWNsPSjTBjS6HGuiNFINTjq4dC8uSaW
y4PYcvxDxUG3eqAWcwdZijEMSno2jqlyHUZhCSSp0s2WMdGvTBh/FlGMA/FQRyBwfG/YUeOpsFaT
pzEioaJH8UUGbtYJv7qEb6ZyReen3JMAIGpPCADmfzcljrCos85oy9bMe24uUnJJekzYWFXNWmTN
EDmMvu+Yb99Q9ftEg1maNMcN8IYWvkcIxd5M6VQ5Bk7RfDp93+Ag4VWWzhNjYRsYfGZ7ICpSc4Hh
0POb1d8quuDGurlBDdUgrv8nnmI90VO8f9/pPXajySNzP1zAC2JLE/RbUx/yWVCsq3KLFglD3hwl
sb9C/8eYIYXM2ragFeN71eBz7JqIl7idq579jWNiBlrpV3yl3LXUfs/dqM8WB9zbm5XH5bAC7iC8
WNWBojWaahu9umKdhAHdNXEAvKDfEnOPRAu/HviW/JH8JhweHocInTUsrCaBWvG4n2CfT9D/E1nP
SwFsqDDJTziv4zkoLUxmrJtG/cKlIkyzJUrar+zl3cwXPsmXcwG2CKsoEAfxY2skJy9dihuusvEU
DglUg+3bb13y60jrvNMXAsith5EYTbvTh00QQuwzbY0cmwVgjS4kLkgBWpDDOgL9Syisz0d0LbkJ
kJrZfd8k4V0t1HwAqRQamfznyA8UzTXguU8kPB/SLKjWiHuTZokfCDKtHgkhlPRoj5KcE6+tgc1R
gSRicmKbVpRlMmvnSm7PtJxS5tie+9inbvFIjSnqntUFrNL6UgfOzaxJTNHf71Js0QSvqjeliA1J
hqn86cLzxWbYZy6MtwvPuLNDRbNvov2jJTT1JSwYjq6tjT1pNWK9muTvQNvylw6el0KWu1iPfWPm
RymOkPu/HQq9e5CcJ4rPLoGv9kEEsWRuPgDEZqbd8ECkcJLVqZLJRyDwbHpl80jkxXzTDPHiP1Nk
7XSQilvisk5ZDoY4tIAYWSEKVOt7XR2Updq+x2ZBG4uE4Y5sIdOF2K5D/vUP6Z2vlCFhNHSNlKXp
IkmN13QgtPX9FZQr0hDdPChMtYLW0YNjS2RwJc/GGuXBB/ViSEcg0qXVG6U8jM7Ayl7G5wG/dOQb
dZ9uTj/sPJwBf7VCRdOOT51YGd0whrldNmZNetHcui5JvMmmrYnmEAiD31zTtRoEx9DxL4ZJDj3S
LNy3bijpXAZK6nIK8tuv8h6RgvQPsKB/KCdqrdeH1Xn9+x6AHdfx1+HraI9imqz/tVjljAHR38wb
lQoMjSP6P81mrJssh9cKsgdDpbtMWqjJZKoZjFKYkZkb544DD/bOxZaQhl15Wye1cAAagXi0uUON
oCc6K/GeLX2d4ULqJS0sTHkZXAhKiDG96oLWsMXWGXeEKthC78dg51nEN3i9l/WS7T0EYz38VTwM
wzKCSLzZfQByM6vpFbgTOYrkKVNmAicJTe33N2GEuxDIJmNSrmTRoIoPpuUEZmOmH5ahsLeiDF3g
jAREAKrcSvnHZJiwukQ9wwe7ab4EgG9LAvooXPYm/Y6PRGd+iktFexjKWLoenuYCIKkMLEZ58UJO
mAgm1dnBYKxzAoyYJXzlYyYJKN+umaU7EncYIoZX5xTHPHDqAcOi5DaZ5aTFlfGLR7E4XN9Gujwo
pSDAFH8TprbaxE065NidTKcIeUQj3QVd9Q9MAGnf666rCuMa7MJqw5WsZtN3fAyHzIO3tnXxaYth
zO0QsQ/KteJldJCeVTwnziMRCBJ6pITi++teHFkxXoTfDADS33eKag12MDCv1wFRk+tB57mqzhWY
8i4ZS8DSekQfjUtHOvGRY6hchIsHyXUPH5kN7yEk2FSLW0rT7RlJdanknO1c+8TFzrIIVMsR3/s3
cwDvpH3R7r2sVBp+Dq66+Wt0YYlI80OKpcw9ZTbXo7NFO9kKgqfXAY/DsZ7Zp0MQ6FC/XZwICEXu
5fdMo5KDYSDdRY7HwBLi2bIyeVI431t2mTcJMckSFtqhnbwZP84GAzuq+unYaNCW5I5BDccRkgqp
waOe03aYZAYd/Jz4acrvBuFoCq8niex/8vpQuNEyhUJ5dcbzh6ztBl88QsQAn/sGC7PZ5uH+Fqkq
ihZNjTJi7xSrA2e/cTqVeckCAfDdlk4b/81c5dpulY61m52blgIXgtnyrZWP+Z7tOdd+umRwIk3y
eVjK9x5zkOoJjUD/9q6DpLBmOGIqseOST6kHLi3I5qmFW7pqZwn1paeSSnQRgJDuyGGW9I449NeH
D7TCDzKzqpF7l0kNyGHYWwjDDN5Jt/MzB461bg44uQXO8XoPV1Wuh45UFIR2gSmT7C07GhA/Qo3R
Z7sxoq9LgGBDjoBIsVoyleBW00nxGaJ7gWG5cLtahQup4L8k5ZWNewfCDafzsIszWrFPRHNVMynW
TaDAhvnpEc/ovqBM3znYV0PiGjbNx2vlLpZPYZTpO3zWO+3csCXFmqClX0cXjMc+lyvQ2SiVR29E
oRqBiXXSLiGjaE3HaudHhs0d+9qAB/bW1vHj9Fs8WHiSFw/BUq0GKF4rhBtt21tDFzeZMhEGts7P
gGW213npJbfXN8hw0TpX8vOsOy2fMRSTuIlnJBX8KJ/yz2u/KRuHzhgvRibpH+uxNB7qhRyj8kow
mDYO+c0VSd0zCNqJ7hBwWqjVlI+/kp48dz5TCSQPDpYmpunA+00abTe3/mKoneBi5yCw8lb5BUtI
9DqcxFIjtsLuEbAeOlIKIL/moaVXCnRF105XD1RT8J+MhXys3zCnheATrV2J4kVFFhqHWSeMGehR
cN9dKM+lzLDCCEMfzk2h59j3iC0GxOrGl29AG0/fseAWpPakIQ0BZFRp9tCRvrpxefM7GGYDXLnt
2aOsv4WGRMVImsiBBqBSmG3EIP/EFAHF1DSbiPmbLQUmgL+h81Dqp7zJEBU0yurOMcoEQkw5H5FV
4ZTdgVT3/bGJ1Vk93OpQOq/5reKO9n85EfDvOCQNvi0BzCHA6BUL8JIXdNqeQBEW3T9+p1EnUlWa
FOR82i0dBtbOvge0bYCTzrhf+lB2aOJ2lJFasL66e1HYCELBPddLbgEea/2cdNGzsObmJ3TVcLUx
Pe2G/ZAMJiA53tC+e5SFJjP89gNuhqDVRtmy7S3Xe5Y9AWmxtqUjAaEE3RAYp0F5XeRd2uCGLzgR
4EFt/Dgk1ru2KT8N/EJpTHXUGMvggjWxctgoc+dJii+gWtN2qjc5E8alWh3e8bGYpQfDiIGNCO0h
cVmSIcvQEFifp6cd856PXZ1IGhOsfq779/GPvh83kTEf8wf3sy0wqLEA1OgJBkCjASSr0lvVTOIN
o4zFTS15adwiucsWYmBcC8cm2gj4TldE/kkEW59ZLkazIEP5RJfJ4F0Cg7o8kSjDPVG8plTcp/1M
XXychXRPyK8l8Sfyyws0TCz0NEDmMKHRuw0r/JX7ZM2O/xpGktZT2eUSJ3Vbq5aFInus34yK98go
YjMzOAI7W/L63UhDojdnM3zNCaPvrUwqWPQ0D8X30KmyIdGPjcrW3J6Xxa3PQJQFFWwS4yEPAGir
9KGY0F2+8DbGmr/Id8O9zQiJPxRgYEPUUeUNWLXeaxZaWeU3GIkwKs4o+rsoqxZkqu7fCfd0+QW+
sKpCPAJxGol9Bj96tq6GJxuvti/U1bJjze9o2cOaPJsR/wqOPD935Gz1WzyuPNh+YYm5g0VxJMw7
HLb7PGqMgMIV8Jzky3nmnVQ69NNcjKkEFYuWR4aL9s9TvVvQDZYeKZwXD+5SVXs+Q4Ha7vdDWqdE
IAOKN+JKZ8a2EExldwaCCfk9AoNzaLxziAVqNd/XxRnT891iznRHAhL+822N86ywrKggff9f8l5R
1OH9U6+zjStmrsnA7XLKxv/YjL/XM/ghiQHnha6Y8YA6vr8rNYpGs0CupE2oLhhG0Vm7nyGQMVZu
Uo5ygeE0RC4jXV2BZAULQJloUlSFd/YzMNPR53B5ukNFh3ayhZwdm1p9hRPJE0M6VcxrNbo/uJgP
aXdYT5aT8ypoIcSdkcC2Fxjy3vtjfEHFyzCYgxVLw8NvoOHQDKdFzAGC6HO4fcSFha3BPv4q0if+
Z63DjEAdYSGUoXzxwt6BxZ5x9fBH8ZMdPix+0COkMl6SI1TzSXVwQKNXbF9fLr5gWNj6ZuTGMkpd
g9ufkBlxntC0eMCSybNWR6B88xVeYN3w5SL3F2D+8BnxNLzzkTDK9NGAaxw/50YbAUR4LzqFYbMg
QVzf6CelIvkY1DC1XOc6Q/w8ZsC/Vd1GkkrQ5fvH4tZnbGgwgQIRRMr+10JjHe+quhzenxNj0kMq
zKT2qKs4O49KDnDxrpsFE8saKjWFdJ89Mv8v5eD3NnQOw4N2G1QcEWjNfg1q2vLE6EeCwRNh/H5Z
VDftvNTb/72wHguxsmtiG+1dpca98l91gqVi1g3e6OgQp6pHPMvnwkQYyaWrkZCjlf5QxuPMLg9d
b1OFIIvtjBCw2/JgKURvrg3kOOBlubV0/tXDkDphrLr+YIz6ILKDO+sjINAVts+J6tPSuw6PrrQ0
Oir+jKdsdg9+HEp8B8BKZesML8TS3P0nRAD60Dkio1sR5IvqBUVBgjl9mJT1RGfOhnROxWroqzvz
Q44foqZEa/8X0SEODPMntPTNKaPQeBqiH+Gwycl/hlGKUQXJSnQGLl1Bb9e9PliGAC7O+1evWyoe
K3v0/h+GqP3/ms0osuk4zmcmkmtCzKYxMA/YYA2H5f6fawpkPXEfGQOKvu07mir1KjMyH1L4pv/z
ClY5A8uYRywYSuf8x0nvY3We+92bpjXN9TLbbU2tgnAhEhNBHSbpzvrqM9g/ZH7plW7RM/Tz4hH6
9DSzX7YOnNJXMMHSjmyp9+TqBFzKWwRhOzp2E72KcmR2CVtcNvsHvBHaFhA6Jt1pFLEVh7FnP9Qm
/ZJ6P2eviXG2+/pumJnv8Oqhihaio9W5e28aAO+fiNF4YHY4XPMTaIQ2q50HRvI9nm0LX1ur4TQD
bthsmVYFujDLHL6xuE8ZlXQQA7Z9AQ3gflP7yu5zt8tssqg2wJmyxQSMbNQusgw8GYtx773QUy5+
v/g6wFHOVnFzKo5yVZgH8xwWMaZYilS+EXp1FIJs2xi8s5PR6j8iEYAiwgJ/PZ/TKStLC4RB16aF
I8lYROS94JL/lpYsQNa98JL658DU9XusydDGmUl2MHFhBIrlT9fO00u51D9YDUV8q3bMO5Ws9QlC
ylnoEhVkxrP8d29gxh/wBmJYwPhcF/9KPetkEQE2ysHLKoMS5K1R1rXbdWITywhHv3obiMHHjggi
dpfbxVOIGOw4o2pA81tq9+DVQijsGmH9AmD/l0OhD/Iao3A8ObjIhCnzqTIPnyAwcQCT5vnvf7ct
4haQN29U01T4+upLQFgR9wXOhk92VaGtEchzs8WZBpH75d+8SYGCUxYbV9Ise1ck8IpTPj3Chw6r
taW0rx22LNHQax4nox2c0pArVNU5hB7KFoy7BVof71vOWuHYD6DBmMtnsA19HT3vfLWZGeveN6oW
sireDqORuX+sJm+fpRfAKoNeV0zkSQ1TiJ1/mb6PYOn59PWE4o+ZvPkmMPr2pym9dChqwtSxaq3H
Li1Rhc3lKvuTqWrnsSjE8VDO/GaPYCHmG9dTwnmhjE/QyQ1+YiXa0ETkBYfalMkGtgajJfackB/J
XO3ZFsDoOncNpUoi2B32AKnpjHFPn5QmwI8caj877NWjhdS2pxmxWiW/9yl+vtfIUylRlsdHBUDr
3xaZ+N2L6OlfriKXdabl+KR3UNBJclwzfNmJMfYc6L86FnI1Rvfg0v2zKUDrg3hSFzBppit/BStU
8O0J3yrIlrNzYpnEC8p7o+Zg6K80p0oXvB7rcT1aE4Nl3uk7zGWykeYjHU4cP3QaB+kBnt6AZrTE
O1xqkZHLSt+l/zhnNSqHGU7L2I+zTLkeREoaDeOgapGlgngn+6fIlWGaPjtSSpKx3Gk46BV3EmlY
YqkKGGf6jp0Uel5HUCVoAVkElVnOcC+Ov9MHoWcBn6uQkZFd0houbYRt1Ji24N6zTQoOQ/szzI9Z
NNNIHRzihAw2Nmd+YTpdT+h3L6smSjUS3txfxjonwXwWUkj+0bICUrbFfUOGKpSOZ//Xi+u3Jxr1
XJ/OplgdyoeKLslF+lowbckWJRqzLpSxQw+go5mJt/1XoMY7wRac0dergkt60i8jW9LpCSfIn/uj
vhSh8rbQhAgnre7CFA7rSMpeAaCdKbadWwc1Xskvhd1lofd1jxKfrlMuoiRBdz+uk0Y0UOjLRNMi
zVx2Tbctthr9ea0CKkBo5rrlFjQ4Ahsav8kSmzrPrwtmvNvmi8+eBD39TNvlBSPGyNUfAW8AGxra
vKFy7K8os/LMPrmEpsrnRnthcM6lqCFnMzJgvkhoAG+3EVCqdqjOvGsW0uIQ+bzQUmc1/p8c8D8o
NI3sUUB1rSfFlf2Qlz27RzBXaok3lnIeNojzBZhN3bcUz/bdIoOR2S7zG4GAFbcZQ6hCkloKLJgs
AtsaEpYA+hjf1WXoBz1j6b25ImjPfz8/NVW4MIpbOTWW8Xgd+Gj7sOMbZCMB8APx2J0psyJl/PNS
sVZvKMNUqDe3vyy/XGvTu0OY1RP/WlMEvND7CjYzP2j4ap4DOW7OK1knExm3rPlV51c1eYvutI0H
jV81mTAvEfVE3nhVR/EVuQfCjnzIKnwwXxx8vId1y697ppLsu7F4pfbaKIdd3BWXQ/QDJ6Y0nVDc
KpyvrZJ+xAfzsdousiiYEZp89pcqjxZyYXAsv0slVSNKxOFBjD3/eK1MfW3EbRadKbbjLjoQ2PVI
4u14U+9znKFnOIBjn+TvNC5vaycYFtgYtDFsUb6CyH0LP8iZpY+n/OCqKvs4cnI4r/xEfNqDITCF
fXL+K7QP7PBcPndOeUJC3quFeogpzMALeGIKyu1nSaCEwJAGlHIygsynyJhs1rTkuPx5OnV/pS8K
3Rx6O8k/a7mu+MFDI8o5NytxShF/tj6fQLJyC+1Fzpzm/M/AjLLIb6qF2n43hQMFmvU0+160ww6D
KUrJLxzH7Fu/y1F3Wf22gCA8UyweB9Hip9cpTVv1JJeiGzW72bXV6q+7J87BhjdeBu6KCwU4rM0G
9MlWS7M0yapT+NVWSrBKLZTh30u7LJ2FLG1Uvx7dyvPLOqkGatBc6qWjWaMNSLFZAxS9McQaeuXs
3wA7u4V/N7FktvHTy16NFUaMEINPGWf62kBNChaqZUCbZ7UyGuuex/7tDcBC8yQlXZatuWNiDruU
j04gl1Y0tiPb9Tf5pAxNS4FR5PZSZagga+KqbYgwor098L7befVxQm/YMHEOlqeUOmTKGcle8ahU
ucxTHNBFC74qm9aRjUHPOjEhYLqwhVBNecWIejgz0MT3y4zbUNY/SgZxi2YV8rUKOu++1TOWFAYz
azdJ0rIfDXMrmM2S90+TZO4PdlatRb7p+xxQARtFnLxO1sG5fnaQiHIAWt5Oxur+/KA57KpJzY0X
QRTlO3Rra5okzxk2ec21tZ2WiUvW9IBIN++VI+6xf0tGdmj578YqdyPzHHyYYN2JX9M75JmyGjA+
x/+RVzYMi/bLx1w7ug5egfHL6tYCrpo8Z03d/UsmzxamoVwyatz4of/EEOLS0Qm0QmYjvvLZBnym
RupLsaMM0+p/R3tEFxms1GjJ9YaswjMlg2DBaSPvfgVsOMSQYgAajGE/DIuDu4bXvAW9ohmj6tPf
EAi4I4Soim5hK+gdJZkTre+mcG7euIJhfjjhpZNqfWKZpNUulvTeJbmBZ9NoobQnE+ZQe2/I2K7e
BvEXyk8MfQjYJOv7R0yQ5BcwvXYIxXWBnumIFD47xmnravhw/KD1ZaxF5pni82Zz87haMQckKCWz
dqyy+mGGq2LWHyZfAfeRQ1c+37EssXh/DyuLIdC3H093h31QM2LVgD1Tc3eKWtih+fLHWG8RvgLr
KkcAiu1MGSGYCM23e1GXFiS6WhlvpHzfB8/nvlHqIR0RW5g5pngfGk+R1Wz8oGdYfHtCIhAzaE0j
xLJ1LF991MfgMB41IaH8j+6GLGNtsIoXWHRDkjif8RlyE8QS3DQ5UptrKTgA89qJPlCQ90aDHQfR
EmEVxZVDhhwMkumAQcYTjw+Nu7Uy1EomjJ0vJ6wwchHPiM8TgDQmFNs7z23cyz1F7z0suS6GNF0/
ux7B3wVBu248m8pg78IYCnEYsrj94Lscs5usDxm/x/2pXqm58BZxszHhxQACjJ7f8jTfV5NqF1CH
zDHZaDhFSAyquCtDYXSgbDyY2hBcE/joWpJ4VkUwrrm5gSAqnwVrpmGgT3WaLyw9puEts0IVtDbI
8kWtLhl91M4aWa40F8Fnmw5sn//W2L2QJKCUW7lwi8XtboQ2rF4IiHkLwoaUigIT6+aoUFf1UuZ7
h4FugzRksJ+ulKTFFXrqNw+R8xuX9PJDLTynlhKZow1aaMQdQyRV78Qj+7hy6/uv+qy/NOqef9DS
Yv6gbYXpZ9+e3WxRcqEuEydRyUYJH/np1aErJ9aTDKd8Ve5rZB+DotSd29giaItCfHxU06SS48pe
WAr1nacj//tg0JYZhEe/38FpYaT6O3/FVzzUwZYFV5i0Bess0BplffitH4tZxO7IEilE2D7OMF7G
2zddZZf7bAmQw1Bsn0AImiFD7az2p2u1e/FhKou1Wq0ZACcKyQ5zZelTC9isnkaAwydfvSH/fBkv
2ki4VDwKGXF5XN1ZYkHhPWCEEBNTz63TNOy2vnR/orBBw0TV5iZqbV2+AtuHZicNDVorvTPpRmCf
V11mWHRKDw8i2wJtWMNM0uQ55MS0jpZJo5/Esmtoi86CsFwV4rRWZmV49tjPYDmRTHVu64TzoAYF
dkzglJaCCbQ1IShwm1VO4KscOzUbnBmAjEo01zJR02ue0tvL7weY86f+ifsa/RJuPwlSj6pjezbq
JSp12wkqqgQUXfO8dknw5tuStmiQ5y0JRfEHUSIqhW3vMqKjZRBrRt5loAOrDATmnt9BEDWe2WGV
p0S56Ggd8mtsws9ZpOgwn57YHUzqByx/8ziTQ4yCuQZGxBQjkuAOqtUni4XdSmflzUtWVKJRKsQb
tEPJjQ1iyx06zpMg6W2wgHFuxiAO4oSCSJnmVx4T6XhwCvntVV893LPmfzFW7Q8LjdMqXyFoCzBs
oW4wrB4Uy1ejw+1x7DAvwlh85O45fX6mDA7oir6tAVuGvWwRdcVjdZnGnsHdOhpxoyowX9CBwad7
RViV1Df2cGqzQ9sM48cVNUbN8HmcwsCPOPqXdrUlDKAnXX71DssA5bqsywNtzAyUuzlgERJO1qio
eq2UYjdYhD17fbsNxFPSkhRh4iMlUbivRlpq7Y+MxYwC3QzNgWMfedTc2/oedozbaYi7i8mPszA5
ZeMAgq7TWOxciFU4mFdXfnY63E4LWQLJa03LS1NT6anBjEL34pOLMoEcwytEdZHTtTWDODPzZ+kZ
1Fkc1VHvCIyTJ6w6eWTGbjH7gr3Y9avUXlASrXoB+eSRy+TfWAczWD/slGs38gaGhR3XgzJaJeHE
HxJpRoMQrOJIvIafIdOqKM9/txI1eid11Xj6HFXF9XSCZt40nxhKutaOx63TExvcDOB7uCz0E5y+
rCTegGrHWKFXnMWK3JFG9OHXMi3UleMhCA6kwjZjUTIXHiVO/elj2fspJYb1fhIxNzX0xcsMZ2v4
7tkijQwW+y8Y9IdsM6sUoVn13FxEP93Jii2p1ijQ52nIod3cLboL+sr2r8zEn2gcaStcoR8vtsHn
EiNZkwc8F+YWTcPMRrAO8yJpaWxLj6Df9G9gYi/wk6upkv3LlLAECiZ9OjtaIgbwzLzdaqrE6Rju
d/uEXrA8VOH3GQ3DFENeluk8ES9HMm+Or1cw760fdGojiIZQjNH+BvQsNb9mNQsg/GgIsO+85Wqd
aQ1h/bb5pzEwMyszNrIsi8RgQ8YTCAgQiCYMj06/AKFForbhAxAZHrWD7+vdy14wUldYgvIRMJBm
WIzt1lFUs3kaTbY/ZsO41MiDrobNaiS584xA86cALms8KkNqjUXwJfttXziYAyaRFtCbn3tayiyU
FDz3LSW/slEvZJ0HW0SQdJIxz0m6UUF8hkGKod3CWs+avQTyJ5yKi3AXHBilCgtGObSczMarQwMH
CMpUHznkYV397lx70pr/NjfXd3grHbijr6KMnI8tRlxD7fm7S7Bh3S71ayJ3oKS8B/tenVDsm3m2
vgE2NFhxbQk2U9MiRG7QZmvAuvJzx5aBMTex4XaB3DdJxZPllGxpF7GH7MIrgP92FHWvMBhKLVhN
TYKUvHbelWrDWO4naPe8MSWS5RoT6bXkgqd4ptV2qU8pk5GtnnHhzql0jOTxlQsu/FLLW+q2Yj0g
gBH5Ao7/VyW6SojzC+X0UBYnZn+I8Au7daxppMJ3kLC8YHmDSamPHCZ9ajyLK+FtVoA3nb35gavL
xOcMknDHUzWIHL8UD3Q4WtQTfpnVXSluA9xmM7U9byYR+oUIcpfPbELnLVhcER5Pw/yVjoSLNxKW
FN4/NCkxmkNq4O+u8OB7L6j6T8VHNyW3qwjDAkntgKwAYk/HxDTxZQzYUsoGMK1omp+P999W0gzZ
tFmWCqEqmgAV+3+/WN00kPSAtsVEuv1KgsncNixjey8UKt/6yMgc4fS8Q8AsPtyXY8Cc9iepNWJ9
+g3wVMos5BjOWhojtR5jBjdtIDdh93IzLH620NexnDoZo+acBWZA4c1xHCYenVMr1eKGQnzlpMAJ
qJaAOak98BYaCLVo15VGJm85c4rAeEvagF1/b6C9gN+r2/7daLBODb3/plDhzdrTtGPaxyA/s0A9
6Au4oZWPFqZsJ5zF9IcWOx32HmPmT3W7DVk5GOdK8GA1dcGQM59tZ5wZP8hoXn4Btc5fFUnt8KYB
rW2qNIQ2P5znvnxJ1eP0IMUIv9QvU6w3x02Hz9+2163As9W8eBFu0JuhxeVY7JaNPr2a+Jljy0RO
TPtMjmxdr1LL+Thrm43sXlIjX8LjktLtNlMVgTQZzgV3EP1TyfRiztKvY+KqlC1uuTygThld7M/O
KTDXD2LeyI3q1akMWRNTYo2Wvs1j0+HPZbYuqcfXm02RhStPfI6Sn/nVCAYQZu6lcRvqHJQdxy15
TUMV+wDq9E2SxVo8ZYmEUOXAwKSe1a4l4Qe56yHZ3n0ic82nbf0qncbWZyasaM7fXkN4TawTXjEQ
fLO4v4ydJYC8R2BZ6zd9eAB4/7clZcVA8zdQ0QuFN8uT4TGwxl+hmG98uZhUagnPTeQen4BsTTrk
2pm+yDuMB1i6p9lWQXRRF8j7ubr7rxM8b3+oSx8MHgF/TEMJswDUGnqUs3Hh9C6VxG+NNwvlJZ/G
7zki9oxs3B+YdkW+/jaerg4uO78va0tSka/T0oV/rb3csv5Dp1oFUBvXbuVo3GXLpQxikSAZZTiZ
BDUEcQXxKvys6k+SYP7rbyNWzpNME10EMz1CwlZe2bBD/DK/C9PLpv+8+AXTjrbj3jKPZ8H+nVzc
mdb6I983cKDP1fyP6W9PmihZ9xLCekBQPOR9tbGizvygmVr+bQPnvAx0S9ksq20UGtyaPQRDp2TQ
i7k9LwKuSpVI5nANm3HGacJmM2xaENBs31XVjR3TJJ5kjKwStL+IRFAp4J82wJQKsdS59QhLmLdM
4BSd3Lymes3XDBvt9JB96BgNRiv0RcaHlp7g7y1/M01WhLrJlpLAS8RSaFR6NoZcFFpf/9kM4VMv
5iy45wyICMADgwAWlfR7iRs22yUynBYqe3M42cRU1OngMJmnucoceCS4r9qvUChvk2cj4jDO/zTg
ByEE2eYrj2lCsBYiFr2X7YsN7PB/bmamHvHwTIl6G9Ue4joi4uZrDkYPl28pI+BUhbcGdFvBmc2f
/fXV/9CTfNsvFOJWg9qD4S0PkLw/LA0HfJ1E0CCJ0IwiJxBEsET8DMm2oKO0G4nAFFz08BBEsqOe
a4WOG9spXedt4o3P3A+EdZywkS1wiK5QQM2tzuYD0L/JIJ4x9yNvjV/CSX1CaSq9wUEpXZtGPBuY
mjDqTHcWkLmiQBhTYxDmaX2xi/Tso7d5Qtz85d4xV3CrHK5MTJ/6D0lQAwf013mCbVwYlAjRCFSw
3Jv06THWsU8zmHPsQZASjnuBd2eLpvaRbd53m8nveYjezHcy06KKRaKw8eEM8sn6xElot73v6ULb
TvmmRsvRGBSPrgJlF41r8VB6sIe4U0U9t3eKj/ISMjPGEktaWayUri02ESZ6ln0Kl1sY/Dme+bVM
jr+9WC5iI862i4ZVJOOrZSCI4H0D+0lmGyohQteWqZngMAsfbP9jwCEw66vtgtzO5Pdgozv1Blnp
ZE+jly6niibABl8509kmVE8Ez2NOoxcfzpM4E8Rtk0lypoAhbhKRggGrb8IT+Bu201i0R8xszfkQ
nYmYufGIz0eIDagaqt/C3+1zzBjrTX0wnF7zHJ2idXHEOXRN7Yea037yU3LOK14Ub4obqozHWqhn
R33AZcnig/DvpXqUg8KXP/fq298mwFBPju3hR4cXDB9jeaL+OZbkKUANCRyWfN1rMOIdjYZok35f
dlwyIyGjRJ7cONji75zAMOtW0lKn97KH0p70k+Jym7M7j21orB01CKUZYVCCgUoaUNYKkmUd6n7T
+4fPAMDDBWK0uxCMvp0y2qp4clJeUuEKxjIccO/0bERNVxp/VbNe4zIMB8RXM608nhyDsyLzz9AV
lcO38o2PpjLmF+BYZpmR7lFsxRuZhS3+9dwkcK/z/5DeLiOIP7rZc6ECe5tY5pkwABLuXjtWprI/
fHhf05/reYXOcQe0EIv4gdUYyrYcX1z/qhMrnN/bcWOcjItHCnRIHSUQZ/SYDenjCqYEH/5hGo2/
vEQwFzh95sWQOl+TX5Yt50wVcNip3y7e4gE6BmXUxeAKI4jns0fNgsGSIkOLpJEBdo3GsnPnYgTR
btU6629r2y2GjaijRO9TZGPsbZ9x+EQCdl7vfAUxBOn+SL8zFf2BdLWWXdrQd08Dm7DqKBwPQo5d
x0y1gFaj/vw4dkkgozNR3Z30sB+mQFWPyfXDKHXOZI+AI/LfbJu+1lw7bEdnk/0SZ+ESesYyt+Ux
C4RPDrO32w1nz0fVmLhB6R9AIGU0AlVl7T073rQ73v8xrF+m0+7Re9kgusF3PaqSeXbZLDLLNYdT
zLN14wkb5tjIVX5dGXueaodyhFXB67XNuekbBNcoVjtqwm6W2hjaRs7JaJUJwex4Yx5Lxp3CvIvB
JaQmbHJVZOHPKGnyI44zDmEPScwmX5D9+F/Vz2XqivaudJ9u0QtF6xkgN3L4sBL/2cYgwrDpzHiR
p2UJ4XfuRaf8qhaxP/PRerVERUBUMDwYjiuPAz90urj7W8+W7+RmGgGCBgEsm8xJs3l1Au/T04mM
T1kP9fpCi/JwWuoaDILISJ95XuZaGePDVZwYq15ZzX27wAKPn332lxIZFfiWtj7vqJDVVJzAPonr
cWW8z5GorIZkI3xhOYy0PbO+poed4vPrwWXUNWN2anfnG5TBWkuMemN5emrTeD4xiM7d8Rdp7ncP
58ZYkIYwIWVMcP1fKgs9maCXSFqTda4TvF38FaT2qaoghMzRyngIJOMscg2lgxooM83E+XtElKrZ
eQlhAhsCdMu52QH2xvJBnxNwwku5E7k04t+9oxWgnpl0zWnEkBmDHmN1FAnuM7cC+1gc0yGjtf7O
lkoyNfs/E9y+MGBrBmoAyLBeAfKJjL2DMc90lr7H/BURD/9OdLuyVpGdWEnLn7X6MJM7ivG/ckX1
tBdDCeozB8/n35w3vHrs9LRLZTBPjdLrLZVTN+NbKYu3IrJmnMmtcv+PUAGyTr2ar65/xMfUwpws
KRsBYrcP0XiMmw3C5zVUF289zzRp2ULtqjWKqo6VJ4aicgs+YoJmCViuJdml5cF6udM8miaEYvvk
xOQO9gxGCwP+v/n+R+clcs43iv9JIKrlAKJ0e9dNQAZmrcygy3dwYYU55jfiJOLG8CxpAQyCzuQg
dWhvLWYeiQOlzn+//A+UwdcDnf/ZhyoVt7xgpd/g/tzX4vlG7qIMudXlZvywhEDLwoqAM9lPGNFK
Muws8es8m4uuazXTKstN8HzU++Sp3MmnL42lSZp6FQNRCcVYQQ0TqD2Q6UFnr1FfWzXodImfRNDm
6gqZQ8bKZ/JxmbPQlpE7fUP0QeajTuf7m527t3lOIaES8SktfXRRM/vfNWe7KvUbFvqjh7qujzXp
l2pW4nDxejN+tlwIJj19/FHPWSPhyeP6Oew4geApsoozNuxU0xe3YdSAHwlHW4DoWBevPv0leWpY
xWjGMDNxrNI1yhxUlQ5lsSnMIMTChEj3AXJHOAV6KNN3LimVtdN4OMxW4XFnzipm7jXpYOG2P8i1
5Ec+byif6vT7e/ovp/KbGrvMDZ2/kgbGPJtsEcVCLHKIMIvdoCnYVG6NfGGzsY8JiHTJS55iWiwX
ziNfVx2ITicdD09qnZTOL4kUNQt96PRXZijtDHYJQmeaIe4NDJAUg42+pV7V4XWAm4cAFW2wLpY2
0SJCWswOKdG2Da+G0sy7qyrCmYiWkdYy3WkMRNC8ldZ2LMPnq+Qu4hMdQbatP78IpM/7CS2sVsXD
AWbHl2krAjcw8btykhw8MG++1cL5z4y0vWLmIFOf7S+z0NNQnHNA6KB7/KUVg8Ht3Q/BgnPRnK6s
ZRPuSOeIiHSpgu0Rtl3vAJh6NjSHmVyklpEE8C5An7haMKXd2KFUPPfib48sxAUYC+VK6RYyaeRw
oABExVCxT2KvnTAdJv5Rpqqp+3+0/yuOW+6wAEKiivK4SAeC+1xQJq4xWQE5/RXgL6ZX46MO86N/
gao7Tlhh+n+tfgTlSzJqWSjosckDETWWiOkzVkFcqzOIothIb2H9I5QF4WtzH/4jvfpLH2ZmjCQs
tfRQhQiQIWfc22XVHPbQZjL6iCtowEu46B3m/01y1O0Z9sju/Xo0aGUfEMyH4hX+VTC5AILh5rxc
B47WG4ezo8p5QYnziOawi5817UfJr9JfrOamP+gHiZbuu2O4NKpv7BV3iy9EHynYjEq29Cj0WVrh
jCpNyPdSKTmYEi7BOZZeMpbuMOcXzjJ/OGGyhCy+kVI/X3FSoh8w2WPZvg5zDtS7YNTSC8Yu1leg
HADLGPNxPVILtXw+0k+K72HALR4MYy2hM3HSRSefQP5CmBiF+OKRDcl8JiVIA2J9duk3hDGEmZ/e
qejKuajXy2GU/LRH/EFfT/e+xg6QTZpBEkWDXnx3roNKmSNC/AhuOtv2yaY6rleKopeT+KTpuGEY
SWBr+z9McUxT7MbLcSqs95TTAuEG5Ce1uMX5CmUchLjuEDaKdkhxSpmgPKFwWi/H4keIPycIz+JU
EGHJiT7kxmcAPZ2maC67aFWWiBQZ2GB1clOgvNcdxI03MOiMFXh3HU8foX0waYebq8yI9pfEMDSJ
jPPvZsUyj7yK4nsS9AFGxuECWZKk09oChEvuQ6vYwQfqrkgrqS9Q8D2jfrSxMF/or9hG+Ih+/Wg+
0q/xrSS1eWrr3BCc09dP5RuWmZjpUOZvt0NiTtfJZrVV0XiDkCCv0HixhEv0GEVq9tBoS/XI5wd4
6V+9xnIkKgkOywI5hbPbHxnMV+TxfttyunKO0gLQtgAWSuEZ9rpFlPrUsYsS3O3kLvTG1M8MZU8+
O4KgoQCtln1zV6S/rddgKs5FLR8EulOYWK3GKw08WdUNmDkgQmV79xFbmGHAWYDrSv/zzV5+w8Nz
mLX3Jza2eMikaeP9RJMIsYB93GCqrOnpKkPWM3VpX8iMtgLahwMuZphYjOAQomF4LUhYD13Hb6mU
B3xvNS/LVRiQ1n+A321urlKe5rxgLdozsko93lU/eW8OG3vQaXV7/NRS5rTXao6C7bawTbqxjUPC
y6hyhq5Env1tf7nquuVx1exAYTk5DdMs7ObU4AAzIfK41pxyAj1JKLMU01qbsasWnKKme+m2XqHy
gdK0RU0h3lKx7AXTC86KNOImDFgh63fBIfT+usEAg031SCffcmgwU7A1vllKhtBjC+HhW+480lSV
QZdPpAUKkYRV0Lw8U4fNc8OwZWe2fmVqeh0bBHUgx5DLV1+iWT+raOMhVOzRJ7vHOnDaG0HltA4K
Bi5l+9ZTsdNNdoPvi92ZIlIDyvAzpBfNrtCdn89B29WXc+pp7WKie5NdR4q3GHIGDyFIA2QGNlaN
JAjAia+JXv4X9+FdgkitFHfZSIRN2W5UwAyrJ5bGFP+So949EkqEwdesSWj08D8+AG/GGskxmh7I
HH2Y/WPxSYE3V2z9BQFh4ndZEglpktaN4F1WTXG8HAn9LSrU3BJpxjd1nIaW6268zCFb0Ro0OJrj
+TrDkpwF78LFH6WkmIYjGWfxj+D/zeeMVQU5WBFI1i2oDrinagdlhZ59mWQUWKvvtz/K0DPCCVAG
M5ZnaXGzamkHxL1wXWY7v8xEpALnU1g9QZDfPGGalD+s7h1fywCWrcFhPnqWSCPCWAQg+6BsX//l
yR89g4MRRAb19oY/ZKMdMLGchqanBikWFG7lo7PWMdWDoitsJ+L6YCd2qND6QBSEGOOqu+quvz12
sFVubXnLpQM3JmO5rcNKbYow7vL8d29iqpy//h7FCS9NGywmetFs6mNS+GU8yu8pgDyFinim+RJ9
Eh5xp0IomP8zoDvgf4DtcwrQpQ+Oq27yT0NMVbVsAZzbUCFkW930PQqiYuFpaanfXB8bTWjmM1rd
5sCFeBDbpD5lNf+HmrqXKM3sJLZwgyzxEjo0kjG8vDksydAkQCkIyIYtW5wkDoqwDL7UYJm1r2kL
QXX+al7TJWVy+1r4raJeKwLGnExSSncSySxFFpUD2vTHC/qJsFBcTegmBVyIDUk8PxmOzvirqotB
bqsl+PbDHjNjXcENlfn3ymQrc3j3uf93S08ySIVmAgqbo1PcSjMirVhBwd5jIOyP5w42PKhT5Zt7
Z83IO5tjj1RcSLOHzer48M/7JiEVSAJzYuGgHc3pUgJyRaTcg8/PUHwrrJP1ROwxw+s8eESpweFZ
clKaGynsan9BYKHCoPd2de7Rio3Z/5BepEaGgUFMZI9jOqeUiPB80dCHMChEKZOip2a8qB8mqmFd
QtC8Wr4s61n1WoOf+6cjtK8wFcWOhQXJb9kKJa+HGcrlO01lSRhncIyPiJsLcKUMTbpdI+BE1RCx
SPf1uB5lDwzzBEO7crIR/9F6SrO/tfC3YGxh+7np+Z0uxKNcCWWnBBdEyjkYFoQpiJOAaUFmff/G
BkdOvlX7RMoIhfXpZRFhpTRkRg/U279XJ8ZJfJ/WjcorVYRUcpLbLOCqLmKC8aLfI5W+WgpHlMmm
V1bfsFEO+762+kuSO7czAkVb9PxUSde0OxQUQqILcLEDYYuW9K6l14Pc2rardFjVUqsAT/FjH1Sl
KzAQm9/+G7JN5IOSr1n5G1qbH1DCOZdpk4FfNi0W6D03W6fH/sNvfJP1Hjl1gmHhHY+QILBeg23R
4aqpNEE5P2RFcQDX3Zi9fJXb+Cvqpjdxylr/RkXPoCAfl5wH2+ls2ew5GEf/YSh4oq5eJRWR7rNt
hAdHx65Fx4sdmL5s/idqioUqWBeJ0hPxoCh8cPvNC9yVQAhpRZheiRPV+bJ40cvNPFaK184Wc80q
UXenRmRosCM8ByzYntHWVzsymAtJ0jtGSR/YaghMrcze7+tXJXa06Z1syxiCeBIY9ANhEff7YiEV
ABO99Yg0F+rosz9mRHkdN1iunoHNglz0Z9jgv85HQKP/mfQDGpbbr84qOfqESg1iF/VGsUU2NYd0
ZkGWnQxJUiCysedXSYTLJ5cKfyPTR+Zf++9rjlR82VBtaLg2IqMPqKZq0UTH+GQLW4yDzxL97mh6
2emw1bVHRRynw8E+arXJsUgj0L7Qqlhf4tr3WQZy8+7MoDna+dmAyz77Mrf07Dix8/MARKFxsnaE
8DmRVVgxZuEv/BS+pVjDzM7prFo/Mp52drxCmHiC8dVt9iOOyw4YK4JB+8DmCDDKERQwPjqBAPwv
bPaypvVwz9a3hLKJ5c6u/j8l/mijfm7xvN1irh92Uckc+o1mmNux3kLkdZ1oQaAA/l6sNb5Vsp23
xZHfeS8j1Ufjz3IsRyL/oXh2LJYn6DiE1zRS9+Z3YLe4gnzZ+Lg9zwL9e7y5bBuE5LGKGSNuQaMg
4MukM91AzoHQf/UW1V053jbca46BDweKcOvc2TN/ZjZWVCjpniZ1rucBnCOIzVC2GeGoXHZxSgb1
JXTa9iTvx71MgJ31cA0LZ6bP4B/4FWQRvUGtPaxmZnSG3+RXarUeSVu9rO61VkM6knQ4YfWB0fZh
MOyfsdIPig/634TIP417H9+il6GRM9X2xoQIhJRBR7E2wUY3miIVSu4ABE9nJgRJ2mzB3R6hHQat
vyyVCIRsQz2nbLBPBFsqtJlSNUqyFYJqms2iDhNSPiHOJjMfTDtzBtmuwKcKuM85r7e1VGvnSEDs
oCOm1FXSwP1Hme18QKWUCSCLPuLa0k3ikZ7RO/753bvQAD0ZV5p0PSTuT4SM4NoH9H33TuTgtwTR
ESPVhm36xqHu1Xb67khTV+yeBbReA68vZClOgDrR7gnWXtC+5wMl4GZFpfDNRhTMgXW7ex2DrfUE
hXfd8yo/vpca182FWbWaw3+V5xDRY3aISgYFMzXPQE7ho2cPfUTYNvIzd6dJmX9aWKFgDyY5eIfr
HBwJgtwOY3snQOssX2E7VqNqLD9XiAFxd7W6e3EAMYczh6NbMzu/ElBpditGMw4OOgOOY9S5qQmE
Y3HeFTJiHpzQ0v2m1oGyUyBEXhp7jJ8zeq2Dm5aAtEP2LgNjoKyedSLXPYurY+BA1Zh1t78B8z/l
6Q2Sca+zStRmI/bTLRwqPUrHmjHVYla6jBwUVjwnxR3qHQEWBOdhdoDVgdoVFgW20gkBLIEko8Jg
elxdEEIASk7vBG7S46Xp7QpgdJgxr+tZFo9GngGxY/cg+YKMP3r28GeAX06w6fysRczmDaYN8M7D
ItkuWwGXkR7QkFxYlz91mCc4SNVFOwd2Mcct9RRyORc87M1/Gij//wqAf1JZMpDwEbxF/I0sz5Qj
xgtiL/gvbhGswg0eq8KCxXcr3nUfCKoFVfP7x8d9k1K/QMnGqG98KTp6fxkYiedFIU/eXWCdfVGZ
vrlNAKGp9nUzxAC1q/K1lm2o/9BnZB0oWj97HNZVWuWxgFlCkmnzprym9S/B+KskJVAEadoc91yL
1FPe3cl/DC3RsPqEWnUGHUkaM6sCXFRXNVhLGYeDvkoK+HteHPp6B2nIvP6E0VLdW85WIzB2GSa1
0x/XmVL0jdwBoEi14VnltXsgFBupibmx2xmhhK5JPWa77s5ypCYUa0ePsP80+16O5DdwpQHc30RN
ECgssqYsmYK232PTVvGNZN1H6/pINytcLQWZOOkJao3cDvnhilLIajoDz+O5JEq4C7OwluknTrdK
izW1oEa9y4fYYP/0m86dAx4BgWOH8c1QGjnbCmoJZ8g8aA4UeHtXMB6eh1NtpXO2NvpfcIwtGviV
o0DtDjFz74l46gytOIxX6yT/lSz/x/XwctL8ASfEyv14wfEDu5ssfVBg2SgneHwGd/ZafqX93YNZ
1McC45L3NH7H4sAGjx32qY8OCzK4lOP47UiNqG00nvt64qNHjXnYkfvw3pMAx6w20TJ5muDQPTT8
Z5oVjLeWfTm1K0PfjaGtyZt+NlN6xJOtGRCJ7tvZ0Ssta/lPBssdIF6VIi4L91cK7GBX0Le0lT/y
nfabI/tcF8cw0QAZ4++6YtTZA/F3XTLez89M+Z6FVwamhibYEZcInDbV0ohsy4/e0HYo2QHOPeyM
KS1gDsXrwYUHUjJhwl9Hltz3BPZGpLONTvka84BK1hiQ1ziApe3SKbgFvGedVbnn0i5itRxJpt+M
DPqdO791VVbCHLCnwLLwPYuqMjZCnRbbTfwLzy6ToHZ9aWhgD+J2CdOlePPXCskCGjjidpi9DpiP
pQDY+eGLu00dqbRbHj+M3d0auytjiuPlb+UiWsC3EmxaDoigSIPNLUw4SEtSWrhtP6gVIUpl813h
egbiypKf3G5pXOdCeYYAvaEahR0YL9j8/hwawGFUAr6sJStNh8LFpVdI0ZOzX6KOktn6fEVQZDOP
Duns76NdEWVaJfnHFqNGM91nSendD7As8q5LdECBQoJ/2Wnkem3thTT66iTLchp6Z60OVYBTX9uA
zHKa6+4qf0DOqsdH2ee1lQkljUuglc5Zl2uPaxtqnj3+ppvTJKYLP5hwBqA9P6Nr3Oxv+PjC+wi1
WfaOKTFkWcULwiQ136sI4zLmn7U246EEXoL+ETHvAqOBbZBGCdNrIUtPrMYgSGAvFzIvRnBOIPWs
jQd0j5ZY8X6UrZzoFByihtach0mIVzxgBuHBNoCI2NL5bOf1oiZ8RVA0SpEKiWJsXPnKSwwK7Gin
pCv9ro6vevsD55HZ1ErdlMUK3Om6H1OcnJWnuje3ENZDgZqkItG+tv1dI80NsfMeATI+gc9aZgXr
6w3okDWezZSTf761G3SP5LsBIMidulLWzLGoeFqqR7hcgg+E6n5HFqW4IsFf0jqWHkS4WzTKLtj3
j3YOholMPlNQvYztFBY0LUD6Ru1O1SGS1LAh3S59n3Sh2j3ykCdZnd0hLls/G+95852RWuMb28wa
inVaXbtv/07Nln+rAwFLTd7ZIeQiJE3Y9OXTyCQB8vv1neYCsLiHvjwGyYTQeA/ng4QKZWAzYLyB
XUtUCiFfPjy8upyf04WUy9EihywlekaBQAORZdOschZJ4HOn0RQtLCp2wo+T6T+lHpYcP2v6CEZJ
1emzwylLpymiUnqeA16pLw6Ik0QcNbkFpU5FRYyhoq7iQWEwGF6mJP9f3DwDN7+WdVfIWPcrwioi
nIjQPb6qjdTcU3AYhrEBQ6W2/GHmLVmtQBlE5LbQZ8bfCC1SbYN1u3OOiAuvJwNsWp+5PZ49M+D9
XWesZ8IYZko6QJeHHGigi6sIvZrwDTAaNzYnmcr+WzHoQFm/X25LnopaVxiIuW33vLubwYJcQG6w
qT+9GlWgM9mDvW3iq3klSOBxbbwEp0kZZYpVlkb3sRJELnoLxHA8K++MfpH9Afi4HegjpMMDoUG+
Q4g7fE7N4Gekyk+HreAZdi3UsOfueUjtVorWaUpi+aFGXYzC4Fa/MafcQJz/JSEf2hr8yusUyUuE
FkFR+TmFHpH/xA2ACHOPFJrt3bfrnh5PXyzaKOjZA85YWoRuRtvDflx7NU1MEAdDRBodgQlgxV0f
BJcgcE1f8w2/EbPJaP1M+MixFr85VsbIFdyKXJQOfkEC0zdy4Vx50pbcSIpN62seAXDOKqqAID+q
5NiqZe1ksW0BiSDA6wN9uCLVe/RoyAYWw+9P0QRocgLho3NP4I2P5MeDBWe/krUBRKGlpmyXGIUM
lN2Gnpop6Xn7aN5UiWPH+Ru69mrt6LVpd9LVd+OKPgggwu7maTVzwgypbot/BXfbF61vRzMvb6jz
P27zbON479l99QTdlMSDwxr9au6n+hTqh86kK+YWNjt85hhg3RLZ/1u0obqL5wwLyWUU3c5/+OFS
NbYlYXo5+an7Gh0j0oYMK3vSpWrecCUPcAj3+rOMI4vw5+sYL66yQ3zZajaOPw0v1hFlaeRVb9wH
8e2W1cAlid2OOtzDJa66LYaAylwOF/FZC/L53XtVP9x6sDwBFDZ+aJkqCRviFrxZJ2lwJk6pE+7L
zCvoMVtfNB2zyWFCKqY27ZpBm0rfTYlmgvl4xpFAQ10PyL1LCeq7DbjY52kcVl9ziN6wcsDuW7iN
p5K4dO5zsanhdXdeHPT+w2+W3Hg9w8G/ngMdOfq1ya49r2TOU457StkhqajTlz9a2itGN7xV/mXg
4i13+7zsvphLnGX8ZzNQWZk3LYc5Xqdh9r6hinT0uFcN9KhE2iahSgRdlbegdLrHKigNCAeKXK91
6hYHMiuEqvbMYCqM0Kg79RBEm7U9nePr+ACsyIcpiyGnYj66YlCO5XQqacLfh8oZXSZ5Sc6SWe6i
q0he6cvmb9411qYa0iWUkcMYtZsLjck0xkkfKPuNJ3VT0bJUBx5vNAN8isivfYqHAvEzPK7k7xrQ
Yjp1Vg5JEOSg4m2veJZ41QJymrtXdHN4VIjnwvAWpQFr4ocvqFPDwigBmg1+oDIYJd5Mad5soAhG
s4ZzuvnSqgUOjZhdmz6u6V+Io+DMav/uEEepuRpvyjAdnAXi7senvqGMI+04hrl17fA65BdjkF7+
dPadDTOKCy20BlErNEhka49u+1RVhmm5+s91qTTpgs65ngpSRNlxAXU10e8DTa9IAS1al1HzkbSU
TQ3ume4oODEBDwkJwwTAyM64G9o24wfBpWOSTbiNaR3iKHS20pHWZ4yyhc4sLTX0XqjGb4UE3rge
bY+ZrG+f2Rkoq9Mf+BsIJ0yucl4mnt5mlCXm8mO27NBpEUvm1Brdu2ytE7cT1JLUYN7TcObxzO9h
5QkkibxJoLb0y/HJJMDU5BCuKs7Oo2h1r2LScehNGdhS7loOHgxzr239A+PwPSnbpHAV55wznywk
FoukQCpC6M2e70IvZBhF/IYcLT9bLeBo/vNpJfUH8BisxiaPDaxRaMUTdC2M+1lIq4vZAbTulpFh
dxZEY4paULVYav/XZ34lUYCTkWZkzX1YJ9I2xA7B/6CdoFHDFDGXnmUIfC9pYC7O2J9FGZSawckC
IGe7oZoVmF4qMpIfmmvIjwdFORjUKt/RSNhXkSPp1s8KELn2fGsx+bwVi0d5rFJlz7KSSmhatwmw
NfPGaCW0kThs+BeW8X2iuDP0l6VT9w4XOCVgbb9IBKfYPtSDWHYsu2WXOJZiYedY8eNB4WtPhxIV
BAh1mQAkvJrXbHjoeLArQbW9OcVx8XtBp9PpkyGJouX6KE0QF3zGxupEusA7p5FiCSrN8hkrD/pS
Vos1JGA7KbUO1tRaieh/oWnqbWu1isxrblDZFNXr8gm88u2nxbCsq0h85GcVbC6tKiBH5Zo84YVh
BkBgD5C9NPXPqk/QpLkv8kLybgjoSXz3As+xhi/FjLeKkgg89KKriu1Bp/7UPfJXOFlJFz5X5peW
ksAr2Z/syNPPclXzPE8pl18U2tt2fxxSrAVdG/uXPcjaw3nJ26bK9gCJglBdyXdSFBp57qesXozc
/h1gREBZzgji1ev3l//i3+SzMCn5ALl/Un25H7cpQBM80BBCD6w6N+jn+onEC5aoS+7r3omW91W0
8Ws21lRItubnmBB8A5SXLyB4Yt9OdYy+QgXj02xQKTI8Smmtsk9MCtdjsdxeOJkQKBTNrZSeZ7Zl
R9bWK0MaOb5TgY2LC/YiI1RAUDOQW5jhaR4Ca7smRoKOLmCXiY04JgyR2gMnNXdJAU4eMfK6f1Ui
x1yuySydoo4tSfMCPbZiZ3xbBBxqMYt1O/tyT+Z4c58ruNmZ/fgXpdvl/KEB00BqwL9Pp454cgyd
O02jbDVfUIze9/I6vLf/8Y90djfK+UEhbfDOlZ1TquJJE7f/aefoVgdGKtfzju/757Bw3CLLudGv
ZHJYjw9YO6lRkRmf1doNA25m9bnls6k0CgDKVo8bbYdyA/6ACMNooQSKY1NZV9JmMH2G9xM/lnfL
KxMEGmKO7k8jhnvq8H1oNnuGpckdAB+uAR0guQRpgP9q8vZN4feRFHIX2pRq/pNM4aeXYYfCpPRo
40NbPwiDwZ4xGqNK7dKaM70eBe7CZ+fivYFe1HcwgjL627cFmM5IwFFzToWUAVqigrfrcW8Ow7AP
l8AoRxh2zuUXM9QjluBY+KMoZpAYZ6jfAsHoWazz/mqjIHIe4vA1bAAQduaX96spTpHLo8JfH50/
RpDxZKB1y7COp38f6C3dMreRW6BaeL/+YINA9rswONdZPZW/C/r+MNjzbjM6XXmthuYuDZbOLddo
EGHL2chLo69FEmCxHrVUWXwXAcaMwTE8igP5ssSLumrLZVyvm/ztvRsODj6nocHfAIJEr4yJHImL
0Nj8E0sgQfx+QGj5j2L6WnYM6QMeEsULuq33pCPQa7S5Qi7ucYQAvIaqkz/UOEwdYFnMEuPiefPR
N6lTuVVW+AbLxixMwXyIbD9lUt9eCAUcBx9YacYCHeL2yGspNYzifzCSlP284hxVAYVofNKtwF42
YdKKVf9nE2Gc1+src9AueU3RGLCi+mPgGnXqpgLGuSUerCijvxdMQVZWb3mFzgk5Ygz4BVkOsetg
eqaWT93JIskaCjy75qKsDYkYFJoMXPIX6roubi9kz1sy9aKcGJXRIAOn0eMKQpOnSwtoeyE3eOar
1EWyiCkVsWS5XOi0mz16vW2fRjIKQU5i1iCzeNr1U0XuRJy6EAGN8fwm1pkc5xiCNkJYtOn0JhrR
OYFV4TH9F4Kd4/HA1UPO+sJI2JFQMz/qfY+uljpZkMtqUundIb7td4gXxK/gGS6q33dc6DANkuTt
pu3xQovFGbpmkoN9hbMAVJWMlWh/r9LS78mMDcqt9V/j33Pk0M24qs8G7QS6p44zNqai0FrI97U1
tzzbgf84T2w1eOdiNcONuYTOEz3KGfc2VUZnXLPEzMClrJJ5UPRIr1mYp28Sth16nNVuvJN6BWl9
dRyEcg9MnVuMWka3ciD7vMAC1ZI1w7eMIbqADpEulGh4NsbxqgV7CKcdKdC23+pngn97QhJ2jzdv
qQX6U58hiZf1muKteKGcEgCaW/VdpbQqv6GxdrIKC0ppnyoovHy5++P6B9JA/F3HhuziTlx2QviS
wgHf5fwbGhi3zDMr9XfafZpqlxnSckpQ1M8xJH0+XYLnXnyibTZWlYQHVXxjVztinXWkUPFxQe2J
HPyGZ8eXKaQdQeG5L+vxdESkGebsuM9hM3Nv/0xo9E3NOm2UC2Wt50yC7R/yh0u9BeRF+E7ilFTN
RSsJTshidKlCoSWIPTOHjiUFxV8YaqJK9MfAWU7Bj5aBTyBR4NY4HhIBAKgYX8ekf4aBc9a01h6f
Q/+99nZWXMC4IqT76NpNJ/bjs6Y+H2FOS1PW+JGGq5c+0/vyPOmuD5tbpQfLJbz7M/WiI4vBqevE
SZN+ik8p096C3WQqjJgALh/mMpyY352/6QYOwXdQvfH6W8s+AkTtCkytaNjKfUTR9XZRwbKVTHIW
qrO9TzaZsD5QC1hK0ggvVV/S+x2MeOdyAwHiQDi3bf0XZCDVa4PLpZ6L2iFdntQcbljIWTD6iA6d
Sf9teDUtJpTrOfSfHGEOslKvfTOAYqBMw5/ZdOpGmPlJvkwjKKCfqwxdiozFrjkX/KL+WuWqbNKk
p5Gr8nGE60g7SGXVq84fR+uMMMFAv3VzPZfCwJMA20Oo/TrgAIg2mqLNxE20KW5p/LZuQ0PdwOZr
WBEsBuZLQVEg8K4xSVe7hCBmNIPOh6ewOZkEqNnn6522OSbObrJUFnwxZLg+dTVp3lIuO32dLlAf
9qN/OFYEAEsFKvC5zhDNZsf/eSMztxz/4IjgwqV7CExyXtX/SkbgIMoNTa4YaB8C6K9pIw19QIjY
Tqqi4xOkdsw1K7wmddD9DGMsaB04bB3+Xdn924X3zpLGG1ms1HqrC0F0JbaK9TCI2wf48a4VbWzm
IW90zaI2n4gXJxLXIPu46d5tlYWKEjNcRooFDJ5q6jDM1Ra1anvPpnquG+qBsp+ANTW7/jYw1VYm
CXaMiwk+IPopL+UFpWEg1RTlaQEjeTdRhbslMl7GlzDQsBy99HZIlDs3/oF6Dg419a2F5Qbk2lr8
xnqO9Grxc7qeoRb8UzWza9JTqBBIkBwip4kBU+KjrjbvGhvncKO/LWYhClu5Dm2UlwDTsLk65IGw
bRLJrmth9Mzs2czaUjzFlCxh2ux37ivgcVoWrktFX4Bdt+TbY3HxQk8pyZUaeOzTX6DqsoGas5zI
6+132yKeTTIRFSQrGKBMYRbzxsblrnZOmZZL9iDy5wCwRHAjJ2G7/klxN+GinIAhWNnQH5ovZwZo
28IZ7KStR/h1XhKjGXyyLCbUphTzaXz293I4nXsJ12dYnr9cZypfExslxIVYeRjhpgUW7+82VE/u
kGU4UbRufA2PcU/tjYU/hwX6G9vKBiF+Xym6wEveDh3GBnA2WI7xZqbthDbslv1yX/8sioznnce4
WhJbHw9nQKlABbZ6qJLv4v3PiGVhnI6si8xiE/w4jDCnGdTSYAiuSxrXbq3zHnZsRXu1cwkzObVM
glul5JjjwoCq4mX3WkrqQdJiMP4lJIuBPXaf5ylNLXwegVj5zJ9wskBHFPumeTHbsqruGlWO0K2R
jRWu9fTIFDmdoumijRml1drVdtv0BPmPyVmnKIoWklrX/cAV4SzWFGOWsIIdH5Z+ccwY5eSMmLyg
psetks0TKJiWg+k4TfpK9xdAxcC2iZTS9IdLfxG1v4o2LJP80g33vPSQ0WJNmRmzcet+heHcv5C/
5XZP1lufP6g1zsu81OUwA0s0/17M/2+quMgspmvxjDEKsz4iUCg+0FmmMxzL8H3w7MSI6to08ZqI
54MZ0yEknsKwbz1BexkLCQZSmch/WMh/fkzouJem7g/n+WHGFrax+UZ/81SM8T3Eo28Y0VLkdybR
DLG/ljNZrIiIVnbo0z7PaCSBXc2171iBwPT/0cnB5PLhcFaRiA2G8A6T250L20Xh19bGn4vOdzrB
ds7LiizibJ/NfTSveO+OBymLwyQESaphitjoBeZxaqL0xFs5vcZ5fkuUjQT/S0ifcrn53BpVXFFp
BJCk0mTb/LFc6vHSij3s+OdfXBVI2YBXGvKQwPlHrf3rfgMdVfE7edquPsbEF6PvWfvTxiKqX0qR
9cGdGZsgg+oI2bZLvILQt3uBUi0NlW3CXkFoZ3WKi1NLSDjxo43z/BTODSKPtPRnrCVyxuG/2h2z
mrwfmAaEb31iEmXIozrlWUC5h7UAXhwS8MkpSbSp4t7oHM++tpsW3LQgkugR7M0/qmiujJ87jF1X
/tGY625sw9pCHt4NkUlexhL11cbZKHzYy+dXrZwuc0kVxe+TP87Nf+hFH/sCk53yMRH7fHtWcVZP
L6qNR7iJEHgsv3JPnDiL8btkAuPZ7pokybSXUYSwpBsHvjzWx1rNNmaErWyvSWzCynOTo+IJ2mDY
ow0/+4TGO8x4Hgrplt4GpPDtuHpnb6qfWgK6lPco4kxe7aWImsF+rwqFKZtkFc+GkTKv0nUi1pc3
Mi1XwIGxuhCGKuzgGbBFxoCAQvijS9OqcU13XPHxtphj1UyfV/9d0sez1HiA/miH/1d1zQLH55iP
11GuSGkEwlIHXxH2VytFjL3CmO5sl8IzVBdxGUUjXdp3tBzbMU5waUThQEeCCdLoSdbRHzHeRvP0
UYYN09yt9N4kzXEYz28L7O/IYk1VFlNqBU1+3AydTPmRrM+RsVDoqOp4ttnjfcmOLTnAdl1cU4ZT
2HJaZCX3uZDzvD7E3gbC7bp43JdTgOMlB2SofGvoNKb90b1w61+cVsyFn+xZDMIfrUcLKLzCG7eP
L6juebGIdnQXXOKfqyIOitTOCH3eti5y/h2RTlANfPmpH7dLIc3thY8sOad04jL7HVshSM/g+cPY
5ZFn4o+drfVKlkHiurF5zcM01r5Zvt6gt6K9b3Bcm7MauWht0UGnrHvIEvzcoDzdpPzDdUc9glXc
MQdmwhiMF1aePeNiv+e1mFT4hwq/d+kzA1QeOce5MIU74Jkj+5HdGxYucR1hZwXz7vDPrWjj2p7Z
FUYHUsQyBXpbNFZBQ2kDarZfq8gSUyQBJqOvQUVtrKNGnBV1SnguehD26XuN/NGJ+9YWoktlNfmW
Ou/nznMZKArSzoHok2fhEHlMS0a16aE3EPMSYsa5yA12jOzWKhaHL/v4DvAW5jFAm9wmIiPM7aiE
RKrnl1ct+rBnZcB3w0ETkxbQQLNSdEjppslBh40UgR758+TugBVEKmjG89DsEk1OruLLazrqudWt
3nCQGGwLI/PmfjmZrAVF/SZRrOEG3E++UpYNH6XFvYS69EZ7Y0Ft3vfBcE3r1ev9TxEe9/HqTeZy
xk6zXpfEHLswbXWmMyiALOGffWo98WTtnOA+AuHukgqkWQxaoi5BHZJ8BWLwT7QminG07atOhhyK
GE3frwYYC506lvoPkP8OSHqCLQ4h+uqoGwWQHE1mrqzgeK1wOKi8tR8wlu1qa1TXtpGsBuF5Mkev
jeirOh6Rdaaxlpc9h14wViZvyDLb88qncnNeO4MsALWgFz2MYdkud/DC2ysCpee4QmUwCiYE6FZn
Hj8+Fy3Hhb1jdD2HQsAumkHqlPxyYtOM/h9hJlaK1TOHBDMxG2N7CcxNj9d1m9Qy9TzjkWTtJ94E
nMOBM41WPQ/43ir2n6B4quZawvSWaAhf1Vf4Ih+ZebCKy2+44zeUUVgkXy7CedJndVWhTSlTJDbQ
WJFbxsQz0QWgbsJkOpsBqJ/YQcNMMPfZdr/v/5PaNmtMULrbQWdapEi+unIPExVIbL7ugqHU+Dvp
KVVMMaeXMq4hpyHnuXgmP9UgTe8hxOzkt4PtTMg2cBAF8ZGh19TnpiWEHvsdlUutUCFedv0r9vbS
MAKrVZpeVGXC2+gBfmJZz8AMJgwNBD7zNgahvqCcOCYSpMbh1giPJa/cYPLfhwWw8H3vR1z1xsf5
6zT/O9ZI2UPSo7yVloFNHT9TmkZxwdvF+XcpKBP6nbdvsvE9RfS6CBNQmQJ7Fj3505Tv+6s5F0mR
0tvo/S3DLOjNiwajJfxkL9pdgSz0bPvGbjuZRvEQN8aUysC+6pGgDXIjP0+KRk+T1Wh9hscDEdVg
KQJS/w0gKY6YTpmfCl3etDuyp8aWhkx3QxVCaI/UXHD+8L0ZxNMk9/VtZKAs2tjQpKD6yNh3VBM5
eC6HrL+3rqwlSjlwHTpBQASpE+Xq0bIPv6TNlRgjPrm6uHbXqq81hRxtm82madZxwsU9ZuER5kvk
Jr/WTsSE9OA6I1eNSLe9xw/KRJaSZrjhbnosbt/Vc2Nnce9LEtCBIf/VgXgVa6Cn83TDEYltBA55
NfW+TG/hzGA5EJBuerYTMJAUN4XPmxhrc81zt1iynO3Zj2BiHFffHe2TeTXAwqJ41sxkk71GHMVq
XfMJezI4QgVb/y8lsTxZPDgJGaJnaRRWo7NwRUOVxHQc1kXAmCXgtcn2MycZU/FC0xZDDHjIB8gj
RMDlrnQUCxdWA+xIUBz6wp5CCjEiFDtcL+6d1j/Q6Q24BhF9JIk4PgKSmT/jzrX+P/ILM85Xt1BA
vDCbUOK1DgXk8IdSlP8l+mG0H83uJHyUbD9MR6m9JRMeVEQL8f/hZbLu4/by03lIuWt9AtO07rvn
KDZ/G+XYe2dcwbRe/4dpffZ3lUeWVq/bPn6c1KPaC0s2QAdYpBNwV+WaTZR1MlroPkO0VgNdAxJG
J+QGlNDQNpMPN2xNV87vxAzVT6lcxR65muvepy5UP57ghHB3bkrYNHmd4WQ4e6+she0paRGNocW2
Doq0oX4JQg4tLKtz4uYxWLaKDG4ySm3NlqJkB1Oj/k4ePB9fqD4xZnRPESgJMc9T7CRlcTedekW5
Ue3lkweNYI4kExa9PY8dJ4bMJgAHGoqUUtgmr2kR35Nokt7zmK/yKFHvbAiW9jSeA42PUH1YzX6Y
j+5RBo23HQc5Uh4TY72MQDTvjeBG+0jMsC3L87S5VLWjiLSQ0T2xQ8etSn456gaHrkCfGxeNAZuy
aTKOnE79Q/jqo8HW7w3KF9sPLjP37HOy/qROdMhGpvgpIEl3WTGj6tgTDEEYmviQE9da4G9jppL0
9WfHR3AdVnfETWujtxbCHzugimFOKXgW5Kbsj+Q8fWiGf4OgF6aWgw1WZtuYU+hCtJCu+a4HOMun
uQfyq4JJv2+DWGupq59m9lcv3cg6/ys4upBGBnUeDBO4Qyuni3Q4ReBtsO1oXgsNrU5FpkB409KN
2uhE9P1rkYOjD8pf/XP2E4rDkkQvsVXclixyyebkml3hp0yJY0HdbivUXZYYiEaUSgfhnXl367xs
suhlsVXPHfDtRoNeiWpCZqx3ud8znCg7PIynV1u5wvFlk3NXthFtRCzoyktADJOePt7cDjciY2aP
5t6W57WWFNkCqFJj3CEeiViOAwaGdPRdAF+HF1tYY2lZ8s/YPm7LmTTLfyyZ/n9Q8st7t7iyMKGH
ohG2xH9cVf05RBThvyxaxhGAlSbvZw24GEGTtKp1aE46MdFTkYDNw2sPEoj3BSEQ0C92BDwBa5OX
4im0p82jnxB9GedhkRKW4XOxF4A19fZzc5nak+l/2Bsmmg6damfSVZnyY0aAc2iyNtHL3TmVdsEl
N63mgHo8Z9g0Ydizgj1EPibutfxmsnjl9lgLCOA8g40OQDzOj344+G6sd40uQkYClaQwD3ZSgc75
d/n1zwcS0vwM3c4BQ2y/8y87ZQM3+D3PYU5Kn3r8n38lZXFCILJRg4pqNdmb258cvuGoKhoMesZ0
TwMKWyMUTRk9qzrLn6YWkrwy7CYs1psyTqf0PXEBxVIDnU+UCEbFHTRZARgy2R7vnGUZho5PPAGu
z/1l+Z77JxPHDJHnjdEP1TXekK8ouaFeJB4JayDyvtOBUM1MqoKAi/rbDuHGigLQ4veua0INvUnm
qq7FPNPrYJ/bGa5Y2rmdwpsBrt3HmQczKxlOqL4X+jzyp31Y9ZVpoP2XfHw79hUXhAQkJmQ1wv8Z
0l2/3GgJpTLgClMl1liPgiwpNlSG0Y6zIWqNxCeTM+vj3NuIYR7WjzyoLtOJieWC3acALAKmXqK4
cxUxDdBT16AxzsRpP6IdXIEndN9t/8z9vpVbx45BPtEjH6tCd1Puv3/P41QUgubehPxdZOIeZEB1
GlnB6t/1T5vRa9ZTAU7gEJqyuvfxU5lxESpR2dAyZ8KEllHG0qx7GcN2x2fR1pL4WeoF0PQIJxla
aAOYdxKr3b/zCDcwzNNlki+Q8ZaYy/4TKQ77w4FCsnmJMhPXsuC78VCnF61EmJBEf+GxhrcX5amW
vSh7SNTaD5eEkUTKEbENCmi5bxcQ7pcSNWeJVTX1jqHzKkL6Cro/NiohjH8ehV7MmRMaH/q2yT+m
zbp9Tm0CAxdq54Ze2LqwfsVAVYj6oGlEUx/e1cUPo2XwpG9zI60HkjCiFkMsjXxPh/9VxneA9vlG
8i67D8cHrnrLVhNzQW8QOXGA0gZbXmdLetWqshxN3No/s3b3xeZcsNY4/Z49Yt3z4N9pKIDtbX+r
Eyys/Hp5v/Hwd47o0qvhJ5pEPOu6v3UcMBDLt9Xhf/ChgXp65ssOFn/9dLYnXe6u6m/WITmvJsL0
cLuqg2PDCb51hP3uok5skgvyB4+n7A0nCz2Jxwt9BcOIeWaeyzAYB6vg78zF/Kn3xAFR2/oOYJuM
ZVdVm0dtdVoNO3wi/MnmU/MvP99Q0BIF7dJZJxYIqu49BzzgX1YvQMNGQ2gqT+eaj0vXBtkR1yc+
X5N+CyG02PZeAJ2AE+TaBsBsd3EYyc9yQNmSClzjcui+RhM1BJOTMUfucGfz5wOLDe4bIAGUu2Pm
FqR0YnQzSBNqT1p1Og0RFKaB/xV+PfXGWyHP0xnlQ78/o23BThy2WHQdVhgGbONrqXa9NA/pmfGE
WvDD+zKvicxjTUt4mPyoyiJrJ1zKJBdZoejAPWKqfHBuNmK8XHGIjlyio3gp/NN6VnJnl8MOrxrN
KlzneQHQ5fikgDKlgzXrP2deS5mH97if0S3ajvUb2SbUynqiNa6IyaYvGOfxuYE0jUOk0pNesgTk
unRWoPJ6jLQ3cu48AnQhR/8WLNGu4ZzDWnarL1zTNRw8W9CzFCCLwOhnT0XoFivKmIuDoJo8aBq6
DCjyyKUB30WmXX37OddkAv72BcNoZ6c8J4DFl0Pdljm4ZA3dp1UPTD0tSLmlsqJAfb1WbNYpkrKk
lqnYwVCwgZLLOSSn+B37b9pPd5H/ok5vjljmf6ED4WutpivuT4AAivL4KJjlLLRBz+h8htQSkrMA
3cIAdTRX+ndhmj5hi2c2XcUxDkVuidu8c3HOXGdkSf+kN/j9Koc+SDGnqdxAaNchmNDRc8TVvbsw
+httWwGCAhW1bcjJ3i+IJPkAilfNoqCPT69OU8AvXK8iGXKUzAnQzbDLLMDkbdYlwhdxIYglnur3
j0+JTw5D81DJ5n0/vOLtZK0V/23VUepFbDsnDRevb4mJStrb8m3y6Rf6bnARPztvA+1YM41KZHkj
EBMB4Qt8vQ/V9sodhRn7HSqnW9v1/fnTmykrTWi68RFKrkqyS2TLI0QanOeMM8cvW42TBtPEHV3f
QBhiV5EuL6JQxlS44h2TxS7QzLNIzM1uas2j5L+7J5gLdst4Qf/UBe+j35/MZrBuprD+IpjZzAhS
OYwYMt5FTEPHhekeoj4B2sdTvCS9vdZJEhDpvI97SxV1R7NCWl8CD1gF434yPMD3CDsybfgZdwjo
30jspg/ec5rFPl9VGkuahsROid0KZIVfjU13WUsQZHWrt7kknfHp2SlNE5VhwMedFjbLgKf2Lx3G
s+DqatKpsHZwLzb3jxei6Dd4LCXntTjjwAkUUOtLBpXTZDBliwK6zXjkOPaWgHgX9BiSZyyDR5Vo
uWX0pPwA02wuQf+yCl0yzveSVVnVB47i4Y6+2/jNDX0JPD8UY/VVHQyuFGCpDANpvoqgBdZF+D6y
yyBBlCDwJV/6W2GqpQJXmtH2vc5TBW7rBc5lxOCHMmXL3pbbcFu9Brx+4pfTCN/3A6Fb7n4dvFj7
C5iV8n7Yrrz2gXJx6x06CJUYsfJKwZLC56mkuHlwBC1JB/T9+U++HjjyR8t5qQrlCwEZJvrMorBD
EYaTqBgy0FwgNVXP7JGxi+QB5I4yC8L2vFW7mtFb7xV3oZzS0/+82hEA/R8w+8bFi5JsOQqciZLs
fiVeYcSq2ZWjhTeO1SVJoyC0WgM+89F+PkmQXfzZq3xWvlcDgsA0F4q+r19qmXkZ10u5A8i8pUr8
XHLIPuQ72CHkvXm/NGpCHJB63Cp5TBYTljPwsPytOQYgVMk6WRrCDH2XfX+6eCFUa18cjltobV3d
DgdKFXZVLRHVBqnH1jwkxhV/3RhxJxSv8jCywhGRtlxXHj1jkZv4i4PxXAVnc8EVfxSGItFbcWdP
3kHRd2wb1ZzRmBdh1VNIgH27NwJFJ2W+HeSgy3yi3KBAYIjbQnCnb+PGlOWf+ryEnijhkEp4Oef5
Zn+prnjGRrQJjseX1312Pum15ZeBJPvzeK7gRUuPEeGaMPHFBigFyr8bMF0shHZ3S18qTkg3IPxZ
hNeXf9NYYFm5f/AwlqQta3g5MEdvxeG808EHZQDTiXlQ7LlnUpNX4V9Sv3x/exc24I7siyxtVpTG
5Sq0/sVdlRnUQC2KVyC4uHvjBkg3KKkxvUZ5kozMVqctf3KBR64BBm5mEKZtVaOJTi+umLHHqmQr
LSlIwce7/QWp2u9DKZ2FDA+8zMnGsZeK3opX5zWbzx2RMqEGVHRz/jQsc1Xt+LCVj/1KPQsBKKVM
2CITrGdN3MYvMXJqErc3Kz8Y+mC0P4aZfuEgNIVOxooOqQo7iIc99GsUOR7sPUYHiLF4eEBc3gcD
LVXXH235Sj9IXI+BEjzI70lcSDQ+4HLs6UzFFa+kHU4GBH7YNVTui+3/UzJr9COUbzbebHP7SnY1
Detdux6JDo/CkuXz7iDctKvkqmdV2lsMzMRirA61PK39R6A8zaBBzjmEvBlgH0yVBOrL1c8rMovE
NMeOEUfRErc6j2wtr8JNwIIuDQvzTsmSrtU1tEK977YiFaGmL5K7bzrTHw/HDmpp0SyCaQ0RlSqd
keP5fPEqn262tsd5fKpgyO6n2pZtmR3d75giYVbt4rqCZIi+8mm5ZlHiv83j6DRf3Cm03Lj5bWje
wbe9aIUDwy+43gya70spgzDpQ5GiPbHb/NmYqnm/lUFDluX2R+52Mg9VeVo5SIss9CLnnoRDEKo/
h2nlVYEV3qbzfPdoljCb3A0+W0NwHsZA5dT1VYu7SAqgigbHnv/fMq3y7KUOwCYpsHZsuQueKJLO
gkYmPdLLr49K0+mXxKR/4k1SwLIlO8GLnyZGbwA8xUm4d9lNmCWxnwNxUy3lVu3WBhMqyrUZy/fr
og9mk8qmj/PD+7qQX6uo+2g5ryQUye1ik3E0KfsMi2vJuE2pVL/JYezWSga93nJZmiQ1BsFhc8W/
iTNr/OAzDYUs5OiKyK5uC20WJgQJLLxyTAV3acSOjQXcJ1AEqu0nGwhrbw9nJAveeqEnVVDa1fCR
amqR3TnzhESHXLXUqmLkLlysJ4it58ZpiZpDhjWkCI3G9FHKng02M7zUHKLCnLVDbU7RG0S2aqIW
WEmzrCnNSpXA7rQbHc/7MNuNlCJetKqeVDG9856Et9+vupvVkP+WwUyGMLFk+Ck/IQBr5jgF0tuX
xh7cCyqcMEHwiz5ju5BX+iUndVGTtIwLPNqfz0vWuW+oY5gXFaC71GdV4dc4oP832N6kumPSwFjP
d/nibL58fjx/HxqVTVdAztqs3/nCRoIhUgItmLjr5IWFol78Bgh+tFf579SuLsb3oqkOXhjwBdU7
XoM1NEbLQKFThzb3qREFoA1OvNTd4lqNtZEzTAGsZkaEuP3bBCeY7FS+TDXDi+5kCVoE20+DC54S
TO9rF8vLk389MPb1cpWO8Kjs4F0GWRn+wtruMqBZx5wLuOESBhRqwjHI6FVuKXVyyLjevpoDCjya
O20XjKwKpDKcB0p1K8K9yW2OSkMFXAldIcsXBrRll797BWkvPE3mTLghQlQBzOv4qvQ1UzOlWddT
2v8XXho+ly01QjTXJn6jsyFJoP6yV5yL8vvvU6TuzPc/vKBU0fvazeg8ePBs47ttm6VshctegeTS
fUiWxODoS7beSz/LRw7AflPXWw3uQja2L9sOqkEVD9K59a7leeTEj3cDiJFSgNdBQnDm0l8na+zW
3Me9aSYq3W0BULbTM1m7L2eLt+agWEdnD6Y8ivLm3zM4lNDbJr1PnqLU+34W5d0AnYfJEwOCXwl3
GoXWyZ+3YkvBBQqkF8GBqmdzXYOcHJyRSRc2qJrjYdEFhD33YkXoVMi2fMfP1yQdWGrcxirxZYjZ
N1gfFnCXRnUBSiCCQjbocZwHKScy6uIp+ncBEaXUHHPTi+yQmUOFWjjaWB8x7zjElxtDPyA1ohZo
GLEwEtfFL1J55w5SlOejtVZwxwjbg3/1yyqZpiqACRh+2bISCDJ89KnD4UKzkhGeNPaoufAOdQae
oPFYgjWozuGPzbEYmXyvXC5qB1qLmRWcBrr86s2hLwo0UP+IU1JZqwasMbNM2rJ/J3t50gCY5snn
OjRsJIvPuR4mVSTwzNuiStSTnBl+71mivrsUsW7lsRf77GMIvUgm19lsTrtivE8puwBIY6AJpIwK
QH4XPh2/FgdhLiWqRz1B+eoV43204GMJasT1jF3AhTStP45xagozoGbWKyoixVyquxHciyR0Co2Y
lI8HLNl2whxteTaDIU+zRHn2q3pBD8Ll1Zb6nfBf6FhaWRX24iHLBqTH33rdr1ppjxTa4OfcUatr
W6B95MYjG4FUocof0xeDlVKSmk6Ktul+tq4R7GOP8NtKP6SLTq2hbXBc2JyWcMEC+sYHmA/ncIXp
ZDj86kmS1ZknaF+mkidBh2bZQKu6qKRodVnh7m90DJCe/3/CNq/Wcr1BENr3/cx8GGBdtNYf4Rl0
H4LVl8P9J202PGxqKFrz+n+K8uNGE7yEqWxmdzx8nKwAUw/7UsjbSUMjIxYCFFODiDamVHDc4jyv
qxa499CEDycuqsvOHgM7kofbsrdhf05RCBIS1V05uQ94gT0QILs7nJAJmBKPZB5x5POdBEDUksCi
fiokkGhmPGBNZyENpZfV+NtHkwo0rYU/kCg6aeL/scf4vcoMOmHQLqItmSv5QXVh98zhgoD71L3Q
Sm8AdaGdyX33g/WsPdfkGxIRlxbWpJTzWZXQGxKapUbXmrqbHqVPiU8Af6wcGmptMNRoi9u5Wk9W
nnPb2SF+a72qTYsGqPeiBBq1SnNZ5uIunVbnSGwP8g96ou/Ynrvb+fTxGw59XeAZfdECrzhkaD8t
vTnvRYjILfXcUmD/WN6U80p9x5uET+w2kGjskf5WBRmF3b892PbeHyfA4q1Zwb9k3vhJJqimID2u
kp0BpU9lj/9NW5iZN0prDBS2Ttshwr+BFgam5TNsX1k2PGEDnQrUt+MN1Nzy7BLLXheF90N6aR/h
/PilEvuFPSY5kr9h2OZm1sTG1+Od7Ik5lAEWaa9HCpboUVP038jYjDmVFpxfGxuNKK9x5qBighuz
pPT6irzEzQ++yDnC4Teb+4ihaWlXvMmZC7daLt+jereuAQidnHEj5HK8IA+5xlD79Pek7MYTHNIj
RlY19ZEuFcrPWJ72UAiXkzGdzMwj401g/TS4moeThPK8CWJmphz7n0lR4guWeb4jHEo5TDm1yeUQ
QdX4jNKjZ/bJQPra4FRGPOZNPEIZlDv3doDWZjB62W4lrN42RaUuIQr9LOe3YwBVWU8oDDJ3cWQD
WOgQHTP049g2HG75Oz3ZBav0E+FJi82toiNeSX/+HbRS1PvT9/QsvpvbAe9tRdpg1+h4tJgIrwcL
X8BTmMvttetWXr0LuCdoOHnf0SPfdrmgN0ixUsC/Zdup72u5CxsGdzK8r9OyP5SElzSqRM5D5jVW
oqGtV4Xu0suPIAB33kpM6AC+kYXM30WqDh2Gt9izQ1eIHsCTo7gCUkl+FOeyhGLWanEl/jms0nAW
B1sEpNataNnOEkDGS66DTdnSO5Ly4vF+CLdUFlat2jnp8iCU3apiJXQn4CSXsJkZKCYoRU3imC7B
5WGBfG89y61jYWnRB1kZwZjvTvwjIZQ/3tixNpURfU7Rlvh2Reytq82HHLsKfEw/mg4ukAAtUvgh
CBbT50ZRqtYiWUFFJYPxROtJ6CxpYiqarTzFzvScLEwL6cp2QxJBq6spDnft4egCTM5NqSrJPQa+
GXQjjKB0YLVNIlhs26QARWqjoVy6n4+VrmWCcYpfbgS0DhTIaGfxFMgFoRuW1UakKQzcO7HwXWFm
6yyVSwb9oKtQuYMQFavuotJ8zEt25tQ3iSd59NG/QQx/xcccTmnOX+NVIluRn6RJaiaLqLsK3xMh
jQtdke3xe4vGnNRb5Oj71NLtaqN/43d9zs7SBX5vYWT55ehJKedYee2eYqabQdl12sangdbvYbRH
EhZM0S6p8TB9af1An+ATPPWO08bNx2W5RRg7N8pCo6d9EW9x/qW46nB5JE/oNyn0g9H3A1ZBy8Dc
38nvVx3LPklA5BsCmPiemZ5nUhNHfZZ2BoexgL7o6MMrVcq6cLeHi3AelfZYTHlLEZjfzOpMEfRV
IN5md9YfPxmnuwkBYU8Fp2y34bN45ETs/RrL8T2D6xffWArUp2c5lE0OboDfWr8vW4XMSBSoHx9r
/ESnAUITjAW5/f0oeM0CWs36v/O60Z/XCIWvYrSvr4XfXxQrxfa5aO2/nFgQ9qSfMP7MGGqn+JQW
mtsAQK0bgdb2aaAbs6HylyvhDhxJWL26z9+/nkDJUdfbGwpREBaEANDd+UAmcr6qUXYB8I4yABzb
bsJVGrgs522LUAo+bs1TLkPvDL/F+W+rnTySSSZDUzptDi2mxjCo1hoO3fLEknl11B03dCPWe8o1
UIlTZtofp8b4gEFAoR3wuf/3jhAvRHKtUlWNjyo8hvy0L7YX+S2Bn0QV8OnmoHq0q9vK37ZTAN8d
uqZXOZVOFCfkb9npXQclOG9tUVAjRW8BUeqDUVr7r1t3ygLr8+6DpqfQFMGuEHevF0A4KzB/J7WF
PQ0ukIQJhwgDxacGCnFrq0G3VZLuauTpUwEgWwran3rKIzSP4UiuOSuHkkt8gPWffdRmiw3rMMdL
mFPZtrIrrdqlaQ2FEVOuDI/l1KN3n1sHh4kBUqakAtLUqNlwQWMZgP+CvjfCfQXSWVaZ4XUaBuBt
5N0of7Cp8WYmD9+gnmyDVyb1m1bUoHColOVAophwLAVd1/mHO7gWXdRhzOdMG+/j5QnSb2bBsioz
FJsrlZxKJsNm0pKLG2fIRvib8NAEITXvhwWhVSf5VzEwkcI1wPXIZ+zpcVv+8bfW/lXAg1MDUzzD
ntjddcd7aKysfZ340U6GuBwmqastCj7zoLsWOmBTq1PzzBk3zWM8lWzZ12JYXI7l5L8lizuKI3SA
vGhSGRX//Lby/qbnEUFeeHXSTXJIjP12eqreVxz0lJ+shYO8Vl9tsneVdoBJYtqLJJJDALPzpc8N
B3OnY3yNYT6OIPLBcUwLZZ2eFoqK7KFaBkf+QstqzH9NAXAbUjyrzX/nMrkHpAeA7TytaG6qceEf
6KrrpoMDyrfbljl/ou0ID5L9/dk3WfWomI42bn5S8TeaHPO4D3Fh02hiIq9D401w4y8bksQb11/T
IpICruNv48tyU4/eBXoZMD/2kIp2yQQhBF37lroYh1dzCpehMEzxRxT4Zz+3h0mUcOz8fhyo7CxH
OLZRFb0gqRgHnEoM5Zwa06KHQP719m/aHXmglbOuDhY433J1iyLGtRjf5f7ufV9lfsMpbujpkTMQ
wsuUYrL/hLk31msF3q3IqRvkowJtH6KSJXhQcLeNEti+7BPjYIznvCHSw78wuPm/EFpBCRUnpb/+
4E8b5v5nWuSYDDHKe6GjwrFgoG/Ru8iYQys/QyQ7AhK1IBlWNSX8qAIQGlHuBc0lWWlB+WowA4aP
jKg8ZxhyPwSLjqcruefpiCM1xQMb2xc8tLVNZg6926VUs4YeXDNzjZ6Xpz7G9DOhUpyJoJ26loB8
Mm708Kuh2zCnd6RojIr3mnV1XvzYUiAbIt3JQhz7vMd+Wm9BpAUhB2EQQbD6yCFg1eYneim6Z8qN
rdw/fGHStTCDc826+wNt/dLN6UDG/oowMKSIIWW80gjMPTBChjakE5BRr4Jec3w5hljs1cyWkn4F
Vq/NDhdDLJ8mYJztYt4g/BTNpXwpK8BO1BnfgiztXFaRn0oqlWU31oTEcxJTuc9T1MfcOTHDLnQR
kVZDAS9uJuQ4PQlUm7oYtZ9dxiDm3M4cgSHQuOBlESrjearGuQNpydVf0PSindEmcUw0VW2h+4Mv
V4f2lT9TJPqUhZaswxYkkrp9bEK05TIkc154wllJhX2wvmsE+1PNgXdrx6znOI5YcRGPoirOUHZk
//374HrbQMFZoKWBJxEoUh8SyQOXhMVXbOBYLEN0gMlqHMAUbhBF7D7j1OM0ujx6mQSDBAVvBMfd
d/Clbb2pefBwnTobP4ZnB7ni2txzgibmmPririBc9ulyrmbyZs7d4Kq6MdqTZLcAsdq5/OTAYzMV
i9evTphV6WHu9YgtpAjk/Wxt4tVX/xkU81FyNZ4fsjI03KwX6GYA4gJKkww/reKgbBkc5OeGXlv9
8r8AcLjDyqosNchQ/HY4CpMbX8t2svt9MOT77JnPPWnet16Cphqbu1P5UW/4Xoy//lgkW5ZxrhE/
NqNRpxSTsyOoLssjHDCkiTcS1Jxl6+tp4OzuUDm1u0bJnLDz/Htbx5BKRiUIEAElwD0cHodcgZam
wUr4MPMUfSjdXpLbuTUu6o29EaAGX1JpvvTfFwx71d08WUCVjxRXQCvUYl3X+0KX3KGJ1buYqOoL
2cIRNC18C1yOlYkbGci3cdUwTSpU1vvyMAUlcKr6Or21M4gklG9BCihLWPGGlqGlcrC6T6ADCbD4
EsCoSJ0XcK6cQt32oUliSzvLtV52QcGh+VN66ZuPInYrW97v3F6sdFtgaMtpbA+ewaNga0uUtF+Z
IBm8BQtrTJHq+BEvJQIn9d2uKb0pTJZCuTyfZB5Y3P1wZBt8zGIFAc7sjpLMXiFWC3L4ZnWXdhin
FFrKBOX5EM8NMvs0u57dO0hhoChIqWFfSymEA+hek8KgLAmv7hVcCMBV9mpslyo1mDLSqc8KkJtU
uCKBJbnv9VvvVY9Ts4fEwfKoGk8T4lCK/fYZnOxJ1NA4E1UZqU75yhYVZUHqKtfc5TT7kXF71u1Z
uk5Y4G24ygcKFW1HYfk7BdkCONXsD+ZbGltckdCqfUYXR+pPkzItaYl71U0IlukUamgKDATiiKr6
pwrvvlR+gGYZHonnqc/yOmYXiGaks6Ry/fCcaWZET4iAghRAz1Gg8y0iCKPWlQ5HPG7HuAQyYnXR
I2r2MTtFT3ENOLLy/0EbFsCZq53A5Bc1cwEULplJ7BQKJK3E7Fv1Ej8Iv2ZuF13rXrKbD+jTIbb0
ZO/rcfQqTiAZ2MTd4RP5zhUmmdiogqWY/2D9HYyzcRZNh4Uw0oN+1WIWZx07j7QfvmJWLRCkdVEj
0LGiAfxCb4p9oHX4VwoGW3ungc2L4yd9YC9/Dokl+FVxIjG1W5pumqCgd7A7SzUOdvwHRhM9w44V
gr7rKP04EkNWPIiok6uzjDTLZ5qx2IAExDgz7jRnRMr8MlM3HoFHIXtcRW956HKp4wDm6i38ENyI
OnmagSxhmJGEzifolYJmdBa2xGd8tY5VT1ikgfD8ZRh47xOTzztljOyj16X3Q5Nbn0B4NZrXu2aI
5YnMBXPKHaTBP5tdvo1JL0nS1nF5WS5dHrmrRkLEd3kJ5TYeF9nBeZef5kD2neawqP9eRXkJhccS
tIJVBO/6VusuNc1r1gWzUN9DRH2jS9cjvd8AoE3PM6qXEVgyd0TifodrJ0/ULE15W8SA+5sD8U5n
WyBcCfiRtBKWqoEgRA0xl1HN0em8vSiXCZ6p6bdxNOu76O2P9bM64bVEY1W3iAoaQ5xjbrDqmgUa
mdDZMTkTBFHsO6lIScIljlK2SclvT9vhvR9EUk9T5wm/wykOCNX9ZN8bP1nWCf0r821aaMNhHXn/
kDMJPvgTRABnWsZl5sgrKq2fFp8KlOARsqG2DzGcPekCsBC39V7VsLl34BgwbGjosdVQsEO7QMyI
kHafqDMg8LvLDsgcvW3BFLSr16EpmJpqTg8Os0EiiQcD2uXo3eEWVIeH0K1Fp5Yey/M/L3nN3XEs
xNYVlBzB/ppwRstfrdUlx0iZc0uckUInwGVTT4kCLEXz2T4yOq/qCv6kZe1y3ja68D+MYfYkxBir
sW7nOW7kN8pLjC2/y7/F8rvqmXNpXLLsGQ4jLbQHRqAKizJvmDCTL+UDYLw360K7S0y62IQTai2U
DlTL/xeHgdC2WAk14bL4EXKA0FZ3RUueIBhPJGJ2Mi4A0ffq3lRAUOylEXSSxKTZ15TdI32APuKB
0E5HQ9nAQqYUPPgAy2czFlwG42hGAKzggv4FsyyU/H6iQ+I0uG4wREc6qP+XtwMtzfmTN3N9O+Jc
kVKwGQRAWFky3z6i8Q+QRIvwAyqH91rnbApdPBKjCCZk+KXouG8e08l0ehv0L/0m8v8ivojsx4d6
m/5uWUwIBSdjdz4JQOPfTG6t7jRGhjsSnSJd4PeBTqe/z6BVYvgYvOzA+kKRX5vIQuJTby8l3D5+
vTY5pjO2LncYgw0ywVAW9YZWZVTfi5/NUsJhuTfaFPHLjajMvOgJrx8iWp1Fwhmdab3+dHKxJtiS
LqIQKnsXlPaJF+jD62cEaWS6fJsn9jsrMgEoeQTAJjx3tbUMXr8rsqxaHW9mXmaxY62KMragWaJG
Crb2agnXl4kHYMUJ/jlwum+uXw4E7IBCMy3PFJ5szeTgM1IwWcGNYicfBsCpF9l4irrv5gvCRY/W
clEESXwp0XviTUNUjDMtKWoFiAHwUoukviRWxm6X59T0AGXcZsF5X/dlY8ExhKM+MBAMsKpscgnV
de4gisM/o0OLVJVr1wTH+Al+pfVB4k5pSB2HE45C5Qq4sA3ToltzeM1GXxg2yaqKEWdodrXoFd9z
sWJStakACK+93YQabD6ywuV3RlDdU1bdpzblpD6uWDlSE4RNWwkGlnwTUoWUPYXU3TgUEwzriuF+
IM6i2VkW8fNhmjZckGo6sQiOqUtlfmumhww9G8v7/ogRvsi++sNbZlrlB6UghobkWxTy82GNAaP9
WAeN5NK+lcTjvSU2OtSOHmMmsGRZH756xC7KVA1qkAqN804Jwu0VuuhkBpjddsvVDLqje3v2m3nL
h5zTS1tgT21VJdHXZUQsvvhz0Wgv78iD1SPk+YR2zahc3rciZpMf52eeFBLM9/SY9DjfqlSjQ6zb
d1LGJW5nUqhFfIg4QuepbkDLdgfpy1S5Kvtq9/iTdlsoXRGEUmFBxihwkGic3/tfXWAUN+MESyRE
t2dk+bNoretijwSIcRpmvDpvOEF+brIqVqNhmBG3zL/us1hCkb8Z14ZhatZQxBes9XlMqXQ7UGTu
rx5Re6SiqGkyVewrQnlFhZl59bZz/PWZuRHC73Jsl4Ys19lPJJQzXIWUTUvQQ98sfOJjGJQDLghM
3CRdRnYgJ0pWSkvZymPAgbVQ6m6EFYNhBWO23WMqrTTA2mmIt0cCC/JheHqvDmKeZaBZLfjZnKL9
xQzTB8jiaQNHniPLowo/DRD0jQ3TSQg7WJKEGm7Q7QEQYqEcbrdZZtBM8wQq+EK7avRAflU61UK1
IM6lBQj45lEm+RUzdg5be0cdoNyXoFrYnHLc0FXSrcZuF9MNGg1m1dVQvUkRd71yiZYH1upFJBPN
pPf+zvy4jzq7qebcZMj3hAcxtCyWTzq3iMvb7eYS9Aug1Ylrr2BEMcFgECSozyc5CZ+1NKh75Iub
2HSM2Mbd7gMpCRgyvlJ6dqXNHduj0+mu/Y6bfkXdLcRnNSa57jCY2xLL+KdUoNwks9oyNwZA5+uk
YqYBlMW16iAQo4yPXAgTb86lsa0+SeP9zns1pE6voXKrT00PvUfocYxu+Xa2FKAtOYAuHdjT66My
FJ553ILSmOPQET+FonJC+SlQZuUC22fgLn7HPb0KYwdSphqJ7EyMNqcoj1iZWREFPOFXwMWs0jie
hCzzye67kiapKNJfJs2li3lCUJNvVjFs1QmnWhqpYQA7UM3GpnEmIiPbTx8EL0TKSzR57Sew9Fvm
YS9UG7afLzBlzsnTKW64SxuXgDBujMiqhxIhwBvayFCawp3R7vG6aZAK1NmPW6A6tOS3J5KGdkle
dGfANek9ommsco7n5BjeQuNCOUdP33PnFHrFxm6hkww3hhS9Ds1SyuhmnFkDcznpxf7rFo8geQ+9
BcxWz0O51qiNrZ69M6d0jL0l5OyIOS+mNTVHx81nq1n40h1aTSW7zIKIT3LVR1jkHPrhA9ysSGS8
eHZvKDgufQOFt5f4uEaVq5ivjAoNQ0QWFeQk6z1JXLtY3xCkTP8Snpt0uQwFviBo9uy0PFvrt9Fu
AevVwX5FJSIiZUnpDDjsXICqGOTLeVklMnxDi/j24mqF24JSmI6HFnyILgntY/yzoL4ypiZeg7sm
+5bSYP9djRUyoReuGM3pHkc+Fqq7YLj0VcQNGce+i0elozLIUPhBlRN6eGrqmUkN2t4uP5QZ+yo2
tadPub+7IwgGPHJNgLceup4Md7kREC+1AemmhcfwiRjBB0hLfaBeebHnpsP+y7d+RDwE3FCgxGOi
/ygy3obeOK7TtPTRBeiigw6i68bzh98/hM3OWgnsxzKV6CMCuYvuI8vOAMYadrcQjxwT9u3FrXdx
xAm6AtNLyfzcIDxet9sixO6w0GC+oAlt4nSqC2yKDEjoVED5gcsEIsmscl0nm0WHis8CTZDfT3da
qBcA+caOUGxFhh/a+RG0tOAWbU/5K8euwRVXrA6vzF44UiyvuNqQwcnkmGgIV2zYpNWUdNBe9M6d
os24SoyHKvbbfNXgY/6W/Ru3lDDCNAk5F0aHoIeow2AHJSNq014oJEnjkhcqEH1xiaD9hcRN0zZr
2fjC92/kkPls/TLk5CPYV+eN3/gnh16SrTx1DRMQ0dNY5eoRWiZGBRuYIHc1n0FhRO3qu2wZF6Ac
4Ks6UWU8DXf+8kN+vjEJW2OqtB+aC+paCZGL+eEHbLx1HC/AA9G0g+zgXccR2D7rzFDMC7A8hruh
59nI/773f1gmNQ2pnihzL3HhPKbStq7HyNoSt7XkX1wbl/YkI/W6ggURSiIOLIkcdOzDysKS7CN7
YcVqn0te96QGHGUFEO7RHwTqA3+A+zhTS/DcybW04Obxy2fZ76gP8wBGUTAIP43VU+SZOuZ/NOn7
7ndIXTUZEyXUnqWOw45mqmCc4HhsDkV7u3tfW205u7d3vSsB0Kk5jyL9seAjT1Y6qfzeqss5GjTS
2E+3ac80iLVA9Eo7wGbdddK/0IYMN3hBT24nqsMDNrwTW1IOFDEOUu85rxQ7Mm7aTzIRg0PHSCVB
DWDxevaBycozp9f6Iq0Nqloq+cXy/aIfvAFQIThqQ4qBMB1wvLee+RhKEt4Sqkk+AROTvaldvph8
uod4rXIjK4BorrkenQysy8m3G2yK7XbpNz+RwN/2ThG56arQ2/13FK8onaNjkqpvUtZ4H2xWCUzF
YixkJH9miotikaYEBIpowzAm+W+Re3siGGOKPpBO4n3L4h/NdRLurlGKBt3ana74o9vBLuPGhQ0K
EIBdrgAdTMz5zA0lVgE5u0eAmlGj+XlYRkq/o9ieqZDYq6Zb01eSuMBW0ZyT6YjW4ltVZIfR61hE
KIqsez3nrIzTC6ONIqId/xxKSTGVbT0xDJRxk/X8J0WLuTUWz8O6PVSC+5fcztehQJZH0c71DpeO
2ck1drUjzMPlt+BlgS+zwkps1zzHrd3D+ClijH0KO8zUvXZZQzG9vC1BcnLPoia5Ml9qN6eq7m1U
q1XAmGf2qx1QTSovT0OKeHR4xZ6HMKW1ugnFnbV5WIb+vrhZ8TOpwsUydyFcgfxQrZqYupcnOaRK
zNgH/J/uCqtVnCHYLURbY4WQD7zAQU4OM7L/uxZOAkH1nJjCK+uQZgt7Fie3eQ/Ek/D4DNEfblr0
JGogvBvkgG//4o9pqBTxmGBqShu+Sz299Fz/LeY4/nANMPYXqy+IREaA1g0CBoRO0HGNNdg88k29
S9z7NxBuIaBdleDr3x0wcdKrc7qmW46thNlUAXfUAZGuTQbi1KZZa28DmP4mZUI44ifesTC7YeCW
kvekL6NsRBgjHSh8Vobwn0Z2uiecNG12UBt7G1jp73IVXHARM5DyHeNrFQ1jRo5nGxAlGqjXM4KX
Bmk18herdi5u9BKNVflIWeG48+hWHscQi9hTTzwMLsPgHK8aIJ1kNLRdoKUCCrIZjEABPkNruJG4
R6a4jr2Ty4Z3XMNjJDiQ9YW3LHAC0BNB5df/oFkQ7DbId7+RSVc1bYtBWpzixtMK0qpE/kCFy/dD
cFoN7lMO30oDNBeFyuxusEhfVOGD15Xo75RhlcwthCBjx1YbF15Vb8uzNIjheHXJ733pUYafXmJw
FKbPek2IHca/foplOqT6SYADvB3yfZH9oxY1xRe5/fsGd5SAsnqs6k4fyqQ9TFvFD972OTupJtIo
UOBA8cQNJMP2x2HWwg47N7iu+V0Qoabg9AP0ImtNbg8VhcD/mmuNFItilfi3X8UyTuWAPO410XBi
pVUka+W93S88Tgfu5sACgc513tbWy/zwfcM4EVLZjdyIEfHTQZ1YY/DFLVEgrNMOPP7CyUfOU2rl
H1tlGL2AH3tUiE+Eizd8eZolMPgdTJwfVyrQqANV3cXK8b+qiNNFw+hIsZ3jxWyR8J9c+tkukkI4
PK2OCPdm8wq0Glg/PnTEEka+39/Q57rL11VJ/JBh24HodHZL2L6ON64RqFXm/ujnm7Lf7yUaWFF5
f0pknLaZ2s9ROxqQT0x9XdUIqPxbo3dNglat77My+2SOYQxiQAcO9aZH2B/nKjMOfbi0zmU/0fNt
nvEB3ZQpPDt1YZMWymKv9+ivtRlUgark+a7rjPHy2DfOYrwrYbaiNrDiCeCyU4upD4dBTVrbrf3p
kq3FqF7HIO+pDRNzEslYUFJxwWDjulSUuB9m8PWfsTOkoM2Q6+gnkZrUP1DSvHSGtYmpcGFp2wgd
I4D0C83bXs7CQ1OSEZWkGKDWjqlwO8CXHGMONO9gei6w0ppSrTwSyKFCvXJPf1d8r2BHP73stII7
Pt5xLwcFXMlVJUq1M2VNwUxkIxoViEG892DE5jccsxmplnR+zDPLRFrYB54iCtH5zz2nZYD1u4Un
CepK298lwI2d3odK13+2q9ivo6PL0tmXGtBVNV2TuE6mv5JXG9dq9YG5rwsTO/wF5FL+il+g4hWE
g1YNw0hOQ9EtMWYLVysjEucg9Cdxgm2d9Wk0eAxc7TcpXSgtFJVGN+1QX947lqOJ+4ApROgF96nQ
GUsv1JdrKCTffbW6p+XjHHDYF+gLOAEJSxEnXXLdttZfowgKvnL2Jylidbd5eZttPz73QY7oNEp7
K7Lhpklj39d73Zl9KXQKH8gn8xnYScOfxcfSAwX762KlkY/qkhfjk3RvY1mXiDKDn90Tkx5mKcq6
YAoBm4o0+iDkS97uCJZ3r+ccihEWPqQDrGkks8CKXwqmE3UmVlSHRPFEQ5oPlUc0OSuwSY5mbdwl
iOwiZjwEQNE7kbnGFTEok66Fxy1D/zpsRvPkKXLF2iTZrx85X57EnSNGBTXQDyncaHl8iB6l561s
foZ/N+Hata2l53y35ee1JQLX9PBYwu+zhncRxFMdweuz957bwdtrbUmKZkmCrTnizN9Kkp0v67F7
gt/stPIcbVf/ttXML7E1YiDaMAz/uTWTK7mfH+zzCbUw8E/kl+ihRygroGkCcAtb3lCvS5t7Niv3
CszpDso8uFsJ2p3m5WWsDUt8ytWF453bcP5M7P87la8xb293ERHKyKLLH/p1aYlc+81nZmVDktw7
RtSb0fVJnyPGemM7mQwyZo8HPqddkTXsyB9qZMZxT2E0MkhSYd40O/nu9+GVLPIlZ19lR4SX77B1
cevnvcp8h6KYa2Se1TbfPxbfpC3fG0QyZcpDiWiHJwxyOZfERuBQs8mYNP5vU1f6ZhAqDLuS76PO
sfElaHQyG8w7SIT0kZtYF0BpqHpW9vDlhmbONJQTMUO3c/AsAtRrHJO8y++4o+wBIOp6jEZGBZ9j
8rblTjsYcUDvnMDrmyVZpsTz+lqmE4F0uP4qRaHMINNyvkcOr9guRgr0m/PH9KA/bgkitRJ3qo0p
GFB3W+nrfWy4ntbd1MXDbSyg1jiT1YfHaZTEGF75shY2IXjF01Vn87bAE8SYIuHRB+1sbZH60qyr
1NOReeiniAt0k5o8WDgERcWUTDKMdZy4IccwU3uIfaEmTxQ9t3cTyq49rHb5cS7dOVelzqx7Cw8i
9lPDbc8MpbUp1OIUgkA1lTeOAoZuaTcKBueR8ERJwBZa5Yh17+fnhVVSVLjvwJ+uYHxD7DIwiSZv
RZmlNXMAXrOYNsc1Q53YQUUgCobGD/0yJ/Y1MhENdMcbhF53Jzz6MrdsOlEPcDuGu6xLTcB6uP5L
alCUZK4I5MJAdFvlAx7ykdgffvKkvs7kztlkfRqrrELy9VPgb10i/TETVEIykKsjLrMZ3F8ygeCS
bI9ow1iDvDa3zJSvmclsk7rHUGbir5lYnkNNNRNCOJ94OpH4M0i2qqrpwWBovrdNlESovFAWhM+Y
HB3zyfnaxA6Wa4f6NIVInE3OMF6Vp/vecw6itGV71RVMVgWucAU8MUOTmeWXCtYXHcLrWeO3fRYk
WhuMJYqblObKooy8EW2Pt8yruDMRMxvK2GteIm9vBiWKiAEHehm+b64bh8kPkYPfsfYLkKmSVJvJ
7OXllb9XTPJnW+VlE/yJbPK5rsZxXhhWoU2NB1eqyJ+aED5AichAodaH2Pw3aR/Cjh6sQsIFSkI9
r+loZwhZBVikOjOpMKQNjKuGj9FkBA0L4tmj7IaBwuwDsyH4GhhdXpty8B6RLdX2nYl4mk5abo30
A+qYVaEWNzYlPX9yqGLvSATn8s+c0PSS6GMdiDRXci6yDOZfh109OyHiNx5yVZ1Kjx0VeyTFVti8
lBoQxoOZPZmQTQQDikLpIIr2LrN5ce3F5J8f1Mhchih6ofuru7Wu0YikQn8RuFYHg75LMYMTo6MY
QQp2PgVGbx0afgY5/FcjtIgAN1yed+0sjFs/Y3eDH7KGbyYeenhX8FQgJVpjpuE4v7E8TA2RuuuP
JjbQ58XK4RgozLXcxIXXBrsF07s2fg6ershV2z/7NWRBdf7CXPetHMlDswL63VQE+ZbcP9+jxN1p
RsTLx6OZ/gsFO4zGC9vlFoAhRTCwLiUSmGelLOj1p1Wx9aS02IgHq9ngHJAXMcJxSJhTSQScITsI
OV2xbz29gI4mnsLX9QMYsursr5x4SRR0zp1IDKYxQKjGaSV70Ko7o6ytu1TJ3nQYNsIq6pbgea55
wZRo3YN5pi9pG7FxhHvfWZmlDgPKK9G7kvVEzPKKj+hpgFMh0huMnUuASZN6v8BFAhNjfxhW9RWC
80edaY4eVte4s+/qhOuZyocmTdbKMjKMpIpjcC39Qk6hFG27g9Dd+CEfl+rt7J+iRFhIcCm0Eyxp
vSgfBe98ej137zAWKlEe/lHs31LYW9OFkGPr0vz41hd9fPpUtr8qbYsICcD0B6UNbYXeGmG+7xVt
bz3f54eESLPYhiK+6HGjlsDjPIOgLUl7d/xnBLW888hV+ON8vZHvBQPypiNVh0WthYf6yROiQnzn
dQEBqJ2iFYUegJjnKRBuwTzI2Er0RkO9HKzg4kKfiMIq974ALC5CuJYNDuAARfSr7lVf7BotS4Wj
MS8lWtsV5yhH05hvY4tFSgXErU69vuAa+YwT0OuUuzsiVfMf0TWw2fUeRaK/1IJKDmKIsa4hOI5e
N47m7lttATBl01b9crfy1JB/z5fNXLgFkQ37EimVx55AH9NczWBpOpw5qPxfjhCRbC9RCZJSQ2pA
w83LffmESFbfNHrOfPwlX3y6DsdaBbIFrYxLzrl7Bgn0dk9Mfj9bIh4PcRRg0BNN+cJ84CIMKj7A
VWw6aJLYvEfR9OAOUJEvTyp6tIYUB37hAqLiaKx55laDi/qMYozxk2UQTI3Kfew7682SpuQ3lGRS
m1N3FR41tuhQZrFBN52eidUA31AzK7IKhNwWX02POZqRbBRCfI9wJTSu7LbaxSrqdZBk/vawF5Vm
Cm3MRcGtXwZuY/tMK8Ao7njCMpFId2RmXnPxK4vUchYzlIJdNUdj/lZFCh0j5VcQ2E1gm7H280UY
FFVXd4oNO9Wnx6T3DWBoUf8gtbmlj1LvHmSyTMfgiukOwEhkxfJlqp1D4RAv4pvhPY8iRNKpEpcR
uYBkMB1oYe24GY0C+PEFpDzzU19oJap8MvPpmVYJId5OuqEQ6Pb+d5RKueu6LcVzTUqizDIf6OxT
EZSau/hcIORa7R4LpFpQY4BmvyWGVRx3to16VwgXywDpGY0A52h2i1Mg9ganKCkTyNExNqSn0aCL
ryhJA2xDG5Zi5UIev9Or28NZXrT3qONKilc9aXROj1YeIKH9Swiy0Ji+J98M6EIE9BM4cxiwoQvy
V2AUdiUlr8tJfdJ09+b3H3Rdl9fcYPEGz1H5Xw7V6IcPcM7QBL2kfR0728pSbGPi5xMncFLdie23
4/uZvkEfcEONFrVsfGm6Aw8Fr6lPvMAsKlGVd2PG5Fpp27WZKV/dwrDji4bm/2zqHZSev7zoINbj
SQ311/78mnVdIbWhklfIb0AmPbyPuEObsE469bqhU5FwojMillWPXi5Cr2gFl9bK5XEMzuvl8gjl
FU1BL2kkV63a1ad/YpUfTlo/lA14Zxl7D1EFLnBSjE0MwOPNuC3mlmECK9dioARqzsSj4vQE17c8
NsD0Jkj5hcwcnK44zPFUhjwjP3AJaZIMhy/UQKiNcLjXvK6oT1FV5ObBIhjV+oCrey8gIdvnrNed
qF5SkTVO1NJojShOAMsfp1dWiylqeMqmQWx8yd22xAZ0O4ynrCMrmWAYwcLkPvJuIvlEPPOE3a7R
q959Gt4T87O7wAo3ctZUE6rLWJbk8D6ua5yfKhMrR2clbgCLlLNVHRCHcyv/HLheCv0j47Iv9HN7
16JZd8oWX4H48YAPHmEIY+tfXL44hZKbVrcIB+n31IIW6CfV9DWrmHMdMimlJ+hnwx+YHFnC3APr
p+uEO647+NuYLxgt8icZ2LwGDRvoDEefF96HaslcNr+0ZpGMPCKCuKZ8qh9zt9IoLdr3vblpkvIE
1a1XdAl4tJ3LLMBYOe3WqmlN/5FOqmAVJXlZa1aSueQRrGunbs+GfM0FAw3uuhu+H7zyRZ0Oh59M
kq36Y6JmsiATZSdYzix8foENvl8Qa9eTDLusi3lTW10cUfeDrxqHhq+yt4J3D6hycEbreMklCkSM
6l03qpklaj2RY7Ar521Tzp1qZ40R/hpIJ+C7e5cU/kFs/U8l4CHzlpy3OGcvwg/Nrml0EwRBqyII
ZBOtzZbCu68vvjuZxggJ7ApLd45+irjGNj06aytIPhbrSI2YH5Ei/JDNLV0UGzipxBHBRyz4Ay4H
ADY4jg+VEz7JUZqzBqm46A1q8hYrhyUfTRspPNY1x6ibXVxih0j3COcCEq9dBA81b80lIddlnyfa
aa8vWSHUkVU0ppdrzvU5Ie+HpjeEnOo8ssaPWu7QRzPlRC9e64EGZja51TUNzlAPS1Dv1s47E8mH
6QlcnCNKKTqqmp3V3N3oI6TEmKz3FocBR8dj/VbWXngrM80ofuxDx1CSVRQyMmttwL7xeGbYNQRq
lwYBl+x18sp7m+QjojJDnjR8engOyouPa2iAJfMCeQWkuzC3oCXwnphow0/ka0LctsLDnmlfvy1P
s/wh9V9n3FLq4ROnetCFiYPS9ifjHMy/qDFI0D+u4UzudM28osIMkum2E+Jg46auPmbc+drRWq1h
Me7RpaJhub4lAm2dEaqH8aR4UhxGmKrfujcDKVC9AbnETjV2tGCZPPeL7UkGqGTJAf5q0SOcaRNN
+rnOlQtw3lquFdAPDy6T0ArXVbBFC6Efj8HKIvs5jr6OIgX551jcOCrNObgpEASRhpq4cRC6YQLJ
4xYgiRJ4N+ZNPvQi+Nz6iR2fysTzh7TudFSucIIG6lWc/wuQH7M/vC9I4KWiEqBZ46CMuXsjY0le
3Y7SVncBZyYYDMt6GXPI16q2p0tYeAuB0OC+v3Bgr6VnaQ7mmQS+6EgxVjz/ThDwPaZBYmuVfG9L
b4YLnIN5U+faWskymjafrG4Gm/8S5uw4/iPDf8yXh2l8uGpUrFCfq66tvAN1uTErKAsPg043C9F3
aevcCzWWvXJQhFj+JMZKjIWFgZzwJdZyXcG/90beJjAaiA+LELP0CRvcJwXEitSmLi3ik56t5zHk
9vYfIwqYvDRPx6qrpMIQEpH4JlGrZwEJx1d1WbH1FJ7daLc0dOFOlxBJImafd2PWGG6Npr7QvyDL
/vsNIM2Io1w3c9pvZDaJ89FFlenTOPuo0gGwCf+NNKir1Tefw+VR/VmbGum/ZDtOa36r7awF1Cqj
Z/H1lj6SsEmDwodT7PDPPB9DRqXWl9yV5fBceKkJX5jGQVxlPnmABhLJGsl6HfVr0FipW8Nw2JkF
6mSFwFbOQXqAkPtU4mAURFVlHD/KpkXobp8PdFu/YjOXC5qKy6gnbdT2/YJ5YMXyzxsmUvmXs9hQ
puuTOIJE8We7xGuKowqebXiGYvGmUpCae6VLETiKok8NF+kl18ytarDOiap9Y7CP1FsyeBqc2VCq
xZIe/LT3aewNxsDuW8gP/u7E12SvIA53b1BUeHluW+MGY0+bzLo7arvETuTS5Hbc7GxYywyQrSTa
o55zRJOB9LZbD1AxB8Y2TveoosJczwhWG0V91aj19+xXqu7IdJBJ0lTPl8xzKLL+9jZPqwAzdwU0
LRufczIQ6jSeS/WnnfXUfgI/Ku519c5sjLnRLncJPf43Z2P9nC3QuIdrc4YTX4aBxAxjbfzsVrqv
wU+5tHCg/uka70o1GgqBi/0k9nSfG9I30DZoTI4QDR2yuz2EsnbeuZUTUeTQUMPLsGAnZ3nJv32B
D1xUltE9V8jQG2rFLueW6Fmlo9NDG8fBxzqb4NyXK4jGigFrUP/gVDBkJfQQ/NzjXoUviu0K5qpL
QMsvEBFKdRwlPYuvYl8Fy877zXS9bAEnvkma/lKgkNaOHbTqxYzZASHzBnxaN2gNW3W4gytCKMSw
n7xQkA1dYcaF66j2RsSpbsl6X2AfsJvz0HZLFkSIqNcsMCcA/LQYl80lQXs7vFYT+ff94PSp7LUV
/esCZaltPdvrNDp3Vzl5Lsga6Tp/m07ja3nz32iTd3rnHth2tzd4mBN7XAljbDZ9PVmNVHqV4pG2
+3Az5f2ueo+KoW0dDj2GrU/aRQTxp5dOB8BRysIzHjnWwO2LTMQYwJzK5npV5pUvHQ1dqUdleBZy
z7IXsfKZ0de0kDaDxBxj8nV4goH1R2IRw/dP5oQai5XWsJnJoYDW0+3bUn+meDYWKECzqnzwUJeY
hADwStoT+ZJtKuwr0KC5/64ntjRVtQUJjcv1WbkviByO4VLPMj0qgFi+NkDr032pgsDXIUvkfoM/
lanPCccRkfjDrcWBIv+ibdAZnZPMU2gt5IuUHLf98buEpvfXckG7Pc0sHFq0My27qezA7XNzizWV
jqILAF2QkpewQ0nJeci3EHs4hM6WNlHZcyIEAbEOSdL7WtVdv2cq8DZwGD+AWpmxccEDKO6hggy5
//XJftGektipJsWSZ/K7xr/y+kCZKN4ixN61KZNUWcDqMsoKh5dbbJSXp1j43lwGbALO825O8Sgo
IQQvxVgk96JWbqXNt7in2UgTB5plYKk0r03fwdkcrlpKxvB2WM5PDQU4NdjtTzpLp4CQqbHNIqbi
4Ci6mypK9MZiM8Qozh1RsmNpMoeVovTSXuqSgad11SPLiud+LXdoFDh0BkoqJiQ8+tjGgnBRwcj+
OnmhysAHqWOfq0ddsRp9uAURP+uP79fzzJTgLl/rb7Jg1x3Ft0bjYVpalBqPWz6s6UWDtGNguuNy
O2pL2TCEH2cvhAo4QzzP3/cUizoE8U+CorIfLeBylvGRItXbn+uKA75Gy/Zu8f1dJUnB8wLbe0wN
UdpTOffJ6GCx3UI2iVTaKzD5G+vnrSAeZgnduo6vSJ81hxRuA5n2x0YExJaDA8wMlFMOc+gvP2V9
5XAOmPJmNLmcHpwqjB0phuDHD7MD6uH1EDJPss3hZRGdMAhIksqkm3++w2FCuemgH26IL8J+4hUy
PVDj2qLKf74SHkJY8shxsX5Mw70nkFd7G+KsglfMczoM4YzyahGuKpYHkG2l7VaSZnzwh9EPj6LO
+duVBfaCXXl9c+qvdKNSBBTiRgOR116FpwDZQYnReOxPMRS4gUK+CVrp0Vl0KpIcHe6KDGtkgNUx
4SDXRkU64FxJE8zVd18XtscPEa8bcKhDRjxG0Cq7RCi7Vy/e2bL1fMe0EsNCd/hwIqKy47Xv/HJ9
FaGkK/0LmvUnUWPlm2oAqzsImycUleY08z/M3Bg91ODqN4Ik1AKHtYKLN9v3TYKyWa/lnEgMy+C6
3/owZA2ppGr7zsQ6XaVpRalIu/qYoYpKOB/DAF1JwONX1hgkF8cpPSL33BF05tGxNNGfrqFJZfSE
Lg1UrEu5LWq41YF1LdsCvvFd22b+8/qf8i25T0S+pv4Gh3wa1oCijaJGpne8UKejjASJtx5NglEO
FD6VOREArfATRg2KvV7Hk5Ruk1HHLymDMDaPmHPOUsPsacqsMj0fZJbLBVw3oMvVkAso49SPRsP+
nJ07J2FAsa4E5X7tA50kUn8uugraNr0zV0Cg2CoZBm7yWlS0SV4GKeIAkN8NqmbizrtQ92ZMKwBj
n2ydFPUeNgR+UOw25auoaeub6N07qlDup9GREwuvgCmk5w1LEZE3tNYVoCss7b5be9xiHxKZrz8W
D6H0HfRAGtIvfZKImW7DfSJP9EKi5bvFOq8lt2ArqPfmHgLjJGbw1NC330M8x2wqNn4CEm9XALQ5
S1sjJKqD/YP1dT8rC/dHwByl3Hh34NrDoyLYFsdcM0CnffNtX2GUR2XijxBkjHqEbDnvkVMKZ1rT
h0HxX3yscUwIq0AZpQT6quVEv9yGFmJ/mE+1wEKJYJiLpm7Xue2UEbDRCbhT4lCeXA+jB2Yaya+S
v964sI2Duxusj8lTvy29PkcReJPZA4XiP3x+u00JBC13CUb42iJk8d7wjRJ9J3zUpSfK6qPz10Lw
ND2+EwXT09pCYph2yHdYjZhDOcw88qbObE9oHBt5iKE9LYheWu34JLRzQQqSnY0fNk3/K0l62Zjf
W/6LLqGarQeqe1HZULW5pVHxsxxr8lddwET3WZ+PWrorN4+e9JiLNtxI/9jRTp9NsbUrz+j85JJ8
w2cZnognBXCcuzg6mv8Hkih96aihniD2Y3Ac0izTAbHw33Wa+QW+Fs5zEMvr9J0SQ/VscIwUuOmC
osLCAfD9nBw7fG3bXwnzi+0iH+NtCEIUhLavCDz9IIV+FMAetKIqDWoY+qfkDbLdQqlDvP/Kh8xA
0ECQgZW1ZrIdFsFQhbGoExenK+0/cOvXYFYVsW/d4eFDNaDMbiJrX6EYoV5nAjs6uppWeBYqEhS4
+7wk0WWMqKn7YS1YIwpRlyRcvwICn3/S6WYV5FaOp0lEkqHgKBzscDomRGQlu1SO1O2BWrhsjsZU
Y/Kowgo/ZDPD9IMbW/gPjY1KeVM7lZFuE+JNTP/KdcKegQzURgkrXcb6OKMpTuf/VX6wTQ0B7Wkc
Qk7NfAi3TJwV8uSNebqtPTzFax1zdW900SfoYftfqcVBJREjuLdenS4CXESO4nk0rzb0LVdeL4AY
WefLN/0JOS/MTt5gEiyO92/fxhBvJD8md5EYk0/9e2rj+1kkZ36GLrjo/CQ2Dy5SUaT0PY2D5AaN
sQ7DiPHANW9kLsURXGVXjhnWi22CPF1olCbnNtJiJCBF3AAtn17RnIeu1vnwOKEdA6ZhcNQzpi8I
LqAhi+0cg2z9LXlZ74FDLaxQf0u+BMqHAVeC2+PuXX1ldNus7yegEpeLA2OnI/Pxa4yuFWTa68hH
uk/OdaWkZ56yavlUmsVDiRytJttTXqRiOKgGy+LxG+CC/AwF+rZAVUdz/6zfVc9r7x1JywEy8mpZ
/Rlfu9JIGBhfFk48EFlZkDRXr/fOpF5U1TUDmXVwcn/u2muHrTJ/ECwOB1vtW02q4wVAlxqfS40E
+/DtDURjGGmVMEu7KVjTHqokS9JT/TWWaZHF/dXnvZ6A9kphQjJ2OIFaxRCzEQ4s8ScTTeeRTPhf
yIcISQUXc7rFOioSc2nxNjnOlXSeqRiVWrMFeX0cRQ/EcDyz+ySaiVLpsk1Sa+5QDLSMFS87VfE6
JS/Kl8qk0onli4COPZEdvLJC95wGo+B0t0KFZJq7xUWdIFIlra50xwtvnb7qsBMRpskzrhNmYBEY
/vamX9joiACJglvN19fceAuHO8T9t3crgPLk8Kk9ewFqTaEKnfuBzpR15kcd7WQBSf5Z+wmXUDHA
oUymWlePWpt8XrpkI9ET+YWqEzw/Tto8UASDBoXSDa22J/MY2RwOXB5Bwv9QWPXPSnOxZQ5EBHAx
LqMVysvJEbFaBTm5avS55OGSxdL1m9sV8yRYVSUaWSJrtqy+VzaiQ//uvH4MZDOQZD13Xs+psG5v
/FnhKP9bdLIUD2ucP8pNGI432GMMwwU4UCd/F3VCaGrhnqlLGHVKF/nPGcunQxZqVPZ3GmWuWXN2
J6WmKLi7UaJgswSdX4Opg5TvVSnQsvCl32vqkOq2G+WxPnuE2H8+EX98NnXigznyZFdmJfS2OlpZ
ozgiQp6tMf3YJYmqs1DvVOa+/xh3UgYPDnn7tbzLpJY0I3yy6tDCJ3R+orOuheBlUpyqTP0PHbzk
Rw/jad1f806Ffyz7p2MAFf2vJbUBldtHrNE4IZhSSVt6gIXHT6qL6OIDkKJam5F7/qwIsGnmpREo
su+JI0GfuUNVXHBlmtbxye2RevdqP+Vg20DKfi6tsisuapGt8RxebM/j3OaF8jZ/MIhKpuJmxZhp
xYIZGudO7DleJMyjbEFgPNprqyVzyS1YsVq524wq2JnqD35GYYZO5Wtk00HZ3UtvAB0XVHCskxSq
Jr777rtMKgDIT0/tsXfuF+UWfST0mWKscAmleOaIOJl0rqYjUeXqOvubO019plNcu9RFw5IivTBe
3iiT/av47/O/7bDCfKPW3ZDDnPO84VFCNXbynX0vJOal3dobLB75HZVxRpZG5aRPrYvfAYjgVs4W
GRyaSSgq8KlSOuv6VvQk1dKLb7GsvcdY6ORG56tVLF/0uLEPcT1uwL32kClRhSsYk8bkmNPWSu1J
qC3ms12KtsSmFHCphu3w+VhGo5besLuLqqvIf392KUbwQ9qOg90mTpcome6Or2+yggKFk8pm5Wh2
gjiwV+oQ9PKq8g17xPkFJ4CyrbAtxdLxAe+VJf+8xD5vKRYiccyfK10Vy2n0g+r09gnAS6CKx/g5
4V4H9pExHeMUUfSJDQGIJHCLGl/AtbdTKr5aOWHcE8dmZ+zfcy7W59hFEM52MllzfJnNXYm3pLbr
L7CQDP8eeRs9z2KIw0RuF5YmPvjHaobpYEAfAmi5Q/KB3xlNU+M+5AnH64tYLngrU1okzo+skN4X
FcbIzcmqDWYIa/hkl70elDkD+1hEXmJn+ZJIlPgap+mhEZbkfX/Av0+hOkLZ3J7Ky3A9arzvEBnt
a4RLHN5I/QQe/DE5F0bz0EnL9O50Af7X8hJur4ccVdnHcasovWxa2cjSBEealmlx8w8sBC/NxOmT
DRNm70y7CstdkIVueX0J7YWlytYRtQhlbbggbj9IFA3x+dfyT1arMWn/lPyt7l7kjCpFjW0DIIwQ
gB8DZ9aNv2DBAVm+tPXeAbYhYOnmW7l6zDciZiqHHRNn6zePuDk4KWUcYdbpfjY89G9XozA+uUGc
Jbdv0XPLJczHrnN1dvBe5Ilp20hCNFS5vtZ4kh9vTlkns/XQTN6MKVC+8LfE7jp/eu2swQt3OgzH
tNsJ53SnoAVTiUeAtpBspI3YC5zmrG0Y8V6tAY/Ea263DdgKqPUfATIjeK6ibY+mS41NuGJtEsAj
RwBKTZzhH1IPcWYrLtQgj2xCzUcj1uL/9Xjqw+L0mlHISe6uSO8rqEjLPCkfObyz1tDzV3aHhbSu
72xOY6Zpjvw2b+5bO2MAkjgPmO538cUy4tqs/8qFwRG4NKX1AcSdWe7pkvMoKiOePzHDvcKuzYqT
4mjIq5Hm/1FvuXN5J7G/5kPVQVG4wLL5rA90LEJHkEJ95mtiQzXHkw9VqiyPJHpN6i407UykD7vP
myZ4WdeMKHCV/elFG13Ownc/oL7m7/+BsvPAP9YAkpgmLm6olQfPcAHAmxMJ9Uoz1NbvvyB6ZRwO
Faj6wEY+gYRk1lAw4DOtpG3atQ48qrRmqJV1rnyrpiqulD9qZGm7Sb+KZEWY+8sDbMjEqMdyTJgS
r7p00nbOexI356AO/UXrwooBRTsNi7hPmXi8g2wTtZyRAYEqItzEh7t7YoHltTZs2RbsOCNiKcj+
Pv+0ot9w/Nhlso6V+XXeNKnmCHTIYT1Oyp5jvZvT/ejSIT1a+QnEd0LYiGkCFMC/jSvMErYJyDk6
Cn0DGCZNIaOnPUwcxtRmvNokNePrsZtRKk0QFw+l3NyqNKt8PYT22jVAq7KzQY4CP8kYqZdbUdaN
p58pBez/j8Kk8z3q179uYTTKGW/fDLlAHB8nJ/s8n8nwrt3qKPMPRbY303dwbMoLsrD8WXwZb7xK
RNSbXc4stZwwQ5QK22iAUZcjjENvL6pI2/QCtwX+2zkCLD8XUb+RqR4vWF/GD5wlyFYG5++U589O
0XS5J02XI2cqPv2A/XyzSH2S6Kp0aBJvwnKiKT7qRyujdFFmVEOsA+TlKj6idl6wACFNqe+tvsfN
Z1iATRTEhoTCl+kKgQijv1jFj9BPfUqPkrUutBR+asZScR0D+c3GE3lm0wJ/FUG+wAeA6fb5f+nt
gXjoyYelE9Y6SxKlNPo/hSWCBlCHgUXKv9+Tqi28wv/sGf/WKqM7WqOn23cBQYBPb6C+o44/dpKT
JiulVBo4T5+qz8lKpONK5ymivF20jhc21moH3ZGnGSR/Oe/1dxcmEW2aCrPTl3OtsAxc9mHMFv/g
UTr32Apu+zb/BvGzeSWGkAI+mAdblQAExO8Hkje6DLzeKPPQazC8aWX6rm8qbHWwAk1th45ZOiSH
taLpppuVYwD0CODZt3DwLb7BNshlwcqpYNAQoPQxTz50H5X3Dl5zJEY5tYFwZhTWsKaFXAA1nvx/
A+1DGezqts3L2Ira4ohuKNcs1O2D90PQMPo4zvFksQHlUebwgOpd17TXxdAbuWUMxbJ+63LxH2Pr
S1GTQyjUqCsPDmeOtjAE9Th3Ohq/EKV8+keXkH0RXFDvyw6oQFIMCSXiL8sVQVVWKqhW6PKKN3Kz
RwApm8D7pVScjQAjHW4evW9VLZBU6XwxAQKjDBFtPUMmi6j/aLEhdWFgMDVT/27ayAViX7Y5L32g
R28VftMeVa5+wEoKxZ/q0X/Vkk1rPVnLUd5U9S9ck+A8sU9mQ0T7Ja1KFQXBaJWNT/RuQrD+hcra
anmcBs/Qi5KcxsNwGTmR5QjShWmr3tMe1MrYvNmF3/r78BqDSJ1Qq3vlEg8NjCJ6/Qmjv9bP6sc2
ue6nvhU7c4eIziHQvKDunpusVwkh7auecWxfVczlSkK/Z6Pf3MJAwNyONhBwXXu3TxfV4SSPWFtR
b86+kp5aDKO+eaHc/w1Qvvik3wbWH0FyxngIfGQwIhEzJECDCRa7rb8nXwjsebXMs18g8qKGlkSw
5+KN3JlONob3cGP1WaaLOE6mo5NDMdHWNIHmOLaDRllJyPbxDdQQykHM37t4Tc19LvnqAOlvN7nS
t0WmhVKNkjzpX2R0RbsIPJ0Y7TJ4uy7WfcI2Ixi+BjX6Q6kvkxSBLRFKcxfNAEI2jKwvpXK+XNsZ
GC3p4h8bSh5sdHqyOkqmKnGsb25FtqEX/TK1p2mxmeieWdn7IAKFBr/vRbHegzg9AdyCYCqEkk2e
kFJ8CDto/2C5HNgg912wcKX4Px5rQPeEmfmAomn4buTKMVqTnuIe+ruIkY9D5B1j+LYi7yBEIEAc
kXnxvRh9yCGdvKVwJnZSVFcuxE/pFUW2TmGmrE9j7Eaw8aJZ/ewDMStRaCNYBxDgW7OzW1EG0/VM
hZricYQBNL7Q+Prcz/mKPywFNozDeDze0AzBBjaYh6jpljaU+V6qI9aOad1nTVT96B0ySaJVxaLg
mzVxVAABaPjzGtxoNPaMp6EIKi42Bh8ebJAiihnndJDk+zesFcaZiAl9kYsk7+s3tf03zF48aDpX
VD7h6hIuvTNMX4gLBudqVknlIkk+5upj2MU1aUzVWHb+GIxGJ9ASR3dWnFUCoqer+T0mJPGdfbm0
LUy45tYTX++6KWlmBZXcjl+HvvBKH+Zl1cYsNVME9ARv8Rk5ZcqTijyMRBM/vYptfAABfpxomf5R
PWBiActd8a3yEibny34ZDfmaQmkqoUNG7Sx8oU4CcZXlKp35/sI7Nyrtgk+QRGHIBNIT5KD7DcIy
YenYszIL+0Zut1naszOOC2ivEIO7U+c1bp9wJ5kOZ5K/BlTWjF2A7kynIZE31XxATJd0SRkH31j6
LxmgJBSB8a7CbYuK1vFwYSbwDH6mahEvzXUKW1toRCji2dJ8pXWwy7QiTYNaCkzZV+VXEageu1Ja
fbDNPCumS42Mty+FrD54oTs7tWplrCdR5uEvCb47YQydQW1sMnWcPYLV8G9cpP44QKk3Gt9o0HRU
HRtgFHDQzyZOMy0Gvdg+WKSMHnwLj9SbWgZuskUQd0ojsK/PMYLlfrnjIh8SBXG+EpMLeOVvECj3
nqbW/55KxQI8AoZ9PCEQ/XVL6bPS1YMVAehDkmPIOTO1hjz4vX0TMDYkNUPCWauewigkQdxe9enT
fldBQjLfTRYZjGbMKh1A/7C3HSBh7iw1jBclOQXl14k3PNfPpCDTa/cx4Bk669Ap75pzU8pNfmeg
tFvhyM6oBa0JaH5y66w3aoaG8AQQzr7kSylXfdRAQmPDfvxOpE1zVDiq87rsBwyS9LByU7BQgp7I
Cu14OTZgWx+38hgb0/4uDbe0qjnvLfLOWWHKPYavG0YweQK0lIvV608p3s3UQuZl15glSXY52Ufh
+UmHsyrBQ37q8JWi5B5Ak4jjY3O49/0D3pEq1C9+l6tUYad7mNBqLB8Sfr01wm+HuINTh9pDNGB/
fZ5FsxaHA7+U5urw5Wvv8Q+LBCsn0CWMm2ARFOgGkt4hfbiK9ioHebCdNu68N9yZZ7a50SyMFRGV
HhbvKK8bJocikAikL2/DrimL+Wgx4yQ4HFzCQjuR8v2H0vMJ93WS90fBjgNwusYQ5oI8oOFf4sK7
OYAFZtXbs47k8ngt4y7/vRComhAD2/AS7rM2YfKTEuCuLqoqW4zLIEzH60zoocchf4yNGH4bA9zZ
Y1W4aFkFzxAQi5bQIyiepT9HneY8vdZC2rQFoieB6LDaM8n/5KukjsFVI6QxLT4kk70VIQN1NihL
MMSHPSdjyQFGeDzp1aUXwD5ofwR5N1TK1A0AD4CuIi4Se/7fgW0WNVJ1UuyaPZO8Vu+zKRlzNVvt
8Zbbz16BL2sK5fh2t4KG73ezec58t7sbKC4vwWs9WGt5dPyPb6GyXMH/DMVW23RrNJHnEgjVg13U
okxBEu3/iSQmBkkOz7AKDdJg59GMZi69EpiHtrHBqgvMEJuj8I73yTSasyiaKGbZeJ+3abGzqZ5m
aQVu9+lv/E2/HsCa5yTGmnwCZrybtPqowCtUZiOn1oqeiVvobODc31ODl/9laOxsGMfx/KdE13/3
Jkm2SHOT8xbFYhs/mU2rEsUbxviOxRTE/nIpznrLDU7aRggTNQOy2ex5ED8kH9mtwMqfAcjCUh+5
NVFwQB3+vWLJjxvww03HnfXZUYaaf5CmNQgTrf8GKh56+Ysupwxvgv3UbzOXUoSfeB47uQ5bxx8p
SBvEutRhV5DPjCuG5E3MOo2o1pTxJgbpoGJndfYDEtYji3iBASTk/OtQRVTRXxKouf75lI2LdnPT
nBEmce1Xv3Nn+qBophA3u/K///Ykf+N1XXhEhauWykaXoxN+RCvjc6rckMgGLJRkjj4W6uyI4R9u
SnMdsCcDGhCEhB1/HrqpN9bLdYDDku0LxtTT6YvVs1TaITQzyoUCSpXw9mn3kMQxCtwtYxi88/Br
1EhxdB394pd5UQyzwUiCesi4FF3HvFQOi7L0eZ490JEC0iyfAmtgzi7rMWAzkZo5Wo4slL8hdK1J
BlkFpQXv4LNerXfZNuSNHnc2RSbAGIZilZOKlsSqBnkv1rUd7FCNi/wrYdPplBt7IjTIH+Lf7vEc
zZ+EfAWWR/ZGsvEh+NspfN383Pyh2AKkeeZW1mYQ3XFC0ilTna9KY4Kv7v8M4dlGBNKjjZic0yNk
rWJHTOIeVR/JqC8SFuYsbgUqzAsbpHNDVkQdt5kQvEVN76qxu8KUZDUNkph7zzoA9F6fHL5rtAm5
v3h80Ir8mJpDdos3TF0tfYrGrXdfekkwBcfz2zW1TKj4YdaJy5YDQt1echb2grbJD8+R7E/w5Yzg
rTkuyhMF390XCQ/SmgmRvwrakNZ5gk8VvYaj489Uz0tdS/cBLX8K7tjix5koFpqW2PDUxVYqZJ0c
DOTHB9lPiqNCZylY+LM8jqmYCtkgczdMpNX1rqSRhBd2JnDavfUror4TYbGH7HBP8IFDSkKSjl9F
5MYJym3NHE7JQf54THmhIALMWYhIR3qNqLuXI4J4N/kCJJaPZzBcHmLKLnBQs/lhJFapMapx1uY9
6Xy57XQRrahMxuYZ6ppY3Cw9LvAj2swJAQKivkjD8V5/J58uVP0wmln4V2WkKe42yRfLU1AEL1KR
sii2v2ArYSXpeGc3of6mQtzrLVP1ndj7G1gZgm1WSEspQgNZTAV8tdxRaf4BEDiYCHvw7Rt2zCUW
i8q1JRJI20PXS6l1+W8aPFuXYb0BeYHQaOcSA9QV8ZGinGUnj6IhI6g4kUoBx1hgdI6kB5ar4Oz/
KY6VCYhtOnY7S5Adm/QilpicvclY1UX3cpfgkyOsHvwI5GRIyUPZF7JvXIpJ+N8WB60v4aUIPQA+
bL9BJ6ynz2IGn9fGTU6UTfddHKHTTqzqvcovCfNfohRBWWX9cPiRMDpPlr8sgeIoT245rPBt9xPV
OioenJoFoGYSDwMm30fARnxUxZ1toyJu9TSb9Qh2kSuvutoBfJIOXdGOlWpWkCmS456UgbCEfd2T
XYRpBmqzjMCB2Nnq/SH5Bfwo2DWTYsI0OyseqFHchsY0/DxOeIVV9TOLE7AfUPZ14zDX/bDwDLE/
6ihRRVLWrjpAQSkBkiv7F2hJnn6uotVO16yDNtTiB2KsG5K96qaquKx6gmBLl08xMfCyW7O4l9fS
EvqVivRJ0RI2snws9LjdA5oblVtL+ERSRO9gPEhgbGy4gm2jqBEDKuPhGVXCaFmu8l8hC33SOYqt
yNt14bZYkid89fM6lDM+UaCwTFzxysW99MbzGhd2x4zSkN7Z0nSFBStnikI1330K4OkwgkpGdlIB
fq3kYjuQY+SPw2xycmEiYEOPr/8/3Am+W1FU9py0MI4G9h1FfCYBgluq89cMAiTCKq0aO7vX6sXt
Tbi6Ghv6V8dBgartmg0o+elTZnpInOitvY3zVxHqa9sLk79yMzzzMVSos/uSAl1VaLb62RkW7n4S
t/ckSrW/S9E44d9YsAxjwWSMB3z+FpUIMZ7eUEiUG2q8DdvdhHFrdRZO2aO3zeYvghcvQfPssZFX
os+QlWHhmEo2WwlfGLddqqH+KW2DdFE5VjyVevDohaRE7RYGKFJVU70mNRoEflEKcTnEd+sCwlvo
dxDPu7X5OAP20o8Yt1tsaJKP4pIYfZnZ7wJ3VU5e7SAYZ8BwfS8mCccql5x9XGI1KrbH3i9x2qdf
WrOISLZe4euRJwFzTO3SQXYF1Yr6kqjU2iUFv3bYuuPX2ATQWQ04FOFgqF5JilEmCoVN6VJFKNs/
/aXGPLKDcZ4hVgZjSMn3QahJ1t+ZpJ0HBWSk6SxcZmnKKqviFcs1x++Ls2AYLJQYhqUphRA/5IVi
ikHaI99Rz9rXwnBpDkYu8byVQDUeNgdjFWdP4jWYMExUkIl8sFT9W0dUEDD9fKCdHSeYeSVGieai
gkSQ+d+UzVUMZYxft5MeJWZYKXMWQtKNclPiZMWU8sfqfb7ChZBSkkNpzfBUpcfEVz+ZZXtJuy3d
y+SsCABMeB1dstrfOqoTnz2XdHuB908pBR5/pGSoakKLifPS29Uyay7XaMdpawPukgrC3x7XY0/Y
TsfPCgEmiCUq6Quh1ejtE5dNtRz5rmKeCE6FtNi0mI6ozAkLQstrmRAnqB+0kzD68iFZkIsYzo8N
9p32osFDtqNdyCBwrQZYYyESoeneqPvmOaKyxpdwHRL/lOF21BYsmDXSA6AYyOZHTS+HskKK6sDt
WtdLGq+BjsYw5vZvzXuOYvh0Z1QG2OkoXR1XnGDMawciga2cqvrKxcuWoPwcy0sZ51zxssyguuFs
nQfiAWaT0TaFCl27G5K4d0dkIAS7OocAjVgT7AgxAhg87Rx3K+26oMf4WO30Q7zq6/cJmTjJWfK6
qwaTXPo62QbS7c20OT1utRlu+LY8mK7TIjVJwkpqcAZJg/NDDocam0Ua23O7LqoqTzgOAtK1MR4K
TNlHAQoa/h81Uk59XJGRn3GcqklqIlifRrQdGSMrO0ethAwaNpYqjHnkKdoizD/3pKp7AYVuggD3
1tRJNqWbBKkYZipHuDWbtA0IB69/WmWeJAss82yvYoGut0lA59J4Xurl5DMD1T59XECy6CEKezPF
feWRjq4XuM0M1rL2nc2jEus/szhjHWzBtFU0lkXd9GWR6rHdEhx8coX+1rPBwQDetcO6+5LJhz7P
DolmZ3pe9X7x48/JNybM66yvuxdvg6xQxmTsphGCsl3FDGTA6G0+9gkldxG8eHMhZ6iK3ZoC2fty
M/8eod8SoleOmiZHthdZB3cmBH/2s0gyYcEB/oZjv70FLQ0SPSSCfKCqoW94UzdiOcFu0AAeDDn3
lc6m3p7R+apPNfDcIpxKnu98d8h0JEhxt4JjfYaNIZ6ghlYkCx/IPIVeIpwh3ep5YGjXuy0VsKFC
QwpxS3/YzpNeA6ZljVspYaS55TbwECHCxjdbhOqgs4C35O9UZkjZDux4QqNnQdjRC/lhNYxlvScH
/wBpYIem85HCKZ0rbrcB9pWIfUEa6/WA1opSJZUv13hnKic7fAY16ln/0/hDe/z642KoLtXfTrik
XTK6intUElN3mxhM2xae8RJY0aQpr/BrnSr4GXUVGlgt++jCs4KnoEA4qdmRnn4C1q5a4uEBZXl9
Jx+DwRnxpmN3qfHIFKzURduWc94NxXkP7leoemPIT+Q+qNlNlXHl1Lk3POnvwoa09gba6QZ8XtdD
1TUJc6YAydPR3RSCoEy809lAOnvpUGplhTPdFCKloqG5o0BX13Z477K4GR1au3C7tXthaDUfyUp8
+REyvNp4vN950CgTOIjxA6ycNCYdrvBoma6I3GeUvwhz/mm7t40zvsASg1jgmxoj8XCOOcA9hNit
pYAUvPhMnasnm4Z6stm9xDpu+LZnlR9r3eh3m84pTbIUv0qTMpSJkFsCyHimUGdfb8Dk65Vc+FRE
RFo1q7qCxOnFLyjzwHF4bwfprnStswyZTj/e+YMQA6znoOpWaSqqlNR+RnAyaSVBWyvaShbSNly3
TFQlsPiZwgBx5S/HiHO8vSZXsb+M1g3b9Ktr9D1Ngxys1qN8xhnjhk7SZujhcbuY654rLnhPIgGf
89vVBgUxbkMHkIxx5rSkdZMy7yClLeymIR47drgLtqONRQT0wwj9zvT+AjFezo7kOcHfn9v+sRN1
V+P7Nz+UPsaTykM5liw1OkJ3R9iO8ms9ghuPFq2bNuGe0PkLvRs1ijcSkWMOcHDQNvmCvg0nN1hy
gEZKS/1QhGpPIpINGlvpLQWAX9IaFCfmQLfh+Y+Jze41ESYp9gF4q14/JrbzaObSCTX9kevrbEqE
+s7FHqFYCRDKNbTP9ZFTtoHikMd+uNsQZhjC8noC39+fzSwRQuFesddpSgiVEGBTz5GQjhppQ6nv
l6nXGzumfqfriZZHsfcddlnEIjtsILngA8mv5kRtT6yHu2MEha5flMX95VrGCWt/T0R6Cp6tCEQr
TIu16uVA7+Wz6eTYEO9AojWsgDr9pdCnUdR3xQ3YuLGdo5Z+iJ58T0UpyNG3L1DaVdEUAsGSFTOT
sFbhkCAXSnpBeaobWai1tasy3XR1/W5zNwQe0mkiJKXes1gbhOx/GtejdkUpKlAHVZptsTbXqPs2
qX+iub7C9J4GkshdkpF+5JkbXckGDJ6T7cycMBvoeQQiZ662PJF9OEoOJE+sqb4JLO4SZWCrmbuj
tYZIbZ/TSA/0I62VyNVNQ9ThhCAZXmr8+Mm7pX87O6TqnvnPJkemCiCyd/9DiOMqvCUB+IdWiH78
uxKWoj9ODNvSrX6x8OU8EFgIRNrhZB582+Q6pnVecgAqGOKfauVoBbNPKlxmtg5JPevuz9XYIsxP
3xC5gZNNm/plTFlyhs2G2frtj4AZngA6Y9LzW1RxNjT2ANX+M3hqLHMIpbI679HLak5gAJixEWdM
i/bjZDzAQ8o2IzP1TNt7aVQgiri71YfxYK/GijazBTWOelw3BENJsW/+YEYtmaXv+QjKmNiCdWjl
NlrqQjrJpEVQzuYXTyS06i00kqgr6UuG5W10TmxBUf1DXteAZYbExyfgLAQKIRgIw6YVX4+E5Ba5
3n4OoLxtORwCf954lTVLellOf+ruGu3uK/hGS6YWKOFXuKvIKk1zIoo0sbzFhgQL30SaJwOdG5qs
MGeh95Uv70aL1hj75rn4v9UjZPnA/3WX0jhq5XXXizXpEjXocF5VUS/ZCj0Btu1m0A6DNA4wsDqk
cLVxFwTMFw+JSF7eIYu/mik9u4PdWt/ccHZ9NsMlvZV6WAZGf1HITG04Sm2ySwQUBYakCrUMBye1
5oa7zdcAlSa5ZrpVzW3dOYIIh0Yn/kIb33TNw9ecCHRmZwN34uMTlTvGHLAvhZ5XOY449cAtzu2g
3tVLVkkmYUwVb5VmwnSA3CoCZX+TAo9YpV6c/zeMe0DK3adWEMVPCu4qmXvPZuBdHgsizm3gKWRa
MCzpWX9bFRlHg1YfglQfoOdNXOc6tZBpU2OQpHuMgYQxqEBAqfCeK8VXFjgSCKR3VWJv8NOqpAuN
ufQ4g+4u66WnRcQ9K94GRPCwE+t7ljQ7r5HZ7cnhKYoIJ31672aqwH7ayfplNULVZzPf7ZWIn9Gd
AkSE770XGdHfw6ZexHrv3UehUtZoKdIPWMsJCDgwk9VBG4NUSrbkJmZSjQq03Dvw4rYynTu2mIDO
91bCkjqEC5CYAOzCFyYucVbgwaeIqPx2yt2bcud2rUs3pfyDJbgAUhOq3c2BC/TjN1LEM06plzfX
vPpTtGpWvic+QAY8K6ZN3gDoRc0bNp6e3Fpk44UdzgZFVFXKEpk8NURoBBAZ4QU69u6jXxLRMJXL
FTu7630UOygaQMecuN+ZABC262RY/gIqcb/4mc883vJm8OAjHy4Cr032Do9EbqU9YdIANaLrwV8j
RmakGzx5JzPO9S6+dcv3nncQuYtDvsatqgwIEe/70iXqoClLpLyx9lPyT5RK1N0GHDeA1T2h6o9e
4ADU6ya0PeOcUTt7nzFp2+GeB/JfaWYih1fJgjgBD3nt6cmpIPI2cCsV4nddcRCVJH4+5l3htFQ/
2kXIACZ6Qb7MxZl+QOQDkGEWHb3NgJuUJeCn7V0NPRwzGWHLkYoOBhuWYMjx3shz768AOg9/uT0D
ADUVQww3httC3saFpgqWxGzT0CUItJRYgaP/m4hMUdFkK0H1ey+NXoZafGcqD8EEULDWi1O/6XL1
Kho3mk4rN2lgu75J98Gr1piRZaar6GlsQQKiyP0Z4qGoeQDsIIyDJ2Q9wWXv7u5sUeIWLdTsrNol
6JGjXlJL+X4g8pvIwrB4VGEr84uQ2J6qqLM5F6SEkY6y1OqTeOgRyllN1wn0L4nkH/PaEXgO3xDq
eY2djh6pyTSrKBJ8r7nduinreD68ccsPx0blVNPpRsWesCVY5cmKqENh178qmthET0N/BG7Ak7O3
I5b0Pd+u+tlT5NkkCozZTcSfleUHh9r8CRxgXom2OwV7QDc23lY7jw850AkxibOtY5FGTUwp39HV
7yUWBz+sSRs35S7l8xyM4GY4JfS+hcgwAc3RddttUpHWK3C9zXEF9WdWRVyoJgJHCf2PeNR0DKBk
Jr5enI8DKt7AlZYZhAELsso4UWLoju/6CLO28SwljbczPpT3UL2eKhojTTu2Qmtgfm0wv3QmYzb1
sf2Vllx/IX9Yxe1v2UhsEwJztIm8IoIajjfgrDKeEu3aZ/5StXzIBv2TmgnyF63BzU5tCqI56UYT
HzwaNOUn9gGL45zsuBY/mIKb2wHb1M7yHWIRzfVK5ktKZHGPBIf3EEsRTbzYTbLgTSMZJ6fZ8QyR
Db9mtihoTPtRWuJJfebDX1vg5VyEu+b3cCb6OEOvSpE/0icnpvtDjDkHZleO+AUtS29mlWewBSNC
fKubFfgDbqeg/VEfD+4UeZGznqUX8qiMxy0tS3Zxl18aj3+BnODzg4dpIv6IVKvCxUkMPiE0i6r9
/SZVY2lYU7BL3L8byXJJvMjGgOI4X9Wdx/I4Mn5QYAASQmVH4JgTE3Zze4hKRFXGDWrNMZEtSB7k
JHVRV5h2i+WtN2/5+5QHoyUptNc6KA9rUY4/zUr5mRqdOpqxXaI4JMTZOqwab6mW4ArlqKIUT8LN
p0u1PoafPFYzAJNlTeNEqVc0nkywSjXGSBy1ana/YHwNekSf00TdcR30SYiHV/vNG1p8+U0H+CvT
V8Bt17gx9VNbDugBxbIV30ecVay0JlcE4/KQ+XVQI17qyHdu6tBBb5SOvrbUQdg/7aY/xF8zUy4W
NbcA9CPtNBL6R8LFMPeR0fotqi/yk7bDFGF30koDWczZRZhKCXNtQNlgPHBiIKAxaud1n1xkx7Z2
kIEBWOUKTLaSeHn+Z+jzGw2XJm6MmMmi/DXlUgxKA1w+yV6lldQ+4enH1zmqSKfsFb85AjA93z/2
7yTkK5OQB0osACiVzRVhHbt3fBkBXb8UlHWtUxKpD0td3sLKGwmN1tikaJbCx73FWOEOvm2mtrqb
S3bB+SKtkpb9E40Ve81ZDgfFvYGO1vKHMDap/EhNxyTktNtRNWe4z7R0R0OEZTrzOtKOQIvPlDMz
CPiWHCZF0EN5HKZlyILELspUeVCiR/lDpYoOzi1Dhpfj38cPQBgVf7Oym7PnPhqyctqeYrRUN5sb
fydt3wEHXyLpK4vxDrFF/mxXtsXz3kyclwI3YP+thaoRc8S2WlG8DK3IZSNHcSWE2gLPdCNaUutk
VC/wJ+21nj2o2N7uhtLHoZ4QsjhmFbFYZeVUGv0K9GKuwQ8wBpx2pBaVKrtuNdOgatYDGi/yBPMS
2xNZYW9nzNYwnYx5V4w9prGehXrq088lBGSda2pyV/bS2HkniUlZVvrrLqh0C9wehLQQSSkh8z1H
cPQ1AoYgHYaPpRUdtHFWZiBL7CUS/8jq4N6ZuVAQw8mtM3W3Dfk3DxE2Him4n0Fk4wWYsX4b1kA8
2BLHIKFVkHnVE/PFpuUtq7Fs4Nm7AsINp/VolbF51Dy/+0Oc/BRmi/E5BfKtT07CCRKOndy7d/ww
qWvVCPSWE/jX0uV45TZRHMzoJrGzrUB08P5k06f9lYodTLmqkFxsRXhivu8JSGpPQEca+i8tB1y2
cFcMYcFHsESjAUcPS09Ruksw+Z6RkM1LTjwU7DATxAaH0A5hIZRUlvaCTV9fpNO1yICwSEVU3QNL
zu6x0spdEt+VaUitGaN6ITRs0+GsXDUQD12O3FVvgwCgl1u+W/Dy2spsUGXCwI4tUQo4/UJEvSP+
POg+d+tRdWJEUsaebIyqEc6r1sZhzbmzKqqC+cCqe4AqYGy2HURIbK5dlkoglGj44bgO8Jm/z7AZ
arE1vFkfFqDYgPuUXf5C/sg0/VxTL6nJd2QZZasPdF1FaLM7+DSOQTK96bEIbVU94W4YgR+i2REm
98rc72dvT3cFThpVKukt5htUz5MVdtbEl4Vre6BHBFbuc/rZ/MUH3Yh2u9pSY6uO7iUIxOjTfXJr
cDgjsI5gShUYTq3nEHciQtLoxlTxa865buBA/vKdlMinj02X8GvAgmpoGF0CPPwypHC7GsjSs5ro
ZeSajb+INXK7U4X9o2OFBuYTfvI9QcW3HwylLYpli78TxJsuHl+DlsmVlOiX0Z9qdWdBqhJrenKi
y1+dVU8jSYpLRIR0b1WvZIer3PQUd1enyRm82dnjy8ULedhd/el3SMkPKYEncEdWEFqmWdwH/Da/
A4ogdonQKpSErzSn+3DKKX1a+umijCI2IOaXYlyhM7fPrC7J8+NcdEXnxSRQ2VgHHEWC0D7LBmah
aNv6JxHpkcGJWkdCUDwRoV0OXp61ooUO5Jjz43aQSERsGWuFu1zV4z83gOs5L+ZCoxwbWaccrwba
ms39eOel06BP1JI3Q8HFWQv9l+lEoA8AjcS5xSgR8hFpXvp1CpbBOg5VkvjCmjFbkGvT10TePx5a
Fw4Y29LzbvaH7Lo+l7BL4+MjEZFEIURGlCYtYK/qO+vW6Cj9BDPJuGdYBANfUDcvuw+9Q6Y8FMFc
GjUqZOJauBtBBI5EkBRWDrRk4fx2pL6CaafxG/mNGtAiRVag8HWUpF/EBwGXUmRkMMlbBRERu7A5
oX5MeyV3CPWjEFXGcYd+iTmebxohi5TIK9y5I/4JvQ2GmCP+vzNug9KMO25xSqlaYXJDkzF/KbQz
dAAYVXR4vfZEyJrx5+obXQRNqHP5/lQNONUaJ+5GnoEoVazKFvklXjS+1UhRDIGX+LuKEifaD940
er3XIln8VnSp6mL05v/USTIrwGoUBme1HrWRNB/8oBSF/JzJFU+AcM8JKJqb/UfTz8J6E09EQ/J5
LuydivrxwaT5WtMTqPtLneOMo0ROYMhuy4tIs4Y4mgoBpGOCeG5lq3FBmiPX/ewc9lv/UsOUFvXx
aesDWoh2675ndCmOIy1HUMmRJmcB4+1hJK0OsBfDhFTCLv6YiTvowVOUlbesJ9bl4qheta4mR73N
SBGphVyIiUpZ07+CUPZuqro7hUaw4UJuOeP09waNpNB0ZDtqPXbQ2LCdSbxFHgQxO6Ujk+WWEaJq
wXNxWcO0wgwhi+yI+WOLGGe1OicmH9MQPdhzYsD9N0rSZL19W0v6SzGigBnlg4f/KqVGmxH6qy/j
brjC2Q9LpPeG0todPABtS0u66MIKS/K23i+exZLigFtJZePw4kR0ym3p2PximNbq8qEs9M3jvt9Y
pcih5UdN78GmTjEK/hbbxamhrSD46s/gRCYv1GyQdJzutgJ8kmOCqvvFTzySlCWiU7pf5yLFQoIX
nwzhQpc2Ghf+kOm2JIP0XXQ2wrvJZi3gZll/IfF2snANC0AL9Ze1iA7huccyBD2gzhS92cyAJHuH
pLfsGp9l/ngjJy1jerCNUWM893Z8EDPcPlH0VcyjsKBwXcXvz4QAyfL+jCCdj+WSWMf7pKC/MYI0
s+a4c9x2CToSQnu5BGnZjK4K59zITbZTPxErz1nigdh1fYABBG8wk4JD1B8rJ8a2v8kScZj8lEjK
itSwfHF6hOHt1GfF9csrACwEjWcOS8LFmf+UQDm0FohNgEF3hqgOpttiggKNXnvJFCeDyQnNLj5E
cQ/QTpVoCwfkvZXh2ewtQswc/mP2uc8OH8NWOU2g5K8QEdOpOaoSOu3wZu3DUpqB8RF2DPirXDG+
5XTpgrYfDbceg7XWnbv/2shiIDxwP9u4Pm+b38IDIMSheKZOAmcObWYSUGceyndGc+9pR4/BbGii
aVqmIJVb1RFWGG9DH3r+D2aeSNvFD4IY3jbkcFRaMf4KWVUnjdLQqSnDNWoJQvPriIF4j31lyW44
mNY797ianPdorc5esozQGLENpxFTQ+CeWwHl66GdyndeqQXQhO+FBPOSvwvreEXof10fvkrOsyFn
2+GcGuXrI6h32i2bur91gVBbHZaXg8pYfQHVzxzu4LHhmkTlYPAL5zxBm4SgvBpYSn1p87VSxmgn
qutOmriSuXy25otmsVzPn2rJKOfr+QYNlcSpqEjZlvZUQIIV93DseugSvKF5j5IZGfVPjihbDg83
abrs7uxeMmbi3yXFeenA//tfbwgRF1KjZG8sEgI3Mbsu9VPrgXKCtALy8t35XN8591/5s86zAkvz
/4dfRrT+gYRLpLuF1UdvDKpDYnL82rbLecNduUPv+3mjO/Nczufy4aE8WqbyKvJuG5c49go17zSy
alQRa0tjhkpqVuTqMZLQeUW3WUvhcNwWvsyEV5S/0XqZVaQmCXUrEU1TZa9Rt4r3mLlZf2Cu54j5
NrDmjLOm/gpckiWQ4bV2XL53rm+of5819/W+nxV3IczAX8+WUqO95/t3mAbBbNHowrwv02YEjBks
URNFO1PczputMydAOnvzsX/ciWHfivUp/LlBrz2+FeDHSMsfkNlKCrGU0YQuB4GYbbqG9nTkh3x4
Cw7wGw6SzNAKShji6I65sVO1B90N3uBcG3rElqewT12MYG89IR8kU+xyVk4c80mvZeEY3tSw4U1T
K/KOGfaggGJsZzxC5ut5KlqkiSyvILdYswRSuuhWuyGddtrIEHaR4InIt4T+98QMYaNXOFtx/MDX
pJxA+B+iD5MiLty+XFqntBa70AxxPDIqbEJole+100b62xfQ3rNyytDHo+kl+2lXxTr0UC4F8t8L
zZzk9dBx2BElMxy4D6KT/M+bScW5nVkz00IHNAkwVvWERl3tuE6gD0jKtfgZ1AJuazyW6luYtE9Q
N8IoZw9mrPVMKb9bHRRbTOzYRlZkWHj5u925gH9iqLbMDYVHv+JeJvE3YerpbW/8D2SnSKrf6Vzt
L/+UYXTAnwVVL2Y74HkFa0dwsfmbu2uthXY3KGc6juz4rLidCH5kld6+6CZBx0pVc9MP5Zip8qr/
anv7U8grhdre/k96kpmD/4QBZEIHBmyV6UO5b/vlbef9QLMkecaDQJhTwyG0KdVxSmL4K245+rK9
uo63R5a3uH5jZ26qXN417VkoygO6XvlNb+uRwuAirVvkE14cwhHzwKf3Z+kmw5yVaSFJbBPHET6Z
aWsfYiUyhnCj/Ruc91c3fjp+icswXMmExLFncxCaNHVIS0gyMQjYHp6OWJiOrDYNzbsHL6pbNqEc
sOQt7R3QSIe1xxJBGDosC3lNwVANdBceHjBPMY/XjpEmTGraGNOKtQx1RJuVl2zTD0rXuQUvU/RR
766CWFnnOjYc0wl/SlFxNIy35wFYjhd6Z3oo6e5dWR6B6Cqf7LoyetWp/Ocmcrh+7p5HATGwT15m
syx2HdlOi6RkSqSRlrTyub1CrEIdw8jXeK7qJJpyhqfFSJ9I+/lmoKfinlIB2VXXE8tTFGAo3VMy
A6lQgsO3KzD7jjhK9a+/c6cm2GzqfMuJaAxlkYjgUpUIz2ZDicJA5q8ORhlpY9mNB/yHzH4arpJk
ITtqe2X77c8oHjlDIkTdF7l50DWPTKeH+wChULp5C9+kfQcvGt5h8N9PlMeLX73RN+1CbOx9Xvii
pcz3HGt0cw6sHRWtGYWLtM2sfuZuM4WPrWnC9Xsh0UAsViDWRGxzbIfmt5virpjs92gBW3NWHYC+
EaWZvOjc5ac9mt7HP4s2TlRhEwDdB4kGhloAKnF45RXEyb6vO1PeLkO7LTHAC9VGMPDfQnKHiZyn
B6lQqMdXVb12OO9MXO56BLZlwnn8Vf2Tsj5tw1ZpAO1i2vHR2JQM0nHAO0phsMuZ1zOzR7Ofe3BO
X7p9PxSIwXpQeiaVMeN7J0PncmdOLBUacp4Rf7RYD7+GybxQCTYRPafPPNRUr3X+eQvX+GmN5LMY
lmitJun7gwwDu2OUb4t+jM7Mx5h3Twza9Aaj0OeZsWrJl6rJKPFbvU769GJQXRTO/HzFjDgMxsXH
fD/rnNlR4MUJ+G7HsE3IPkzRVgKMmHTLoy26j14HYVZA7/tMWygMCmPuTOdyuB1qMMjD1cF2DanC
WnMjnuB6r005BcQYYw3JgkV4LdhIenblix3L8Ut6OMpxaaumkyVShLU24cOBFHhWkyB87yLXyeHX
8GhidTZ+6jUmvnagv8RVzBQ/sZtr3//rNxqbnFFwMn7yAmjHoVn23Xn+SsiZd/1Rp27m6yOnh9a5
2ypJ04txYknrvli7GIAsanYksPiMz6VTSlxHQtvobFehiL7E018uavAefBreMmQveQq3hL5cW+q3
uAyjWmXI/IQl0Jh0pccf2H44KwGtrm5wpDKhftuOTKo6p8abTJZvSr7/e04V7aAt6rpGR4PaZY5p
heuPHjCZvTpQapjRzMnX4iUJb01KZCi8neEwKvk2UG6DZ6UBxFeP/Xk2SEGZ3aKJkBT/BIGiRlr0
y/OQQ3seajtoqxrIGTFGrrrMziOtPZCoJOFIao9UAKh6Nf1qBvWJb5VJqImDX5zEbMym8Dun353d
QJ0riLmAXJTRFXGacw6+Twd90q7uDaYn3no2Sw+/lJk8itB/7ypycrUM0Zt+3LF05jBwkyPNCXX/
afPwEPRUjaHDJbSPKbXRhmw+MCK1nYDT9DyCYWBrCUXUdxo0qDe9BSbcx/q3USJSfWPpNAvgVfVK
xvU/r1KQSZ3FHo+b+LSvxh7BidoU392iIDIn/rBgCLJLNAAviTGi4cJx0DN03weyZMOkaxFlVQpZ
OU6g1/v5dPvvfHE35gCEw+Pk0dUuF+IO/zbY98Jm++ybGOaOHwTq0Ai0fWQaVXJtwKGm4LzyQCUl
T5bekzy80lG1geK8K7+YeOuWxNBuG0oiF/1IludYnUtZnpJfk6cjc7tgBf1IPcbJ4pc3Gh9r9n+W
83jcnjrh0PeAlj0QyrU8GN4zpLVKM5ITCfAmcisFDULAQg3rt0PKYOWrwipGzn1s8P0kf1gEZlWQ
piFfrrMAm24dRamVl6IVo85n/YnT8NzQGbh2A1O4OR/oj2iCj+/cKa6luQp1vk+tZnP+2bF/HKKi
jYvL8o0oTyQZ52snzSRhV+hmLFW9QSsM7+8HQlvnBWvO+lQ0+IZg/q9I/iAgjonhGXYjKrHjL8Hf
ndd1XXRk7LVDKxQELhviWrDM6BxyvNSrZXjn+CvFfTO7IxHearhcOARzk+Q9OflAD2swdfvbeiGF
ERy16T0OfyWhCUD9dwBgPn1evxkwXKLlrB6vUNS/Q+ImrjtOYLfNrqaQFvyBYA4YJD0RvIMnz94u
AwbgeQNvVSp+gr5aq3liyFWLMsivPbERULJfaMFI0w/e0OyjMBwe22B16HMXH+1maEc/5SaCaIH/
ScX77ETigNZMWGE8B5KILh5ts9ygDKRtIpYsjYtzsBTuD4mkBwoDoO/hkmdIuptay5LRtDTlnsl8
IYsTLlIyU4IYIQKHCKicCIZP9fVS/ZA+k2h9nz0sQF0zOVse7rRPUMPqcO/R6zmAGYUD9W73AS2k
MCaU9FGmQrGDU1tCYiex0mnVuFc1rJkzbnplGd/gfxcnY+zloath/8RpzQoRT8JWm3WGwJmJW6TR
BHQP33TdY6PsM1rdiDC3BPHCLA9DQN8NSVpG1PBnNHlZ0vapomhTyWJMKBoR4xPnzPwsXm3k4zR7
Tnzm/AQWnWrFOT7Wj9/hvrOnB3CKMp6YwA/bPhUcTFTigJXfN2Jv59JfJfnn29XrI+AesDbDqX60
+qQzb8UocHdrJv0UsCBxg2K5djExQf81AYNhnLlXvZNpPEPTHtA8+VxccUnQ/DKmkcyqnpHAa0Wy
6I047DveeLUDftVF+IMNlSw3Lru0TxrCk+xLU0pzIUwIsHryX0ysYuV8p48Fogdm9msMi1pPpByj
tEOIXfEed2it/9PSnf4Jz7dZVOZqro1u+aoSe9uB+PDuY0DM5SDaSfQR7T2evVXVcK+Z0uxLTKCg
HRQB8YaLszIQAffURVKHsnN3ieqqRQckZSdHeEboiYKwd+I+nM+0IHlRSKkLzqEINZzIIR5Z+Muq
pEoEA3wRyAJPgiJWLtGPXb2CgcRADjbISmVCiwUK8wMIVZ/6uByYFBno7eANVmP8fH7YX0Z4wlZM
qs8sNr14bd+SYXv1iXTCYvpHNd43hBsVMXrYeOWQH+jX/RhYrb03JzrSj3Y0OMQNKFhJMbPdn3lv
mx0OpAG0gBroOtfZC/nno5Vd5DwFpMRNsmJK9z9ggfpMo0jCiw4/dnrVkHFEOkScJPI+XfVLGp04
2HOq5DrGntU30EGMkysZpIE4YBPUp1gDV6B5BPC4nmGplcpytzviGJ7xYjoHfbV02SycWPsT592V
SyIaP8qJbxcAhFLZjBpFxHDfd+hSkvBm1EoqhHAMPtGD69foGXHrqrQ8R2tyfB4lN9ip7aSZk5hG
NjQKPsbi9CjTUwEQ4x8l2qpk5i9li9T42NsC5IHct47IincU1QyeG7pz+55qGWkGIqAjNK1d9QAL
uJwHcTBIUMH2R6F36fzQu+E67gm353EI/XtpqNkHfT2kjNOtuf0WKMFdujpXxIeAudRDGxybEraz
G9X4rCQ/GRQMearzd7tVGkUJdeOxVpsQaRfwuScbyOLGDWLG/TEwQiPD5t03gLWHnAog3zT5Tnhm
wZmBSV11TAKZ6eZ7RbbwTj7Ao892+kJCKRthShE14uhI68rWvtcLryClQU1TULgLOccL/U2LRh5V
lthB9MgzmxegO528hFjwwupjBVkzOqHVUcgQqXvRHlq4SiUkYsxvo/JJ+7B0m++nY4TYIstlNf85
7EDQyuDnr2Qd1FHPzXX18Vt/XkV6zrybULhtxbZMqfSu5HmJFuS3lgKRD0NC4V0OxIn+cyYvVqeQ
U91/FmMZg8vlu8frNaE5NuX62u8epS0b/dZggbeqbNhn4LGhx/YvD2DNaxudC5DJ5cWaKmA/wFqS
gIJcT8sBMAbfo/cTiExIIfzu41rqdTeu22qVRhpFDaIPi3k799AbfZ8Wze4U2hTmpXuH6e7/wXk+
5dyxZ/R6se7dNnImpPGtJMf4vIe/1PV19i91DRjciQkvihsVeXWxWpVXwfZVUmA22ZZSgRykBI/3
EjnLpZ19CRCIy3Bv0wFUjEafi61NQfxVroxH88B8+1ZurMghiXcjFb1PgGRNaOWGaset2wUVjHA0
c6pT0Oj5+yIqYRHJp6GKetgu/1gWPR87TM+HX7tzBz6OlfEjCyMXyzPr4H2DdAunmZwGtYO7Iqkd
oHe4MwZ8A+P9/GeedsfpwGbS5805RNFQenDhPbhRRFayYvGHJKhVAYhFDY5ymTha1q8zsRvJtwkJ
Ngy6B7S+XEO50sFRzlWguGfC6ndANRzCVyinPQdHubief/rDO9rv8JhVt/QzCSvdlN0MWws4BXBZ
bA2KgAN2L2u2ey8WLRFLdwGiJJ/c/unIWsl0n263SPP6Wr4KYI3uyrQqN86+j04zB8amf4Q84Y72
C6SAxW5tZob9JxrZHZPGhdAOfOPisHoC9HMuLl6mMC8xZN+GwfKV2T6YGN3DB0Y84ZINMyvs6F3/
Rhb4F4uC+KpC1TiDhnGrlHKw6bWFoSDKOY5XQRHVmXOstmFuhHQSjlYlNHwA/UUfr2K0Ibjxmqag
bynqu5aF0Ldquut1jyLnqwhGqAipP3zHCH/L1kwf/roh+fAYx52eSEjGp5uzmmhyQlbkaSSVZN1b
5av/msBhqq4QxPnN03E2nPXRxzn/nntOVoZc4aVc3oyKcFszZwGfv0Z63rfeBrFzWMsq3vHSCe2e
WyjqubYCV2FmKgX6ZfqUu0my1V0DhNMP4l9PIT28D1w0BwGPewsFCqnKPkjeqbjY3frWqnlfud3J
56qDPhJ8ewjr/nwADpDyxLSy0h/cYxT/rY7pr8Y+f7uxNqh3E7IOk77UNoM7cQXGx1o6S27zojSj
zUqZ0Yyx7CddCSi1YSJCyIGps91Fhag6CBrdwGjnx35mXJFC9WA8KiooErNVtWnx9NPR32QFwSl3
xhPSvljv9Nnp0b2hNKveC1ixe60RyRGMDWdma0ndTMb1NhUCKmSskAkHN2iSNePI0wwEnorBHp27
gZrWqICL58wfZgHWktkS3wXFgYT2V7GHGPNXw7M6HSV8ktY96TzqE/t8Hn7A32Fuc3g+cwQulFUy
h3+RLoENO+NEzopJLrZqVEVadbOROyUC/ahmFrOOrvMXYL+inygIcYpK2frLg29WbbaavOX51gw+
3izhOkYo/7NfrNV9wX88kZWUWrc0pXbpjqhpdd/osGx8DRbQva0iKFjFyTITLCOp+8SudpJmiwin
dVAG73OkUoFIV5Gxdq+dk9tRXiN/WtNqhkMqQCE4ZbcUHQhrPP3wFQiVNtxcqg9EyTw+5ak4LECk
yp7/DsCiCimoV3q3Swk7AcSei37cyGqiGRXTI3+Wm0suKEkHUEE70Lops49gj4jDohgo5zs1+gqv
1lFBotNS+wjklo3FWPoGKWLF2oMMQvz7zRL0PszZwk49AgZ7h4hzbxdgDaimS9455mS6dSj7oonB
DaBiJm7jhSfhrXuyiEU2FQOuK0lj9povW5gZhNABPblKVFwmq9sYdmKwSb8qtPIX5IGPd00ekt2B
cAeat79hDng94+E2655o+Vand85xkoX0MZf7VM1wURBCydka6u6tSQ8wM/O3f4Aqouxe27Au6QtH
xtTMFnjGbk/Hv50ZCTcORloXnGH64V8O9fKlT34NMKJhqweWIL5xEaPkLXzxnqC9dH82XcRp6Eva
27xO3vO1T/AuXgsv+0aZOjHx9OR0x0lx6isDjd3nK+T+nnhgjba8zeBUZ8ZV54Zc9hExHsr5DQTb
2koOMsustbbJ/diN5+thhAVKRCNNRm+wts2Bb+YH4d+DT7WOqGqRNgN9JBGeMDUkAhuPYl624Rrg
+0E2AsQoHxQt85Ez9ozN8JM5vfwMy03anoA6iRypqGFw1Oq6qR7belFjouWAotymOTEJ2iyLDSLO
qSIOvoUCZ5Mm1Mv3t48XklaszK84/2xkws4tqiHud1P/r4JmI59AC7KaEtb4DR7r3rl7w4lBhSgA
yTodRc3x7v/qUsuKM5k3STlCOwDzz6XdYWQuG6YOmP903bnKUHESspZJ+o95NwR6lBi/HQCQPB2N
FhQXQqA4VqAttPIS40tUR7nwD9t+CHHx6Pfrl8ujjPNBV7L9HcjHCbgmB3/061+VbAIqvTWXlz5t
8upNEy5iBJlBT0p3cKjnXWgCFjkWYOzWIdBHXsGOGpCjFYwTtLvBDg+tWqBM48zvcvl0CMEpmIan
a7v2xme3N+ageAc4b1KUcKdhigXhjmwAicQVh4O9ho7QmgC1q5YzNPzuvKD9N0swt9jVusSpmcNK
QrJdLlROu0j4I8x561fyH9Glx91EpqL/jqhNqhlOB/nin5GK6X+8xEGBfXMOBgzr3jg25P4RO1YY
gm69dNh9x9LHMuYXXJ88F8NwLE+T/SvVMuP/12gtKSoyIxsXVFfMr0IDDdemETvhsHGvZkgPtTBx
9YqvLFnhBrlXOlugJ1Wn3WSjvCZCnWH44fAJma3tQC73V87We1BulWvBfG46ZsZ+HcaEXK8UzH7W
QRLtOsCtrhz+KCLJD9Hu1CVByleE+fSSbPjrGskiikJAlIcOeWch0dcxv3txG4FsD6AXLov1nwJL
ACf4ILYqO6iu/5Wi1pv7M0A815/mjfs9ZACjFjlOW18/6OyEJ3huT3FggTBmPXaRq+KlVZXk72kK
Aok+E1gTmiBEZ0KVxyyTl+O0nNCb8nVTjLywP5FTUMsMrioDPlZ8au02bmsSvGBlDs1Iz7q4XAkA
Be4c8RJ2nXfVDQgei0D4SkrBrFNlMj41gUrxYHvT7ysX5EUq0uH48fvpzG5n6JlFukfi6ZywTCN9
ESZymHtunrU75I4dJenmLYlpd5flYpyWPVwuaj2sucZ7G+kKW8zTHO6hNiLCtZPvvovzzTXFkwc3
18Ihaa5fldluIZ7+/AItvALHRBxTgW7fJmvYfkkhSxMcsLTgZBBakiAfBkZ3nlRsEovq56sUXIDf
6PpJLzs85Tok+Mit1I6rZdCEr2UwuPtc4yNOMh9Z/zOiNrClhRhse0HdeXAUDfZnFDGtaR3qDJQP
V9LwVh3TCdNHTaBCukphTAUOZ2fLPhV++22HudiijJM5EJbwTjclbXiWXi2hk0NRzmlgue910HhN
EaDkbNzR0yyIRNn9j0Ni+WYTnEwf7P7/7YGPnylGSonZJ01sZpHKKhyUhJjdJQYx4K0Uqc5OrKTa
F1OfLJ5TWge/d9Apd+BDwLnCJMVvMSHvUDtztx3gXys/iWrt1GpUKrgownLVF5IVrvzZ1LISA3sQ
wGoZI8URevAqKXQRxCbQwW0P+LokTKg2OHSmk996DOpxcd3lsLUsMz2Q8b51IulcBlUB9DLSvovQ
CE8JjC8p2/owbSqWz8KmOFqwLxwEvtL1d7Jt0oLUfy/7GrtxQpqQ7xUayv9hzOPwXs+KhnZDTKLM
/KRr/5V7ZcEsAzbG9xZ0SQIse56pv5R6hG2gi430tLpq/IFdEe9kar/7JiozyaRnDzebHL8XBroW
gApKWs0+WdtTgYifDuJGH7d/nTwyBxmmlrLmg9NFzWxzpj81mBvWiQtLs62GrY+QNuoEzIBINEwN
d3Ek5nVF2+unDesln14gDrc9zg+xnw61Z48MNSfxUsq756GlPkTLwbEBjqlDi2MRNQyYqvRRPHeQ
B6HuQ/AsRhN4tTtV0l//xCmTTA7IFamaylNx758tImjs+mdUiR44Yi6OWBbFnUsVjWXcdgB4kbXZ
itxq4mp9upZRor8DEALdogIZXbxTMfY5G/rg1zhUB/ku4fac3ExS/HA94FS0SpSM4/IvpmLEVOkX
svVJDWl9JuCy68lIX6FGIpNs0aN6tcbQscpavE2tSKotDJlvuTZw4zZno68vq8Waa8b4SvZARVJk
gDvgNXSW1PXNn/9uet+kZYPu9b73gvQYuNlHc15AjhUYcHc/SFP923H+kJfYA9OggnWq6i/R4huN
Yh/3+F6RLD5w3C3pLpt8ilvYfyEzqP3jcuOnluZRPt5stXydn5tC6b0myWcymGE94bWT1ZQN25Hf
L2mtBRWwljAigbx46xq02l04ZJINUGS65t7gN9TgvRryauWB4mni1DIybA1t1K/gtqcyJTV5xTOp
vJ3HU1Wd9DEnQegcm9pmZfCjsdyho5/dEu7VEwdZO2wcVpQEsY1jEqxXDmi2OO4dyNZjF9HqRKMi
JSNUocSzZHLNMAjSi0QxXUxvkFqYrjCtQcnCdsDlwoUKNJ5cx2yoParWhOgTdIj6AAXIW3VdHIUg
jkBZ6hYt/G2YHJEqfWZLBKehxW8TO4JqEw158Fih9vn9akwu+j3k/mMLZr6puSjQnOhPtsf0/uNJ
jtqMxDwr4ztRjv1C1GG/j06z1Ge6pF1tvJ8huVxioaX/p3T/BBJ/y8GoVN/mkoFEec7jnImiOav6
fLrDF8BK8UbweBAM3nAaN2Tat7D83YIs67oNsmBsoL3htAAbJJ3dnM0FWF6Q++5N6Hk9xnUbfa0/
Wr2m3NZ7vEjNg6SQBnZYgq5hM/0QRdBYo+t1ehgSzHuz8sP7mDU/xOvTwZU5G809bq5eCC7raau/
oOtfU24pvzrHto8FNvAiWvchVSLH2QPj41ZQkrbVNsngGPvUQaOzyHpfd3JUFkUh7bbW+PAe4fc+
5uiE0SNGCTkuGCDh5rc/n4CzoFJgJC3tL6vU3YqTf1osymqTsBLIJWhDt1zxaybUZO+tWczoKlU4
dr7NcxEQS4ektYc0pEUy6fsFgDpgxX5iqYmYTB+Xj5+ovx7BKi9g4a7gQPUl+g5SY9K8dif55oFz
QKMi5JlIP1ADtMF/P8rI4FtSpvdkSJr4Wfe6lSlRfQ46drK/C1DfoF38y3/JvBTS+yY2DkMC20tm
IJ61BVcZZaBtmWsW9S8lotEJ2qtr2sumRQDPgATQIFvHj0raQJR79iOf0KNN2KbR8abV5E0Te6tC
YC2bvIXAHhGdSb6JGygjWbDPiN/D++aY0ihiS+xjfeL3QVUgcE5viaPGbYjTE6OWaQ0EgA10CQC7
SUb+k2DTkwMLz7JNoyqBWOMpu6Rg716lOE82M+wNK3Ck0RL2WUCqSwW41D0bekcSUk0xq2Yb6+vH
jGC7s94lWOKTjhbw5hopbS9QqO9xjYqBNSMeJclYs41HqhGsZxay5eVDAGjtrQGcoxGva15R95k7
6OhFwQTL0D8KmJQIYtwqkmzEKWy85nc7/SUelH9LDCYWE8SgZGyG4o/iyPIg3EPgMN7Dx7bZtMZ6
268q14IarKhP3p0u2xeXI+47MfkPXHsFYnlk1KLHnivEuQHejuzv/50N/hTvwZ+9qOhCAMTcJGsy
T9lb6oQZlVAwaYYOFafyQ8l4f6q7xj43+qJH24W0ZKyozKhAsMU3bQfGw96JENPsubYj70uBqoQw
JgFMyuyL82PA+7HOkDMl5iVRifK0a/vMnSuhgrW0br75jMpBzdXQKIIQOSyd9yYgVQH31DbJq4Ld
AkUaiO441SHDLzdA8PV+SEm8dh5CbOaFL4hsSNi5JzW/CGnGdjznp6u1TRk1B1Yhzjg7Ki0fAoIi
+SB52WLXD/Dtw3zmUJ+UvBgBvp2JBRBRCl2r36NizQ+Lt8xlRYN73AshGxfClnCP6mS/p7vduu5O
A4IDmGOZ4yaIFhdTLyCWmAWgcvXBOPY/t2evFnYHucWII7aY616hJ3YxdYfqsrSwt8xS+cXWNFaE
RrSCP+uGGU3456gq2oyOQ7b77dPYMAOxMW2CsazMQEdkbbwujWyEubCFWw/jFDA1xJY21ATAu0kS
QEDeGjlN/Ccz+2hehIIlKgqNAc+6RaCefNa3ComiqLXjfsRD//dtNpHK7NHg5pQYIYuOa/Wfl2RY
Tu8BwNw5gu4HZwYKjkM4JpYZiMzyoG/u6MKJjUugMPz4Nfie6ce0wyXFo6cWlHp+4CWmp2GlVSsq
GPj2IFt2baxJlLTUqDyB0IJO0pmC2/OE9Ehqe8KdyFejXL+HFhD7rvqsKQfjtL7IQXOc0m1JiPVM
6H5C+/wva7QvvzrGnmbBMpRqYkIPeP0YS9G++aB5mx+PKqG4MxiqLdBEaCubl6v0M97YCT7QHV7E
i3QnZAc16AD8h/33ahad6k7OVDPyqgnZw/vLVrLdhx+dp5jGi+FENf+98uX7pOkUFKT5oKvs0Ig7
dDA8dyFethSmPK/q2ZP4JV2RRzhudb9+usSJlvOGX4Adh4pv8mLyyO6f2tGiZsTLvFTX7NePRJN2
JlCuKyloEK7xOIFwATG5TuLv2JukQLMQNgQzii+BUzaCUOItAgsLU/MJu5G9PzaTHquyEFSZYgRt
CMjR25Zyf4rea+zR03Ycgf2ywutxZWMIpaeOa9Og6/5dRbz6EF2UPupE6S4GsqWDMjNEeM81BZEq
yA1OzlRffMwYWwhzu+tfTyetUTVYG0/abbf3Hua0zLCLgJEixa8MPM49u+JIm9MHp5nJJU5h4eTm
BuOBzkeW8XOfhi9w/EbCYPrnNWrpXZvWr8UywpPDzWkICh1t8dYlNy53jL8sfn/6vKP+r9UHFs5/
K7krItBf868in1+3KYXdmjsNSNf3Hv4HESlRNiOgXrec8FLzTGIVLjALlkDDKST41OnvPXwGD+38
gzxlD9ynk3szvGAu82+hRFjxMbxd9N5Jkw6hXdOVYWLewQWvmAGlRJkSpuwqdNL+Y6r4w7vq5jNu
e8Ewk7z685eNi7pcplzYYeNDWKG5xMzsIdzjacrlYPJmIAsPgRWmz8onTZ+qE9yhCL8Mrni/qdc5
ECrmD7HA7pq3Sz9/vmPhVSBHBTy4k1RN+dOhhFFdPKed9iF9yiVWQX7jlYvbbvokt88iOSNZm1ok
Y1yOVm9UpEK+laPjYmUk5NZk/yFdQxOHNiinR/zWSLr2nVCS3P6Hqe8hdfr7vxD5lh2gVmoplolm
j7YatOhdCoIgtjzCJLbeu35brEZKZ7BxejnrfVASwJlewFO5M9q8coValLxR8XTuMbQR3l8wFgvO
1jSHH04a+SAHWIr2s94D+040aJBIqSsBRyzbbtLPktvl8eRuqYVuERLB7TYdOywABW5+MAGnaL8v
q31kI85qQzMrPf33rxdNbhe8crNBIhBMiAJbYZ9/nAxSCjrfT/a0MH8Eo+4kZ/eaovPVv9jU/elm
Z8NkscAEtXN81TRiGOnquEftVOqQQ6JgC3LyqyZSSi9exhmTBIENoqGQkCAupO8INKWYmFbD8giW
AOJ4T7ufLsitwSndgxKY/uWBvtkY2HRBEXh4YsV9lcRmLn1Z9V82oeMHX/QrSPl3StvxgieA4OEZ
gBl4PK6v3P/R/h0YCIdiW6BlwA+OobFowtO5TnMqfGTIruqqCZrCXXDFm/GKagXqefn496w0V0lM
+T23gMVuoZ9JZ4kycCp8WWXsYmBfgJ38SsSXwtvQtikp45Hng9UfXMngY/jPmnOGWtcqd6+ZYRFm
RPvseBDz/bkeDhZGD7O8r3BGcaI2yJpPSJrr/ioc9Dlc6XP4D5YKI77MscWKFyoa3IwzjNHFZY4J
EJgZ0pJi6edAc0PpurPmOQg8FPGh1czOPN6kjZ5UhyUONdRN+oiKwlYZ9E9Sn4+W/Cl4aFzj5CFQ
OzjF4oNs1vgFjJ54e3lR7WPbAT778ERmn1QUTsoZtDpsCkmNCGP5Y/DxjM7CpWoOPI++eBUc7hkW
9Dd5H6QHVGRm7uup0IyBfAMUkmRiuGMkH9XdGGEyUqpCZSBnqQB9tvXJQ+WEtp4Y0veggD/lnZAj
aq33HV+nV1vugzGHtmu3LIUUlJ/ia0bmklvzkvWHkOu/UZ+4W/vjg0Rgi6nCizkSWHFHfgo7lPEZ
gidJmQA7lzwo2tjYBH0s9bVOyDQkgahhMnqSGko7bTeQZ9RWvgl0QEPI/z/3Ts+BHkIYukikGEoq
jeRhUP2F7TpoBvUKeJPxWCB+xXQYQzwa0ZR59QzWbOcbXan7GoqZkt1AluUo6LUvKt8TmvmGlaJA
qlKAM45ufWnNRACFTUnhjASqRuVrHPQWkVExRpxiLsbLe9Z4FJiu5n6U1BkalNDDVhLHERWG4Ypy
ZoZtBoiZaO2sozTjOaeeaPz2BRneWA2HYcqP4iw3+/dTVo5KTCWICgs2dTlUoMyEvsOiil98G7wC
kA05Oulka3mrQyxnKIjgoN+uDwGWouH+Vq3GGUOPK/Sq9ZgVGHSv6AZpaLdNxZvGJ9aWvxFx63lF
8mYI2larO2jRdR6mCo4QE9W2SRrfnx+voT1uW+9VRvSSEr43x8AP29ReqyPyqpmXNGAI9jnSQ6Ap
Z/9sHtEcOmjDLzKZCDMp2GebWskYveBzx2QUJEnnVKKglZtSEU7KEcqR8HG4mGkmJPviTUOC5x6z
vOgjnPqIjGSRaLHN+cjdhQEhvEuFRqsoleXOeu3isybOSKWDqtesQOHtdVYtR8lxY9x84jdFRP3C
c85k6dz+55pvCZvCd+H446vT+h1VWrY6ODEQfFNS5d+dT+jfTzy7ouz5mEV9Aun3m5ssd6y2+vzH
3KrKAjUdEtyJGVAmEI5uMyjmHZnLWU35Wniw+TbWK0QaIZWJJpuBMrijurBwGlzsek+rg0BnFezV
3rl2WXK6k2UKWWKoYseUVI+Vl4B1D1tkkRuPnM8/d0cBlYds7yVgVMnWqHwcCthEZ1ayC07uel5k
bmtuXNRbVzMjAh3Utm7cKMv4ywemHsfjEnAS7PfEq+rhfV7veZ22GHGGBd5S9/FXTRFkABcwpcyZ
Pu2F5eEnohMlV393yy/9WDYxLXl7+O7dY4K1Rz3LQsUyS5otKYA0Krnqf+wrtOcgTggmhjnqspbO
y9hKKRJnKS+tQGiHByDzMCP32cWkhCevVJVoOmj8xtBHyqWjDvn55D4t7hO7/hLvnL2SEwsqNoai
SDO/B5ppz0EFAVIiX6cQGcqIHOHpuII1FYYKSDiAt9hvynPAjq9buXtw+6sv3g+EixRfoVg/hPtc
5B/8NAh4E6wAuCCVdG9v+Jy0MLiuzyt6D/3S0olJKEEh9y9b7okS2GhlH8knXMHRG7RwoKBn3VHt
pkMjcmTNFrQ2Wh9E4iObhNtIAyaNNjHrxJxJ/UbgOkJMhy8komS6k/JHx7PwXmSaYePZe3nBkm9w
hKCDtQJr+jOXO1ltScqGMk54lSKk4C/XCHASsAC/GY2NbiVTMEhub+QL9PYBnobM5+2+ccOx7l3v
Dthccw/d7CHkBIkz2r6NFIQuCpdX3Vm0wBTumehA4xKY1C09iZQbVhE4icOqaQ/5KXDzvaYXLgo9
3pPI5ikCAV+E3Da89SAUiRgX0dQdTGLEcRhvgx61SLXxODKLDLlCIoM7yzhOSAvcUbPBflIp97cu
JVWqZUbzDxxTgOGQWzXOZT34r7tOxvRvogUrM/Q5GM6gK6fw0P3+EEvDgSXFu/5CYUi/N177lwvy
UfsYqCHMSKbgoXfOJJ/LPGM1kVq1NCfcv41J0jFk1bP+JoK8yfXlaK7h/cYQeQqVhUA/8bBQOfJc
1EUy5hLKn0JOMNrE8XdFi9GPivjQgkjxh3UL+JO8mhTBexcqXDha82BQWm1EhNSnvIh9zYqMaL3T
I5eJHnaIqU5FUh4e/pmJ+w6mfZPzC83aHaVemhqPfZJuROft1JO5+EifO+ctF3Wew7r41sDvLI21
SyL/Z549+AtVo77sb1279n4KCohhoZUNotp4RBj8t//RITdNcdNAbwXkQBjmcUSJ2wafY0gFX0NX
61FVU2hfIrcCFkGbxawCsJ/A2vWSuAWXwVCfLyevI+RGrU6oA3SH0VPkLbt22To3704BasxtMdxt
L67HhtmfdiDxSIViZAsTAojvizsNCIei1nQ+YZmNc3uXrvjLG0bNn49Vg5qkWGxEzDLX3sLIOiKv
xCrs9WeM8NlJXFJjS0haNHIJ51HqY2SHcmclskF4ZGNkfyZGs4dAX5GpdffuM7EnxzKWUMSDxyPo
kG29ORuKREnp/tgPofZQOWYylSyOQEAUttbooWTIIaSN62c0xFOiXbTA/BuuOo9QXGsJ3vii706p
dtGxRHmsIZTyu4SlHSa0oxF9GPi1pP+Iwlf5d3leXuESSKBj94an38sJykhlGrksZAIrZT64aYSG
97VzCaYHxgAc9d3eTgbMAvSq3HrNxpTB1GzVEkGfzlQGW1hv883/7dQqcqekP6ZI3bAocI9h/0h9
P8oReCLDvahAeaUtGnGIHduGbFSDuBGORRlX8N1Vz6W8U9jZDxicOKZS893ZkUhOQBpWMAuAS+qf
IXzxQUQ5lwUVRsWiONPA3xRXK27UbzAerLdlC2x8NeBX5xcrYCi1ZeQK0OppMC2kY+WLZ1NV7DJy
va9wdC7ak2A9cw8WlKGzNf9UXvtTGkO4yWFL2ybliQXcmTJVjFzkDeKnyumHU5KFcoNcTm7xbct9
hct6VepRn+k9kDm6D+a/MGcrqw8TBC5CS0RTuViZM8r8lLpSyfWvnu09+AduTjbiCSFUu9Kbyvg/
Gct2cCjmBcrcsb7KiXdfe89b/Ij1+yha31T6o48ommKGA1oU9xcKPlMAocDjiQHcuNAs8tFig3Mc
LtFpF7gViG6kSKCRQdAWc2bu/TLiwqbOvHjYLHE325WFrc2nMHBw9Zu5Kiunc8/PMG0lGKC3x92C
sMcmzbsGrowociFxruDS1h+k+QoMmiwsehn2cs3obPL9D3a/wgvKUehbQzZxajvzOJmuY9td3GAi
Xi5ix9FeSfdihXIiZo0gWWhDq220WVbYKguLat6ke5qJyV962KN4dbL2RO83HqBSAN5htf9u2+kb
ll6ip9uhqBnkoBbGhNOVhFZLyp5aROQqV+9yqlCAmxPSsgIybmlFL/RxXpSTpZO4zImi2cp8YMJ6
ly0yAPZB556S+0Oupt0s8NciDf38Wc1Sb/HpGQdlHJLPF+2xlScE5NqnwE/kqKspcoE0Z5XQEJOj
uNDzANLk429SkPECHd4G+RUm+o5tGNTtv4Wi/8R74nsXJhILZ9k8lJ47KiyZUwrMjlFWcP75Wh4h
2uAtEJeK5yD2uTVdmTpBYMAGzuJk0/265sGfGGzQuuZNy6miu1OyswmK6HKIGQgd13AfV95PStvU
oU6w0cXDLtBwELHARyKSvHE7mDEAKshLwOQJZ8RMYVCYbaGhVjCt3K1MBuW8dfVXo3NC8r9B4KJR
uw2Tdd7OH4cEIoOeC0xU37aHheEgedgz8blXiAR5TUNOtk+i2g3IwBRBAH4fO1mlrSZPrObecuwN
VYmjcIdaWJp7txDsqI5R9lRZSHmmt4WfEQ30tIpiSQRi0D7wQ5Ql8y3Al+SyWGBRWIg/uVg2/WGJ
CPEy/gvNXA1uoke3418piHSOhJjKRkq67EfQkvO0jCZUoWlKo9dyHEdN9ZPV6+qjdhJ+AhAxJqI7
g0j9Zrzy5+hPHEKCKqwoGTSB8/Y6v+7tgstSX35DPDE4S2z/biMTJ8Y3taLfGlxcHifD40N1t6q1
Wy9oKgO78ShiAK0ZAXexHbCtUq+y7i5V+7BMjijx4x7Tr1zIWtTn7kpAO2N/+CFZ7DEEvjrCIH0R
SpcLydTB4wCXKuuizG2BGAF7AnMdSAF5d5/vtydYtOcIwbKt1/v/R/xTb0oAamBrfgzKeecaAXwT
7eE6mljsRo6F1EYFnZ9pLRZD73/0W/FWN5SXOdVssORrt8XEv8qvGIkAHuFHYK/VSt6iSnW6SW+d
Os/5yJDVwWbmCNAS/6SHpPZEGlddT0M1Y+lLUu791wG9ivGldofSHkFuPjgxltkRjz10oI0HNyNX
t/iShBIbkLhJ5VVCLLP/D/j3PhxcotdGtL7Kl1uZP5k5Ed/yfSAMfxO+qEWMjGSKhCwqV9x1g9ki
KuCwGkAPliDJ1pQObq/DvjU33yO78lzgczVYW7/HhSeqWh+1OU4lwDVpt92fbAtEOvA5Oho4zEOu
zBpu23SM/jwKUkr/bZee0LA9zJI9VPvPU9t8cHv5mYzXQZUvB8LIu3YYDJgCd9yXNOtkeht07aeI
rQtjbeMRaXQbSO4gcu7vyvb+5Ru8RvJFeXrQW957dPqu+n+MRi5wW7Ngyvcal0pShsmkwuDh7Ync
5LVRhgXSIMLY28/r1OhLxCby2KpYG9tvbJhVicF1/z+DLtbavG5lNIGdfqWcQCLWIOrNQ/z5SbTd
CwOKxQWqZDI1sPpeVaP3PnF7ieUNFAX9GI286BfCRAG6AUdHf7ADghjdx5QKIvmeZcb5IM8x1eh1
hSLHZ/pEskFg7u/f6JSrur8NqFbGFuHwLzWcZHjnAQkJ0XOGOq3Xj15iozC0Kp8igMedJ/yu2KiO
Yut2DFaFfPowJapVlJqx2E/xzjxMu07J4Gr/lAQFXILNoPYBZE29PkAehhXO97Qb553ztPt5rn6G
HIw8OHdNtD1DrYQeBmjIWinqfkIyQ+ClyhK/wiBZB901DFPOHvhv0SA6JkHpIIxac0eH7Q9YhgpE
SpUCckNvDxUMHfdAwKvUoT8QJGfeRtWPtZdlDPqeBpiQl3qWJqUL9GO/h2Jhw1wev/9RUX/REOrn
G2CGiqBsXHY87tLQZge/sxFxQakmfDkS1fTuav+ZVwEN2wqRdEFwvplZ1QP5gEi+4MmECbPPDwXp
77UhTLKS0QJ0GJybSk7/DOjGD3Ef158j2fCVPWFaFkm/6Is0f1d9KPdYmiMiaWKlFMD5hHzvNIrx
UQsZv7T3iNPwcU5WqbGdZftFJ4YaM1pOBQ6ECEzFgOIwtVYNJEGhvysretnBpnjcyjftDdkrA0pI
5b4m/BOUO6wASFrM8IAjju9tFYmy8SUaxlUgltSOETWRZjHFuLoJ+YiOshAqVwX8c5s/dHLkMyXg
af5/3KMvoZEIOWtbZZQu3lzK6fnpUXe9+M/xAUTAEIj2IPg3JIgs8BUK9C7zXu0x/iEOMz/PHeru
ymRUMtJtCJsOE78BnCwX+RFds4OIb9YuuhRXF7zQFUfM32d+psDLcVtkGArJtRX17t+Ov4a9fGxi
XrKgvdBLclAK0OdNJja52LhaWPy32rJcM+hSQnsXeVRvMZFWPoop8CEBF37ajLcL6a8WMCwCZQoT
I1JYYxpAURbKloABeYDt23g0/lsbPOvJiH5ZVgWZQRh/wJ2eJcAbD8VQPzyPOlWwl4AUcS8yyV0U
E5Y6G15gJ4P4xT9MWWvmczzoLwlCvYDPKJG3K0ptvZplgjrXVB6r9U5BRO517R/bBJ9C0Eio/8j1
RlZI33ZtaSIVZRNDVKevOLQKV2YauS/XUj+iKQ8mCwaHCxwLPw2WTX+mm7NI4NcoH1GAj5zcF19l
9APYI8mZpYicVH1Y9CKkNTgdlg2HsEdt5HuwCDV37j7FqbcCOf9auXsTpOiFROC42VtHM2AZffZ1
8NbIwbiqh7DV+1a5H3qJTCbVjcRQ4BI+OClBPgeKPqjUe8Fpt3YP7isNgft4kFPihXsxmcrWSAns
hpXWbsYeYdBHIMI//RzYwOUlxM/g4kxAgt5FANAV146i300ohyzb/lrcvEUw7Uz/1SsszmgzexhC
U6Isdl5nsTRthCtO+mo8Hjnt/Y6CyMzFztgPHZHUQ4tYekpWM6yPzBpVQr68qJQU9uda4jKhE2jO
m4Vz+Zlivz6yjUJr5+CcIy03OzqyWPDGPhhUiPd8ZANGQ04kp4/q2jnzEu1G4y7YkvCQdQS/C6Rw
/QtI8ul0TDfy0zpkCeF9Y0ra+fxuTKuaN00MUdTqr/kn5rQ8I86yOqtkARuIi2LxBUFGNpqu6cAp
puKIYQvgmrdhIr163YgmJzq1fxhjf5BokGUF5wNwrLRqr/bFHMGkSYfOvMG9Xl+BkaCcFhV3tDli
F11/LpK4IoLXJN/NbS+J9vOQMQT/V/5LyDJAeFaAHybWpmbzGbA01ysN0vONcfiDR0Ngngi5pwl9
a0/Bq9lY4MsMaVh/Mxz0dQVnvHrranCqMyxQJ+1fIJvzvpmLnh1wnqrF+vilDyIdbjZ7azNFTqL1
hjGCW2rMoyISJLz1ZgAk6/Z3Js/INSP2JVnTOckNw1TWUHKXEP+ltf9yfrl/cikJK+bg+6qYGTAR
gGfVndKKFzuG3j9uppYBmwoM/fw998zrxIRm4eP466o9BwdMCQ8WD9bkqn6kMGWo0HF9Cfn5uNDw
/mAtcaMSGXdYH49Xyk1IkOC0ofl33ame1D3/ZGCQdnp/fu5EO+AKMguGGduGVycsY4yZfJViOndK
XrjZ4bJOYeCYG2KtUI6xhTrXCMMLakAdT8V71XBwkeeoF4IbkgyQZ4FFc0I+xi9d2hxn+UeYwsnQ
vum208OPAgojwT+n9kfOkxfSiyO8DnzIladCvctQaIjriNUyQkX8RUbBYvO0AMxFIbcEtnLhl54J
H1QsnyZjXxKoCNgoI8kF0M67RkXexZ3OU1fylfE0nsYJUPe18WK8J6fOrhEikmdpP8/lTKznJJLC
SCvIOKqn8Qh5DcHeAyQg6Cl9Fsi5AXaBQ0FHHbzXJuY4YyU4H0caDUJVeeH0EW7gqyv8a8bl7kfb
d0laKUZ8Y6bpa1YJ60OHxNJ9iTusD6cJgOWDpI6/j9nPq/WmRZqV7mfSLWiDzzc2Kl160bSaMfGK
zUOikrmxmrMOcd2W5q1GHwVtV4xhoYC+Tihihl6Z5aORKb5xpZmMxyCFyFQfLpiIlknhWfg2mim8
sJ16bAFDSNlC4BLRDt6zVWfh2xFsmboYv63COZWodznWjfN4u/ctsGScahA7T06XblMqE/Ir6y2F
v/5qP7r6Cw7B/jCDW2dThvYmezGhVqqtJPekWfi9uMiESCdHCSnGJLv0UIS23MUg6u2ENFzjIvC0
SP/vkxYANaUDr18mXaba8S2bUnpaRHNxlntIb304gE8HxF4gNQTrVAeHRkWLp9kveMD6E7UucRfM
UfjS0iiwBWI0Ez2T7/7mfzxRYEk96be/ce1P6ifCAB0hF0bkFKvQDsBQt8EkMuxvkG+AdQgd/rCP
oTGsb9a5rHznlfY4wrxVmuxcROdVk0wb0apM/rv8nDI0r8kjTNDOIF5hqIMZWuikDCpsr9LDzuCe
2wQUSc8dgHFLKxkYd6QDWZ9D8TOzIU++UhqM8FlWbNrxf2dUnjue7B1/yTULjWbF0NPla5z0+Zci
+w6tvREOpEc9be712gNxLulg9bNm3BWxHvihU9+OYb5MLh+Tj8cJZdyRWyxOIGMtr26C1HTeqZMc
+FzsPPSc16xSYTd1Zf05Z2zqcMyGju+n4rZ46a9SCaw+s2QDq5oaSEMQaZXWGLilUDM4rhnMp4K2
YxyX+r6EGTiT5wx8E6KNhkiSidJRXVfL5wXB0FBAGsiQwDIO3lXa1rPOuZRYqL2LZ2D//6JJ67jC
zUjyEvMy/VqphrYmJdsGPVThbluNKJ7LgXoV/SQecvkSc9NGaJufROxczi7knYiN9vN5a+zZkHOw
sURgGJ9lYAXHMj7WPXd3Yyczzg1TePP/0aF+wVfrZljq2x7L2k3HSfBtbTgvuTEUHtf53FxGUTG9
b1crxmOQAY4BcQZ7ibFP1Y6d1ZGKLUPY7i/GAUhQXGlCtJ7duxAOeOK20Eeehto8QEYv2swFnsPZ
Emr088lcxNbkwepQovAh0BhHwAil82pkyc+E/b2opVpBx0gKC5PzgTtC+nV4Sk4MBgY8AszbiPOi
KjhUbLfvkViJPph9qOy6VDEr4vmKMXJ5yiBCkFKAX0j5POc27A4nTpkDSpsl83EgWNM1F1SLhfbY
NybXfOyTF41O58nZ5gtACMUgDeZ+Mk3j7kK+vX6ugkPwMrgCTTho056bFoi6KX6lbgUyjW8h+GRJ
UMTSSuobliZyJRY6Rrl/vqAlHm8+DbdappS/TmT7zdyK20vXcExWhRB8aXzcGEdGjzAoWIYyazCk
KrFpH4/+MYOeMmSp3ulm3Bk9w1A5cxN+/il0CGwYJMqiIZk0OMyoqHSt8ac+2kfqqa/MA23LEALY
JoLhSmib5n8kT2wntnpgLHC7Xb4/vM2ZVtCPGyXd7IWqmtVdmy16iLex9cCFNJGuaKDIgUdpQYqP
aPiYBuARJ86vLWBuVlKv1MIZuvzc+F1Qw66vTvPrs5DAu/sY0FNKaPPGuISeFx7ybi4NpROXwU6f
8ThWnKOuM5m8EAS2Vtlv7VWS7zgC+EV58tkQA5vIv/KTLR7vRssMKYIkNVq0Oq52+UAkQbhIa2Wg
3bkpQ9nzzhzpA5OPQtq2+1Alt6s3+8d4oAmF2oSEy8FgNaJb0JR/NSFEODJWydD3afdToq1nJ4L2
wFI2yNIkPWbBh89jNHwCSSWHLn6tBH2u94SFFOzbkXCxCyByq9QMftv9pvtbphDU0ABumJlHD95g
CIRHhK5rKitKwLKVR59soCwO04kwM1Yr8QCaf6k79xHEdYdixWB+WIsHmp8FIqb53WKcMznd9LEZ
NQqiuRlZCv6Gaju9Ui/r8MHisc9aWji1DFPKkbf0nffyyUtEUyCyd+xrJSpZf/H7lH9BZWjlX4HV
meC7R5T4fM6sR7MCvC04/VH7PPE4l5cYtAGCIrWtx96QKGeAud4fUm3Mad3IoK1ySJduWYOXHHJe
8a2tR//+BAy7RCHVhmKu3iDEMi1WDU4fA1n11zfb7Y3AP10UEreoJWik6ypjAzayNzOBCu8bmQoq
GMGab2QF8mSfyAhRYMehDNCzaRHvHOHdRJewDdVCToCb1kAto5wB8jBkfLgjbESuRjt1+9u39CzU
EXIeSVZUtBnBNZO9hO4wfLCZjnJg9haKnYeFrUttwegHTyZaS81pNP/ZjCYGCKNB5u1dL4YWrYnB
X2Q9Qse5gOhkew/EU3vnb7fvnUuT6TRLlhIga548vvqMQB7mhQgsMhhfBIdEP6cLxgeidWIaN7zk
T8hJXrl3zXonpyMlD1GqeTlN0aOFr+IhC9N9j43GALG349ebtMuQi9GN8EVic1zpaqsi17PcMRMO
Wbnl2SRvPEuTXnt9+XGY2BTg+LaFgRkz26BNkPQkjTxwV2BDJ3IgCmmxbPcmrYSjxNPVpACgbxjy
jVv1JLZIP1RTJYylnP+3BVwlOg79zVd6yqAKgHPmXEJoEG77bgYHfyuWAqFwpUyUh+U3lx49kXpW
dJwKPw6uStAA6Lgy37AVN6sdtN7HJ5e4gtAQK/PVEU2C6ZPjPbPb4ZAj+fQtCyIZx03RX51xg5Jh
O9ciUtRca6ARujs9Ntls2ptM2jz163q8xcc5PG1xJ7+3Z7FCzHQ4x4Jz5IVWAV7lElFoSv3SGLbs
b+MBZHDNOFHWfmEURY020msX60N/tG23YwaoxvKKMtkk/SvHLQ9bSsMwXHtSsjR1sp++By5mwFL1
sF8UIV0Qkb7TfYEwRk8dotwXaBON9Ww2wMR7O0u6zhQee5+teAHAhYaojCFxK6o9S+/0h/7cVlb0
22jSm9SnXHrNTnlTE4RGlxmS1ZIONJeC+VtWWgBeu9stKES8aCzS8z+ib/w0jFuykLGtOtW0C/sj
Jlqc2Y9l1XMILPcOQ4iLOdR2qs+ro1lTJVpGLOa6aPXo3BOdt8KaSzDwr6Yy8oUaRKQDzg6DeXlz
t/VIZtwNPDXYqTaqtGU/jWttlPrpTBko53Gnc2qW0Sl6DrSwU5R314cHCM4NjRyIEh9nbbwHN6cQ
KF+itFjsLyy2qhnKy0kzIfIfXrpCR/ee0VYTbxGu72xRnSGmlAxTmX9NR22f59nghalpR38vXLnj
OCkrTfy8vH7tAzI122VT9a1tWWXhRmmCm5MnOQcQwzONZP13D67ei44QJ9uUoy8CJZNtWBvnAk6s
8/VHQf447Y55v9RiypS9gB+duwYQy1lpAzfSwTGTdKAPtvCRS+HGgagvJFPyoclME+alkUrwlQn8
DnmTgJxzWSfRzDpZaUgqUe4T4FrZhVlYXcx+PDWznHSD7X8qYEErpHReq0GihyUv+tz9GbysppWX
uhWH+94FHIQnNFOFdHX0KBQOx9F9i1VlR353HTxUMhBSKK96sN5ovINlPGQGHQy3TqPiLQJJJIWx
HhojmLUuHeA4dheEAUuZ2/ez4A6htbLXcaPswTbXERrBePfmKPImVDfdWXgsa8hvlbcbtUUZ666o
YV7i9Ou/LXryQ2jAseSny59EWNoh+vQ2KC+rRn+0Zjt4Hih/fzccVINTzM2DrYMQTQJhZdeV2Zyk
j37PQs+RZfCkPDFt3JJWHQqe5BZeKJn2z8b+sg9S+PaO+7BLCcAIUtdPNEeFsynPDJAR/IjbN0dc
JDtljKF2P7HvGBOVJMPnVqd4OchCfeudsF3jCQh1Lqj+Z3+RetqsvhyKP6SKbINH5V80u/xpIQfh
ng0fHjTM/C1BsTRTtDZLUdyAKg8sZlgFq3/QFVSExlp+QUiyrUqBASkLJYwUB2XHi0BmdRB7z8F/
NUVqkkh1mFonTEDY02DUcb0cVl2ae8dlyPU8P+J2SKrLC1pz8yXOjOo4HUyGgEVrq+4ro7674445
LDEBPy93q/L0mltOsQM230ENUZIj/uPICgsED6dnF39QNgvY5cyS0YXLKnqKg9Sk5yaTj8zfdgHd
wa4Xdh8iezLJkeVE1AKjtnttoNdRU+T1r1xcjxetCRnVwgfevvmj7A/a8P6cZ/QEHAx5cIpfDQgl
vBZPXb2JNFPjr/NGwgBPdUeah1BBXG2gnloq98IcNPvMybAKNHrC1SFFd3txC9ArPKaNc1MJ95Wo
h5YGm8m6bL/uzmzmHBfnibNb9R/qhJhc4D/RZy7mvTs0F8+LSOwqHu5GJMNpipS2Gmrtu4T1OXOo
Q3RhWM0ocaKWQFnXqzU+ymLkT4fSsGutAfwn2oD1ENsrPIVaErLnpe6I9WzwzJKKHE1V+yYdfdvB
AFk1REqcVLcHgBGR1ccmEsYoBBoMSQDLsAsf47hwrxGLCBo97UUyOCxPt5awpqq5PfXeH4VIG+ic
DiSU3HrHlUrPUWlms/xKzEmAHBdKGaUOct5tHLDwfz5gzDw8S4nKBeS9sMIz+s2FAigU/uuTNnKW
0vl6PyLYiT5JOJEQMrzdK48hPz4Z3jMgWjK3G7kTHWKLdFTOSX5nOCJUKDvbMXxY+eeGfL1dTdhm
iCjFknlQw8o8BZrbIsUGEdS6EzbBO6wP8CoJZOLHccArTuadeqW8NjU6Wq9WvMFik6gHlpvtnLc6
0F/7L2Moo8HHXyir0xmhf56YdLyVF0jmjW0MFmKBwpA1WTiQql+ztc/1vgDQi699gfQE5HU7WU+l
bUbfmY+/gyKPD3f8ifoCMDHGz+qvCItZfeIB0NPHOU4YncGtqlabeS1XjIP8ICwVlvaTnS/bLWNg
Vj96Ts9agArce+kspzdueh2VCbVkAA0oo2yKsNCvXPcnbJuKUY9F8B/XhJTTZ6toNdNc3G075zyX
iPKy3pyRVZuj2qKnEW+QHRLiWwbwwfdSKWdAHkdGi/nujFmY5YL1Ay7PgXL1EVAaTfM0XeZpO0tw
AZjywGKjlF7erBET5lIO2C4MskYZuVDdg8TJIlFkgyJEEeDRC5egd1tXI8ug4QAwulpm7PGUe/vr
Q6Bl8xh1wbblAdh6Wps8j1Hge7u9541A1SigjjrzUqVdBo1tXRDxVq+mjq2O75KkyWPh30AgkNxj
Y8xazxj+ddCFA+kvBIaJeWdMIZ0CPmdUezaH8EofNw4JXidiy1GpFz8jaMyorfnYq5cagAdkC9UV
+PYPCU6ZmkSkcy47//RdWKCWeTm3jVNeSEsoG0HH9VDScUyZztcBTZXnvhK9qGMgWldBg1tQl/5X
2pnPyem2uopOXNLrlCXi7rFKGzRhAYZATAlgFd2RcunZ4ljdQXXlhd3QHFyhWw+EPfldZbwjP6qp
wkoMqB0UstOmLk2TALW30yvZGg+Xwp1aPlhpMBWc4MEdgr0jB1N7pSESH/ckKUuJcFJES7Xar1nx
afyjuJRS+S4j8KwUN1pqfAxGHwxh4Y+H35bKHIHtcFXFSf0Dzf+tXYdJw//62SNc9z/yhaMLTgdx
QXm9aozcmqk8RD0SFAmISK4d8G7SBxxnOWSus6YDkPS+ZjAa6/wYGM1vvBLWdVQacgL0fi6pjQ9X
IPZzkr2NpTIMQd0A2pgvv2RO7gfqNMp9NEXhQX3Rdy1Mdox0sUfhedMSiuDWRH8LPVvIcKfy/DLY
1FYfttbDw/Y/53O9OSmHq9XN+KLJg0ObWKPoslf5v9Atyy0+LjqsCq1na3b4zXyVmTv3M1AZoR0W
FZtTulRANqmPY0dJnUAz0dMo1zbGKnI1GsEjdnBHDPk2huQ/uDof2P7r39q5UKUrSodXnvM8rhJ7
lgp3jqXmQ9OBOCrZ+nOZSm4Zq/HChAQXoYwmeHkCmRhMCLo89mRRfEhwKHqvoqpVg3+wG0LOOu2t
/MddaG1JPwy8ziWffYGjHIo2RTEed7OekSYckWx3YKd3u4VO4p10B7k3rDPaVh2b9IUlpjq5qhg+
oweI30t/QoPM3CVg/XfrhwHeoNdvseIao0f570ZR3mP2faJIx2Rhwqt8zG5Ru8t/Z1hkBgXvj+oh
kkw6irG246z6qJ5pmhcYbgYMQpsL1p84HnOLkIzz/xXLzOGFAfGsBehihp3czBSSrPPOOapNqYXR
B9XvFdM74oXZZ8ff0PlAkwQ3UvOga3bGANUi3BGapWcqrDUDpBnCRQSJCQ1gapsJxN8AyDU6Oyf/
rtpL7g92AfgFK+jFmAipgWVXOLP94U8Dkb//rf9SLCbY8ETSuk6I24HNO51OQLdsO4sRXOSlyfBr
UO08LUoIIMQ82mdD/bmoDnUDFgBcPFhC6PftafyeLuQXQ0Apo99E2KibmlQef1wZL6bAc7a/rfgW
9gB8vyOc4kD3OmRFGSE6RcwwGTfmFE2Pthn8bfQs13bYTaLTGsRW8slFKk/A+ScfhIDNawc0bldd
ATpkN4Kld7pyzRlHXWVaTdJdhupnOPWK2dNeYjUisIVHYPWeRzbqi6mHpO1mtmI4PXZBhmvIm1ZF
mJowVFvk2zxzHemswXwkwZ3wumd3UZBt/AWR3YYJazYltfFOqPHbv7ORYCjlhXst2233i4STZE7W
KrX0kwtVSZEdiGlGAUIpLbM30Q5uW2um6qoTWZkT6qSMFyok7xdBn/uONVJT3PX/fXed4FylOe5k
00w8MJ4aCwR8Hw2FBWPHkLDU0tN/TPJlgog1rGY2B8bywzyZzLwzhjjUPWEpNt0ZI4yNgvfJCF/D
OZ/NvBYWe0Su+RjMzj8awak5H1yPW/p7LBAS3vIieOcn4+jNAf/oTdROf2DryGHU9UN1VtqvvWVe
NarV+kukK8fSud3j2afuhRSaQEcQifiK2pIoG5tWq3R4QuDkmclxYwA6i5gU3XUS5K5GFmECQEzP
tY3FZ3KPQjdYdWY8ThbJqshGxi9cQ8g95Lx5XVGSZXyYa/rICGo+TIYYYZWm7nturna+8y7AB6Bg
XVQNzpvtl/lRKj/jYFOr+roe4FV1FPFIKHQnTB12QXYP15OwMC+eceQAKA6LfF4zauA0e6lONkie
su/jyx9tmmcQsONbhd+5mU2u7wyq3ILaXt6KzZ16YrfLrn5fzzeaIIl2P6mfRDdoqFsX1HHUr0Bp
0vIbgxeMWP8wakbIYL82aw59frxoWfj+ANFTeIF38gXga+05I7VAw5m8mGREvUaOnHuRBmUpSLgB
R3Magk/ZMWPtLr/6m98y8ffpNmnk5TojoU6Z5kKwqgl1Lh2PJI56A7qmArvyxPQqst3kk1jDQLxw
s8bP5z4mNlowTCXFfpbZmp076qpc7iuykDfBke8w/sOG0NTcwZ0GpliRdUgpqdonj8TIvpZmKqUp
a2wEZTPH3Hj/CgBhtOY+NHG5t7kIzhmsjV7CjOduLyQW/aCA+LHFQ1qHhtqRLRofizFw727gm8EW
r1a/biGx1mOOCFD8QcC+eWaARjRZPEh9wghmvcrswP22/4rgPoHBBGkTtx1/hzOrRdRE/4hPO33v
sSGnGfVR/31aY5W0wXqs44zwP0TnjMxC9taXO9CrEg1jj5NX5nVsyjesUYgNaIHIDIi3DfP2uJ/l
q/7m4MLsDBgrQ/IijqeMbnOkrNVRMWgVzpqSECZylDpdajal/FAU1GR944MALIBMT/Qx0Io/1zaJ
iQJ9e98GGQ3F9Iw6KDmhgnJP+++EBU+eTx6hFVOvpcIh49M4nbRTZXIAfDdFoOEMiVlgRChfllMr
MYWdGk3Qsx0k2ttVv63gSClLPDHjbPuP+Ae+LFtTmdw3bMRm3yT9y/l2tKSmIMuz7qWtjOTbqqFP
iNfSkdhn+e9Z1UqxMUH/C741yaU/m6fPX75V7ZqzCnxQ4R0MLeLw1FWUfSr5OKLPzW6HnYaMYwhf
797bEi/sw92GCNinGF8FFptWhPWoiPIge51zYd2m0Zxxgd56VMyaWCs6AAWeO5vwOLp9DAzaL1+L
ImfiQmSE/E9dz67XZzLtTkf4GvuPDrG0QssrcCMsz+kT/JB/S937c20O9sauCvSRY+s1SHR7qwH9
36xRClUsNekXH3BkrtH3/dokFUQQsQGow3Oro2u5oX7moOPDNLUo8gX3U8FJlbmGfkAJFyCVXtbz
eCQ9+0m5SCCUmcpa3hfHjjS70XlLMultn9MYJNksXeD0GKmQm6L3G8dVBlfhSwyZyMjcbnZE/pjM
8k3QhWDbsHvgaNA+603VKFoPuh/Ym1qpVzoeVo3DK39LxiE0yH4jiclQNLzBnpvz9ne9Tkowehv9
8dxhiit74ZA/1x33/Vl1cs79TJPxqfYwNtACV2iDjIhZ5IqVmBVu8xCLPjQOptYtc16GBfGXLqkx
pzTWVFBcYjFLVFm1fTG6k+4qcAOkZ719oni0Y/nTxp2k6vmDxBQX4TeLM6vMKnViB7bnGLKLRMN9
tA9JH1gcWmbNqNoc3/s992QwpksNkdMcCf4ruK+bhPNMJv0MrPCEn+IqvmqnBMdPWvGD0pyJJ+XC
gtJlomvvlUrWoG/Lj6ga3uBN/QrbhVd3+vdpvEZEhCiLxTLJ3MRLwmWhudxIi8Sks3ch3HGZh6kw
m/oFbIAQsWvfLJuKoRtMuCcPODCldTdB0dvXnnJ7ix3gStPGdEj9K4PTIBkQY0OhYsMFOU8uzIxC
VQZEANCMVXv7rjUigSQWL0j+09xiDg5MC4bzRYfAdLRfIDDR62nEewMxlzg5ocK0gxa7nsPVr9hA
pFQmgogqiZbNk5YGHDWYOPJjexyo8Jr4OkySMCeQ7hedh75AbhWXzpDq4oDCfJk10lXKi/Aa22nO
NI6yJy1o9avh3H7HqkoJXXOIIEdj+mt9cZSX+MWbdzFcE2j5cXZmSg19CNg42DW1stV4/veISsv+
HFR6KuUfaSgdeQKbJ6QgqkYZpaRFovkLtgEmv2uSeKR+JjtWoYM4dH/5wYhfvRq52Qhfu1p1X4RG
h7njMFecvWgUc5gu9IwijYfyA+lew956WMFuj1nPIbXmb4eIbQYerML4pne9HfoX/aSdd6UAirmG
rBV6d7xqiGN6uD3fvxMGBDq105r//bcnfms3N1NAa7CnHk46LukL+7w5LxughtmKCgL7BuvTZaPe
2zknCBA1LPFJ9T85Lfehin9sxMNmxMjMCd7KO7AP6JXNfeTu/aAWzf9KFIkD57D9QI3eXjfr06p6
kruU7R+5GvxQVKhUFpMSNzHuEDbyOifsgZeieynrdGHzdacWhsDpL5NDTbXxDDGY/zUWj+/mOeJy
AAXUn7HvlBgDUmwztAX1KqvmX4jm4OSl4WyeDQAcHGXG+btVCdsaagRx8muSz9KItGN4TnLfdht4
6P12VbEz2B8JRdz/kRx+1U2gI4T7ORbYEkJwQ+VqMSVqJaRZmg9aIFMKJWB/6hF+/RxXMV30vqVB
nthRf0Io9FQUkbpY1p4QEM1oYoKZKgCcW4HONmiAKlNhWCbMMyJn/ScjYBSLQqcBGKlmqCqF14k3
E6V2yhObgZtAlOhXjCUFz2QUbBu8jW3VMWZvggO+gxg+9AwHLCfMZY5cosINO4chcJKFU9k8b0k7
mvlsbPPYnvB3/xYuaX13T5jrmdVWGsr91Gu4clcG34hErqtWpRSs7FYK1IzY8I2m3hv9hLJWZQRv
0/cgul1f1MhEcQUBe5Y8qCSTRI2UbvL2k34QQWsQrdd9inypDJTDBxrNvA1Fk3irXna0Cj/CMpJM
mmzHpsqPHhhC3jIV4sm/GN5Ens5zcNGuINx/3Wxk9xojt/7hsbXed29urGo6+W0bdjUs5xoIupPg
vSHMEoGuqoY82Y86ieFi7+M7bxu6u8lpSD8cD6bskTweLDj8j0GpwicgM+M4pI92e4RkFhv7Ccib
ebG6vQokf/7fTjd+CgCSvcu2nhcped0Wd3zUfV4dX27hx/bkRJ3xXI4d8VPWnVpFkEEOBpyRGvm0
dz5p942scAdtoQ1KlrHBiGm/m0Xz2KWUpNfwiBCvzt+C9uw1sUDw3O4Ukc2dV3my6Y1HiTRx3tof
4ZnF9zgGeIP5f3Sf1qtUKG5CrFxtIclWlmDTGXqTzh0Jp7dwEJJs0qIxVFd/bzaX4Ri0SsCMNvJu
N0F63krTRaFIdo2TpwIPrWrEMLdMicBWEtJSEX22jQlnB+fUrr4dmCuXfgow7L9O7LP7lKcbvRPA
VFovyHccTx1CMv5satyx2taxiy4A3uV+hpCIZfkq3WS7zx2++Bv3bjeC97rXyy45Z9mHPyneFNot
wVCxIHLopuw6ab/vxTFAu6vsqIsAYFTuL6m698TogjSqEaYq7ykX3oc/mIQCShxZnLIpvq9yUXfK
7EKC8VktCHLu4yoTaFwO7hDWasCGeNVNNnkpAwKFafO9fKCAZ9/Gp5ZVQrrcIoyIOPQoOJJFzAnk
FuegWEExp8qaQPe9Xi2TVPm+sGSVy0A19Fi0OfxiqHreUhPtEFLLCF+GKTRQAH25LeVSpq9PJXbR
U+m/ev9DDuTpGsz4opVeAcj6OaZsrqwccqI1qVmP02Gp7NzXX6qWV6Ay8Ykg1aQFPwKIvKlZzk/g
fVsxt0EqBFMiP/2FIACQCEdp93nXnkcKKyyNR1Yop1kDhQpwRa7kcehVbw+z6UMR4C8ImWzdPcUC
ox9VopmPCwdS/fZ0NXDsl0y1jdXJ+c417JU1uWyOpFpcEdreK1nFcvSu5sbAoXith9+8C+wGhXGk
6JXlrQ1eN3BEU9ZE9CNs14ZI7qTX3CosB5uYPlmSx4IaST6KuAEIDxMTuJs0B+B3FGIYdrh5yomx
2APLhmoXtMqilqmNlqtpFMQFmxdkP0vUTQZmYRuGRoSSmRtHWkKa+PLfPYxvuHTlECX9c+bh0Qgc
1O34xwUyEbcKov7dlWIrInbByXLR+4V+PEePEOec/7/nWZP154gbnRXZG9/XAT5sNw21nqVzivSF
ibYnlcm1pz/is6rqlPDsse3J5gG0+XoK4/myuoPC7hOtgLTKpmz8YDfaoPbOdssgiE1NUZZrinEe
FfizIhU1ufOfajRznUgkLkUOtfIv5VeRQXbt6csWLfrOBycjRM8AKhAumA7Hea6i+Gs7V5FqGKV9
RyJ/jm+xccIO81fuESQh0Vp98668BjtZ/r/DsxOCtUzZ/0aSmpMAwsj29wKAadq4PLR2Vk6dwpIy
inNdT2UsNYGQbdkrlaTqvqiXbgA77GLFp/2D9i8sUqmKCChq3fQhESiCsts8MeneyVaC4iiWDILp
/FlJi4r0hlksSCn1Y3BZdDvUbJufbkFEoUvwGYWzJsZOjH3zUN8tXrSBYoflt0ydSkj+mdkJplIl
Hf89/mAb3QHM/oXZ1LsG5z9Qns1WCrsZLYbMWQKt789QO6G5JONQ0+wPvHRZi8mfKQ9E8jFCOw9a
PVFp8UvN/1vPEMpjZxmfMixk7C2yuYwHDNSyESOSTP6z0e6MwKPC4R2kXqDo1ZCpIJSDa/LdIaQB
H1VxHAlyVLJHS/E58k/eCwBcMPGhvciOVsWS4Stntf5QjcVgF5iyx96kdooVoms16OvRpotA5NHg
X/ht4Byv75/d+c8D7w5o/LD3ZtaNV3S6YBaFlGbcNYlRAsaLTOcbowdpWcWyB5xd5+zyi8/yDHHt
ppG62YRmlwA3BX8wZ07U6ueI4GoTKlO0tSPBF343s3ZykMihdt/48SI3jY75/SJDMZJnHKHYoO2+
FqIlFemoDajVvUr6P7QS8LD/hEj8H/KDXsBdIovU2TxBHs/ReSatWNR/MSvGY1S0p65gRLxZ+yfl
uDboc+1vg3AueyUASL8VXbarp0UCnAT5zSVzyLhNTB+8Wa4jVI35uoTrFRsIcWrDKH/KFYU3eUc6
kAXxqvLs90zVwn01UNsPJLHqjFemJKNajnRmykRRxvrRRI7iAhpeDK7QFeC4ZQHI7YTKeHOCzy/p
5hdfhmM0++yIuIqxN+hixFYNFXJAM7JnhOjHVdLeHZPimfhqrKR/4aG6kMcKiWg5qEcRaDQeEhXc
48VEihSku363XlNyrQ/je3iqdt4BYHTPbEweuKO5ClTJDWf/MhmoJetQCpmuXX1Vip2kTJi5PEYu
saOQ0re6/YkwZwL98gAd2rE6wh1jWF09eAyH6YDVtArO5UsyJD4Abj1HSO6W0cdgpMqtJHHWIMCN
s5SmqHk2GnVB7jyMkbGgMjr4tx7/LJW+vgQf7s8/OxKUoBlFe3dXw0hAyeuXt26zjPssyJQ+WnM4
IYILuH0Rfy3xfGe1Avsels8UpsXcdx0ju7UtvvQ0RLM7Ozc+i+grqK2FCGh260wvDYBSvpKJ6wfF
VAiE8ltkSeFQnz8u3Kk1/jpC1tpKGbh36JROsdHeRUd0091PKGIRjk5IRGWHZq0hNyGgi+itLST0
B6ukmKfG1b1W6GnrNjXNNkPA0NWAowPi1gVEnV5EuqYTOCyWdF8VrZ567O7NV5qtYgtehC9ryurH
8SgqSVsbB2QWhq1PBrar9ED6TFLPhqAMqZPUYHjmf53XTKAzmUr7ZboPtZRtAXyudqRnjh1NH8Ku
P5yq/4/XZ4PvRIF91/COIxOHOeUQT2IZe3BFPJYETC81GzaennFyNUhqWzo8h0phqb93E72IyttO
CBZdE9bP/LLKiiz1fcsXRl9sGB9sRDQhn5rLwydxg2NKyeZ4KCMJ5jn7WPvTMThnRf0K6//CqKeE
kFIARk0rQj0PnbRz/IpG2uDFfJwBkFHaijNDLPw0IA3S+M08e2a5cfYX2uq5g9hjY7De7E/f+72K
MhDSm1HBEpgAPPUSCsn8ReVkpOlzPju82xtQxAEzB4cVHDIXTbE9CSafR/GJ/AwOSJ+PR5W/TlJq
znqbv4PO6kOv2LdUK04RRUVzdKG8WGMtlxTR2H9s09Ktvckg7uhYcWPLqTFwcPBcwSpeIygdU8yt
QxxWkg9KHVXAo8bDtUE0dPMLCOPMzKOcKTZweXZkAkrSwGoc60e6smePKXNX8QN0RTFpknO475OU
rayYvdM9wpH19d0NeN6+86ytqXnsKey68INF9T7XsLP20l65t79+DwsnMyHLhwSXuSv6W6IfmI3U
DAiGFL0gyw3NxIxe7v9M1SI+H8ISZkJHcd35hjA7yAToMi0FSAKA4j+rfK68Bx+yn4nCyJ86PWXy
VRuziZ4Wwud/Ltfjc5Fal9CDtIiIcsHsSP9jdAT2oFR31p2XYV4B/0VRTCpJIiWJhjEZcex5d3Ki
iG5H8/Sx8N2DYWHQbaIZ+2aj75DbXup2dlWLnvIFxDhgVW+ELVgt1zfaWsSHS84A+tACE+DsWE+A
jLnnnnQ4LoaxC7pFNBJV4g7INOSBclXCwDHJK0aivw3bymhjQXesrAQb9J7xObcli7tuO9peGqDH
i/nnlEBszTnMn8A9Oajj7fnjBua/sW1g/XErh4/RiQmEQWwZdUX8jQ2C9EfMZzSyji2HsvVcxtvT
Qm91p4Kn//lBXVfD9bdwy0+f24f9qDQ06eXAypUsUdJnyxvjyslKHuxb6UUZllIVGFU6w4CIgnBT
7dy3B23PLIor7dVRZz7BPh67ezn51sYtVyNeZu1t30y9VRISkAYYhrCKHy07GVVdCYQAXU0TlkV7
r26fV6mYDYNpI805R0YwJXCajWIVftVr3+Ud/9ybc1n8lL2KTQuPUnnEQTjaS/QOdaXutgXnrA/R
KlCMzlAOyE6GGSjdthwvjyoWFEOEVi45InBltzQ7bDsGluHfLU4ZGJ3gYq6fZIoblko+GcONctB8
pJEii4oy/mJSDIVlz5GPtwi3nMOhm8y/hVv7iE+hfY1/ZHSM6w4ecQaXqzoc5d5wrlXIEBvQB1IB
SmRgJY3DTIuyR4INtt5Wu0eIsfW8Qh2ZlnJaQKxmHn5byGMmplQ8p0d5DfgEsPcPot503FbbW1lN
rUZtkwjlXpzaHIVU+QfZnc3hZYbxoRqyOSaGwiNlAEgRvbbJtUM2D6s1iTPxtcukLBIu71VwYQh2
jWZgIU9eH7UWDINqW6EX0aeFlSgQqRLI6+sQS2PklN8vSaxEcZq3+i0w97gwywYRfSMZrDtPGJ8c
iiKTSYCuFaJ7r1C6xhiCtS94TKy0Qh/pcCZ5VET2T902NqqDOKzSbLGEnQ1IfZi9GxqsDas3jSt7
nAOgm+TQwtg8l5yoq7jHI8Je4gQb/IdXajZKEVcCiIdUStGHTkMfovFCMo79xA13ShZbzVCkcE8Z
Je4baas/iRRjzp7H0Zvb6/33aF60+M+/GRKhKor+p23dcnUYW18OiJ3NobbHIVjDhMTYiWY5KqKj
X1ETsmrn9V+oLl/1Ch0vKYwskdXAP9UPjL+mqJze1vkU5pnpKAkP1s5s6+X39B6kCo24sIAsUrdB
owCXY36gAj0/zhb+z90BXZFk9TFlOJZ93hFYgG0WdKtakax0TnUlx9utoOlalu5oITmsCuhSY+69
Npdg3VkaPjpcjxAz7MpqcH0/MSmf/Aeu+QS+gV/MuJFdlUh2UKbFbjfJW6YLdY/6rN0nPdVMN53m
3BgzqEBMsiRvhjOpCtlvQ+v9yoHcasIMRXvktDEgCnqu6dI4jI5ZGsX1cup7C/snyZN87yQaJuXs
ltxDnQLBfIhGP5Oi9eFASWMB064CI95ucJ1CJRrJMMWZgA8yjO9N6Yw/GhXHZhS+T/pZt7FpptY2
TE/6WsVHMx7SjYa3rmZC8eMKSUcq0L+C6RaPa2lYWwTvwTIZsqOdH0H7Cl46L7lGAK6G3F5/9DkK
RoBNc6lhEUX+2o2jGugM+ugIkIw7jviAV3ia8bCI5HqG2cftQEaes2conVLDTavfIh65LkyI2tK0
N+G9twI6ZDbYy3qc85goKQaLyWZooHmuc39yel/gv4H7zbLGYF1u9e0n5m09BSgDj+EI9U1fmtPc
Z5tGvb9ijBebxMW3uF9Z+MdoQzDqxoNu9vwyAfOY1AcxoKWhFu4m/QC3+TXHtZ+bUUwC/QzucWk0
Cuc8SWiGhLNI0/EH0hEhpBxfWDNRtbLKy4aC61lkZrD1W/Hk0OSqpVKPe/+g5ivaes72MAZ2Dm2O
7xr4Yy6hZyJjCx7Hwrcr0+uKInwHb24N3Vk8MZSezItD3wxVQD9+BAjN5SLVaKe/OMB85HCKBY0+
t+SJFj8qni+GFwUzruyZjSC+QVbqDqE5SPbLtt7MVkQDvLJHyD6B+8IHYFglHmUdvjrImj/tpzOr
KFM2nRF5EY+r27BA36GmtuJihz4NO6xX3s9WrB/vgNBlsZeuEPjkBck9+y4LBkWauYjjVpNpF3gH
KW/YKyJQWBtGOcXNmYQuXWlj/IULdJkDB1dMQ4wnKTCM62jxbMQQtS1iebjG/kUa8EqbRB1KrMr2
VOWNwk9q47Wv8YwA1yOJML6K1PsHjks0ZDHbaOWSq5MQ8KdI5ddcj8/GH2Aty/AP1I27T5W2oxrt
2m49SOlsjXxKTHEp2W9zakTKvxZEUiCikoGK6y7mrP2UsOHTStIrgIvL5O7mGul8awKUuUp0qIAm
H5bukKfFU4LB+XVqFexOIJE1qtDYb1indN3uiy8P4NdoamaItldmcuQTU/AmcBJSk8SX5Ib7zWKW
ie1gMZBNMifCe0x62T1HhYQJ3A7+AngK9qJIZDWHjogljbK5Zv8Vj3iursX3IE1nruJW9iZVpw4P
iJrkEq1UxznT9GjiAygNIV+gmDR25zHniK1ZNKG1TYc+WmKbmQn2mJotDtPtkCrojKtZu9aNcygf
Zuy/V12XNijqx1rH9RrgHAILzMmthsFmLCrrFs+5UbxLsEnHcjEMQpO0hLNtV3nEGv0Yufj4jXkX
/b2xXn0ZHAgudwNRTnE1durwdlMuL0Bo8qJcMJXtWGyhNEvbYZRnUEUk5ta0JPtnwoC/w2s5Pwr7
3Us6XqUgnUx/L7fbNK8u8f7gurkDa8BaYyX2fmHi56JtxS6xtjMv394HQo78GzcZlZvDHkyakC1P
fbUhUjOP9RoEj1lvuQ/gjbOj/WEZlQyNl5HgbCKIf6H+c71DbEMdrg3WmmZvpf5zigu9Ke+pgn/a
SKGlrUYuuqNXIDPf3xFWbI2NMLNFpwB2cJqUelY2A2Lpisrc9VP5LSUmoLc6hxaI0x7pgZHGbVD0
0JVTXkVNn4p/yyKzbQb9mxTSQO5LjHqE0ED5xgXiy2TpAzyQubwkHIyHlVCHHx3VbkcTo+FkOPAd
o2MZiOqOx+Zjy4UhYVj8LaVPV+0Tjqk2DaimJwgo3lvw7Ix6s8Etkw7yfphtvijeXm0EGs9QFaJ6
wX7Ri4Ff5fLJEYOyWIeKC2bZXV6EqNhAKZCzcfNkY2FurYQmPow/xgbcXMRJyQdaqt5ZV+zP3YMs
5JQJqXpsnl++HT3+jmJzk1vWr7g0qX9U/5j1fNET/ixnMwNtsHKV/mX2a6xJ5ZbNRPrz5Et4wcaY
PbcKuAiC8aVPkaG0phXqJks7Tkj6k2gnUxqmkkap3aAyKOQkIC2nfHvObc1vaMCFOBgSLs5RSoI9
UIecHxZ/55jET8ouXHdGwBekMOVsUNITe13DM2rr1bnm4HfcZaWnREw1Oib0s5sf35WGQpOl0S1e
7LIr1G6bT3+7zHgkrYxL1k7cFxIRxoElaJRWtRExtAd9Q/NetxhK4GJYDkph9Rm/t/goTXJjSKCt
+uUI3cQjeoITpRv5r0VSo3/SdE7wEwFfRyqZvxFjoY/tMX9S3pArk3y8Z4J+Km1I5YcfMnCQcE9S
vNuBZfLEP1wdczbLM4QpyI2aB45kp1eXP5TvF6POfeeYK2XfFwNXWzkqGKoUHUlTBtCKJowakPAM
zbBUwEMwa+Vmz0PX/MfTNn1sogb86ZMX508MiCQTc9M9ytDbVyD8pGVFXaPaQSQfQAzbYHu8IIDd
EPZHGhtMLgLTqEJw14V3C/l/4kc/PeYEr0Tagj4Pt0fOS9LSY9s7/qkspuQrutH8/dLhJt1076SO
vaAXnmAnwB5i0Q/gFCIE5DJ5ZLsm7Z2I3Ak5kC+If7XS3h2vdkJiHj3IqZ2eONBnx/gQeInkHzlL
6ZE8XZGaGa3l8GJ6Ziz0BH1RLIR4M6tTMePvgUbWKFc2IA8GBFx/bpd+kS+JggusP5GzNtb7r8Mi
Q3NMcJCCU5185Xfclis/zU3Uid2xw+9DrA6NAMP8vNZX+l3cjdtE54wMs1WPm6+qPthfuUvhvanH
W4lN8o0KaL7PIqPbzPX2A7aFWN7tGf1hS7CSnF5y3Kdq3MHEoIm6pcuLqTxRYYFWcDx8sHA3oWEi
tK5HqsNKiSoqcF33fAlx5hyGDLulDIDsZdh3s9f3YrYFikZC2QzABS1AxINXUqGR35e5m3IK0mox
Oiz3sbpbcagBRwIkA8meT/IatYNCmfq62a0Na5sGIS6M018V0Wq+43ihJ/KqEhQegK09CFqyoFTY
wwVZJQ7S8nFREqQKhfhZaYqTmi8OcXeB1SvU01VyU7txvBVmF83NrmJWDIr9gzZ7aZ9FM8pyvaXA
iICGXvNvLmsfQ4eUMH/hx5F1iQvbKN5bVJCem07YywD5poq+3F3QxutepDG83CjG8tbxrwMXkqW1
vj1/UrOmpvug5Kdf+m5f4mmsmfUIdhE7X87yc0UNGoRvjslOdwBcYjHBihoEtu/tFQWsk66MGSlb
wzOMp6QfUImCzFM1JWvbd6DGp67+TWb/G+PDuhWvYwGk0RrdzbvQdhS7tGQojsRW1/HBeJwLp8nQ
ITVhUt4rJLhQuXDrE6wtj2prdZWocpbGSK3gXJiysoaze8nWne5xKFsIDqOhswJyVLDtyMOcI0ni
S7f4hPfEBGevVR3Ka7DQFzKnfaevezs+m+Db8ez5AOvD6O6Qeng3PvTYIQekc0FRKjUF8R0QJikK
i5xKbkB3lxIqvwMwO5rSQ8agTWKzfmr1ucmf5XU0Nb9NJXnkfs7HwNoJHGivnESzheGXdBvdQOE5
3J53Ca1FxzSbZTazg/AIICGbnsOFZ5P+SYhiRSmv5QxuBKd0va5EuBLfRfjArfWGCtKibZYmLAOx
ENGn9TB5LanQsUWdtUtwez3wT6xecNPqPkd6oEc8qP1DUMM7b5H64n8dplWPGVvfORhzWbPxBJ7i
cqwJkksWi4UmpcDhOg7ZMtj2kURz+m+fWDP+mds7k/3D3dO7bmsZCfnAr27Htgsdo8oL7pPtBdJD
2Xs70RapCjVhdv2AL69DQ4eLrRxIxjUlFo5NQo2Twb9SH8uKPPhcMB0u9zM73wGNcG3GXfcQwsuC
kQ8069NKkV45/9YadRJhOFc6lUDjSEOmllRIkCaQ//dlXC+VkAVToLubuRt9PXV/WvTazGo4rlRk
U/KtzzDl4acMXN9V7GDPxHOwZCdXDTP9e7TKg5x4twDxpSL6++fzPukcqc9lytaoYpdCysfsxQPp
tHhMsjtk4fAZphlQ17Jsa8oOSkNCYF/CkCwtNnpiRK/xS3dN7UnDgXZlmenlOY7+GxjRB4Cpm2t+
qP1mjYNGssubAzZKLjwOWjZbbvgfIok9290GbRlfvBFZhPVapVXDGkGhNOz1MNHj70IoMF1cwBeG
tv3yJWn3XSsDxWqmXndLtfNQlgvKzcNj/y9S8uljrJ/Q5TDBorqPEDLLXy1FMQ01VJ1LWyX9YBIT
000KlH+L6FgmnNXooqKxyeTHsmzZpZ3MgKbhyiajqx3+cEDLJofLLDgXIl06BCkOXo3A9yUFJ1IS
e5aU+GBIxl+keaDHYbhN39aKjP1h4+8p1h7qc7aQg2xAIY6XA4ZMAlEqYavqcJrzFPTMx7sqFokE
M8Xn6yOi8PKwwVyRVfjxlc7LQoPw56Ah2U0FIETQOZmK1TkIquyDg9hFjavQyGelQ3Do1R23yLH+
pwTN72HbfPPBLXW12wBRrXR61GMXDDgTrhFZTRqOSyEpZj8NDIa2f5KBIeKo3GNo6eBI57GzM27L
kpgHX8VwwMdipJwqZOEGvtTl/s2i1jCjc9aQ9w02xlP52Of8y/GodqiZsbXvfzrt/LP3XM3+DU3Z
jGsCAcmDoULhzeS7ObYLZEW0JHMl6JaryOove3QBIg5XKvN2t5rJ90GyrR+1VJvQcBiIJ/UI42xf
jUsahn5cnqch3KAbVczKqV5cq/awzWi2PWWOzsfk3uAmFEFNaT3QrE4m0t5Fso2Z0CDFpwThYTSU
62gqT3QWqYK0edlw62k31He8RFXR3q+899Vn3Kc/P3dkcGhnks4+UKTDFwKl9LnyN4tpUw8OUmld
enQlvZ7QSammm1Pr0NgveiCzNiDVDiTmG5knDZkjb6fBHVaEGVHeWBmHgGWbPXCCpP5mfixg6IPv
aiCmIVkd4vfF/D7/EvbcygGhl4CFbMn0TWUu291Obos5lhynookAoWpD0h7aPRjG0lEUHi5m5quq
FsR+1d5EoOpP68J0dngCMucr/Z4O6mrGYStGRzJkS5jFWhL5y3nOw50kyRDsDfYcu8WP1hqtZLFX
SPnGO44f0SB5eBitlaiQ7nNdqRmKmgrY2wIfs0zYS0Myu1+qDZhZNEaBmWh06Km54N3zQ26I6qVh
nUYCmblwefXvXh4EBhuZqBIezmfOj5MOUdlgu0RBw5QU8YFsj0+sCPkvg3bg1jkjkGuLLzieAYMl
SC3aWl/pH/iCwK63Grqics2qwwXWS1yy89+5FtWusEUITVQEzydx81p4Qj4O4SuRxNzUnAP2s6Xs
Mv4O4QMuT51+3y/p5UFDSW5lmMbxtzWmYk5/kv9NGWTJAb5spms4ODv6aYdm/YNmHdgvUjGl228X
QgiiibuVPNRStobbbzhjQj1O77t2oLHBuJsDRro6+7TL5tKV61RlPS6YEsClCoT1CQpR8B2PImFU
hTZaZ6p2HPcmfTLA7hZp5PBCksa38aRVdgKxTvIhPbP4j3zuRbUfgSlq6qk6+Md9qkm4CDqR5A9H
jKfAtV4/6bnnzxFr/EBt4qX6MgtAIBu+03N77DVM7UFKyFYkod8FDEX46LHOE06DqmVEHfvj45oP
5vKT4FYidMI7uVU9C3WWHq3mBU7r5BtTPDijtNzCLX43hkpKbuRU2chIGNmbabrAhBI0+WeI1wBt
0zpfLXQDhrJpOzujS+eqLYB74n5Im4YNJLR2W/Uj7yYawVb8EXBUFbj1oF2ezXQTy9KqhrtN19te
9P7p29SX8sg9vQr0kBN9NhjEiGLiFHcMfbCO6zQETf8DpQ0XmqtY4ZBETwqn4Ky1tGa4XJMpeQf+
xBQaG1XAO6I9WN247/+KJT6W5UKG6aMgiq9uHwVUyXI+105K/LKa5UC5kQzcAHsdHgbD4N1OANBd
uSuYdDTKpFrucX38sbk0UdplkvSqTC2ZlHlyQWUYU+BHkoyZeViAx0/RXZjRTYrAnGjLwKjT28py
sk6s74sdx7wGCh7IWIW3zk5sE6GSsIdnvg0ddL3MJMy0+ktZuWdW8QSjh03JJU+SbWsQeo0k7Tw9
1wljKP9eCP3tDdZAYblR5RAHh17VnYOzDPA3ISsQOBRJiGA2+eXy0UB0oNVenzpDfYHHjNrOanno
436iZQogh0rd0HeXAZN5K1GQ/4d551X2cNPMXtANGojLuxg44do5x1ojVBGwbG9lA/u01UiQsvHs
9CiHld1e576nskmpN1x0eUUxrujfH1uwb/Aag8EZe4wAezX6/XtdB0ODnMIZHqXZqzpCClml001O
7aKdVL/8+9Nw/omrHJJK3fpH3TTgJNBAUAvWviRAeNqURj1J5ilHHkFDkYXtofIQimDK9d2i2lbW
hl81fR1XB82X+/FtHbZ/PMORbSbfbMiD4QHU3ne2u1lU8thV5nyszNuuNtU37H8wDmsqH9z3RY7L
YmovQ+/KTn5+YproUMsy/2MFXbEhRYFe7xCPdgu/Cibsk8+tDnCvp/0ncxcyJsZzGPp1MyI+mfqp
UQCS7oda2GAQryxywSQiFHwZ1UZ6pTF325hPv3RtzHYDxJAQCiOrWSgGa4Z7mv9/Jf1NQwvJLwUq
d3rgiTEONqOjwAaK155FbjKnd5RuKy8iGiDluddbzyx5xTdBNfjGLdW1D1OPQ6UOs18565D7Nit1
Noc8shGZuX+IR9g9eUVhV4Ku2du/voJJSYwZUDa3vgvx7uZUsWzeTgXDuZbzFQLg/9twzz8VimM+
0iOthnw8AK+0UPF914c1wMbfnMnWrRIW7mXoNHJrXZy52sINNKJhJtlnh1HF01jDydyvxQp0GHIh
wDeQUbboh1XKOtX4uhldLmtjjRJv88uNflj1qAF/gSV/1Iv1rAFzxRxdGfJ4gGbptZguwKSZg7MX
juk2hoIsqnYWBydLXvoWJeXnzYhJmf2F5L8spmaHAh9sj8xuMSHgk41GzEx71GEyBtwZhLqvkvqD
kKq2AGcR7+dzmUDJLehpcxLmcxiZuMrICSpPuoqUkfyNoqFaiP8R0OzX+EeGD7crqGGeT1l86joO
osWyrRvQpsv6T8ig2RfuqMFAF5WEri3BbbnnNKcGS0zIQ61euUW2a8RFuDcbqt1hTaaD04LdRMEn
qWQucXjTggT/HlTCbm1mapYGsCjP3sOndqXjgKIVOjtWJL4okCz0fSCgX/+lqQLJ5s3wzBrFDBZx
yDHslO6cuEQMTo1ACBD7huZvnyKzoWqPeHviX29EBtvfdFtKaetBEfF42J3z2thD2d8OmTqOR+K8
//G6tUMsiHngbHGS3E+/agIaOiHUyQKhzIMMSTGcM8RNlCroDTIsrp/sv3oXDIfMqAwrUoe+FFrV
Q505XhcboqnifDE7I2AnUSlK6CWHDbwe+Oo7Nii59VzlZJjc8Vagyd7sSBaG5eH86GpmXDhuZV2Y
BKAK1U+JyDVSUzxR0ByKNf8Gqsg9aplhOYuvSMQ/8Ks8mvwzHHC5s0Onz/CYHAPsZuXarcaJ+ksa
JjkIzSIasqSka3Ita/SkW0+ybgtYJL15YDdu+alrWOsO7WMl7ZZS0GtEZ1jKTXJGupt3ApPzbdk4
G2xSUY/Am+Sm0eZgZ+yFkgzRlkxsYTuKJyrzLShvj8q3LYpCktx3x7lP9ERuWFmc2L7vPFCwUdNA
VPSTRenpi+Q5DfunRBDGG98fuEw/tGQl7owOJuodqM4NaD032qYx2SVPG799UJE75LrYB2v0jLOa
LzJPAgU+OP+ZJ2M5LNvu1IA/vqGNarfHOiPHw8A3ydQEavjb2mPw3HfURufl2wCAS4VYlbjPzEDb
m7UVa5OmtuyjfnQfnHIwmOunbKZLtOCp/MbjLk0va2JyCE7xD9RrS1+gkouyr2RbBh2bW+AU6Ala
fVBwOP29zGfOgb35GW70Y9TbHd5v3XZBT83pGRH8S7KOHCNkBERxe24aUzEUgk2A1UerNDnDak6d
mdcDZY0X7dMvSgmJm68LpdHpd4XNF2i+lhA+QRySB/6xxuCX+R14w+Acy5y0jK+Jz9IlLxgEGXOd
tvN0wE4ljA6m8ij3fnnMsq879frQtXKD2i+DDz9xLSfaGHcVP8JtnD+UXNy5uDItpVXfLh5dt/Dy
gzxW9khbE7emD7MSGZXLuNmNWxOa849yAKO7qoQTc/KGcSZgVHm9cbAsZ8E+/NS1nvofNLEZeUf9
NEOWmJz8C3tbj8oSrBxCQho0eat85jt+z2qm8Z7fOxcGQtk4Jl7HWKg7ZbcetjVFrR+xVw+EPQc9
N994iqu6OTSMGlTvF4+Rf/pUoJ3cVzsg5Kl6w6OF30VsnZ4AKLHetvxk6LdksrRUlaPyenQhFwjL
//m+7mZsIT87VO5QglBfaiLX+tkcmuj4Iv00c3HthpY78ylhp+C2m5Zmf1prI1dL0ApXNo9SqIhu
nikmE1VQys38RIu43GSRpzZ9kD4jzTqmGF0aYzVJ+RAXRZMPPS31Si+uW7ZNyH5SQuVHKu+iSNv5
9zflk9LfGWa7ulz6V5iLF56j3SpvIILKccCiOFEA5Adxt3sUSj3dUh+s+h2lH+wlLNYCFvj8dq/B
P6671z6wh0T5aS66CUD8YpVAUTVXulbRWzFXjtBhdLDfPzVexcQZ2VXBmE72dP0sHBohgyIgxOSY
SAli9RuRaOSWgSB+wKXKwlaRIkc7duCkKOAN4MGIQBdhKhDPFOiRdW5JGODKdWZklwvdWdiwXbTC
FIP2cmlqJlI49i1BpmTizAksd6quF4zPYEJR6mj+kCW7l3z38RB9gEABVS1+6vcPLKHc362Ow07y
+4NdpeU7lViuJJYvH1zYy4Q2RkQfa8OJVI9os1yDQYOtKDMRiZRkAs51EyR8Ogzegamkayh/w1A+
g++BLWxOXlVA8Q0bTqeSeu7io72VP2+bqBchWUMFho/iaac79b67IT9SUZN8xByJy2MLM+UyGisC
ZTmWck2KAsH3Mdww2rOgbswPS6U3yhLgyKTxlLOnY6rHv/objS300at/JdPQrVBlhITiFHC1y3B9
7en1s3pAHNTpkp5JILB8CT3B2bs42NSN5zHfuVBGwB/iwWvZ76wmxiL4k3Qgvjb2eFVHBgNwF7zX
xMcWVQStY3vdro6KTMNeSdPn4PCHIT3I/spPuP6KMImQ+2Z2ZYH6KqjN7DI6raA14zSbUGybxSZP
H3J6DNBT3/0AcaWCv54jFfzkvPuW4jUG0JSmDSG4GUScotMIFnn2cH/OYa8dT8B/diy7n1BdbG7H
x/D606FjSSZzt/DNdwxAk/1WakZ7GvQcaCjOF/WiP1ldTRke1a+zznRTzltj8VW1cFVq5gGOQZaT
Oc8c1k4+d9OCaX9bxnyht2J9GpwJ9fbUZiM0C2f55SpgcJJm6JtWMDl12JxCGR7748vQeQmZ5LZl
1QQ49/IBW0LnOcb60kGsrCXPtq/+d5woS/oyzfLfN+l9pVc4BPs0Wwa9gCHpT8vVz/8C4GK5dnyQ
9H3LxNsSivhz63boYXIjcyPk4ijz7dtaoe11oHVmPIEXX58Xcq2jvHp7T2KaSjqlwUJTQaNm+j8B
Wg7Frut7cY6oM9SQtylv+ZF5rjy9++mKQXVm1Z9/QsxsSEYYm4mH09wUPYFdpAKCg6+Zy3x+H/a4
WJDieneKYxN0sb8jsyCPJwcrd4UiZD5NBPMQ3cdSIGrWkwIf9CDtPZQFdNd+XSST+IWF9ntzPqBe
LrfUBWIvqIB93noMNUKdF9Xe9qV1UasPrx3uxpIq2AQAJnlu7H+sSVhY5Kj8ijZOV2GVmp4DUENM
b3jkML0AvJ8XLX9yRIBGqPKkL3jNCV5Xc7OvVMdP36pSa9qAOZ5WsxnasvbGKYdgSgsdAlTK/pQ8
u5QGYDNLNZbr+z6tmDBqXKLNEjOgKT45TD0hsYWkAtJeRoaOrSGZ/r81PozRQAfJxQSs5RgQuI4s
yLJQHk6MaFormDaPzFsGkCMQg9TmF1xfzDx6a58mOovP8GuimxEVi4eDwoFAobyAVTmnILmMiB/n
xOHhHsBQuYhGhl+BakCnCSiU7zQGsrR4JkU2JqOIlgp9g/YPMYmbKkaRyoF3UlHKyrLmhA/Mxop1
bFG47O223CVJ+VRt2l5LTeR/AOBfOMe5ETZlK8G8ur5m+7ZT2RrY4/Odo/1mhncz/41EYgJ177YJ
3JltT8V8XJP68JYMPq63eojM+xe+TTEX7/DrU8fcS6/R3Rr/fFgd52dTc2g4TUthrxnJxSZFjf2e
9XJwSbJfXZynZvCiN8p7H5gpJVqvvQBeSXbuNWsoOqiCKii6WJPCzCtYOMyg3/Wj8fb53nZnjTAd
rKQ5TVwIfFBBMNhOuG77AeYa8wjakLGfgRiDCH/d3XNW6Zo8Whi3N7cXP7o//GQJBaHZ6qFreGRX
B7mq99NSc9+jud/uCViS+5nErRsJpzsr9kNZ6xUJBBTZKZfoNlL+n/UkLuvCqDuir6MTqXJ+hnSD
Z0bm5adR3Q+PndZaPvCHbJiTTVN/GpY26sxoQlgefav8/DQl62oD3o6MFuXJHShDr6j4g7kiGMjb
lgggGftKJcfVrkdmyQ2IVcvwTaeoO25wCCK9dsCHhbcTFL8dTWUaSKtY64MjVqShdm0PR6vCDod+
+MnayDRuFfrRif8hydtlq0VXL9WZWjecmeLZsvuV5NlGc0NurYAkdU+yxrdJkms7OwIvBozyjTVb
JbpmuttUIKew/99MpkZ65Ab0kuoE4+8Ykw5TO2tA9ZwS7vgxZMXcMCJNkpGWWJLXf2My5zol8BnT
S/ivMRzpNMHqnsakiAM7QvCOpJ/17ZK52rOORzffMYBBeet32nhbZoo0tOpMYW83//Y4h6JzHy8b
7z9aeon+io0ZXBaLYbclTstwVG8O9eM9kw2x1EX0ZUye9zOmuch+6unNHwTvqsw6mmoRVzMeVzAF
98rqSflPQzXtyuFypBfw2U4WuOa4p4z//diKzmB9vPITAM2T3AsLPk0hchYoDnKzxkSkL9WOKO24
zGXdC7LnqFpAzogwKCDnf8jDOuaC0dzrsR9bpP2tkEE9dxa/4lt0rAHpprVKCVFkHFXqyRvmuCHQ
ZG+XIxz/1WEiljXOQ2kvfazpgKAKNDsVMkxhCd88djw6sR8eTlLTdihpH7CCFUOTH5bVWnFL23Bw
v1QP95OC3g1g14hBOU2O027F7q3kyFoi3Ma1CHTXOt4kBpCSOsIafum1xlgqiWh8Xg3pebUqqK/2
oM8QJBG0lDNDsqaecCZEzAvOETMc0zLS87yl74flG+zghh4MKxtAfj8IVdw7C6YPwDPaV7aob+wx
Anz+6iWVaxhm/9G4BAW1oIKU/xZZOzKMhdCgrjIcNtOhXUkcO74CT1VRueEBdim4wcIPV3MOv+3I
fBF/C7of5tZoTmv25eRYE/0A3612VphSQehtxvlFB6P+0NOH9shIUipGg9vQaKpb6HmxMFoM3SNh
p5hAdXwp+WiJNkCahDkeY5ijbu3EtwJVRoIzP4xqMysBSSaqb0cslPlXsFdEUTW5vlpCACP6vZ+a
pSuoEgqQp1aWrrban731oQ2+yjO8+8LNbDrwDVKO3MFs43dgBtDDI5/A8iuHY6rXqAqeHGc5HoNd
elFJCMq1H5yNlF7h4W5hzdS+PWhISaOfgTxnCOzU538CSoZfOHqO+7rcFu1IJuq32eX8gg5qVgai
Ay1oSgsOYKwUH1cOH032ZHMbuQIkRiZuNHEZgjJR+IwMgI2jrNOKd2m4FSwKk0GjzToRe7B4TFvS
odaSE34Tx2pY6TU+/1Cctswxei7UmomhXeLt7WUaTc2hUerEOqQZuLVwh+TizGBddDeby+x+hl65
YpTzKaHJ0TXz7RwOYBXfZWRyXxINIW6hmPUbGEUAyUcwz0SazplpAAJYdzHnr3eU9epDEWsdy5Nc
yb4j4V/zD2VkefSbzv1F0gueMZETzt0FqvAhbn2HurMETwsFjdQKwgpiTyDB0623gL8eEBR4V1ie
D21pP1y725uzHitIP4MKXjasSJz1+bfRHgUogeNOzOcWjT+Kp0o5zTXfKp1eJq3zyTDnqElBCpMh
iog/DneMk0+F6YpuMvj5zPHdXMIY+K7Osux+9kVMK20iiVZGiVZGvRGXQw7H9eDPKmseDi3tsDjx
CJ2yQG/NrlEFoQwKjSsFElko90TzjKe5uYMWvBsOcnHDmxbJGjNetxV2Ga7tSxhGMqhRVXeEi96a
orSGNfq1Tl15O8e5VebhG394+HyWtBfVu7Gw9T/785mTix8Dw6Na3l6Us1MRXFtyqGyRugQWjvqk
9+7tDjjaiQyDFz5XaqSyF0yhH/OKbRcMt0txpOEuiRTGaN9CC+Y2p29xjd7qC3xpCVKOM+CEUbu7
74LB2B1OP7t8iQVWSlRREvUoHL3TS0tacOEuGDCot8MDg3zW85VOA79eEgHVrivxDDA25ak+Yw5P
CflQZn13DauqdKp/EpVoOX6ZlJ4W+dCA5eXCtWD5qBj3heD4q7zhJHglAjbS8fmrIG36xa9qRoA+
lmkBDfvfPRsD8n7msvHyNGBOgPn2aPzXpf/HDabVwAM8bla4ffqHqsD8+4cnjN60lUcjYZfVs+KG
mtd81I/Ho7IavreJoXOsAIE4UVgUORtoodVgsZp53KTOgeMMVRJmqPac6wyQ5IC8nFglmrigjlld
vN6IOu2QIUmVJW9YBGWd9uHelwDWVeCVAPzBcMYv2KXr7zKIPvIyp6OLO/zMF2O5Urm8e8YBqlxf
24MLhoElEU58BJr8GssD+z2GbXhODzLC1mbSwEYa9jHRA2A2Qs2yM8qMLjWkUBeEdOnZablTn3UE
xFJEibEg5ywMIgcVlqLB4Or05nUWC4RpcgyrgyMJJOVzgFLiO8rga4onxinQB72DeZ3BL3SScJzt
QyhhDrQ5HLmmAaCnEKwHTwvQWvw1otbAUn5v48mPniV1+j8wJ2Xxa8ANu6+l9yLZKtllnKnIycop
buZGWUSGkmVHuuP24Y5/kwsuRjcQsE/A+LecNLbInsuiktneZ9qlhufOxcGpbex9EbqaqTlQJru/
RrFfrapTLkKnqRvehY1mX1QNTF2wesFbsA33WWbUyiCfLXeIiArrmPJR65YzkwuPELtjXa956GC+
DSiSJNO6Is/xRv7CCgbUf33YyzfT4rXqIYuMG0fbZ4Hexb6eOVm0eEH1p2gUwh2TjnRvW4VE86Zk
30f9JOPrTAxhEIJYCEw5Cr2av84I/WNezeePI7qYJWSpNsJG+4TCL6ic87t7HZjp7BOQ9A8fddOz
tLNpen0/F87tmTi41KXtCeKCckhYKwc6LYAMLrZsbDnJqfEb8cDKYTEQYJSTU49/xhlAakQ4ss8Z
fNErTgh7bu/PIVaxHxHM6U28BXwqiNLMCdmmuQ4689eonGT3+Bsrncs0pD+jDQmT0HPiTX9ut/1p
5yVKR64K08pw2stIVBTJrA4+DgwYcRlV9ttgmVoHobGBBJYpdmNgsIkzoEvq6aIVkRuq6WX73gME
qtJJZEdZkDv5JRpkA4OQ7IXNHwZN/jO5VaA6/tw04Ywpjka3Y67BnIsIGJlCtvxbVxza5oyO5A7T
VsKL96jl4c1vpuCJVKsJsClQ/qxWNjxngHy9P6UltWGU7/NkpauHLvPYjJSn2x0zY/yFLrOsQhwz
CGp3L6MAYfHIug6m9RY7wdpPazI/xKayh4/QpJaalBDq+4octcOOfJqw3h8ut3Liuq9SDj+JClDo
puyPDx8ixC/gIKFsBFy0cs2CnDUqz/IJ2rjd6dnK4HJYXqvI98L+VbnZGrb56MYSDGBxVV6hgIXp
XtJCC4kjTN3tt5Uu76miOYvdwbnT7R/+PkwktYCXhZJQ/LrNps8q6JcZggwWAxrzAjNs2RspnqMN
2YoQBkZ07BFG8O+gXqvPqj+6niouqqVUSll1GnNyk3ZmgMJIIem0PlZceeSnvFx4NVEnhL9xUGM7
3/ylaItB69RGyazZLnVEymtwJF7fiuwHcc+0yuwZHVJPm5GTfNJ1TBPQzlrXI+wh1DMvydN6nM/r
0Feieo3wY+7+a76r4RVirqx5UxP19a7LdSmyXK+PxLhwIaAYEk1NUucB/tFhduOxaRx1mEnTjMzf
K0N2jYUagMj5b14uDGJvjoeCNegy6XFgegEhOSZCVk96s0hbb1uDYIoazkhlDSrNtr2fO+8oUE43
kJiJle+OlhqNul5eNHdmjiiJ/J2ygFqvQkdokjMtlqqteil0kIfxmaJLS+LooFGORhB/uy5an61x
jQShK0mBOFe1pvvfksxJT9UCkP0cXoqdifZEybgZhwLQ2HaT9wM8zaHLoRtGfp33lLa/CtA4v73j
cU2rIJWlml/+g8hCntvCPbPzM6Rr1vVcFKqVhhpd1DwtUYo1IOrIknltO4ws2xcMcD2XDRaFVeRI
gRtKa99jxtp8iTQXNNVVt8Fyl/OQ+25oNOGq8K/P6z9cuMS33ZGl4TsZh1E2/z+MlHu05ckQPr8a
AqSW89wZhU/68UrAP+ynwAQZc4d11M4Ijx8q9RGEuda4DHqCNhRSioNKl0YXTgWJDuM+OLazEhIM
1ZaooiwEMBzIQ70Bl4S8YjaVF8u+DUItBOf0D+03MNZIT1wzX9xfm0VrHCgwh1L2Wf/ATwZV0Zaa
khk38KM4gmeyWRI+iqX0/ObD6UKVzXL70WP1a2cwUKzyTOpJ9iyiIUhJfjZmCq2fbwG5FHnqIqxO
WDgum39YAohYSySFGmmCXNHBtlEuoe8UD2M++AP7M1ThHzCaqf0QydUE2tUvIwy0M3JkhcBmyWrT
JkzbpMmRqRzFxrlfez3s1TKm82P1290PutxFldbkpRO7YGAF688/xbTSzq0yC9vs/MX+ygRzzL0A
PO0G3C5XJtYztoL5wmNm3He+jtDQz3rF55l72QvbTgOlQReJXbd7/SDV3qMILDd9I+IoTToUcAjR
L4KUQqujlUY81mgg0/p/QyrSs6bhzgDcXsg0gnQ8csHQfxAc/Yq475NTsY98xmNMM3z5HYMPhZcF
Pcj9Nvqs0JOic5jkfDsfBSd/xBbQhTkYWYFOa1I+EtJiOq4Mw7pio51dTt4OANlrntddvNzgWn1t
cIUfjVJQeNEUQP/hc4rkb/C26m1fi39hgT14vL0odjjKDov01qMGKEc8ud/opNYtzBFTWFkukXqf
EkgBz/YtF6V0cksgWL8ulmHBT2+StGKR2HDU+ND2Z6yzfq8aR3Mkv9EASsG5I0gXrYrXZtB7jy92
2uUxBj9lUMuAANH0TjIYzZswbQmTiCB9DWIw0M1Xqk+Cij+x0cBO4XdQRoBmtCvZlku3qqbAqomU
Y5FI5IYRNVU61pxX2bv5Hz3mT0sEQ7U71j7JqijWB/XaGGMlBAcxAMGtAH1kfFuMF+T3cWkMuc+h
pvorZji52/C5HgcV1JAiscIiqMSksZnaxmMNIheUSPEkF0INV/9FUVZmsXm3bBl3kJk2kXQRNFlW
NzVn4vN4kGvDgw7kwYfZLwK70eYFHCp8heBwLTO11P/IBHm2tWMk26aDJbUuzUsDmPqD4zHZw7Gt
97M5Cbtp2mCIkkV+uLfdYHTotvoWawVAIn8t/vh68SooGT+ghb0NQFjXTNg3LqvJ+69BhfiQ9lZB
PbBZjivBfC0f38rW7OafPWv2+hrEGzvoJyX7hK0Ny6IGxRSgETrWlRwlqIUJhUehHlZv2tvY29G6
k6PpmSfxlJZe+sqcNjYVE96V6B/fDw7JjxS1LlJvx+oiICJI2at45U31Dp++yPlgDiyD4SIo5nnL
Sc6vT7/9CSWObSYpFuMmbjv+u9FRT8GtU5VDsrRk/8S1jkEfJIMUbw5c3ibE6qtOymH/I64SRS5v
V7C8EZ4d7gDHGga4aDffJAJpssDKpycZa4ZwUESKXF3iav12r7qTkOH8fUsK7LB9fzzvNr0NNtjG
JLW5ln3KTjjKZPAY0oAe1umSdNZU+xVsGkMSyg/9240qdTuSXwYFAJSITGfXGguAjuHpMrrWrRIb
F96LCALWtHEo8QeoAYGpqaxmKIC7Ac9dm76NBwltGBsrslbyNO7fU3Qpwxi+c56obXBKv/2if2E/
TIyeqNNxtlBq3AA2Ljd7JCGdQkcS2CU4i9gmkVmeodE6hCXnbFZRAkjvyWprS6P7plB46vl8lnaC
DfckrxxsTyIvT0NJnK+hH+gUc4caj3Sqx3i33HJ/lp2JFF85om31GYvYzWAalETbZ7+qpvkhL0QJ
BPxDC1e9q9zlZ5g5rLYXgOCQgrt/i6n5v70xkWlHk4C/LvpD7aX3gmiqHCHine5PFybwTf74gPHM
fbRUCTMfCxl8SpTUV4E7wQ6M0zXwFk6MnraFu3qpMe1gturysd1K6CjLoC+Jjmy27RFXgapyn/sZ
oLmvgCQ3gFPYbeiSLgihsN0is1hN9eMgPCMc4fhUNse2FPoEKsAIREOYL25xX+SGqQ4it/67SD/h
atC7Ol4YRU72bJ6F5bRja+05tm31WKxK2vl3a+8Yn1zhbU/XhEd3DMQBeQfEK8HWMP9ebEFWyfBD
mpv9KexIax7YK3BCUmZd4QO154jq7mtULw86wlnLH4XklVox+CdaUNVUzSzozwu99sJQz3rhSyaV
3syWQfL/kIFWZRlZllFGNAcEeApxKMQw2GJaKb2MuM9ayJeyUBytvdeCR18iEeCfhaZKlzU9AfSY
lYFndQAq2V9XxZ3Slt8FX1EsoJAkl3LwhzhSxXXTIFsetVvTJ/V62vE/n8g8DvgtSRNb3AP/2th4
0SwG7jXfmhfILMLZNimDfGUh+nO7KnHP5L3RP6xqXwFROm3ahRhCOjIIVLV6TGwQKZCTq7Ekh1DC
wNgv8Sp8RdVpv4yy/XIXvYbdFOhNPiWRX2HbHFPLdSUilLkPMbWe1DU0iHfxpBTXzFrwPc9xL0k2
1tsOsVCF26uYFGucl15m5MgLKNnM03fJyd/mYhAxAG2bvJx8zhOLHnfh1csG4WIOu/f3ylMWN5/j
63LyXFEX/9y+1s4ZAsENTfjMeTsyeU6gdmTh+gC4wNhLnCMDBWjVLMFJ278pcyIzNhJMLDirhOlQ
Rpb9bAmrYo/b3mOAHR+WEQZd3JH7Ihgh3fyhhMKvQq0BEAc5x0isUR0e5RzzSsglUIPF+193p7V3
m1YFM3edyvmSZ8AGb+Zkyb/yccrffQFaSd4sdeFlis6JqeWBU3ju4oBA+zKoGKdHAS8PR0k4bTR4
7ymvJsCDx/3ZjkCp6hQRVFTygg/eW50TVaQhH6xO+uemVFFkKmzJhVGjW1zglce8l4n2CNWuLZw2
4afrxo6BrFUmbfyy71KcITz2o3uDdO7gqEOxWaubTDcZZjYWlduxHEY5DfIz7J8WGKwddPxrtfZR
3Kl8owhE0kT0wNgbMBBEiiYHojBxzkKIbEo2ijBHfglqNW+STpC45tU13h0Ta9QpuZ8do6IYhVb6
aOXjXdw+69ojK5P2zQtF4MmL/vreZuh47BKtmvmr8espTv7gHTKkJDAmENTCHj2tm4Tx3MyRAPTf
rD0F5PQ19mMhivKzAzpBLZX80Yn/k6UZ2S4VFVK3H9oq+9BjdXM8LNwSX/CqNTMBWlhitQhLVNfr
8KENdyhfJkZs1d6tUe6Xrl6O9tSMCY1zsr2M6fss9GEtxE6I+C9EJBOQp6qoebIEDU9xUR13Cdmj
8lqJuFIrDlBqDFQi8awrR8LnOz7juIlJcg12F0yEL/HkZXo8vee9tqRPUZ/duiTWNNI1kZRPtXLW
ckspqNOojl81sunQ1B/9eHoz0NlDCk5/Fsos0F5bD96BtpIr7YjT6NQT2O9xj0RlReFcrhzXeo3Y
1unT9Fg21DYQqtIeysDO2wLURoRSGSNtHyotU0ZvqwBoVQ/sDP7eS0kfnk8l6ZINpEEtsnJCBjaV
gaqCSUJT0KFtrAEqgFOi4ubIbnPqzdv8IBoMeKBNhRd7qMAUMcVj3VqaIpB8ND+64i1zcquJ96yd
WzfV5hMwKrRqRHTTUM8d8KPUwtKqEZ71vq3Iyk8RvbIIVTIyd0onVJ8fmh/HqeKm/MMt6pAcL7R0
y5+wXUlC8/kAyBErU0jpoI87LdT8polN9NaQyRRJSmCT+5skQm3p05qsRKirZPbSu4p9Y04YwMG9
bpQDWD1D24kfkE/9J5CXMXsCogROPZkRdCtOdfZRGv3yQw4F1dkHaAcs36kbPm+cA5FGctm8ue7D
5Sfd9NosnYK696vTY6g76j/Aqz20uWbpDxFS46ZVucfPxKdxVGSgiv+KhB5XKNbDS8bDYdkeLPiS
BPg7PY1a4MT2LQejEg5sNH84LNGSDynzlTjWTu2HeYpFz89NLePrzllrqf/zyqSjCvi5P6iWEPMZ
7iz8xoqYNC9DttVjX/gbLkS9Z2zfTrTKPzalF3sgzjEEQStoDpM5z30Fyp4Vipf6m7/FRhIilfOl
+YoaHWxF0m6R//5IL1cYwmf211fdM2+Y8Mi3OFbN4gnxc3d4LNJ4VPlSAqTcJ6DfncA47RkX7/8h
Fuy4nEOQYVAutdrCzgmx0zqhOYIlh4HPb91CMUFqHNAhqZZVoZUpoKI/EXckBR5lCVNZQJv9mBFR
ZRnDbJ3zs8QptDUjHFyHcOIUGo5RbPIgxRRA0oipduNefsP+vPOXp9GWQO8e1ctTRD9xCwIpMXy2
q+mAp3xFS9u4C0ghOdSZ1rgty84CbmPzV5ToRlmeh/xgxszvviURzBxActL3OmjDfzeumGJTtpRs
K4LSuwPwEvrDn5TSM1BOU3Q3rcjXVm/CTY1Xncbiz/f1CzIi+YVV/jZFRG6WCVFIxtt1Jdvo5eMz
UvdGDuDi/aa/quXzGvY7Yxbx4llU5IMMEsfC7dAhGlmgcv6PUGJMfzFEtk8GRzIQpZgRoxoMYqkM
yAb2t50L9KIULNpArqqQpznmeSsFvHh/1vT4jdk0fqrFOefypS1XArhG9vW5WsU2DrrWxjobdkVU
rrpqiY9OD+MAMGlJfKkAtuFL8g08w12p5ioBf+iLHLP/E3rMSpjR3R/iCpY+CJ1z/d6/aiQA4Zp2
5CjMEoj4Ru7F1SA+N/6Cpk0CRCPXB1dr5TDq3oQQ4Iz6tPzCyqLnUzvKrChwwEt7pggbUpKQbA4f
d60Zp8LwmFssZn5V6Ulut88p2aGpxnWSwG9jIDiOEu7xXS/Fqdc5xNLtUBkFTX4ARexQcZDyE1Eh
8WBgDlhmKHNvPCQBT7dQanCeCpiHLWnBTlHM05LaoR9oKHtx/vahly7C1gmtUGPS4YJ+KLSthF46
phW225bgooN3I81QZVDBloOa9z27ppIoaP0eb1yZopgI9fGRwuoCvHcAfPbmV3Yk5MYEAYeQvxlv
aoZ8Cf2V5rb1nYUk7wBU33vYH1f49WurqNHFSYEGx8Lr4J0cXpEsaLAlfGoc1PkJfBjOr0aKRc/P
rkYT4XpGzGo6Vg47rJ4hij0kGL57SGxNbzHtPOfFrwyH17okR8HgUBtQGj5J1HAtFEKkCBIsqU5H
EIu0PkXwMCiU+5FJYE8Y3NB/r3kHFFLYk980fyLqv60oCpugMWZx5ZylJjbaHVrtF1klW+a3AL6M
7RUd95peSKFNr8Nj9lS/iP0i5JiVQfnkw6aHVuXDeLlnmbxrGnqNUsjh7j/c+vkJi6A98Vp4vtCf
b7OMXEvpYglOaLHe/U+1hXopTIgI6PrRN1zACctiZIKjjdYL7K/sLPVabFwM+PbkXS05L1Tuz+9b
Z2ZYO5kS8dlSna/4D+G9bzrLt9goNQbilN2JOQEmWY2G+oULU8Xm56QqeSL3ioTPrYj5Fas076Ok
B3pIdlzMoKVJ+e/GmzH3dyy5nxNSnXs3nC4mygO18jBq1320Lp/2hnnnJo0/f3jYjoCmerhBe0F7
+dKA1s0LqJ473OX3sgRqrgEvFih8iTFuI9E1OssX0cwiG31bVKPvSGsnTAsJl4RA62vWTyQNPjW9
NcPyHFQ05hTQFfWpRQBi5C2FCSyOlcXzcoqPKyr/MiUGZET27zh8ErA5mMlG90X5QQ5L1YFhHjVf
MJR6SA2ICTP0co1SZwVz0bvhLS4Q1uuTeD9Q8h8v8WohAhLK/OU2Gqx822FiA7efbJiY7J6bVDyL
oA9I48myeqZ1TH0f9Fc2nPYjg9RmdGKdtgAZWWCqpFtsx2TDeQd9OUiOYq53pgekWowfDOPxWjb5
o00VJcGT4rHER55iFNuZtPag7IrQqqByIgj6wEgZ96mx76gzXg4L7y5+MEgB/brCkeAavXZ1ypau
bb9+e3pc+iJ7Wb4pJXQmByVZCwo9ltobtyVD9t9deg0N6OiUIaaZapShCl4iWadUv16w/dBxmpDN
9BPw3GCS7yr/TEG5ErgquxQhLCHmcwJu0CSNH5VY+mZB08vutDd9YyBMmDLZ4RTRUea1lx9YpLAD
a6At0bikBvohHizszhxH3Mf51Z05LKFh9rstTvjuCFvGviN4BTLuHY8oTPYd4lX2A0VdOGKiajeB
A+hwSqcS9nMkN+e/dlaLOSvpHsCYSWOaTvIHmFxmxgAfwVt4/lzMOMMys24xSnMUiZcFrEiMnMOS
YUZBS96QAsbfEqVzILLdZujm5WRh6JL19KFmzHfCQMaCWcSMka7oXmze+oCJYzztsZRBKdAT2scd
5jw/2TBJ4jde87ZUdnfAEdLbc4kvuKyJNaRfx5dVqL9iHV5COvjDKBv8QAGS4vPxISFaf+L5rMO0
zssJCGG3mmnhaqoz4tBL3CUJRXyzlaL/IjVbg69uPJZ0yPIaLOWhBs64Bl4L6IGntDZMfFKNQsgX
HUYpRSLp3hu5oRvbklEn27e8WImHTjsoAv52TORPhJHDfLbbbxTaCmwxZSr/Ej9l4Z+XLUbXVV1x
n7fCAMLv9Txn50FW7MtOZIXR4i6EkH7K+NVoyoBlzj7wZIr8OEEmNJIIRdnqPSZmABQMyV3n4R0w
Z23FNC+vwvawkVqZCOoS9T/5TGJBYvvlrPfVv+uF0tCz2WNq0XOp/+RukurZUExRhROT3Q1eDCVu
I4Aq+G8x/lE0cBmim0eEcmu7uRZ9UCEHZYlX/cytlScF6Ly/LyUOKtQjL70wLMXjWtlnsyMoe8E+
bMcdTUwFtTuVATokM5R61XR84LqCNJVLDgCIIRoYJ4E9HBoDRzGA8jMiq+lrgl4UM+XZwShXf+3a
w87/A1Ojx69B++R/XDuGbfVlITwVOyobSumtaMYZ2Dtl05tY+5HM8dNBf8b2CrEnvcww/pHUTBzQ
SrWfXIwBiZQPH2tRYgha/MM0iv53nD6ROK3lKnt2mMZVo5wTMpJWEhSvJNNLiY0L/d9m9+EFn4zw
ERIWrhTqmjShDXZZUe6jvk8E6zcPQDVTAL7ehc2/8wq8ok7ssKXdBcOJZtBh/saGdIcTUSrMyuT0
MkeOz5RY24XNQSub/KtSCw1nCD9/l67L/rPCeFc1uwDccmPkZLkuClzjMVvqVcSiuFW1i6rShJpf
zvLTnNj862snlNAndVn10llNgc2XeUI1bjqJZRSGRjoofvJApwk/GNY1sXSzFQvhA96lnxjfHLVy
0QoFR1u6jbeVGjHlbQ894uTt+DX06RyIxQxbxADypT79qmrRVT0Y120IJeq83Q6PZNE62ebdpGA1
hEfqO0tex19lNy5tade0KSdczj8O65JOkW5lWtuQmv+lpesAP1GmFBAJeLHwWJc6yI2Aw+xPmprF
jhP6wdw6aK7Yl3NdEptsjYHb0J6M/omvToCpyRm63z2MPpDiZ+kKpMGHNTPMZO3QtefOvpC15tJU
7trJq6gWXHATDTdmmQbv/QF83X5gjnbvVDUjaWhSIyJgFBJRySK0moqM/UOJx/DhxcBS3j6eD0jt
72dlKW8oMxzYYA48P3XpCBCqk6s8Q1i5COlhK587wlQpvfx0ijRA/3qoArgqu74/X8uHHvKKtu1I
EnIxICnUlPuQU8Z38PNoWbZBojnq3XUGDAfKrZVGVjKWcwwITYbohTZ5L12KqT+8/KOMBMgXY04v
xUstzvpYG7qppHyRjbhbkPWw7yascg9Epjucb/fnV+POH3roUK421OUUEY9werqbzc4icBdt9VYj
4nOYkoFP/spVGlvZWRIS7bJLfPXXqoHptKsPGPmIDIt5UGF6S30iWXMdHwwvQx2BK+hdsQXYozY/
23PsASX8iBtaujuHTmCNSgdKWKnkUFsRJGycv+lrOR/hUmQKUpSkQ6vd//vEV7E4EB9PVoMuvl/F
LnI+EbiglLzR1HgVy6Zn3QuGsDYMq5e/dqWkIMPaTQivn9m31X/8Z8BO+88SyORQ0Sc++eAUNj+a
4INCa9Y7Ep7w1M/BUs62J58DyNQy6dyT0NUzZjueH/MRwjboma9cMj76mY/oTk9R7QB0hl/DHr5m
cjSmnAH9pJ4vIm6gLFqBbr5u4EwM24gO0KN1/R+zhD51g6nIo+zzygjBlx/UgtDghKU/Uto/9k8Q
I7+Kzj0QXUQhbZjeRtxNT0DHLRtK/+B815+k+W1uaDAZGkz7m/SY9AO6Lw7D0c9Is8l1ceKgMxqh
ZW8pXIXNdmRe06yUk2EbdKcy3F6+1u+aikN9Uzl0nGY60BjgYtiN/QZDazEsWSO2r9Dies4fbwPS
lrtv+UVMvVuZxCo4fe8lThrz/R1Np/pvIMVnmlNcc33JMWDjqd/0WmMon7RbVq8fQfrg0T/MBXV7
302OM2Fc2Te3jsnbpoJP6P27YZtLrP/eqIu2/BBwg2JRng98FIWi7TKdIk7qUPCTxEIAjAjHllJX
HjRaNmoBpwrao4miINrgM7ZtiTQlaLr5ruYXK5uPJ8N8W2U8GjIO4AqWV4Of5VW8pJPqfGPM8aYV
UKjbn7G+05L+Ok4nph/y14W+y+sGTA6ZnsYkTo2ncWqC9mCOjIrZ11tIpzlwLcacrk8r9D/Cxr+z
7uM6Ofz6p7KBRUiWKGz/bOpgF+0dR3gJ1xRz3Qmy12dzVC0Ucqn/ptAGTtayWwGSPPLutQOymhX+
scgAfrTkFuEjeXrKjiibUOCuaOPdwVWG/IxV/HeP8zCNCrLlsXjM1pqiTTdKElZi48X+uP41ltue
Ubffj3vkUAOcFAUgmp5M1HVV9jcslLgVOl449dScdVlNqEZvQoAbCZSh9Vecb617wc3l/2I4wNGj
SHhIYE19BarHqL8nWzjIWZTHZiQMNUreQseZm/UTmVHgRkhlwn5+u+uoUowqTCyQ8+3+RKzhE+Gj
U8TB2IcDe7IbFWOgtRLgPXzF+3MN9CUmYRw/TvSZvqsQ0BD2Cm3QdnSaog8TvlmOu41RFOKdBFzF
lEz714AVESO6hyZYlnN0uX47iMfo+usTU8mumNh8dgWk286x4B/vNOU75yAORRpEBkaxY0/C0imk
zoSsnCwcJxUIwCFUoiA7akIQRETh9jwWCB955EF5y5SwUhRw5snB4krdAew1uOoSlB8rvRgPR935
JGZmjtL33oB8ycgvZANP0n/kppEWDD+4D8XZgvSNi5Nvmn7bJxZ6VoMHFHYXHLzoh7uGVupwWpAN
/qoH/YhpmmkgFPoxbuQDH/1y/jbzypbD0pSPL7QSvN2S7BV/V6Sfn11UVdQK3srxBY1IRYEeLirh
BRf5kDAJlnbcH5F9tGjM0/Q8WpnYIP+zs3paB21AIlcxjWcdK/QB/pze/XaqFsGMlRLOMc61bGuh
z3gDA9N4/H8Yc/jljUjZYnjaKmfKauHYrCTgBnU/e8L1+qbIPbTQHbm0ptlRxIFEdnA/YPbpAKmc
BYda6F3vByOr4+HdnoE/G4Wr6YZxKl9j/Imb3ihsYI57h0gMLCnYBQyraty2hhBpF68FHY04c9gY
x+exWcGZwsXWOT886XCrg2rhXPAbdLxkGGNvdaOMebGQj0p7gsHsBxl+6uTgpbiiT4RW5IOu2pG3
tYd6s8YZKv4r+UZ9Am3ur5N7JMkHpuYD044rOsHusHylMqNP1iMQhwu4TOt1sZGzc2DZESsnxo9e
IOAYVEErpll8h572TpTqD7ZjUHUZ1xN7gZvo0xnFOt6A7a+0YhMYrUNOeKPTA1x2yvji8ID9ytIM
wbtAgu+BCb+BpAWtcZVVRQ9PUR/VoP5jGbaXQZfVwT85c+YxWEJV1BkyG8XWWN0bwbKE9bgxVWDC
+5vOrqGhHlv0OnFsbPWf/EQrRJOkoOnjLYx9TBd0tAX4aen7f93Xp4Q9wr2u8dlVt7ybZmBREofh
XCi7aR71IcpX57v8bGWYS9hfVzuSZDsT/b8QMR06X4AQOWeKBTZPBd2bJoRytdniDq2ldM0gbd4t
cbL2EPetqaPT2uPA+n9kq3Uhe/vOXb9D+kKqO3psD40lpoAFZFALO9gAG5hWegCho6EWIwSx5ONm
gWEbuwq0kTvyd4dLgcZZ7+BAuvIfe68hFh/llZv4dmBfq3y5pDA8mDw5VaqZF6NxcKA1FBNvHsmA
t+/hV1k53IKzOXlWj+k3TKbHmtVzL5Q7uVzgssS/Qd4hXkGvvEQq3QeLBO6O2gu7zBUizZYJey6F
UhtLMqNuDtHvCOlvkBA90soY9B6cF9WEzmnWDtwxLACX2IUYXr4IgW3TdLlMiuwq7S3oCDcO9kyI
35oV+uAe/ykglhzidSqmj/6ZM1Q4JzQht5rY7TGuHtaZiQZdknJsahG5KLJDRx4/AArQQg5I2CWV
vZb2JSsEAgA9Sxtv3qec84X/v2gQTJ/i71n5EiSiuxOhJUrd3n1aDzRTxEw0c9Y3K17IsJf6lodx
+FJfe51EVmdMJQJ4if1vylKxr7m6beikgiOhym9nP7xgMtjuxFN+to+3yguxG+W0s7kPXGuTNsoG
X/BiIB5qISLUJBAYjhlntTR9OGQIzw+4N50AdG0Km6x/LIQnTNiD/pY2xBuJ6MeMoNP6XGuKfWM8
R4n4PWwPrRUEA14kZrG6m4ySFVZZrn3w4+oFjTQ+BvMw3U6I5B5GiHO8twdBx1Dy9RZbYrofkEVB
QBLx1LwzDeBRcEujCK+yL27K63aoWH1Vr6rofvtptkIDAKSIWxemwsu71bkh/HR7Kzag41O6t1AA
RguwcnwyI3cWYcOxePK6YXhkzVgIXkk9b/Wf6KtYXvQ1XTrF+yhz5ZfZXMNE6ivGhtUj7yT/8QMt
lhoyxgbv/Urx+epKj4Vi/ErAYwFuZfPcFG/fAnzSTOu2ej3qrs8ZSbUKxSP7QcGMypKyYrmN+G1I
X6ntjxQWpnapYK0h211vIbkHQywSPu9rdnWHVpP7XLIEHNrVBg/qv2+7Plqfbh2eDp2MOI8xpzDi
oSOqNtdltfKhy2uJ+N5vJ9NY4KUEEAr18x5/knqqnq8h8AWoxK1QjeBiY/pWDYDe9+Mdj7q9rMgp
8bS/GA2ZYyJcV7nWvAwSqniwjsCcsUOwmaHN1xDzTKI2xemBLsL01PIkxaI1m8Vg/67DjCZ0XeIp
bg5J6i2izk8YmcHx0U6d9MokrH5CEySe97+WtTR/bN6aC6xBtMaWbY9AjK80fOAYKA/rYfjI4ouN
cN57upQ00p91wcN6j0JfVSDPYzOQtf+0WfNU81vIGjd4XixRFvEkgKmsHTEgELi4QbRwIC+kJN8H
UiTVybxPYPuSi5gh36DPl2yqNohYZwtRnWAmAJ+BrLQWsJyh66tjRB5WO3oq8RlTlzP5KXMiTCcK
UzxDPLLe+b4J2iATOeaqMIXTUMQ3zZ1n/UbQ+uHYDvE37bEiAX+JXeINlyX1Wy6olbJo1c4UOrBg
JUawXuQSujlyXv6UkVEy6YdUR6aLnNOF+tKVtTwZJHAolM12YlRfvzwSfdDbn+21VHCY726nVNL4
M2Dwg5pjO3zaJwIF39DdREdrIfqZcZhRrXjcjOqQ3k84FAEo5K4vCZB/0Bsrg7eePusiWkXWthCB
9JccEIeCKamk8ZhU7v5fEFqrwxotthn23gec3EgndHHPEhskOMfLmfdk3mgyYEiaiZ/h5cbSfJTj
LsZNV7vKO5+KENwHH0gyE4WJrfdwq+YkjCUBaV7+mgjtlJ+yrOsoYXXWkAvnuVh2CLthp203HPOz
2u5l5pWUYOIDqWPY2rt/TabDnfNSm86MmgmwItHM/bJsilMklpnuj8pDUi/dNIL6BgNSPQyIEE7l
qN7uREYy+GMWaNSdN3AkI26tKxzyz5ABHIROqKJrDjWUx7R0rf2o7zJ+t0/5cIE6s95/iYOTXHtJ
Hc03W1GEhmjkQ/EDEBw25EJpYS72/VKoNsfSiAeSfUmr+y3ZbQx94AXUTky6bpVYQSm2oobHRkDg
Q+BHWafjP7xSxcAE+dPJo6i9Uah/MyARg/lHqX4N3mgo9v+EbKS7zjQsBYwd3LSfqoWGQat/DoLh
zFDvO2M+zBt7JAAab+HVtCNynhQM9HJIzMbkW+byl0t4yf/uq+WszNrQkScDPK3zrIrNfGghb5Xy
PXnO9Qu6yme6BT+n42fZMEflTWwvRRkCnokUl8Xt+AkZgiAu819z2vBgFm0sSje1ihrU8vAjXrf1
e3stg4dKLnTQLfjM2t1YQgoRUKkdDz9kZEH1ZN7FPkbku/6bAUIPoXiT/TNHiM1czV4XrJMdYl5m
dHqLYmaqurxpxvc6BCYcqaA6U+FCVnBXViLRtqusb9ILfhh15z0cAJzqikKXSteRHNyTEaAyEFWn
i39cBrSkms1tVFh286jWUp55MRnwh5IsFcg5klgMFWLDvJDFko7Tn7ssCb6o/rM/5cBwgjsF3F7V
cFTpMK5MvNzGd1WsP1OSYzo/uJf8sLN/chtmOwIWlopUVW+bf/9U47YhoU3qGqm2eo3gxtRfUiYS
Sy2XOOoQlOiBNAbA3+4Dor+ecVp8YIjQwX8yT1PUN6Kja96uFZ6tPX9dmwbJ++YomyjU7b11BHEb
uSGD0+hJWcuX5T1KXHGvUoszy6aZcF+1PFxjJ0TiAXe/k22EO2TnrPi6vz8Lg1acz4JqAPQNxQnm
HfKRzE3YQmUA7bNh2o29/XLGKChT+ptrhUANk7bpokUY++hioC4o+xx+dZFgr7M4qyDpklu7wuLK
WAn00yeP5pUU7YqZwSExZ6qSamCzmjZw0GZCxNj8QMDFaM/GeD6wGFXQ2ycC4a/8mRtm4wCMN8kT
fcOaZUDxpeMxjMfsJSpMGzVM54uamqT134/sP9D+w494ISM+10zBzOZKDJV+kPAIB2SlvMeWxeIX
oIX6MpdzRDy5+fUYIfADfvXVql+Nhue03Jfv35wmRHljd+uH8/T4TadMJMWvGZA4wtF+7DB1bFnD
Qw3D0psxWzJKL+GWt8PHHL1aE6QTh1PnsxzDbManGi1k0OGP4TH+81srbXosQtFYDceP2vxQ0t8l
RbE9PlGMxYEPGnKmLqUPmWNRhshOzhXWyICnKemAWhLoqk9O2vSH/QAGyYzdiRM3kLccQJlyj0L5
2vtTCPH9BEDQRWPlH68fvXBaWBHHFmNWO3EmqTsLFc2iBlRETmwzjdyhtGc6Mai9EBBkuGdMG3Lh
pC7Ng8Macl4r5zd+E0X7Tms1vgnRmEIU6OYJ8Kiz4+/VuSkw/fAmWpiXP4P1R9/hL4tXTlkKlval
GVZifN2A13wYg/qkyRv3aAQfmNHWDj81EPlmmep4BFlbq6FpsTkYFSYNUWHFvneGSkRzxcav1glN
by0QXajMpUi4gA+SuTbPbZ0Qi7H6u5o6vNaNtd27ExpA8fogQdxGX6e+I16XIr14RFUTWukXOKA7
5spzOpJ2ZJFkc4CeAZBIPtSnp8pQLRBCriI7DW28zMIjT1xUozXU6gZXx1GZH93G2BccAloyVHOj
qBQbm22JK/ZdKGczDxkmJQZkscmZM98OVpMMGl/kxldg1svnxVTCHE1On8KRwUlQPvycVU+5mG0R
asRxAWqQKx8fncQ06oYrtjhEVUfyd+tg/qLQDsKVxD5J98qHRaSr5deGJzSoaTEC9V8PwhdbGwEH
OwsacpBjTn6tUPV/UEtHUQrIs2yijFvgqRylKWRKZVsCWZVAtrFDJaicoze+BQaFwVRnQZwhco1c
y6YZaO9qGuCJYE/Is3MNpZJ2oE3j7bxS46Fwa32YjvT7L9KnHmnEOkZHKlUNNh45WYowxcQjfUZZ
Xe+KI0wfwELspYOUzpMuYrde9rJnU7kjXhqFHeMfEBM9GEURa9ZWefEO17N7B3thP6p4iWtos9iu
ZpiIArjcFiWJfigtrN/eTfAsYDD8UPAy1j9IgAv0HemnBfKWTdo9XwWtxNj1wDNFd9/zrg9pEpw2
oiYTHiFKu5DB5Hhshupr+hmce1wGpFypGTz1AAh5YSDOnkuDnpuBU2DfkL/XPKtNI5GwB88oWFnA
YZUje/ykVX0NP8qba1rTHDmMyShHT0mjPb0s5CtAFMadX2+oZ9OQemQAa/Z+FmHGQ12g0Zlaxrbb
fCdOO7iZTdchc5n589qw7i29rWdAElPQYcIprz09d8flFpAXqMFJK3hThJuKE9Mi20rVHvWQrQYa
0yZyZ49evAvrCTykPjqU1i7aQ5VGd+15SE43itiDR/fe7lRrKssX7pAhKwpoJ4zptCiotqkFUqsm
IuJX98sxH34S/wV+QY8kIqdFAlRJSVdIAm6IZgoBTxx1qEP6Y+sZ7nAKZU32qInlVswiQeJZf1hd
2UnLgkz3cZheXah0CoHVV3I70PszNCBzDeBaH/KQccnc9RaWDNxe0jO0ndUot3gMdhDAqaXjZAay
jUGaqZqNJtrHVVaxCu1zhQ/OewfCEfumi53oNzKzM6JvoUpnnhyy9T5/jWGj5zgmyoXFV81gpW+5
kY2Rbs7RK++hat01vXhpjpeYprSpLRujuz67f/J5Iugm9s/KLoxBHTRJFnB+iiIt6zQSy74MwhNo
8J/zXPrtA79NJgkoFqvkk32JmmAmbKni51QbIPIE3B2GS+j0ANV0N57Ju3cosQcabyKdiJhoB0Cg
+AHqCE5W2G35fpieVHfA4myaZ1PVaaF4wBO582ftgZaooO4Mk0Dz5Cp9Rn6KBWlLjKS5YjjKrtqb
Ju9Ox2WM7+RdXbVdC8fZtm8wCOYWAJikhmkEw5Gp7UCpxtUCxO5/jptv7zASdY1VEOLIx7sh2zZw
tzNpO6B8yr26i3c0n8Y1lJQ92ACFeELl7ITGbOaYBwl3oHnXnvNSiJt56PwbF+A1PZxauva2TrdI
dARBUEiW0ef3UR3hkyatUU6VYdP/x04YEuhQN4fvYyiCMBdEMMidH6xjYNrDk8gz22ZgeB2wxaE3
T/uSUtpjgJaLqs28zgd+RocpL3plx8f8dgKjBtbbc5EINic2cXpJpxjybRy8hevlyRqaCxa6N9Dn
oK+F+AZItgQMrsDBlt++h1wTulbIdkck36/G9JlIcSplGzEuwCMtq8dA6RjZLFS1aESzrW1gTau2
yz5CaoCNgwA4qwBQo/YESaPPFMOxVEYutXykwH+riFEBsbNit/TcNSu7oDYseSmvhNRcYenzMIjA
lP0XqulZw0b1fwcsKv1W5bSSJXQyH2+ZY5TXFnZxKiSiVrbvve/iTXWZ3zXJSFuYxQU7lpTzEUVO
ZuYSj+ueOdEfel1hzK2AkDfsNRfPsDjJRudsa7uwiPQ9MXCP7LbCE3I3Vsn0zGcE4UvvWn7p2Ws4
qyXn2oaIN0+ARtl3aX8eZ1qciTmHH8O4hdb7G41lVZ8w8um1tZrnPeHyeD8iZG4zfCA6jwczrr5p
X/6hZFb69ulhjPxlcP7Nhd5kdnhxPCAXzrFbLVaC+7OlixnEMxMv/+EH2J5HO68h0TzQNUZ+udK0
QX84xHyhJPxotNfYu17waY2EYflBYenEInhTUVVcYIAYksiXzSuVr3x2dyw5VmRqGK/RK6d2n3L/
cPV+WmoTV88rvRxZlQBUtrXro3SC5n1Ildfm5It4HFMciWH4ge8sVPipnXOhPl0bhbgxEuc68S1B
lC+oe1qbjZLnkqwQTW6BeJq2HyjJKoUIgN/x1uh4z49IJGGNgORuq/uQ5rheBVINhU9UU/A+hWNY
QTL+/cAixc6Sgp7cNBMdGDg4szayGpwJwf0DkQQ0D6WTLX00S+RHOSaUJQ2AN+Y/wKclXg4B/vyh
/Q2D70wdZzAOPQt0Qp6s4pWcAFMc4mYiqmC1MHYReY2U3BozAaNjr2RxfXD+vpyuTMgdW6G3o1Q0
4/9u6eQxp81L4GL7+acFN+atcGEavFZ0zVrpzBhbCW3o5K0DFzIrGIMUw9TC+Gg+Y04hC3+X56jv
kTPZ2LLlknQbjgy6unQajPh85qXAQl1sX3ho5LjOajT8Gydsxu9RhsaX9GuOzfb9dROH5chvr7xU
jOzhaTEZZqagIINQSIKCaO9dAUsS2a7vJwfAXdLXvC9gm5jAgcbUr+MlGBbXedy5+9tAbtwgiZSO
8RTGRlElGGNOZfz3rsNahmhJq93/LXJOREQUnI2ejND6MbyjjCX2bEF7BkeMG3S8w6Wf6Huji/Rl
gna0P+R2ZxRX73Z4MzukL4F0IQuMD0LlG2oD9LzuoPxCVHHUx8I32Madwtfweevc7gZkLV5fZ9Mj
aTY645q16yRXT/cBhcotjNDVI8cwxW9zh0M2TipP/HXhozObGEkwtny5hYRDYnZWy+1M+wdG6MI8
RjCEqr6qAKPRThch1l+1kp0tFyj18T3I/Mzw533vzOiJtn591wsjJLFz67HhZwucVday6KBYsUaf
MHYprizi5M/u8ZlvGkZcB3t8ooPHXRN7zyq7oQFTljBOzOVYE9szp9agUT6gPMbN5Grc2m35UoYM
WIxNPRP4FqH/uQIaIn32vJiLe2flx5+mlc6GZPIAH8oCgJoCyibPl+M68/j7M1c7TNvsTqnf+CgE
/KAjH4k/1zJBu0aIbpN1o4ZEbYUbn+Q1QUEduj5YwjfcD1He47HpYP7NGTxDL2iiuFTq8D6Vaozs
UQyxONVmHxpjYRtSCfAXP+7Tbnw6zNAg/y7b8nL30sivYhRL3cO+7VwrcwAnSUh4Hyw1IHN2Z2Ox
dxJ0nflSFLmBGxV5OBlkbbT0/pXhxbCFqWH9jJrxi24KEiuNHP7FZZphEVe1g/hy95hXaQoipjan
JMm3dJvxrR4j3CM5bGvyou40zDSiGc+D10TMU2SfjAeB+yRpTy8uTa/ka8+rUp0E1iSu1pViLsIr
QqaONaUWyGw43rQJaKVNmz0Rp1edgclczJbDC8FAY4nhxirPnHdDPvRdKDNpPSAMTDQTXj/94GAJ
j3kn0Ss5giFDHq4wh3GF5rWviqxKJ9wRwUFRbvKz1/SGIIjc5FNofI/wvz383x0TSheIotVEtSZj
5XJdOGKhA8yVe9guxnETP9ACgYCmQmlROyd10TzFy3J8HTGG986FIn/otWY6ddCbBTfe+IP66Qc9
YwNzjsT68RytdVQPFFpMFLC3YHyZsXKkTrHb4Qtpk6DV/gQNyizXLcJKvKsci16YQB54d0Auhypi
GWLMwIrSrolAO3nsqvySQPYTD2wYxmAZJCucUglLS8j4N34cM1m84aOijGXmIqVcUP8xzEsLtoWR
107YW7mEAeVj5RCm9yOnbFyxf3AIZOA19Hk0k9PNm3CKgVff7QmPZNpNcR5H68sZz6hS/3Jd9epk
qxWkromqnt+UCwq4hP123KvkQWym3Gw5sLlPO2BGZx+u1IM7W6Z6/rr2fZ37yT3DTBKefizQN1we
Uk+SfZH/rrGnwU0JUy8clhgDhVLaQIUvttww9rv6jTIrmm9tqQquFeb55MlegN+GKbb1u23FQTUl
ao4ro59KIme/yMjtJNSxLp5LwkYObx/IF94wwPWxCvfyZ03A/2kELb4V/Tp8Vj7ESAFUuXBVsz8g
sJQP9zsBlT7t5bv6JUOnhylKkCf7gehR6msAwznMy23NMsec3MUK+9o6iGq543mn+0h7dE0V3PdA
rmPnUcC8+xR9kpkB0oL+0aI6S7q1kHLY6eVVNidGlZXvzO1AaXwvPb0k/+caqvIpvqYvEYJY3MAF
krP/QoHL9NJn2Ij+dlDU4NaswTOUnOFE2KND6fP0P42EO93PqFFy19tkB17JonXREZXZBdJQPMKz
VWn95V/xWVug5xeg4PgGsXUIy/HpI0/IfXaN1IllJ75JdOnElDPGlFxwTDTP7UKteIhC0TW8+G+u
dYkzeTDt88TDtE4gbvWAC+EvLFqIlE5uFNs2sBBeBfm1mgFDfqSIJsMV08swsJMmB24MTXb5zBb+
QNParjhAg0PK/aMdERZtaQrchGjhJ+n9LghinHfqNBrjhJh5eLhv8I23AFhxFtV8VrI8HtowVf16
OcQ+cIdNlZAjTwDhFUyof1YCnAQZhFAtkKIKzZBVgReWxpq0locGxfjHP/UrMsgP/fjAdFAS/6E3
cURs7XOUAkVhiwDage4adbQ6pybwfNPeoL9VQ71rhe0bdtlkiiB2/3gh64gilPgKJRCwYTN0EgfB
Vl4E4jmxUIQfpfxL1jNiB2BW/yR5hAfVI0nyXsJDxyORKvTKaSnaMoXZ291pJYEFwbnf02YDdAeq
fCOTH2UZgCEhtK53yrLvbUDSujQO7DeuZ81dZobylSSfgWemhgO4vo1eGN3Y8R5iTan7WE5aPm1x
t16ufNWIT+WuG7XppbSEqna7aTHDQts0cS3Rm5OA0D2BLF93U6w2qAHx8aqcmfrqj5l3zVSABKu0
Mz5HW6YMBCwquT9ZXIp4PM38z9eyCieeXkyIvFAfd1cQmulS7ftA0mumZ0vI2SY5+VeA66zP0Uyd
h8E6ZW/EsE1RNJ/46bKNSvJ/WUKH62mBeqxX2Y+bE/0u4xyDY/sKK/1nLBfgVlxEKhGtV/ihNFeS
6X3CIKy9qZ3IWdnm22chUIbRO5MB2WrDiBS9+Je3eLVgkMsn6an/4Vu3UO7ZtRFThOozpp5anBpb
/TCy9sgsmiKqgcTMmJXNkCQ6XLW1FQKiiHg6y4H0jCL0oy61peQIuSJTh4bZirz+yzVDfllGFBRs
ThZGGXihY12j8t1BEbHU5PdZgn/Ja1DanjOemBsVzFHKKFa0ZmYqgZx9j2jWA+3FakZuFT/jclcx
sOmSfvS3Zp8gm6WiYA7iANQbCuf5leaqOJhLwNQitSk5j27vWrj6omMXEVzxB8iOo2EiNokE/j/d
vrjDFHcwSCDpOKyfMMWSNOSD4nSc0OJHfc8rsweVLyx76WMphLug13nRWmwUu6UkfBkI9GNvutKq
biZ3MmA1c5E97z3GxGedUQZdPpGV04dUHGrXYjkrhoe+ZbVJx7tFi02m7+NZna63P4QV588zQKXd
OtBnFUxsxorPoxm1DqeJOLaqmgDnLwWKPV1nmCJLQSBJMDCcEcZo7E6EgNPACY1Im8IpybQvmd4d
s/ZAjyA8GmkJ06P+V1lYHYfHFQk8KYPNY4a/p94ea5LpvtD2luhCNQ2VF5IC/iiCER2LAXpejyps
xG5yxzikiZLDQQhjNWepH9t/pvKYX6vTNg4v1P2cGh9ciNUynIvbPKTlMN3Auh4FhXc9XWb1Hsa+
pPJ+JqPR+yWLLKwnVXsdFD/3EPp09KSue4LGVP6YLBx31AK4x1C6lecqD/6PYWxkYOyeUz9P9Cib
A6wFhwfhYqUNwULGEZQbmunVYQ2UqxR8iX3+dmNEFaCu8uC97Cy4vQWGHtRWEuuJtRe3tD+AVBhh
cTGdzFh4FYNVcSH9Bu7CAwwQug3ZUcCVl1ZQ0wV5sczK0hOvsRD6NlE0my5u8zMblPhAS4VqDznC
cQi/pcMJ3/vD070qqNvi+VObMT03alnDJqN4eaab9aVxOBHq3AJzcUM6Ap4OQk8wt6eaGuMj37N5
7vZPINiHBOuCh8Ry/RERYbJB0Kyjh913gRtxwHrxKjwnK6/oVq3cX7nHYD/Gb0N8Kh0h6qsYGf6C
bjsqh7F6rXE0zAYP/G2iQWQa01zHgNY7A8oUOH97kvj97BY2Hd1BNp62AmsX5TnWgLnGUFTQquj8
fRCcxKhy2TARdEkXuSVuGruTk0qWY90rx2ULPqWUTq6P2NU9d9Rj9F3XePTP04WGuQFRkbWZawd+
DUMaJcxpgzGjNoKFL5SpHV2oiJr0vgRkrd7Wtv/M7g9n7aOXThH9ViBNC1LbnNt3A9Fnh3TspZ0a
kKtQrZ23POCEhgnn+WGAk0XnNG7eFWBfpAOlUtv12aPrTg8iK3Km1hXftso8VJMSR84KyaZ6dMst
aRsqqaNIlxLxW7HUVoAy/76uoDhXzpco3y4Sxdp/LhCFSjXdnAdE2aHyFhcyz37Im3yMH5PcBtRC
8GtDFJAutCx8sUZdltlyf68XW/ox0WeM9qZ+9KD5b5jGHjfllBmJIqnyaVufPimB8zvcFv+RaZ+G
VqoI019oVi4AEzr0FZQfdW1KJEFtVfpxRN37SqUg2B6b6Ppj0DwL747khT5t6msmOAbtAutqWssr
TARXHvxHA9IRebqfPSU8Pc6to5ffg10RaGsZ0STH58Z4GDIYyhFIpyY+xdNoBKD7rFQWytDNwjZB
Xun+oMkJ66dQdKyPZdeA3qqAvZtH26zuZ/jNJLfrGI9msPP0ElaRWf2M/K3EXDI27+krm2U9AEt2
AbgckAmXkTIkaZ5eIqwJ3EwgmkxUnkLwrwDB9mqOPPte5jmDGabVuN8z27H6sn8rMUzKM9bM5irC
qblW93zLECnebKsNDPT5fWF5L4mMFt2QOFgICnuakHQFLI9jO04WGHQT37NjjXQBisyvcF17/l4h
7pydNuk2+4TDvHktYfDnYUxycF42/chhq1TyLQXMJ3dX/H/vqnTRSjft+YvYDKrluYSWttU579Pf
7HgNYjy3v3qOdCXZDJ20fib77kjvw4n+eMBYBmi8C06d721kRBHEgOP6Zw5K35gQGoWbbIxVVk8J
pI9f3ZMqDPZjqzJUB+ZSBbC7fS/5beNpkFJfxDlS0iaXVzxnTa3p+aG0jmBPkvliYnBPTOB5SccT
pPA2g7fCCWshAia0nvTuLTzwcpnIAn9hX5H1IsXDCCrM+Z+5AmSlUTuuZDWINCKb5TLlCUyzAA1n
pAS9eqFB4+6zXQOGEV37OXzo2FyMf7B/ixwpdu0MqP4UVDe+Wu15FLNwujG6mLEF85b8m2BP5OYn
BSVC7ALygjZlT0SxhbuTcz8NH+jVI0XVxvS6wqeWou3CgEFNpU4gzeGX2QFTiRVAY/grj5yytojy
pCY+x4GyMcJ4i8SP+CwzKGrBzGM7Paylf4cdYVMC5ID4hhjPM2qSOPtDVEM1/Mcww40mlg9RiVxg
VSJf2ZMTsAeb5flzm+9y2N/9HR5hdtGL9KhWvdwkR5/eIz0R4QhyXQX821NxWj0g+kXmTdbtLpDx
9crB7R9v+yKNW0EzOzkpVrZgixtYFh+yBdacullAnlM3HnxYAH9OSNGMUxQNbrAsW599I8NcyEIx
nUGRCrKMSz1FSTTQPMIgzV1IwvRQeoF1xV0498mnzi4/BZz4eIdp7TOvoxpeczrecht75GAK2NEA
+MdlaaMdsBxqy/nnhrwC08VA1gIpf3FwhZkNXun6gNEMDX5z0ihOUOCqbLMWQco46pkKBh10L1af
s5w2c2jWc9EkpYJ9KLUQEdWy5hBuXjhue+TK2OTyP581nIC6stDsMejJOXZ91PEo4XAUiokehSNB
g0uuNaAxIMxtYGUuMuYH1k54uAy5MssuIcd1BPPUNgCmAmuGJKKAGDiV6LDnlhWoo7R4SmyEWicf
dvw24yl5+XtfuxJbhqoyDb0NjQUNcuTazWwG5C6Xwdgg/2WJxAK5tkxVp/gwlqGKLmVGRpBXB1hU
efL0NPqOtXhWFNJK3Dlg8X08O0WK0MprIWcR/NkF+gXeLQd0LiVT+QNK0eA4LK/wMc5LguXKk5Ox
kgd6joWR3Z/PB8d1TqtRJQitMTxFuQgOikdA6G6WNesLjcSq6gEG4rlMOSWuIxNW+ZQ0OU1hcJiY
eDDu/yloWL6jRe7B2bOOUhwYJ9lakeu5Y3UPckTGdGatOzCXWA+uqMgH+dbpsLYa0XSA9uOvBBAb
C5Fw/gfMJtkNBZWmesh9CPu3psZHCganaz2je1HMtKHBhstYyh2RcFQqzp1H6q+TdP9RXL7Oy3El
/Obb5X1zpE+XnR1oN0yeqxeVg23skuKPek/SFUfuRZ8BG2UVZpoAsX42OXmKatJh9pOYkrOijWY3
TBvDtmE448sZ2olp8/zKPRxEbONbNCeTIGH83qh6030cyeC2/FfypsaGv9yxrKaSyXHTiZAcBY5F
mWVSdDowAO6QFk2GbJTlL2M+NLeUOudxYVStKfycBntiOcpRnhwDOMxykquud3hx6qoTilhU1BtN
RiCycevR8oTm5splvVKZBDCCXAFvhMnkX8D9p1GjqmwisUYGFKSZ0ei4O/o8J+b49yvPVgSpMc3T
4VCEHXH9XVf/n7kHf83UJFzkLyG53tF4GTFqsr4e9uhxOMaX72gej0F9rtH0T26V+KUZHqqM1kz1
90n9/0BUj/Ti5FNXmzctInKwNoQ5lLAtEdwn+ptcHw94HajhKFjYiLGdK2v4/ol/W9eETkPDJ3x5
wy38zoxAdunuoqp3A8YY8fYzd6+vNUr0UJ5m5DuR7c5FpkJyHXfFrIG24Y1Mpi05iSISOGMhSAH4
rRQxd6k0OPToVqoSCVXQlAEToMQOuQPj2QsNwJ28Q8wXr2QBS+QlYrykUAD+vgtYmQesHTbRtFya
UQYUkJCFGlLSGAVpppG4XOzdpJ5imKM8p69VWLIAwYv4ns30D1TbXXyrjpOGjTHYubLzlo+Lbklr
FAFeSyP9kzgBYKaWH5iIhIe6VdllL2w9krJg3d+Pr00a1rFpeRlzStr9Qt5JLVK6BkBgdH9RGr1C
MTXPDKUBdXq+fwaIUuTG7aCRpUj2eskCxMiLkJ2L8hqSCfzsXTh76nO+Sa64AWvfpmPeUs6T5Ypv
92GoIbtj3teEzdMs6g+1GbJY+YbSb357tWpwXFh5XmHIOWxIVYuwp//3DFyaHoHKwjAYhBPZGDXK
endyytCbRVhVSkAWmuxtIHtnRp8zbMT1lxtojULeF1W3NTg7WbSBGuGtDQvboCf+6bJrVYCrY8bI
ph6NA7lUsT+aS84SYQ7+w1CKjWNEJ28oi12Kdjrq5wzR+STCBU28vc7eiNRfmAVIffFwMTambBOa
rxQTED4L0n2jQErVpt+Wn/0JggMZUK85uvoY+rkB0EEApB1z+cYYHoJGNZGqCflL7Jkr6CKgGwyA
tkvyZ1Ljd9fHwWc5e/s2TJEFNiHvjoKBs7p15dndjgyJZbpRTImhiuE+Qv6M4tQA3m33/e0c22Um
q/GtsRnzOcsx3tj8iKuTuOomgxHPgoElWYPgR5Kg1+9c3DClRFOCJ8iTjTgaV0DHIgcLEs3yjm8s
mchKJl39RFCPOnTnkBXsu4iWwiUP/hpRp7Fl0HgSekwfTeVkrvSXS6CsQzu2J4bJuOg8ci015rAx
nYd21874hC0g1+j/k4jaecUsuXmz9kLMoirgbJhxUsnQa0V7BfP/y+09pYUf/vKbOWZsWaUlGgEm
fO+aOfaA6lYuGF59LU6bt/YqZjyZ1Wm/FYX2cAZz4FfIb5LxkN0wsFrhcXW+wu6fV5IwhEOQ7r6A
J2OQOouXOI4Codq1cZhQtrjpmgRBMew3KJp+ekKGN97FXUg1YN7xGM52V2g17j8E/rcicdKqMlVk
sMPZjkNYOipXytvuqcqKG5T8z4Y+YQ3n/VYfroeLmH/7iuwkx13AQpsKFEzZXe10c5WxOHdoumHa
BbNvbrI4zmRCnar+SJMSksVzT38IdQfH5c/u+7GBoslBhIToJaN3WM1CsP/c+r/T/kGmga55653w
L3T6NWUoih61NQrJ7rEYtcQQB8/61vQrEXQFue5x3rInilrT3B2fWjgmcSYIN9LwD7bSeC9wKyDJ
Kxhj6z91/THODhMDOnY9na2mE2ZQV1Y84RIhZ/NVF8jciwsouFVnboX3Ovr0j+i1a77BsWkHwMUn
RxY0XLm6kLTClHZDXd1AM3EdgvxwiHKz16qA69oQgrunSX8rw0VX8GrIvTLp4Kv3hFCfgvGgMqp9
zMr0MarrbPjv+vdPOejEmAi975FHqh15igncrrzf6u4s1u4tAvAw3WXLLCMM6zjqKHgZdBOk/g2/
7OepsqxSv7YWrI/BVU5MMi7d3a0qQsEDv14k/ScUI/CTOj5MjRjz51OxI6XSPGOnSUE/yPY9+Rnw
DD8yF1hmgVVwi6xvkh9gEGse1fDaE22w7WiMHguOnW7VuSHYfAxfjOO3toujtCjb0wgIbPI4jt6p
sU6rB1opiSd4qExu/PtrzmmN3V5ITW/2J5GGGltwSpQmvuA7RU7ThxNegkqW0X+0QbFeVieyaa+7
U4Que1o7iw0tcZKrqy+B+ew99k8Lka+QDWPHPsdmCLLd2T2HnpxDuSI5dVZLDkafEYMjDbMOASGl
zQVB92ds+xv6BhJIIbvi9RvRZspHRb2TQ5rq5ZWpcPbelpk3LO9YH5AeF0PQsXvDwtE9uClMrunW
uxqV0ddQ6cjdsafEFcJvSvfj+wQDrDneJ8Nm8Br3jXYgVd0uMahFw8PDLTgDnWL+95P9Px7/1h0g
QbhB0OnlPC2C04l1vn3Uet+O7GFlnt/CgOdTXU4Oj0pRReqG8f3NJsvvlIfA4eBprg0BtOKMYjRv
i1iQR1xdaCofo0zmo06sAKoD9awTu5/yswEvn5ewWEtAkUyYINsKJPlGtNFn2nhhyt0A9NG9rAiB
1aq59JWfBitXEL+FiR05OCcJ4GiNAWpLiDrKik23PvmWB8OG/temlKy2XWonTVuro66r9sXRMKss
qNqhr/pqESCWl3xOhJyWjbv203LkGEvHnG/4x1mzVUtX2WLUxipUIfm6B3clyl/KHNEBd8TOB8pl
Xw7aTvRyOAwCtZMdiWH+IOZpwfao4tgthEf+ZEhV6BNGMPhbessMApx9GN3QEjNTHcqBsAxVzJiu
7ssrn+ljekuoBMZsObUVhWc9wFjwGI2H44XMAeCM684HjoNekMVpif8JPNAcOVFSAQapZ5fdG9AV
QAWHqKgPIw+8OsJT+4vhnCcqUmdVZ/ZkZ4fO4NrMX13lWlBr4fQNGFDaFMaclbxtyIcRZlqC/884
WiIgUMAOa5aAf7l//TpOrNw8oEhGjPr+h5iHMUQjHZsbgvLIwahcCYz+v/dH/Ijb67/hcYLO0p1k
mpYKmUKo6HHnMdkAFcXwzDrY5Lek3SYJxL6+83NaUr0sGagrdTA9cwrWmY4UgfezKqpy6gizRr+s
Vkwgv1fRCOcWaW88voB/bsk1MLDKCDK4GVdTHaAPFR+G8rUCn+85tRXj5FSMXD0Lex6n6t6Wv/pi
7L8NEjBmL3N2CgBcCqipNqisy5w78637fpydCni8KAOiErVsqJ/L4uiTOMalOA93tkhC5hCGfkTm
2Vujh8fms4dtkLktLHtgb877XVQDLFo6Dv03qQTE+dbfUu2cbi/JLQhSCp95i7iGkgoD9VhgzZPe
JD4Lf1UOlRuwEDQpWjfcKD0xdyBrTC/CNZFP3oUhqFfPzhMB390l2fo2mqGCC35vYpmZ21lkrYXG
NgCbfYNqXkCsMeQmJfT3Kz0R8wzHGSw3sfMPfeURbp4WJg9xnFzHC1eXUHQ8oe97ZYjR51Rk6HXx
SFnzyNbhlfJhlnswrLZ5dqHckW7tRSiCTQpg1so6P4tfgr+NpVCZZrIupsxx8jR6mvxDUuCD5rTx
7ypaKa1xd+x3lfvlI1G77gsGZ7A2++/O8eGj2D7F+mpZdhyg3nPp4JDjl0nCddUFcWfb/g0O07d8
UpXBlRKAiOuqIdM9ZAkxaulH/7n/9MIDptYjLCWvNEKuBW0VZe5asrCf1eWp93R+q85uwyeewlm8
hXZqWOowooiF9z24W1tjsGOVM4+4UD8eTm01mYWEbQvnxiZcLVbIAaQ4q685Xlj12ZwmbxlrRxvH
jj29ygbe2yerWlKaDn5h6V6iddL/Q5+voqVSPmEy61i9dFM75HEU3WXFRshD2++Jwb0AyzG4YZhB
J1LnLbDjUgn5LWBVD9bC4EQMW7dk2TG9JPJKt28bMIHBRE0G15IWIw6TbJmFKwjaK+1hs/k+mrwj
WTSwtaudlrcuXAl+XbewPsX9LJebBs5d5TLJ8ga5psDQrHiSzE5ulpKbF4WZpmu9H0HZIjaBCu75
IlfONEsrg2pcryWorG7s1VsTHyNWZ1XIahTXl1Z4NW5/ssowyORhfkHP4FoGNOibLaatYF/Kyimv
0zHXWPNBf0H214fNbgsrIAj1vhn9k1z+1QOydycPhuz7OVFHRpJLgUVRP+EgM3B22repS88emujh
b+223ZN/3erMr2gEQwVCsP7nYLZvUY6bz1jSDXEXS24NY+b6Ug9YUL+8m71mbAkg9V0CpWY0xTNf
qrxn2jGIefPOy7zJWofdfHoveCAPir4bqUiMqu44JfJSWWv/etP14r4zTVTcSzlSmAyplamlObfa
pTGLvonkv6MWBpcUziDH9M3pOqndjOcvevzepRGQ98qOETnwA5IvjskX8wwPqHiuFYhpYpJCIbDk
Zs9SSBBLxDitVWNY4UabJfiILYA8RpBolOyL6RmodoUVdp2jtsC6qOD7sF39+4CzrW65HfM8QGhD
W62h+wQXeLFc1ms37w8Hf7Z7CbqzNScZavelqFDgyvgIyt8lUo+itlaaCANC66clVW1j+AW9uGav
qu5JvKs2bNTiGt2SfI3HkPlqnCT/xmCtwn6kjPGERu5JM+7Tl5bTJD0EbXh9m1utHDRxJg3ax6Xp
H9IYQJdAUJEZwXiTPUyZdl4Y1ZPn/97K7iw7kxCH6CVnX0WzsxwsemQB6PVhB9am5jmp3XpqC2Ka
w3S+LZ4tGaxJQ8a7ivXHR6DUO8267cyKaOzDWv3x2VhQvmnjXj2mGPCsXBvX4XoFYJRnsGbPRRw8
u++sT+ojbEJ+IZ2nKpOtcb38wV4x/x0x4m+R+BUDGzAJ4lCs0zyR1+3lUzM9nOysVXACou5/VSlh
Z8Ky48STCGND4eJmpCZ0hcC8ODbFYzAjCWVSd/JVTUPY4VUI0PWn4NyJZ1eULkSJCyjCBQYND2Rr
T9hwkMPAfqARB0n4vzTTdq0wl2qv1tmaM1cjgJduV2XqUu4YujDDwZX0jvCNKrl1W6HnpKcgRAT2
+1p/bbwPGGCrF+udPthavQp+6pv27b7vD6dsO9U9pWATg8dSDP8wf3M9+JYJSJuLAGrukFrcO5f0
iBxdthmEh1iW6NweR6BXq6XNcZVmir9qaFa2Z3GlUxtwWtlAzZluzlhNY3DUh5wpIk2BJKX4CMBC
HeXrzc6doXzHdgK4Fdaa6DNadUtQsVMYjN0m63iUz7Agk3J1+KgFOtKOpWa1g8xBUivUvnHIJOka
C6JqkBGfnKgQtgM4uXdv5JhjMzGsTWZusDPn8Kzi4siro5d2RxGdgQidjxHTe44UC/Ta02lMSOI3
v/VXnHUNDrlKL7bdsaLMvTcSTWKQiI71qLt9M72OomEVlR5GvK6G6mfOvAwKfapS5bFjFrNV50N2
+uVC5+51NzPBS8nQW2M5RVWYBTZeVZvvKG8VhBF6i+fGlXN0GsoLukproWEjA7tDwLUYyRwJfFC9
YCfNODKKV1Tck5Mw/pzftwxajmZwWo/RtdINyuxVBru0R0vgUXZGM/2anZM0w5+DpOKIlF7ODrn8
5SZUxrEUZ6/C9lOmrIHJqaB6SzBGY9QluY5zT7hasHWBk+ibA9veyXsxIaRnn3grsy3jPCG1MC3U
AJP6vzC/Cc/uRkuQVCC1GCgaG48Sl8Gye8YRwqPX0Z+3UhsbLjI2HZ1Ay3evB7wTj216nRFITZiI
lJ9J1yLRvVGE1FkdGqflnQ0JOKqacW+OmLmBrR4CRbz7K941cnfdDO03K+z82jKc/9QRLuzFmdSD
OL+P9jOBiQS0aNRwd79GRo3U4z5vxoxK1TkDei73gbFBCsykMKn6KJ8LwpuOVD/ERcJWHfMw1Qx+
8l+xI4JrgXDrG8UX/j8NllWalERww322gfUQX3mt2+6/lGE0f4bcQK2kHOv+AeY250LuxPS3cS6k
cPe0KA+0T8CMZE6j22IKFLCATVpKCAXb6lCMYTdJRUMwzK42Q6XGItPSAhXOrvTMujbFGSbzHq5n
niHpKyGQHjMZI/1zP7LOhUCOgSBwUz8Fk+F94dRa/oP9xEOSOMBKvjCwNnNy1eqgqvd81Z1kUllt
gQ+EzehB+pmnPxz78X3XcHyvGIWMmSLCIXBoPIYcGRrqDjFNfHNq9YY5PuGBcN+Y6NtIuOO4VfP4
zTYKJIUBTZ3+7HevRhhZZAu6KBrj+JKBGoWk2ZMonMLIeirHjptkjFF7JhecF2iZV6xzgiz8bT1i
zXX5VUbdwGRSgN33/IR1+FOmWOFm7vXeLrZ9wdz1WKhH/Vlsjiou0BzSbyXLzFSOQ+YZiBjeCHWn
+Tjl7bNSiGRfPJRP36fetKHbRY7vrjGbJjxe5G6E71q5LCIdDzCP7l0ZeDtiP0P5FLpD75P/TvpD
+6O3aQ9kwUcU3wtOOuwHrrSCqMqRLrkqWmXNLIOz9Lpj8JAlVGYmnFzKNtg1oU4rAZHq0s8DfMcz
zdGhZTGh6150a+PGRjMiRMcAcGpGVSwBMkWHPjdoUlPJXlJPtNyg5Y8+KJeD2SGvzUdq7NmwKppx
9LwpeMEiDTOi5lNzOqGweH6T2bCJnhJbkzgmRiBnaASgnlyAvWQttiArO5x2hakMVh5v8V0goSvt
XL599zU5M1EQHhlhJdvpycN9KWw3gsix7O5enjd0jN68FSLJ2eF50yx1pQiq4xKpI6DyklCKaeY0
xpTLcd9uYkDmgN7Lg4cMM0Dih3FrSQJdSZ9mJ+Iq8WiHvle1kOlocdDt0BxbcuUlNB+eGYnJYvoC
O+gJzdUFZAAbGH/buuvSYVlkI3r6QTzr8K0AMdwfTm83Oauvju7k2oDbEPo/mq3L6Cbs+7yo8flQ
pT/1F2n+nOQag3BrbB8bclh0npdmqiWLFgDhZOYcC7brmUV1NSMCbpnv5lW99loiU/oRa2CbKbZG
bEYbcxIYKhyrCtC8PfcjrmEGs+RNiUnj0HAWB7OAot8ySx5yTOgHrL/eG7dsdi6SNZGPqzKNc0FM
pudXknn2PAqpP4b8bI5WyrIaSN8FubKIL5P48jTXWy9Ft+MJ7b+O6qcMVtqEiY0uyu3r1GlLttmC
NYgVrymtdlmDreMSKiFxEX15y53+smb+8HAm5LDyHIFDha681/9IuJK59M6pyKwAS4s5HUVgDqiu
87gbaWGm9t2iJfJIemEYkLYUFalST79CZtYwizkythToas5/qLqm1UuNPNPt6VQ/KAGaCeZ2t8jo
L0zTovae4E8PoYdm8AUaT//VeUX7AS5gIArLpWsuEltbTRm+EjNJaXlvvwD9Av/SYzhQyl9sJgJB
6d44SXPraFphibgr/1kNxLy/fR2LBxK0wgl1xqGSlL18ZlvvX0+Zq75ZqvO0dus2IPALpa5/sMJV
OXO9qNDR8GD3/7b81hwgo0Lxbu0F2iULMbsDGGxFFpv9D8RrpICwsIgMAruujYfvuxuLbuDTaCuZ
VrkaJ4xOuj1G92D1UDDSDdy4mfyA2zlFNSCkK7TC9hedlxsLuNSKTfYfbHYzkwZ5RyUfrL2/aBB4
0eZYt+EC5F9OxEGX9SNepvx9d/nf/yPL7sI85T4ivNmfIs9eHxhJVTjeTq60AKlK9nAOvzVfDoJT
wDzCfMwIz7SwF8oYWxsgsj+vBeQ1nb8/bDxai9UZUhhcsQZUFo8Rrg+Zd3sAYb5eUUOaFlWqhWZL
XefSi7Iiut4UcNXMdr+3qsxFhIZuWCSkZ7PFOUhPzof0farZSo7hvZyUxLS2YyzUVy2ZbmyR5kJi
+uozUnY9RJ3RjUuYiTZFV16A19l/JnQ21T2zHZCKPYBBT3kOsNyUQxrqvi4hPMtZECcx2y0G/UDs
I3/ZMo/iZniUaRPJ1jOTswipodX3NFrjebKx9pMRQfVOKHffQ1lD5/oSOixRZ9maqmaUb+WEfplJ
8Ax66LMcNXpMG/HFfu2HvuBc84WKkrNqlJLSh0jZaEHOf547n7FOJFtNNvol5btxgQkMEycvu0AD
0TE5SatGbPyPlv0++dzv6FP1qYWSV805WrCt0pr6fKfrLd0AmQZD2YDt0XZck5a39kKTWrzD69xz
wxebC0Tgcn5YFUhA3ltrd2kipIRxXog6UGWL/z87+kLzKEik6JNOInAWcLgDP/H7+TlgN2X8BNPq
5wgRMEa+ogS6YaOPaTg0ahQK2bOEbXCqet1Zh9klEhXdpZOLkwqY6ohXLu/Fm844KLnIitCQStIM
a3lhsqBMOumxo+EnJ2CTgOX7RKI0/j5/hgAezNcvpXX7B1xw4PkuuxDkq/J9Nx9t0aZGCtBreFEA
VIfshnCpoj3OWyj15RM7iiKcvCYypMn4Oj06CZsPXHFmgQKAUL+Y/NatrV4wTmg5PcJz4pHgvjxh
BUQIW1Tk2qFwVqI+V94cYK28WhuUmhIJ5YSNyAjhndhYXbD3/aRUNCNix0qQVe1HzXgRUrGDAjaS
BefwdxEHQk7QT0TX/ap26U7o7yRUITqGg34aOuFMyODIwxZ0XP4Wf/TNkF3adIrKgo2JMCIFl2eQ
NT21dWT9CbfOrtmsIP0lx/cXj1qVF0Azlp7k5GoyPqGJah7LJ50/wc30d1BaPenMmg2tMtyJJjDA
Q6OPFIvuDditXawqXEXva3iNpi4VZZNW/iVU6EvsOAHjMAHzXINrmtC+12mgTXXZCMJ2aKjiUpgy
CmXmiZb+0rkzhbyVgUd49c5+5lsAj+Wh86my0uekTdV9jLKkmipNpI2MUPN+fIsvqVR/wlmsn5le
hiOAIzhaGJctpb9mziTaR9cb6s5wWne/IItlFCGaHfFGuSCSOkNSqztTUmwQPHq5QGSSunvDci9R
zHwDL/MzKOI36yleIq7mlNPZ/qjbdNW/mK7FYfngB9chZe9HZxwdHnMPOltHkQFem+EG0wSYk9gz
p9TZ33VqyMTpC6oayTh777XJGs8s1qtWvoHnQVZ0ICmgQ8KcC2jU2hmOIg1zKR3+p/9Z11a0JANg
pXKzhsBwy/m5bY8NBgPvgDBeUD6kRV+FG9dNOheel/J+aRpDH5ccYf4uq+ksSiXCgZzqDn/nkFnz
lwLFwC4pJlr2EVbw559W7cj1KHVBs8oQqpsNg883YzT54Ge21EJHZCMNQ95FuCfPpKpfpVAke2TN
sN0CyXyvQcS6pyV4Hjg6JGBelEbhoj46yalj/Zf/VaKWoeW/bDq0vMArgN6S/1PrXmxDEzQZp7Yq
u+2dA+wU+mDdTWCMqh5jd0XC67jOBfuhLpWkvLkS4k76SBpv5L6pN5Ev5UXJROqIHTfLJxkKd8j6
fUp8QlYEF6SdqAb0Oy7bocuL2IQKSMqRqWauGZidqoYumhNifTHqhv5SZdg7sDhNsSZCUhjUgH9x
1OiXeEjaHIlM+wWCrvDSdgJ3jDfSZ5S5AoeX5hWlJqBlexu4wVzlc622stodlTJRbHciOrKmUSyM
MBJIsEu40OA88y25CXG3KxXdE5YIjJjz3PAkub1t+deC219Herm8kEAXXd+jVHqjAVnxGw62Nul7
v713QwGf3PSBk6hUpVCP55SQhlA7OB8t8CJql9s9preLsUsezehZ8PQI1Ogo4nSFfYppq6KgubyO
ntClPtoyib/oD9Up+AU5ul+/2N5pEEMJp8IPwXdLY9bSnbMlAZGgZ7MA3UwwWnhHqJgYJTgZOUmu
H36NI9euE1LTskt0X8hJxMAxt0QcZph3CkkD6X6ZJxvgsGyOQ4uvBrZ1O0dBprhiDQerJimUmbFo
tXmlVh6WX+40cyQfAKMtrVFFj8OC0yuQ4rI+njLFqXLvVYjswwhDJZQ87gLh1mQVqnqXgFqO/TIo
8ifvrXmOjDNa9V3EAsRSAmthhFLFElwcJxgAoNfAveYxNcx/orx897VWxY+nSSS+lGoRXq/OO4qY
pDPnSvpObnKRuWbhcb8801ecJYkXLZw07NDo7VsJWBmrxkVjZMWnbeQrK+R8HQyphi2Sjgxj4X7y
G3Nue0ZbZSdPs9jwC8K7NSfiFt7SwFz3IFSP8ldGc00fQuSFOwNFglpUVhKYnfDQcCPuQOCpA8rx
R+aCbLPfysNbjfSaXGVTYtHunG9Ixd5uEqpdBSYLmE8DVDduvb+w0pNL/4XIO8UkIfpsK0i0JI3O
8r4++H8y8zJVh48lYHn3+PDd81LJR1EwHtpLhol+bPKwV/VSxjLiVwWa+ky5gexZqHUQOPps5jN5
ZjXa3bQDVFOskW43z8u2fvOhPJ2pjPkDT2zYCZA+lT9ly85+VtcGx+QIi3dKIYrYOaK3t14FdkY1
G41cc0/8SpEqdxwbO82ndH8KEpef/k4BPbDyROE6XmjwClhXJVdtdeQCokd6+ur07pi7IjFipbsS
7rm5L0sw1UvR9PV9IVPsLiejaHk4ewOmzk82vNLyqeGEcJyrBqeBwNpKH6HBV/59XZ8iIl94VSPe
rQpPcRTEkMtoCsTkDK6mlFp3YwR2z8rNG8iPIb52eAxHt1lBAVOJTR2LNawEoL/pGCi7l/Yt/lmr
HkuziDa535kQ75yfd2pXpbJcLF3N6pXkgEVziFpE2sAio8g6WfF7pGxMF6+pJkiIuz+JG+aJa95K
QeVhDgCzTWWqpdeQ2Fwipa1ymwqWU7wTHDrC16wJewnLf0KF3ldl2qPTpkq9n6TqgVEgGsFXiMUh
RAFOEG/SOdsK7w+WJRuRVAEL13K1Ucg1Zosw0TZ9zD88Pg0pdb2MK+nOJNYIvpp4o3hWtmi1rrPF
bwHRXCmaUcLu1bM4YPrDXFf+Ahm0Tfyz/QqwsksbJQHWehaeKpHLmfp/LHfLVA7IkAHLq75JI8cg
rceg0qRl+GTKA6EscA/AuGtqsAmBRuUL2DIwyftbGp3MypfWKYx0Kon4YiyHTg+3e3wKswh6v9wQ
gDadp5ZTmKRXKcRGZ5Dyup5Bb4BpPmbXqrg/9QohXdoasxQwsPhQ4v9T0kp8qB0xP4cJMTGiqUBt
iVul7nr+aCVNt9GWf9QxYNi1nPRMKgGYWSxPJK4/IAce3IlJdDZOPKv+6UG+vwYpbJmWVmpi3N61
LiRZaqnrLKokOsoD6cfOBwOOEkIU6Wkyu6RgKzRWcjeBbC6A9zLZB87QQWCZuLfs9s2hDfr1CDF1
irqWGRYSGZtrdpddyKlYopQh42OfvxbNdkhBKrJCdRdrqIyNoZE7IdQ4forbb70oh6F9hvd3DB3r
I8g9av1id82nteM4JE7nuUi7ocYHijZ9MyffW146t+z6EgXlYmjHHgMZ9hAWW+wucB3OCzMkYnqm
iheQzJlFTwFoHzvTPZ+N4g0yuOqNaafPRfETr+DDX0nEDzqj98CZohp+vRmYYsxsLkpG1jIVRw3h
wIdtq0zOjpPtBar5K+oVbVT2cbfzitzLe7tHI7d5DLXgzOLDjeIo/RiEZibkuOcDAt1ehDow38+R
m01QKYbLGWoPJrAh75WBTT+fltoYywgd5nnTE7QI4cpoMT+Fv6o5re+mbv3xMwZJCkvskTPU3ypt
wGdZgryhX4pBno59+tZzwY6OY9EZc1qxF4srhXVfc75K3/g8vVtiO3XTIBedOzZnVVLWENP24X4J
XrFwWevZFhO8wooLYt32QWy1sAKVfsAgMKg291es0+YjKG4EMC1rRxCFZmaALjDBrYfpwBeDrVVX
NVIg5OlL/Nz1uZDkgBh/0ZUYWbyeCithv8NpPigiOhAlsaUvBbPnpO0aKg3OsAtROBcb25+nqatx
tukVOb36SsOL9KTZxOAcPEWHu/AiFq4H74tyQYCRHvv9/pCsuNVwk1eq3C7cvkIho/Wb2y0zu2o4
Bxs9z+KrDGVkX5BaIBSl5+rQDGgKfiqgb0F30RhSdU6PZFCgHkkSFGcqvGP3xl/H1QOCkHzNGOzh
h77K+xb5KRD0IFrfwKE8WpeknK4nxg5ZcdgDvLfhN8U/MPPAAJ2p7UAsVTn4MCxU/xan/jFMaTMW
UYBOA6MWII/Hu/J54cVMKoTe/Go1pEf2kHzoRpwcaRSquvafRxrKn+mqU9nQblkyAa93wsr/q9id
IQmBsnup2DLYFiH86iVOV+wJSOk97meSixVULllrDsQBwW8K2UFgj8L8TsMS7TyvJgxA+bVpuiv7
8caND6R7o6DlU/O3pEnqnzXmEwil7QpwVUYAoamG4sknT/NTDJURTySVo5GZ2gKcafFtXPRoEkmF
pKy/0v0aloFrQ6Lw7aC+qfwxQY0cB2/IMVowQz3yvGaK7ukx/PF5VVMk74yyzK3dKYcp8dTKcKHl
zqNbDSZPMynq0OG/vSwU9/wkNwyc1XAYk9ySbPxaNNvET2FAGRUy6nLld/oyRrZHNAfsM/70VLj0
LWjtWRxIar3EUHdI46LXVaXHYnBReuqjqq6LQCCyCpXApks4WdOdVxhDtjGdVYctksbhG0+baaRc
yLtc74ba1S2lGLpxjHA2vZBhoMoGTOC04oMbsaluKkwN1NP5DtBVCmGsBW+ggFKqPUO7Oaik357O
amNblAFoPONUsjAQNvuVnRPkfVVFwhVg0S6SkXiq0jgewfeFaoZaHDtVTypa2kdkkDdmEgW72Y6O
xxmr58inlq4M5yw/a0BE4TTtZSMVHDufOLKMYEXr8DIa/6BK0qgT3XTtSWWeh7gODAdZlCtiLsmg
FDNqq2p0WoLukVsDd544gsge0mr7vc3yTDyJ2ui8T2EYJaT/6Oy6DwgW7tTXuD/GJq7B+LaSdkqw
KZSBejbTtqb0M7KVONb+YK4m8YMwtLxVY71ZSENmTvEcqVK1Ox82di7awym/QtmSNvNqB8sloKGp
+HtVGdQIJyW7rXVNnWowMG2019LMo0x2gmzK5AAXcHuaDcYQqay/3eDooEZ9y0L+dtmivq1dE/nh
p86Q6gKom20sTugaJhrECX1JEjWEDzUirIkeJXUaFI8k6gOFPT7vkcv2PMt9yOvUpaheSWd/ImZ7
2Q+jECemX3Ljo1ATISBLEjGXoO19npi91CdyHOdEZJ5NrZDpuQWF5WTAO7PNfBZzaKOTKdnIwcdH
wq/jUxTesOXT1lydN2ffE25LqgO+PFYiiLm1dsOVFrNTWl7Qk8aQpVYV6uAphiWQtfZ0IPhCewhc
ACYZ9rzm+ANfvnLCYU/KQVqN3IV7M604dcZ/SqJVROtZcEgbV7IqboKIkqL/0+AP5c0ddFGooMCq
wwZ3chem9bKPhLLlFPdlVe4xQHQXhb2xNVuNlxAmMM+ZmEiLJpO0C8ycQyFw0dMgu09xfs8w3DGO
srp5PM/eY5eIuBrOkK7d1QwxwVW0opBBXVfqkCxlbahuLwyJVCrCwuMxbQC+1Knf4H04STuPFRsk
thTzMWtgimc1BZEF9S3owhcSTACuxLPnWsvAPjaNilk3KxlAsN+/9GM5gT7s3Wu8n6BXW4Cquzst
aJyQ+CHFyVcIrznEqG+OSmFaIcm+4imEnseFKsmqb+IEGbOSiEX6EbTyHuibFd2ILmiaIl1drkp1
vhMX3MTz4zHH2V5NOAGBfrWG+7kK/GdeobnGJIF/II8gEf6iu4dCPzzxajnOJpeawHmUaBPPDAKt
0Z0ROzaeOdf/+2uEwNDV+4B833r2BefqadKNeI2hL1znjpNVl3hdtWckyDXALjJXQ8mBLA2IVbaz
G7s9ERlVBOfbZkhB387jApb6XPgia2uFhxNCmodiaxjyHSnVfbKCb4By3chCZRHcvsJpiDPJF0Vu
wJ4458iUC47ug0FYPxs8f05SvgowvB0OQKBkqaEphcaGyn3iVfP5+PeggL3P67Z874r5Z2OPZ6kv
GpLIBwrBCgMDsk2hW0LCnHz3sXyN6ijqzB+TBtbv5F7fsiFoYEmnM7qXv61E80cNUB6EKESGHPu1
ZcNohjm4XVhbbmj47zRdSn/96M/aKu18C7WOw42S0RExOot3KpR3w0HSWEoruJP697dwfY9nPvb4
2WAkdPpc8ihpasZw3hBTsbigWzEaCZapE0LkI5c2grPq3H6kEg4rVKnhE5hE4tavxgJun9cMiH9I
ldlIV9S+PDpyS/fDlu4xoX9YtBmRjzTy8j+xHwe9ZZKyWPo9DJdm4shKZaYVo+yNJW8O7O0BTZ8x
KDnnqZ1h0J8B6g1Bq2BNW4UeOtr82ScBn+Cp0+docrISzy0CrblqfD/Vkg878VQujxuXVODm6yrv
FXqGtckqwLOWYPQmFvntBSQbTiXF9TR2EEB97nZrC8DW7d7ZBZyobSAxj2AWk3ZeDOhccSF+f0PB
MV1Yb2Bh8idymzSXMO7X/Po3n4xJyUavr+QeletajOMFGkuW6yTbraAULjp+AEA8liUP7XinkI9L
Q6Mq+Q3IhuB4RPooNi33WmUb8csMOcdU5QpBxKrpsK5kNbJEDbSAEJYCfJxFmjPDR0P24wxz2nIT
Pa074twB3fWhefFyYWhiKE6W1nt4USIgMQ+w35cSD0WP+VcYFYOQh4MxQDQ6/9uEYqNZ9Um2/GSG
7RZEFii9BYwa5/4k4dEGrqLfKAddwbVMwfjTbyBDLs5b3j/LWTDeyFLpj/70/gyMAirUxfPZNiBO
RxImtItR9HkVe2EbWyWWHTMuPpuFAFdMJUthg26zuSgdgkak9sLq7DbeoeHAyAWctMybx7Egzfmx
ek2Bwhsr/kUEXpnPjOjW8cJ5l91HRYT82upEu6MwTNH7u+oia7jS+Xi8Kc+y8jVD7qq0W1sdPeIA
id2xPIacfo4HPRTjeMjr8nC050fGkCSaA+UMFy8nMWHS9yhGgtaPto7QYKNV5AQ+JfHNO/KQNP8H
Ek7/pktwkZL3qaXA0cbifpJDNUsNbUcT28tnLUQyfo15VPDxY6YPtzIVq2kqPs2ZDoSwAFwferRY
eQIc36XkGmQI2rf+f7VvG668d2yiQAjr5JC9zcLz/qkZ4TG+s2r3A5/kucFrS3+j2CskcGYQtkzc
7QNUIMa8vcSchTmsxOni5aPI5W43jrtz/JQLwD0ImYXRvoIbUbFqI2D8tEH54KvWTnPIalF44bev
0tTcoHCL6fpEoOkJy1cL/gekD5aMPAJWNlKxLjFaXsgRszeUvTSSzBBy9UOVhaTClvQe9h8CEMQp
+yZu5xUtMihYvuQwpUCo+GjTdBXbLtx6lmA3fdwMZuTmzGoEC/FI8XewP3h5maFmx7TMv3vr/rad
cyDV5TvQrerGZeioKx3tacdUv4zq/l+9HSILnlixKpuzHj5nT9NoAgAYuHQbShNNl/1c2lkYWKjD
4FsLcR9/kz5dtjcPHix2TM1YWC628ALNGpcEnlYncvQatzog9KbLrpJbd7fYMIseHSMQc+m6DK/d
aiDf0YXLgYbYl+RFrTq3MpT/lJB/t3KgsO8hLaXxoSd5FzEeDYuLZDLvgoy4ME9jUy3Jd3u9mhKS
ZUwVzsHKPSwlyRZt996sNzNHj8+E0EW2aHyuNfGxwrTLxZeTQ6uXRUlpqyWDhbzQc5TzYM6ZBJa5
yYbEyqTFPi0HzyrUrtNjEXICeUbC2eVpDWXsB4t3EKseeBOljV6ghxTh2jyAIKVBFv3qWH5+FNNE
p/GpOGtIiE1N0HKo5ri/c3364KZbZ1qjrH3zHBnuYf4x+p5e5P9Y4u58U2DK7u14YXVxRmSRuuYz
7NNaKGpB5gpRLTnWAHbG/Hlj1+rbd09ZXvUtotDj6gzoHTYXuLgjPTrHCqFnyMN7naK9Bau3eQ4p
jN90KW9tqPFkZS60YfMaTuWrigypWesKgd33ZatAkKI2+dWcKVVJApaCUDd3tr1m4Wp/w8btNeAe
qiyP6X7vMgNI2DNsAaQBtMIsHNqRNvs2bFKRPqyusgPmMQpiXN0Mn0TPHYJnvR6L8CS6Pt7PFUWb
3PeCDJnUiYnUKss/ammSO7TV9zjt2hDDEUAX2DY1LZ9lqlsRkoGNJXGnaRrceiN+lPSPhrHXYLII
4Qe4EMnedC2cpq1y5I61qiWml40IpmFOBSWROk/5BTuyPmPrGnxP3XDfFtUbFaFDh4A7RyxYJ8zF
A0wQ8jbD3LQO07/zhTxcMz8+0EKd2qUqwm0I9fHY3IeVrzCAIhze8q4t6AT2lyL23bK+ASa7bSzF
dyhvV6QZ1FZPytpAK35+CwMF4mWHAcfVHEObOqIkJTI4gsiF4JasheuAvnzfqj4EXiJuxWQNS+TY
vFhjqITt6e50rjPnFoWZGMtd2L/fXeFdzKx1xvi/M6EH8qnQX88UtomxD+140A9MkMVwDgdYaYM5
67YR4HNv1Cx6pEyKL7ujIRjMo6uKHc39wtATUJUdZbNlg3UK9cHTA4gS7C8tcod9m8TsrA6tRAJ/
sFqcZuPMR7yaM1zKKMsyntrPKpOLsBUPzCh7jA4KcoTzOhOeW0IxMKNDHokCIoy/2wmqxAbbRIox
+rsJNjacbgxv8MrU6wYUZTLVQ6vqAonQJFTibeVwyUp4cgO2S2erAv7XU4xyi1jgMqaCndzFfpHN
5dTIFHIJ3xFbeRmnSveSXMmApZ1GcSFGi4ElCq4VSf7Ah8qEU6OebhEGk1f2dAPgM2N9dfUPEWtE
hg69JN3u2SbJu4+hrJo0U4El64dJDXm8F9LP9QxFbLkDwdkw3f8wp6Lbw37teqzE6xweK9Gcu80N
Z7xfgr4ueHQ9lO0oO+C3xUBWJCCAyEvNB0i9udhppdlWFDqWCLbW/EBv5vqkKRcOeGIqgBqSUj9n
D/N+Rn80rGwECV1YNh8i8NDVZEitHVZ39+jBBLkrddlSfsxPFq52ipBKomyT9gr/dE/3sm0li+4y
yOLlUUXVBnrWojP2ZLtaGrz9KYQm7PFfg8eyHeAIkqwRXcybyAiyJ2fnivpmXQBGHmJwKVpWHDnx
IXP/vEjYTRCDddjt2v6Ef4Oo+Y5E6egQqtmRaFX95Fk3Imb5EU2YFBTT39Ndl7JOpPLcJ+m5Frku
qEZTqKJnbq4nelXDczjCis/owgmH++3Ey3TXakJwSVznog9ZB3HeThKxFNqEaUGx7fJEvHF8Kkl2
rYgrdiVzV9nJjCx/LqPtTuXduwjCr1V1DBD0qZQdSbXdHg9AVED8dyE92Mv584myM85EVAiZIlGz
8QLWFrVfZOdknI86BYG7UW55QX8lT3FyZ8u7107WPIXWaRP2cRCIgfv3aLwauvOlAJtDb2olrOpR
0NTxhcbouWZXkSkzJtgCpCLisiA6CSr31PTcd39Zkn2ZGZe//hUHr2++3TSXOBeHU+TenLwCoe9L
YUt8XxO0X793ACvYUuWmv5Q2G9ibKH9AavOrVokMbvBwzK8fwDaxoijo0MUQ7fM5pcHEh8oRt1E0
V3PB/S7rXkUh6sIgI4vDTFxaXaZxDolWVI1zPdrRjQxtBVoJt3iBAj9d71630C4vWhYz63XBvKXQ
dyYVw91Kt5cF/F64viMk5pdnY+izoB5B+dYNkEZVcnb39RrsJfJySZMlYpJFrShRle2YvHFG5ucJ
15yFoH2siwJPblNtyucAhuJLQPyH64RQl5+n2YXmV8xuRL1Sa/guxCyp7hI5F8lxmyVggEhnOUrW
G+SPpXAmQguMfDAm4DqFBH0V9Gd2vBdzPO+uBkjNAhtX1Zk79Y4Ifq94l1plbAKCTFPVlQskZIrm
zVa+L8K8hwG+X4A6+ySC+z0dHyWwTF/lki+vWT0nBLSPL2GdiayuHxlWcWz60kS8TsASQkQE9P42
ZqUelEgag4ryKmu6XaJhzlSEfmMnvPX5ILeY8d54PlTedwXIw+LdL5k8o5Iqs9Vk0MygRjzs6ZZO
PSaKV4zvS6Oj5FYsomwLRyZxHDQRIfmpPZM5CpbDXBDndwWnvrHgP+PZqIyo6Oxv4p5Tivl203MD
l7b/gU8T+WBCUGNpKvrxyGXK7X4JGLKQIKPLKPEtB+YiRluRCUhHYTdal2aR7YZAkZSWDNcz7CR6
vAfk/bpg5YeidjXALNxe9QPG5+2QCB1AqgwaTSaeiAe+ANIqiE5h/ORImBHskAhHykQgr53c/bF7
TnB46N7p6jprBlu7K9zGneirKtBg1yiPZ2B/lHMfBK3HvEig7ITTUyuYFaKbn6d0AiK6UdsjO01A
dumj49rBzgCptqbURP2EKXTVkg1fPXr8z4EpeCb/vbsvgfLZfqh+mVDB25Y5+UJGbg4aHlmyeHk7
fFXweWckpAPdaS3EqiO+podzxBA/QFmTpLf+nPH/TPbos2CqvWX94RSUdAbdBl0vn1cSs6UNW8Tq
cmOCpn/XQj09plwmfRBH01CaPJ7358eiLk+JvKGe2NAHi9zjdq8tlyV7gQRVJd3sGIW3Ur3TjMJn
Xv+NWhgJR6HW4ZJzHLC7vBnbWYj18LWM5zawMR2Lxa6bodvm5EgS5qlK+ikh2dmFAczw/fHT403z
ao67XOs1Q2ZHu4rhEwYcSj8jis/RCR633JyhirqhZRtPwTmWF+xo6o4r4K+W5KB2bK/KwBhYLm9R
nJvtk/tXaVVtxZD5ItMWO3ReLIZx6mL1zrTciLyUwuBXc2zXpcCZnMgeHuB99lQAialwbgNXkbz4
4ylCEdK+NNxEZaPGWD640lIHLRz92XGfwa9YybURpWMoX4cZOYLnlCRAUE9gsMyLMZiY9YBr7sFH
IN5ryIdYlkq4UrkiJgPSqK5ynwduGz1e8RfXuUqmrtskIfEpGV/OjyX3gmBXJUN4VAzs7MpJTldY
i2IyF0gEjtj7l4zJZi7U9xlHFHm2Wx+DTOr2JsXN+WqtalbA82qy6TMyhPpzSo9IAJvcHNL6/oaW
n/ylSuAhbSX1AJ3gW+D4cRrRTyza9J4eQKNmZiTyl0s3Hqj9ynu5Lh3dIYjGp0qo0iNfwb1ogcai
XcJBqwbOjba+e6POqh9QZus7C2GzjWQPgZC2jtd17vCLOx3601ReG1rI9KJC0JopLVY7aB97CBEc
fT0EWulYcOmAGRivfUlbBH350d4hlRRR6iCw+bvKrUDJQm83RZPnBO8i8ESmw+/tSKYrl2FF8nmB
Wo45Y1UpfdD301J+15g0rVwXO1y18UWJgIUWP1RNeYhL2lCmIayoMPlR1ZkiQwTox09oRGA3P8oe
pK8jtZmrJMGEc3ijaY31VEQ9dUrYY4JugPHiAspN77FScHaeblGD+/A8bDQdZIbsRgPxD5QzBXpa
gLjKSvoc1iq4jHC//9t+j72cyB0JJAGva+yI+OqvPcm5TkoPDspzBOc0qU9Yc5MtfDeYxCji/k2J
Xl4E0Qn4kb2AruWkZjORRIe9h5K2rSh+O35nkA5B3WbVWEiLb9E8nr6Uo/CCCwwiT5LV7bv6ZLt0
7RWyZRr4wDC0UgtUTuBgDGIdrQo4A4txAIv5kJQaf+aeRvEX532fN37oUbWyNpAWUlD/4zsVaVJ6
bLADITwwmBFYi7I73feopLu5WjeM23iIQalaBFb1fN39w/XKS81CcEdT1tIvpCFmBih1xtKwqcs2
JPTtnoXJNFJb2e0L0YOnd9QSeRyAdj29tHlfgs1bCcG+uc6ZiysuTF9Q7nV88W17D+wLQxpQaF+G
/aACELqXc8JOc+ynCzCN2xc2Fp6fWdpL+DnbIMGwB4iKcz3UR3dlF9y368/zwIaL+zIcQkdHTw5Y
LhK82L3dKdkciWlgAEwPBfXxVu4VvpW7EWcIkPf2w7XItj7txdeZ2otP5h6pLHdhNbal/fGS0xnM
vSXsTR+/LRINC6vXupg66VnwD8Rb/bZkHSY9JFDLUqq1SoLLS1aD2QqSBi57KsXuu4a3oA+dnayF
RK/VUHVnRICY3DFwTj7GKVoRqGKZhIukjLwp8HEzoMwyJrXFHMWkL3sTikLgZv4mmCWjpwLkC59a
zWHtuYVlPJkm4hUqxxs0LpYZGuYJKkOwuVvuO0MB0Z1/7fBcpSInqT7R4h5kNsqavtiO0dYnVfbu
BUIBr+bvpo8hUmaDaxXkLNVXcQqjBS8daZhApC75bG0MM4cRd/QFhTRrH6pNGjNlK5kE81X9ZDYm
hOv6kp2p182bUVpPSb/Lwiy0Fv/mP0eI4aJZn0RZ3He228Cvt67kl81QSKBvRut7w0//+mvmiVDi
vAd1/Rqpj16f1YhaJ0K5bUPFJqO1lfuC9/V0JUX1pDGx4tlsNDOGXSD3p1X5TGRZQfbj5AV7FUdW
5pgvXsKPA35UZjFaizmfINI8Nh5+dBkkumLbjV2q8/2xciOBZzw6++acIYpXZSV6yZ/G3tZG1aEp
sPJV5N3V7bLMoE9OWgAGEXzX5UmQCEbXZaF2Okyni5gU9kUb2QXLBZvIkl3RzaYGjRAY+RoHFJlz
GUdV4i1hW9SLEyuwhfgoDME3p2RZYnTTZVDXb/XOSaWB/+WzGV2LU9XKvtI2E9b2JCMSWxd3U2M4
m112EQ7gfQ4fSDHv7igtjKDySs6oIn5vzFJFkJRGpwnC0rdeYQJKT914S+nEKFRTzemic46e3n/F
nRlUfKTaIzXck2xtuLr/JVtGOx8R8oRg8GSCtZAQi3hE7wTM0pCq7q2pb9F2QYoN4AtiEJZommtt
wH0wVss/k3RPu6EAYbgtE1MXuB5E+g0UbyVSeDyyxJdSIKr4T6mPOwD18+am/vRQw1WMJE4c/8TS
46AuhYWw13tsSeWUOULJw0ETcJUqxHkKQx2yOKpsXnoz+G7/flSBR1B2jOMsNganxaH7K3j/XcNU
RqCUEQSz9taQ+V8MV8PEX9S/0jF2ZMGDye2rFHIM4YqhFPDD5MgE0RYIq3kQEB5xGAqwW31hhLKq
tVBRitwdx7ysGTZCee+XdoWbv6S1xido9l4bwm+pP5K2bwuVUMumnLaOnty3yBKjnsifeXHsumxu
zCL8lXjjQ9OdpzKj4GJlFYg1vnKgYkBT4NsMuK+EpbKn8ByKKj8OfQU/gXnsUNWcOVBQKh9SfK0T
G3Agu8jqsgmgeyfc8LIk+cNn17qDYUs6zU4ySa3R88j+qSAlpkoA/xiBSmVsI8yMo8tHHDNZew9V
k6JbgIr4SwxvEQg38K/vZnNmPDNyiCvb2lWYknuc/MSyz7iJgd5ZNx9rMwqLi2jfQMTPP8B0e7FX
pVVfsARmXpJ1YtzTtmCcgOyRyVk5eGrsfkyETAZhPBplg2fe3TnG2QrKdCLj/rA3u/FTRtPMQ/Dp
iqjS74ea7OK/fe7oVIAVM0UpuXKR0rvdPAA8Hjvvy+uLoE3ZGetluxFSdbHIRwrF9enY8KHKwmjt
L3PpwcKv4vdmgKyFJDWle6NPXqazHucrIRaH2I31FZ6WLBSOKK4VR9T2zgVCR9cPweUavz9MN6GV
WDPdK/tCAqLgZ3O5J9KuSJmdTKKLBWK/VfpxJe+PzEKVYadZBBlomyBIiMtvWopB8KOFfX8lJCCk
pIobX8Vh8KPZrtX09zZuyEMOG+3HfKJl2+33MoraANaVsnJ9GLMfSpfHzFR2MkjKWas1icGAJO9i
7wCvFBeqqS53OqguJAGMjzWfW2uCIqDoq3a5y7ZJGbkmNO2uDWKZPEt+6KnVqoTyBYQIOhTudGZH
7pBPXEbm6C0kVg+yZLZV8kSyrMuDKk5zI7xvqjq1IKVK3vFsxP8Mr9Gy4jsmbn5SuwxMEZ9zvdsp
MLiPikYDe5oBdUrvf+XUYHbXlgvpC7aprkmRhu4TJdNu0FE53tG7jiyJqc4jdcuOkiGqpq1lhkSH
ul5t9o/IaPR0wl5Awghb3GSAAKj77XTHtQuJI/DdxPIJtzsPYNB/JljAAM+LoBTy7kH9TanjVBvz
HK4tx20Ljw9IL1hWjoBllKQBsM73x42JOpxUW0Ewq7DjEEBvbO4glpRmVLPc4JwlRAbz3F5f5KfT
m9k1sjhfdVu9o9KbmpTTl782k3r1P9x51/butBQDbL3LzrlesKusaP24AB7YwqJxG2hpaIRCOxjI
xdjV9RPoOClhLNkhI0YTr1GKMfMfSI010ghRv+n3c+tC+4+v0ndi9zwF42RmEaZoHm8svSBCVw7c
OwhlsSz9N+4bEjiZZMsLIxaNlHHPV0gflbZkb6+t0wXza0MzmyqSo3zrom35edf9lw1QFWlD+5p5
COunHsTGcEMGTUNlQ6BeUluU3sPP7Ql4FavN3IDXhnOJ8q2/QhKYPbbMpVilW0prMTFDLjJQbpcu
9SQ39ugqVLbqhSe2qYx6f64yqtMG4VR/BSOwJUHh3RAOK79pS3o8zNhjagczD656K2BZOMtvaIDZ
HP1HQluHsuJvNgmHSVft0ZgKAA+dRiDJCDMIXISL8SmTpI8cR8KHgeHy0fBXXRb71Iq7NvlqDiQT
WJemXYlauF53Jf/J4wRMAOaRa/s3KiiX78f+GP4R0iaAAMqXVvmEbXmtd2TCTeU8DqHoF5leRPob
z43qSe1rqV7cF+jNDn499emWjf4YBFfUUCLScK97SHbThRBesLFS5jAd/DCNF8JzBrjwgTKFG8YM
p8FM+il/um6aMt/o7HXbitF8VjJOuMCrXSMQlAo+okVlIasyxUO+RT+eDrlrwD8GGx2JBvU1xUau
U60oms8mIN2nM97zAUoN3k2A3kY6wVvUkPEn12nXhhkg4wJHnWvC4pOkKUVLoUzdwLXnUlebmhxe
Fniweh7sbOuJWF/gYBvDHwx1afDKqQ9kdVAlsn8ozD/+HHEBN4oeWThgH9u38kBcZ/49SlkD14hG
DZGxRdzCEKbuj3Cvi6H9a+ASF/3aflQr5iKeMxvxgqcXG77k9Fh2wyeJ3Qb/AUz4ifMKFIQ19NLp
4kbHPAdBM5ThKBUmAWgc2N1B/yXj4n4J5lAn3/hfjjHkPJYwjEP0DwtBPOUi9ndzqx6lOaDpOAiZ
9FRpvlYnKfZu0rDPhlFjS9ZOXK9O+1Wj4FCDh9aaBR6M7F8mNfJw9Xxf5rVDV3IgLOtSdaakN2FI
mrmPQuYZMJ98OpSZKlOVDVE2mrtrBBI3aKHrZz/WV2dv7qFErNzkybMWvZhnCTSouo/4pGmNWXXR
9rL8qx0K/UAKMBqmqiJ3X9xUF2xTCuueY6m+jRqOPockz/Bf5vwO0OH2hspm+Lhc4sq7QHhVup4e
njFPEUlQb+9hL61ti62B9txNnuiN2vsmJBkxOZ6t5U3vpvyxOYtzJlEXbLnOkqWL0ffYJaR+Q1WP
9IWg7W7Ai0+9nhzzpc6OXPSketecJj2yVpzCC00koq7WI1RJ8Rl1aGZQ8dao7RWG9OXYVDPZx1aN
RuremHeFEiMOhAns1ngr+4buPFV8ivONK3adc/V5K352GLZM9Pw0WouS1L+aBxI8K4TwUbl0l3ng
WoQek9HYJCq8Ks1idRuAwrpDP9ztAiqeetxqOYspyGS2LSkieGJw7XJEH+HxLwdcbTYQdTz41PRk
apvy/VltD07D5TaNVSv121FSYigB2O+q3h0NSgbqrQc1gjQUDXyN6sv4oG1hOp4y2+mwXXgHhVat
uUIvKYyPU7pK2BQ7i8OqGCMJM+4QJXguNGnXvs4+dQqOzTu66XoQRcCHqTjwnQ747P06I65KuUjr
H4owwIksnNv3SN7/LYJCSzLNZOIQmxmJTMvNchd/p19K5qM9VfUP98Je4Nyj7+vqLjUcTIUOUKvG
rJfaByURcAJDL1K7oihhwxGDkDcWMvvvh6DyTk5aLGkRxIlUXv3glVn9aph8okEXnrm9EEXpVs7m
+8rp+a/YGkyjh5Q4v0vgGnqsHVEJPRuUSj9RjxzYuczk/zqx7DpMKmMpLIGMcCZLVahWsfeAYNpc
ylDYGL1YQpb5QGj2Lx59ki4+ytQ9n54vkLc9gyTGD6PZyq7SAHALqSLc3G4C1OSn2+wm54hO+FR2
1V1l/iBvtK6i4/S3bGqqi/LvFVWWuy4zjbcPfvHD1Vqy2CxkwyGJP+F/xncrvyAAcZbk6CYPtTAd
DtAVBqMShixWG5UjpNOASjJUGEIykZ+KiACOGe67ttwIK3Vaj6GLL0hp5dE7ETMKWus4E6KgOA9t
FoQH7WOPOHx2jjObMIgy2zmep6kONWiRqaD6/4J2hMcot0psiWZbRlYH+pKRxSZ8KyKzz3vyX1QZ
YXT5uuLXwtSvcNxI/c1nEOQgmDBNT7zvsaJTmTkGuL6m5DgqYO5P7DancBlnTqZkJxezc649Kdo7
24t+JXcDo5bxTxft/d4DkbnqgNBolkvX+56WlcOJdYjTJkDHZY3/PjS0u7NwFpscgHfkSkTcN+Ga
RP1ouDn+Wg7iAOjGLg8JWsOc6R+jZ+qWSVhPHXVoOTBAC4nvdMHmMU14VNeCwZRUCCQHBrme2gKJ
p4S4bPgdV7T9PlkbVt427Zy6tE+YxeeJaLhUGC9QLBISSMR4/SDrJJMG/Qv6lyWpLndI1rJjL10A
yH6VuL8oA5qJn1FmNiP6Ggd4gp4MxTZejT7IoBRqrftC884+VyYEKAnO1WYi1T08Tf65LoVDkwMG
WsIswl9pqtkRcFBqgQ5v+eVZDUkAQHFEH9tbdlQvz28FdnibAFz9y7I+TCYmg3DTEZfkCmrMg9XL
AXDgh5BZJlQG3cg9xB9GfU0uhZBFT6W0V8NIs1IxYhLsokqhuf1BJSu5DNrxj56l6/C45nQAW/5x
kRJXqv+P1lZ+7phiaFgRUGtfdZ+wHcu430uMISOvgoGSaDDq6DlH3OtLLzrvFGUfLOvuO2MMiPCP
dvyyCFKRpPxDZPWffOG4HUGHTq+PhXhRSbAm5+xHuj62rur/QVemGmrodUKXr/84thChwum9wEeA
oSu47O5PAF9Sb9gzc9hMpZNe06bfuf4vdNSGqNbgNN6LTXpOpmkgS2JzVk+qCBOoiszEo2dMBW4h
zpvbm310LO1iznStan84EhY6Ijx+cCrvbYDHeQMQuBwhODmayXabhjgd1P7iEz/LFU+msDocTrpa
b8exScXNT/ytXrVoe67aUQf2ZRyVINw+pnIQyBrLJ4nr6w7KJra2YKz4jEOYEqG5NCImKCmUMG58
iRU6qvtPLyQrVYrMaRkbl7Ih8kcVUUi3vwnN2hS1hV3yULasGaq31UwaGXNntR8XCwSpgwDLZXSZ
G5mruD8m+JRiph13GeqeyNFWkCzFBX09D1MFOlWpmrsAkQoosvnWIEi4ZGnGXIoVnFNRwE1Hu52c
U+0GqDdjQnBLerkueEJVGxS+V1+SQ687NSe7BYgIRVic8Zeuns4nxderijVGIrRj0ywpHAESAive
9oCI0O1WFyMvQO9WgIB7sWGJenaBWpqMtIrsCUeEIfUoR6PnS+wscDlhYVeCc4EpWPf5shIKP+XH
5v1yjiU901/tj3XecMxcvw3OS7SUw/qIukkAsDomHQ4uDcV4rBav7LC2m8641LHQzuQLnIDoyoXN
8RbPkdurVoHRG/0cCZEMcar/xHw2y1uQZEbqw23a8XWIZfbljWIz9wo3HuggUIymSY6QaQx7jzMY
mPPHsZtB4RMwPYIycU2eHXCwMncJT3ZBeqJiDCyQ5Nz1iUzJJ6M+c7sG0t7NCfuiW0CR+wEW5o49
TOaYN4crOacQIDe3yzaT/jJw6Jly8/qTu75q+uk4U/WvAjNzdxx5ckv7L0DsqLc8GecYZQUtB1EV
HFIATZdcC6cIof9wdJeDu+Ni5JXTlPZxKohUQDz1kB6nWgOvXI13YU1veg1LpZupLaH3tjAOJcJE
Ow135jJ/7ay99SroJ6+WrAu26H/+47sjdt62HANWjUzfjT5jy8y7ORamNZa67APQMlbOCmZmvnaq
4sI0TDHUg5NCC9xB0lyaGesYbSd+shFB+UJv+3PXV32XlpGqruKxaayxQTizH2bxA46HYY+VEjsO
lodbbg65iU7236vH7xE/HiMnqkCHhf8FBsWqnXLIIJqKPiOJBP7trho4Ro3YoMbEHczx1y7tUROj
lGEYtnLefUm3dJsfCU0/ggvwb8xuQY+Fpc7J3PBo65FkaN2G5+eATw6GyePDKpPL2soEN3vqckc9
3mwy5GjoJ0aDZbAeJ6iSyw8fQBCQd/utRadJ4vPlJ7n6kGc6cY39JhGMtozu5PXOI9/4Gm3bJPXN
R/2F1rywWg6LAZvqGkfObmzfT4fR5NTiLjivNIihZZFtAMKnKenoD0dRQWavTJ0bvdfxIkoIsak7
EskJVfdFnmn/g7j+EPz8UhMeI6oYqdpaaOTjA4iQBMvmFHX6zJeJIf6aue3LO4d+kHMBzFbnBSV/
6RBgR/GqcCZ413W+dbVn4HQ3j7E9UX99V7gFCk0BY41xKpjChMN/JHjl7CR/8YXH4FySTIuuaJpj
TJghGzSfVVqeIFFo0ap7xn4n5Sg23PFXICmfms6EMHj4exehYfgdyZap8Pea2R2yqpsatawqJe6k
wmYqdk4TcK/OT7tcG6qBBZdsKzH2DwUbyqlDpFFFrd5AHOw4HQ88BLCntF6MA7W2VuqmGUsf357O
EqA+l91cTJBxS9cpUIGE4dtXfmnHUIKTAcIfXgOOG2HrrUFtWTRbkxQH3qtOZe2k4LnjCxOZCLTt
8U9rU3j2/VriZwX1WCUrAK/YejwGxdrpIR5jWeVYSjWBB4ceN4zS0NziDboPVZsY+ymTHrmYfhSD
/aRSEpLKrkpcu/+S47D1LSI0yT3yL7KU22nR0vvXP7I8BSUhJcx0tC/YTfDB+T1/klzjhE4bw1aW
mv8nliFf0dvCmvas55hPUn0SPuO4ZiDlfuaXEiSuh9E203DdBrfQeoofTaIVXn0pKIzVgDaXJ8T1
3mRfXd9WPCn9vS5Dj7aVJC4xJ7PFft6R2g6rb5u1nh+FDrnfjdtj4S6nsPK7PtCIVq+yNkEVGz4U
zEug38UDYvUvGoPnTrog/emOOa53T6h9koJAnnZmLls6x+X+NALicUvdtKHM6UFkUL5vn2XZvfR+
hN9vN/Ivtw9Yl81PccEKkicz3ACndrZOY2suOIqcvpLTJeAqSD1NS17z2DVCgkT3NTn2QZ2M2Lph
4tM7rgZoX4FwmRftXtGH0EQqkJEJFZ6AwoHdxa/+mAYvRENGq767tS1rFlWhuawzJymPeY4ZR3Ti
M7KTsa38m7f99ztKuaBibX1/fhb6Tsmz7yHW09UKlhU4KLA4T7KU4XWXP+DzcGvm7z39aXtCc32C
zXAKZo5uQPRqUukTSL3EU9z7WVRa1cizgUFXB+1YN4bQAg7JEgCnWPxpxUkkZeDFkih8mxxBMty7
AjwpwM+TEgD7zU3/w2ApBRcs30Bi3PRX3Z4vvlaWpUNr94wX5p2cm6wQIh1udcUbsSQiQuZuM6Zj
wUxoSO0dVWYRdlC2X/TA6ej1zbpTZvXJh0AmXkoS/5w8fVSjzDMvDILFPAvSVZBXACT8yRvPk8AA
Bf07m/1+ev8/2uGRnr0L2uojTaRYs+0+0d0iS2MLvKTj39C+GruKhuqsUtBLBuAe6uCsAlj1iRYN
YTk6aRO2/ziw155TWnmsQYZxeBFHvXvNPbUFHw371xmAod4oUKrXhJPoEy1k9p9LAzOSoBwiZpwd
kyZTfa4A9Hj6zj4SNukOi7k77shrnYmENeqihtNFFKCZfNDWCRlBXAr3zVEf2kSlo+1Vz2ygFAkc
+Sitghs83pf4cobpMSnHH19koQTk6CAk2Anysn2TCmtBFm/EApz5JcaUJag00uLlyH70ZqbDu1/X
lBCCFhzVS5Z4d7Ha/BwK/bmqUSrUg66215Aa0qCJCXrFkpPTUXOc6yplLtTQydZNEYTFI2iCH2qV
SV1V1DZ4Tnp/SkkqsuRvSR4P11IJqomArYqV+rvE9Y1BhjgROgTdyrK0KEyLQgD3gQr3hsP3+u5b
NLFTuBdoKArx58+spth19GphGiuiJD9uwWzf3FLAFT7bWGOG/Ub2Id7i7wB07iW1yeL6QQtMmIFU
jgRNFgw2G6urCskR2jFUHBXkPlFFAtaerDeq62N1CpuDnP3RH8x4yiiMJJd7SOpGn5mqIpcQh8lY
pFwE9orjXq3j3mwJtUQR/0rr1JwtX587lHT7ycEmAupVxfSTQP9YSnhFB1lORrlHlS9oCk2vWhzy
HRmPqMboRJ/ZgWcaNl0WQt2bQpe1w7B1YkHSr6rRsdUJpNRVYpn4Y3mbg89oroVQ8WlMH+TlwciQ
d42COUiwxaRCt1SbRXgIZnHguWYRf2bvNmhSBJOB4gH1P2x0tqL9q9roO/qsYREfyJwnqu99Qgt7
haEp5Rr9nEyHDYkkG6GoSuXhZDbToNvzJ5biaADMNpQqVvES/khnOZVep74IJ6L1zEIVZ+I959ok
G7PgPtN0PPWdzl1vyFFCS3Pb14x/7fD75WOhaCj2yPRVoxi5oSYk+dLUUpv63clyF8m+ZH3kwc0e
bq5r9vezuEIOrHWsldTKGqYvezEgUTrvAlEiHmSPK1nmFNzSfzSAMn56RvOIGshIWLZ78QcItxsR
4W4O9FZDILmB5GJG4DoGv+CJbR3n3jQnX9jnCbMytmy8pKLEEc9GaycacYUBA+Uq9i9aFf238Vkz
L2UbgqE4qsehcSDXpXyUdE6osmre2HAgHvkseCs3djr/g4XeYKZauGZeOm4/Atohd3AnE0jvSPH7
IML1LdmPXaRz6XjQBj6931FdHO8Yu9TfeWOn2WY6HzYBpIias3OhPJv8LbYYojvDSndsR2axxjZJ
Gz724Gt/h6RCaaxCIrnpOEqm0veW+NaFNufeS8MQYQN0YwH3n7Fv0iSK7OQY+qFxAqw2/Z0zrYwp
nmZGxeKZ+p3xEd3XNZgy4424VDcUs609KasZHfVM1HFlKLoOyXbudH6BEOLqejjxSNcaBqLGy8Rd
N9yWuBEhawzwddFYb2GJIsA7ZCTsvMLlCv4Y11L/P6rDj1aQBsm7NVoQQC0ePBOBJ4txpLMYrbdg
H99wovctxnKZ4Ui41HSFZtaZRn1pHOddhd11rXi2l00uA5N0rXr1GfsFp1APVOlIqHWk9vSoSm2c
bqfKJrStQdWh4MvErOs58MUoeFTdpbPy0ORa1AkHtzEcoMXwZ5btEVNtCpjRnqcpf34HKVmxrsXR
nKrALGn9EC3/2XBMsmc/o9moabtx5Z3kHPec7Dt5aohNM22tANfNXOhCa7DiZnUUMfJF3eDZdxsi
B6T/NLqr+w0f/9na9h5Y4KmrJBoOyCIkOP4+4cPYcR1QFnxNMmcy0OjzAgxGN141zcIaa2rXVoW1
r+eckqvX848oSHSUvjHtKW2ZTxLj+ve/VW0M6zhFBN5nz9sZ+Df5L1G2CatxqHewDj+RAujAru9O
mtuCgfwcVJJjTORN7xDkgAYZRxYNsLLc+L8kfAaztBLYJ+B8ySMQotRwIRAXHz+0M0LJ/AMoghl4
IpfM9FdhmW+sXKb2Es15nHMQQezZHQkYZQjOWCShhiFpW8OxcF/07waQRRo1NvrPlUjQHCX5fnFC
0dq2KSolYdZdmEF3i8d3bnWtgrdusiYttZ7+NWN2MCobW+0qG5E5gJELr9rX5314iCIQ2AGKfFXV
NtXnsN0iJldCSrvCGvhazxc2ZECpyDC5Jf2kA3unyKAtAVH+uUiAPQpQXCtFDHsDCGM08j5FYCSz
52nWsJ45paGX+w//wv+okasqCuHVB5QaebuO6ROPj0YDMMPxQcoY7Tav0jg0Um+N3D1sFYyKmmOA
QejfM4BctPOalHcOVXnLMkRrE2Qzcxv08rUDOOEDuYZeO6i7rHLCTt8Zaqop/WNLytcpnRRarhzf
tFIldiPmFstToAhr/TQs5DZLlfc25AyNpuXJgLvQgGkWIxzWa8OdFFmE743dFC/0nbeppi8ZVLTw
EE/+rPLQkve0eritymtzUji/abTUFir8sZUv+hF3i0RMHXVfy8Apyb4A+oows95I7fdY0bQ2lQd6
aBMqrcsEmlFed1XCupabOMtnB3AKV4ZjtRdtMG6l424/d5UctbycQ4H1qF9SXYb5jq0SLCwTZerI
UqxSuc/kcZ/hOoaTSVh797qWDA55+WkCam/EBygwDRT4AgXkNs06TjgQZSh5JkrNQ6dxMNnjAJOD
78jzo+L/iR79G/XfLfECSdxXKwaMsM7v+khyvHdk64yEBLhXnmvfO+jDQv+JKIanAdEdHPUF1DjR
jDk38u8cBPiLVQxsBuUM+htqrf+nBXzG3zFBNc7luAANxnyU8qSmqmHiYiBXLCblo6JZ52h85Ktv
C1RqW8n4e6Pli/eSVXC+a+OVVhK4cdUqMigy38eYRJdU419fPCgDf8bHhW5PAjisLqC6TXivsNNy
0evjrEslsF+JVMynLfzucePYA3kJwWobyhgTvjPC18bSExeKb+pSeDNLmmEixaimE1XosLMkjwnu
pYyCYHjOSOxbDGmiP27UB5FOselRZnJlyXKXu+JGPKMDSF0wdlmh4CMkPwZvbbfFP03nfu0wocfE
J+7q3ynvN6juZYecTyAby2gGnr9iEZCj17qG+l5venaeUyrr2hUrRyTGsrKcJuOLqsFc6LyIt3TX
KjiptjJT2ITPinMGzaA58khyWLOAjAd+f+CdUXfuOfCAlChNaOHapFgXq/j6aY0g5AN+rDqjiaBt
ARn2VcCv/tklY9raTm/Fn7BpBqQmj2bBxbySpxmWywwCGdQJUZfs628/X8XX9jjFkhbOXDkmeMfq
KccrEh/xixbVr0GID3pNNyMHwg7ww3/ZOPpikvludS01XYDjbbPb+GZYc97VBg69YrbjqesPmeaz
e94gPkt969XQslB+6s0OAS7b7MFycjT1IM3E0Bafj7kKL5QCNqlEyq4CrRbC2O67e/ycch0aFPLL
P4yXXj8v/kx4AfBZA5jFTmntuokLiS/qwiSYBPGXmNTvK11GrscqRZwldZKAG9yIp5ujP0MRATmL
dqeDMBCPLNroyG9Qd1bSbh1Ve2yD8QyYXCtzP8fbmdWPql4Dzn1kv+6lcEQIka2zjgd+zBlhLADJ
JImoHd4dmcqa+IL+WEjNsUYVt6RTe/y32HJ8W7a9zF3NzWX/Exb48Rem1/HglQgsujTN+3tm917x
uzNsW0YgeCqM/5vrSlNhK/lhL04hTVDJpbH1SO869cdh510InEozAmmOMxZVcM2MMPq8iyKOYOFQ
x0ns7WADjllPRP4Qntm7Qc8aX59iBnuCCdpRH+K5fwuTbi6dOQveSiQaImk+KmyWCEbEW0ns/ryc
cpXzh9mWK1nC67YHFBOJJhX+8hBnlL/7bTkbwICwS6K1NnlRyrBVwCBjS7i3R8EXbk6ruTJNckic
8qLF3mtDksN3HUtclOJmULZJE12ukYZ03erug50cOo3Kbbq2zwRl/CKJiXblHsHCuNzpC6Swu5fL
MevhFMgePbPmxbfhm6DVj+jt08DyRapXJLx9cA4cAI57VNXJe3ADf635rbT7ws0WOEx3kZDukZVN
jWDQ4k1nXPbq/ATKpHUM/6pdW/mtZjY1kBn+yBSUQP8erXxjmOCfvh3lfqEYU3IaTVqBy9k2DskW
LsxoMcioZr7udaRTCQv8S5oa88eswWaT2Z5HebeHeAWA4q0GpRJWZI0bBwvyJEWPr4NdQuzAyfwO
87Dqo8EwYjKvlqm68f7GEZ5Ir2vTcRcXsqUCLB1gsxCIcg0UXZJ8Ho5Kp+wSm/duQynVGg7PWUBy
LasTPC1KtL2ZIqrZzg9vuU/EdyETDAj1m6Ae47kRxXRTfXg1WERNjcXly9JFNH+7Wre6Fuo6iv8R
IminFa2hvjRpXAvJ5CiObfeHkstjdx8ujwUx8/i6fewGOjtv0GJuPp6X/61RcxwCvsB2KjVKkfha
2MMBzvciGGlnwbDFraSR+bXUEIcgtNy9m4QNH1/Sqc2mzlnRtFFBtOyDiseVzB6pne0sojrslJAs
xdyO/lpyS7KMRcY5Ic1k9oo1AUoQYVEHqc2wUMJmkBjO4oOD0veD8Jc3C5EW2NpuobdqtqC8zw6K
BEvKjb4894hrjsq3B2wfghN187bOIwTdLrxn0ieXn/73l45yvjB8VjU3Rd0gpHi7CIojbieScmeT
ivi+VON143mw1pUY5ZrAmhj7uiKmCYskPinPXaCWYN0neYWlwO8Hc4nOxIPP3cwuTSMP+Gck8d+b
7f4tlgO3tNgyKkj4dr5z09ZjTFvx39kD80KS+PZ7BT9l1dk0/l50ax43QUeAD8VJbQvY1l4QoiZU
e5zbDD/l60ja5pjCEKMk4w7ejsHhFVtTncNXVf93epAtvxYR1RsY6RdifJgIKx0QsPBbd7a0lrNP
1CD6MaNidsSXKnQJhXL3VYAQi18leXhRGzBkXmxR/a2nz3xdm0SYvHNmg72478NFnXGfGshHVifd
cYcKxaUiWWp5vhtvWzmEym5ImTYZSTQ266XdKdzR7Zihqt/S9pXL2W5UO3Agyi0pKWwxx1Clgq0d
S0UlFNYPT4O+koY+4PEhl0HEcIAah63xMhZnnqJ9W8NLSmwGv4xZfqB055vnVpbmvCJz6bDNFezw
JzJ4GYLb8rPEYn9z0X9YoJGI7T5PNAuI4ZrppJssKWhlFIFCndAzJ5qtPpT4LIQq4q0cTtHItoVd
SV/+cqm3h55as8LrOgGo8AwaT6usEHBzdFxlXIjxTn8XN9pOPFQyVPmRtRyIOxLOHwnjzc6i698e
ojlHMh1/Pk5l/nmoTPYMXrGpgF4LewZ4dntcO3V7HQnhtN8rGSDuVyEg++pxiC2qkM6Jh5DW7Lc7
FjBJwwE1EuK+79suYzyLnW5recKj70Y8HOrzcpA3fseBFZYMiKeQQYSJr4RBAeEqpoUCnuAsNL8m
cEKotII3b8pQvCbrK7xNXFl5C408eGK0itgmXgeiuv5YrpfJidf0pktdiMrz2mxdglqTMwuQjmVV
55FEpAGYdv49TJ+v1jts2aZ4xGzMGpkUyqeY0alLufbHlxRyI7PwHC34LePBy66Rnp/JxZKfX6qO
nCS94lpOP2H+hS60hKOf0P2d59FvkMQiFlWO50q5vEg0Je/wy7dyoJRco4Wp8avtb04fVgMhwNnp
mSDEkHXWJ+f7GZeg4bT3+zlQPZzX/u++bgHo8+w+GzTn9jYFPKSea8HlZwIM748/pW7gR1wnBYWg
bq9kQkfygWgGR4w3zOAGAb35kyNhm6eWzODNhJlH2Q9Xx5raQ92Y0qjteN92inL4FVT48UEWjRR6
cMcI12ybV8edU5HuvOTmtJ/qHFQq/2L4eU/NQiRw3J5X612GPtxzLMV9FyvPGbQly+Lp1V79BuBB
Z+tuFpl6QeflODUlqlw1zBA3KPsxh5pFY1l1x/tjrK8e6B5kN16+DQ14nUS7Yv4d1tR8yQThIIfH
EW4v6Xly7T2OwOjm/K8CSFDI/Uwg9unsfRIxOrQ9LOguX5NL3qABDGB4fh+MSnhF9b4MX424muv/
qT9GaZSLhzXKvxXxOJrqZnMPCek249y+Vj4+ZwC8UDoXJDRdtAkQ1q55+FeKRfMPknNkyOBddVU2
DOge88Zo0zDyZjqQ2j7YDNkounoVDewcco7Uejrx8srEVGPE8dyZ9nNNQwgrSwB+AkhpHT5cNeZs
MbDpCh8NBhK8/vbrv/MkveFDR4Kx7Dnugu/mS0eRouoJlFui4kcnnCiF6ObxT8JK+Szz+p3hqm0U
aRMOBuym1vfTx1V3E6A7QZYdOMmo2/BxhuFW6o+HG0UWejFog3m3vPib7rgoIDGy1fIPzdfK6Ayy
2zksPocqj/6vwmdDTaX9GFugrpIOfdFfPaugNq6k7I0yWkHWK13ZM++0i2fDaTA02GLTP2KIb1Tj
5RrOS5DHnvfaZslJ2Z0BRsURACmC7UhttQZXzR1AKFhNm+ZAUwc93yA+4Do9M0fY3g/BwvO8iP49
qxOZGWYzVthO92rMTw8Ldyuw/XcOW87Sz9HXHxyRcuyJidCPFUBIsFiJhfvBQNHR5NZ6XISrk8lF
oQTDnepav6Rw2HmllP0JubG5Q8LUA3zRMqUwwKx2TD0HsJVgpWvF2z1T0ErRZXGuc3hnzhgY+3KC
Oyyf7OqKhZPvDdwdHAlhhWZkLWY7f9eQG72yjALbhHMW9XFByKA2izqm59EIfjOP+RThqvXg0y4l
dqyN1tJqFHGPzlbHjQsRRIZKrdcg7UGKGP4f+djQY23m26BxDih+8zlWovlsG0tNtAtAc5FjsmQn
fXoYC4JIjes7OZ/V09oyyw2QvMDyVKfUlJ3jS4M+wJCc8ZRHlwL61wE8x8K84BZWVTdSVHGKjNKu
r5w7ULRak8360SXDx8p+YRQreWlracjyPDxLF7r6Sf5gSNAL85gKp4bPUfmV08kCVlhKnKsgzqeZ
7VBOJ5b/KgHodi7afnGHCxxzMOo5Ftxgr4LdGY55cTn3noBZpc16b24XygVsZ8RSrKEdED3qjJYW
qm3S2ee0VcgMuUosXljXSGMBHni8YXAZolA9l+N8Qvv4YQpn7WBL7Um/JH3qnGjBTJYOIhNTEcNk
4dCDc4ucSvSWxPTp0pebAWObl15YljFpgkAaaVV/aHewGZ7heYHrwH3h1nPxLz3yYXPVwN144rjn
ytmOUeS/atwuzaHVVNdGr1yuRBrOgwGhv6plsagFbbtIwj26Gl3S83rSYPccytYVHEeYzLJQgpMg
2fe0vTlyDvTIkybo1RYj6wYNwZ5mTzOVbgmfQduC8mCPnfRoBXbED15RhFlEL8g7249LMVGPVKTF
lWmZF0s09mbVYT9oFhGFij6U1XQhs+bp3arWQQIZ3VUrrHERf0P+HJWMfTsxS6aJOxWWIpjLc+9O
vQCQyNyWEqNwp7Oor7e06nIIGl25FhWzuIx7VKPYqDv9SGJ6TshYrr+5fh4X683FprHgahTYJaWn
w9lVszaIM1Z2LiDX0XwXgW7dZ45IR0APKYJHCA4cVGWHbHpqgMtfTYhkJ14zpAIlzAnfVZ453Hkn
YOUwqHb6MfUm/JyIXdRAhtiQyZILji4pkp96z9rXW8Am9Z0zf1bWxcO1w6FUsj+3hU5txdb984Si
T01LQABMpsDuHzpDmWGB9+PByGNv9nMIq/ETqz6HviHQ09cd6RFwrmSpCkjz0NpddHlgV0zExgUm
8BTZmKMjOolCtXkIsRbDWAFdaPx6alPMxfueHaAQEjTeN/TtGI4Ws5Du80dqHYDG2KqOwK6t8D+F
NMlPlEy6gz876U9lK4R0LElUDrZxwKC+CZ4Ng7fbvFBLNsnxzuKgTMIaezrUKoSbZuz+Kbu5bdU7
SMnXVzJ9h1tq0Ak+9nbmkA7O6qAKWyhmK4SIqochGdvZGERw2P1b/vYNutYQwwhTjC6srTXsXRMZ
k4lajiA3hSFHnvRqqTO+/xrYIzqlz6O8T3M6YWJetFNaoU713Xi4dpb5cST+v/sFkT1LyF0NIPYa
y9aOlS/F5WkmM97NIfz27Mhp6ke12EUZacfrlSoe0wbFneX6CQ9dof3qLCtV58JHUcQtKc5Igefc
yawGqDbhwYIUsLI4BTXExGCJvGVsn5/Fil9q3Vv7IxUsJtAZ4fApxkBf4ZwlrlTlhlzbrKu4a4ZH
JUViuC2UVp89fmswuF74BmpSMdb6YHwNUTFOC6C32pH6d/iCqaMEoKTtF9speX7EBOyGm9/c2uYA
EqJOvheZbwoL/r2kx5IQKnZS6K9Pthk7GjXu8TkRIFDPOO8VNjNcLnXPcl9HfBS3WgRwarIPR4rQ
Xf7MzITj3IoxJ1RpS/iAUJVb/9HZziwrafpo4yTDT5PcbuhyvTvNa9ZI6I9qhE3sHgx2JTYcHh9a
lsY8W2uL38MVzm/FMAvjoQlF6T/Lta75JuiJX668taPv9gHqASDYVfavNv+V3LdQ4NGtZWeRk0na
ZaKxX99xnA76GVSyGzXq/96IxDhEEJSgtZqHNsjIZohGkXkc78TO1PvQnrziTIHTcEnVl4Pn55Hx
Ul5TdjU2m+2BKouc4wRLdaiJm85gBIDBtdUTCmUmyrShMZB/uujsLPf4NkELTWiXeZ1KQl1vUCCB
BXiN69dQvnLEy5iDrYbUAh1o2g2Dn/OdthqqJMSxffZGgZU868gNLZpzDkBZt9bxnEYu9FITpT3X
K34pEjGitmA83HsEfHz4xCiX2bg01ODWhvzPhM4G67cTBuwhxW0HMtDbS4emdYH7mGrnSQD/JuEZ
1WZIxfe6LX1W+/jsz5unJMnNpxniYhcU9DfuRyyoo9ev61ZsTR9LhNrZ7kZvtqXFWW8xt/zegeed
3mQpKiyot3cq9EBozmu2cxJN0ik/8nSf8wI1y7tneogl0EDags/ZDsnBcUoewyYNotTPLkXoqZ+W
fR8ZV9MMIT4U7gJghdw2gf3Bw1PdL+YmWm56Wl7/ohljFF4PifbX2rbTI9JMgckp97+PY0OKPuER
Qb2bTta93NZWlJk8heeZLpUEE5Iu9czdVN7whBPVUfN9x5HS11eNjzMtG0nr+6dVbpano8ZiCjlm
PGbNW2+l0CX8hBsmYwVWLt/nLqO0qiYYswAnl/jVsmDCHIIXJxBNmmyFAbqH1i6p7QqVQvzfOJGl
pJj1cqYMVukVXepuWVk5shKfZ9mEfsW2whcNno4D7I95FAskTNR56FyhYtOYtTohoVigYDbGciPA
wvb3876Wg0Fncw6eCHBJrKvzdW0PlHaX5C60OwHO3J2nhXOnyGZPG3qncTLqY7M3Y2UTr4f9p+uY
TjNJVz0Hw2lrPAncUg3zZHZHtkG6KX5mVMj2MSMKcQLGnPB2cl+Z6hb7ZBSuCNOVaAzs4GHR+HQr
XhHR6oXZRcpxbXWNsxnfHWQOAwS6f+yjWUPd8hOuyrRODmMJzMLk3W4XUemfGkT7UmwZpsPuDSZ5
nXNr6tej2JElekKQM1psiRkrq8Eoyv9CeQhFnornUsV1C+8Xqzf8lT7Is2++MfkLkmixP+++G6Mb
5QWGH36Z9RAtRQEbfXnSvTr+fudIyMvFPLKQml59EdGwF/PKTWCi6Yrw0MFLIsLwvqGOXn7YYx7Y
JCalkcGKAAu42ezCZqdXV9DZhvQdb8NS4I6zcgc5bRjI2JIDSdTIChQ4UGAxZZ6sJP8qGI4sInwA
253r6E7fkpbbkdI/G8Mq063CN+NwoSZo6AHha67TB0MXv+REH4Q5gtzszvHb5MgvPU9+Ru0ELKLj
RT/BpjE80AxJfi4FUHop2pPErRXkhlVX4frPMBlriv8eJ1AqeVIaRJ/NBfK0EH2y9lNwlBMolzfP
mARkGxf0iDlxfuX5Mu7wnawZicwvbp+Hr13iWzU1tyEjyCouKFPFwtRcEa61cYm6QxvUeJyF1Xg6
ncSNp0Dw/kX+tVtRFzZM7xi3Xon9rIcKFy+Pf3XXArQ5uMkI0GQ9TgFV9mJjKu6pC8vwQFlg5Xjq
0uzGgKaf/ANMPHwwugWgXC0VgIBosu9ArMXAJ6vF83ikubBrJ/M0GDON39aP8pS5js/IgsAmIwHn
5A0By+6fwzB/xX8Xrjb7PGeTBkOjQNlSacEJiDkQp0inNywc1g959l9ARGeEi5MpgVi/sKp8pUux
fxfOrxbcrHZHAs2r4HHDpcd+Cci4e5gA6sysZ6AKf20vd8bpZ8V0qmLTjJVk7EzNZWMMv2rodAoi
65b6GjFR52SuyzgJz+sMnOVVGo4dYvri1jepqLlk3nyXMSoAaZHXbsCnfE7LUV8cfuSiYnLMgQV9
ZBm6RgKKrZvQnDDsJfWV/nPGR8F46ZoVc3s6PTkoPFnQQfHBGz6abLSsA3dj9icjfehBauF0qLzl
Xv2aU2IdnGAUcvvDYx2Jj3o9W1uL06bfh1OKMfKtWddgqORXR+n8XOVsVel/IEEwcsZHuVZ+AKts
WKWbrLLiHMg6DEFppnOm3LyaJMNT5vgBHG4snUh6Kbl888f44NLRfh410lv1ZtlH8uDNwunnUp5s
Sba81T6nVWhO23ndZD7lUm7MU6tKUB+r3LzronCqx77g3wKbReDE5/6DnIvnLWNSRmXw/Jmk9jiC
6r616SukQKCGdcIkOBam7+QY+Ml1VCEfwGmO7yx67zOq3ad1Zebb9ZGk5y7F+ivmIC5cHQZP6NGV
RaGWuXcDVLpsOFczSKvpQ3TWIiHHIJwsiMczCLvubk98a7BZ1ak5ueIld4HlXg6CG2PImwVNkCyY
r9ogKqamKLr+2WnLR0Pz5ClUoHc8BnV+mX1/6LBC9rXMnI3/nwxO309XiOW3SO5N695otjVcUOVt
lxJdlABuCVa1vb++ed6WQM687Q8rpC3GtD0el9KiZ2ZfEIAfGkcUy/Lhj6wZa0wz8gcu1vQTYGBx
hGzx4C88kfhbWG/HcwCiGGUok1LX2/hwdbyD9/Du6Gza48RTqA2/StBlfUaveIYxQDyW1vGLiUh/
Vth6vgL+knB/yO+EfSRmlGNgZhQGafnOuNVLuKEtJl6TScYSHsWqm3KW2jzcZWArZ/QBrj59qc6n
ozOFUpko8TnyP+2pMZAscIJwjq0zQJPbJX/Dh8sQewu0d7AvdK13Q7KazWJXJVF70zdiMHzJxodW
E58HfRIp+9O7YByuXvy2VGIPSXMmQmTdGvhPjAnA7742F0gCjK4Rc/yr2RvwrFYg/vYb9HtF6D6R
DJgHp2jkpixzqlzn9+yHOBQZfUONOsEmHxa8UubCczb083Bz6hBfFqna3818chwi1+ZiXcz7f6BC
MZd9Hk1QHkoAw3EbxiX5kluJwExqTmY3ibysfKfcS2lJNfTwvTy1K1gGUXQEcFuRJuyWVu6FGDCq
uFQe5BiKanHnetWOEqoUD/wHvjKe3fLHO3vvNq8z6quwPqV/FI9kOEwCGCO2n3IgVu3n1mYgDxnC
6Uepbb5YTlanfovAf6T9tX6FHpdkJkh+/IngorETHVjPSY0hnwEJIJzo+Umeh+InoMl2jq/t9spV
NtJaBsZJOi8LlqAygV32K+rg1V0K3u+51yLIn570BQzA6NfBKZPE5g4j/jfBAnTFF9raLz0J8ZLt
paPGfXpOS+LiPE3yVZNn5fN55Dm1yMGbhcgsrvzC7kWV/sBjLsskgbQPQkizcBS1ZxVUe8J9dMKy
xqJxvTiNZZtNvnIDFIVb75PDawSVXweBSw7L5R22fei3XJgHR6s4Rh9MI66zf9XKq4zH8m+LJJkb
eF5lHB5B2vVcrCPh+kXtf2u0ckNSbgxmqFDZXuDv4zn6HvVuM4+rpHd++X353WtaFyU3AcQ1D0HV
KrxSAiK60aymzY4yW9SfiqrUPTBaqZFj0MIAHSQm+zSkzsPgMy7aq9vr9Hqy4ZdO1lzZ2Nt7fOhA
O70DsmgqeQh7l9x1ejrCViLW1I/6AdhsYH3tHHc4lL5AT3c3WKtJgypJguhvE9Jc1VgA/EPmcr4f
ITVTLjPU7j6LgTYGzt55FHWdxJ2ohUUxf5Mp04q5OJ/T1g0GsJxEkkJuk2vS2JGmRdfF314safDb
+R4fi4OujXUIhTrOUbA5NZef8n50VE8z8eZG1lw4rZiixMdeAsIN7rwhJr0fjtNhvdY1wMUdQQnn
MNzWtMViwHwIXnQuUN3MBKRgJAiy/OUcZ5TyyJTifeb5FWQ13BjF3ebm/+2dCtxNKXrukgcg6MPu
Rl+5MzQC6LR8sMDYpCsDaTrAwvVLbUuWhN0nt58fIlG2GdClBVRjxoE2J5C6qCjMBa7cSasvyDmg
ThOQBDCX4oRqf3AlJ+ATgzye8z03urt0rqFHjSfbCUVbnojUINlOyIGXgRRoU+GtyQ7B00B11oh0
IJCJHa4X2EcvjKsm1fWdHa7hPxkJmluazSizf4cOVfHr5Uj0GRtzRKNaEkDXk9+65DIy59CTwGon
696moMQmtLkAGZalp+1pYftutQTXb1BPE9XAKXRxedr8kBZOVUtp8CLFewU2uQgpKycTWkqQRw2I
98BR3DP2vIlsH2XtyzFBkCNQTAy1GMvCrbAsTSQA9yDt4wG/SwjLJpxHV5TU/iijwo3DZkxyz0mE
RZjA8muHDRH13QtsLS8gicMAQKkGSjhwyBkz2r3AgaHzlLB4zE9IgL9s7m9UDUbqZ30Opns7KvAF
MQcKvPhMtSJjGvYN5FfgLKbRD8hZT4WnWmAE4+EedhI0t8/JigQCJJW/En/V6RqEZC/x+5medy4w
yZrXPUhrEeD7b36JTxkutn2qQaKswJCuGLEOuQHfXxXC5C6+1TatCwcDYtmYpgn+LKbCjIpngDf3
c6jSHOp9LT7bBTigCO5EJCmw8KHdnF+9No1ILJ0LaDO/RHPgsBA25MUDCShfdQcuknF9SvM2CExA
AeAj2VjDHiv54zHD24fGSlKDpBzYd94P4r9j+D/5Ln7woBi96NQHffrJTLzW/2i4fZWmCT0YivLJ
S9yUqQDTLFcavyPHvWTQXNt5gmXEXdMR5XZjTBkjV6ez7LUwXMZYAsirp4CN9rUlVfHrU/9ndFHf
jHWM9KG60loVyBm05KYnpmuky5m8td+KG1ZP7o5+jwboX8UD1tnYPcwyPdaucZ4mM4I3Ha5wOSaP
iKFYKSngnPnR7ZTBhpXoMWUnrp/A67nfWVTbSbpTfrVVdgTsXt2HHgWhHeN4Ji2v1Y1/DC39a5KL
N2L26KAlCaLC9VsAHFDdAo5qt/T8N6z0qMImWC1gchzpzJuFknuYj40GjhB61b8YA9sDIWEQGg0p
MyKOQSjwubL0r1dNBwKnGcYZFx3ikYgmsmIQt500IcYsq3tw2FfQki+0xRyBlaG0oTkuNvq3Fjw1
ukruEUJcXdoVmj0v3+9px1TYrNf9yY1uROtkFv8iHuNk/ycNxrejGD3MZluAmsSTaXznkoFF4fpg
L9NsGM7lpmoqZlrb01HHflSe/VCUTx+Vs1uGPY1u5XkDXvp0QXjOUZalNlCIas2vbELCXCNn2PJ0
VSoPtj1WHrpFhzG6MrKP24AaiYXfCFG1f23vauJ7AzArBabOboq7KT65Y4DH6+Z49b34rxo0GEDt
6Pt8R+AUp+PfgGA5DvCuaVDUs+aR50ffyjSEWSYv8oFstSg0Ser7rIvcKPrS7UZonAuW+gvT+efp
s7ZL5Ghy9yHQXc255HD1fp+bFeFQPmuxKFYDxKT0vvkbmIybaXgXws8Yfg2jcR7FUKDXAWVUOSeM
dQOw/dV4HSNTViAKM1njKvus/kcUyqDqx4CdfG8Yo8CWnUauYcaHHQiyHPSKur/B5AdeuuPqovC4
+KnNmfUJnkLQ8N2SIZic2mlw9MveW/uYPcRqVy/O1QWTtUbP4rx2laHdoahkP/3GeNPIyrUU98aa
Adg+aT5tz2d4M1Wxkrm5banfwnDyPiXGrjZRdOX6X3Mk15TQLPOpakBVfZ97ZtGAcFGshRxpoOOp
lefdw4tUUIIXHuV0x+oB0l6AzraC55hLXv5QTJYuM4EZCXCpq9fbypK5gx8SNjBAsLjMBXn9TRxg
gqAV2tehGWU/+S6CBoNviRBu43bw/Ia6Ke+DBGdo0P90fmt43Q+IDMPtdcGK4gxeBeEd/bB8Yb8y
hYxQZyY1Oxm+WXb7JdGh+GPXZwX9YdYfhFUjELo1EnCSAEVo9NaJ1rwYJzGP8v4pIyCRPV2ugCJd
r5kkFVLbHgX3X0Pbf3gIDGh1y9+R0dWGVgQkdCcCl7cSOX3MZZrFdTu4YnAAMouD4K9Gxl+lAjoE
E9FsKfC7R96Ef49Dj9il1HUc7ZVlHcnTMMI4QoT3ddMPVLwosvcQRq3E162dnBloaVBFECmKYDRO
R3N/lS1QEf+mota9zsNPiiEJBZ4qnQgQBpV/yimVvybr5wVvFUuFEsZ2JaKyMy5CQ6dAI570D4IO
b9D2foQQDxjAYO8f6dimleo9tRuBJujTgkrETZSgKhg4/G7c1O0dnhswSIy7efAM8XCDq0ZxCHAP
j6E/jURXNL0UtaAz1DzVQSHhtUfHD2eIfdMxlSMidNsmyXjyY91WYupurJJcMaOcGHjABhh1OQzP
1Cpdyww7GOb/EtOWq02AVygx6YaVvxRirUm8QTOXHkvb7iIrr0Y2fbwJwDOUwq0yLi1IPG4lPcDi
PdPzr2GE7DIc+GMRXKkebMoLoIdCJZhLDa6XE7ZN6OQz6HfbhxVxmSVMVP/nxWZ4jFtTEJmWdunj
ylImnmDjVrDFChXyAVHW9rUpCJqAU7WLKzH2BQikc1Xq6RC+UDi+mlk4jL9CdvMaaKmkvhrucx/Q
DLWOEI5R1ZKk1tvdBKMApohCAkhp7uq8Fwn03YzCNOL02LMgLmipuu91pUSvSVktK8/cSW9oo26o
4kjsIZOIPnGfhGGSN/k6W/d3QHHRZkoag5fsCJPKcTr9HCIXi6ViDeMjCIvyihJpRcibYVOXpR/g
WZMt90+gjKVZPgI3aFkQa1eu/RU/pQin/DjCLRpQlTssAl8dXYcRwweHaLtz1/AzYdVvm51TXBIM
ynABSmDu7wMPdGOlXYiZ7L4JqeaEJIzIov9WkkF6raMhC4PGSwxx4MH21lYMaFem5GZS7LypIrWv
PxZhrRyODUsYQHnn0Lvu5vsjYRf++Jo+9zRgMC9nZerYXpYl8oGR7jshbz10Nye4Zj7tVoZ7lRl4
QfJ2zPPfGrBiMhMxMIiziaRKpzai2fb1mR+2bvl1oSoQJqGtrna3mjj5qaz8WPrAiPFBvkjwDf9t
II5Hmp6y92qjLOEdttK1+3Rkt+06Hy+IeILVqNli2rUGB0o3+QeuNHITztAO16YWPQ97K99E4RZI
pS5i5AlUbnFJacAGW6/oJ1H+e8+RaZ1bKXcWqvBsl6+riYk1vIFaoyeFBHInQwX04slHyW4FILFE
0DtNOrfcscqChH62PC+pF30kHxAZcIXDtLuHfz1T5JbQX9xb21Zoye0JEks5tCf2zn0uXwJWOlKM
y0/IUQ3Qs3mj/6yIUsHlWc7nEM+oNIwxRyzjSMBa6Y1oadkMe4iWNO9b7A7AY/gKD845g2pJqNMO
oVW2oHhYuaOZUfzDbg6HcebLOV0BDPSAyg/cI3JFyaJA0V5tb1uGtT+FXxkXQdiyh4znQKQ3vLAx
IA8KsLjqio/8GUJ9AMpKF//QSSu+borN9K/NNb/t93HCgFgad9f7sgPzGmgYG3hfnZ9C96V6PHZ+
8h/5xcz2TxOvsALbRX/NF18Y89wTn/KxkOxxhAnt2yt5hFoRD+k7KYDBrZjoqHybb3d7AUx1kawZ
5nK0iXQJaR5Gfkq89dv3v1HK/YzMF1j0YjWgvbCHFjM8WtzVVHKoum6uZpLbNtYaBRT3iwljC7p6
8TsIEOz/bxP7lE+lIQddVwnj41zUAjzYiLg3WlK0UX2OQhDyp6aeTIvmNCkXrorioF4hetvt74+P
yiuPACkGvUczi7WN9UNMM7ZMuu5CYUBVqJBiysAugMAtOa/eETmBuy9qMn2YuNJDXVbMmm9yMMHG
jKvMj5t8nibBQKboaO6OzAFhdChgIoxmoSGXGFarCyIsmhhH9QhiUt7WUsLKB8UT+/awKu56Yiq9
54G3s+damaTgJkEoVZhAqx178Qq0Lqjre3RvOUmMFyQgwJa/r4RAl/a6PlaIyLVT3xdZJmsjJgPG
NOwM2J0H+KMMyjIMd84Xq8ZlG0uTi6wLMFX8Nfme+pshpzynZ3llufqbkOju3f3j6/ZDGf1LU77W
K0I1do14O8qKvl1UMjiOcaClDH22l/r4XV6n4xpoLB+odnuja2kZiClqEnnINg9aQzZ/C/71Xv6s
UnFdf8czRrRZY2EIj+dfuIr1EBu2uYKvsZ5EC8jxCTg+IMU2VUq5SS6OS+aNVWa6YZa602qLufMK
C+Dseuum3tVI8rjlCGvjsmEM6avpTrJ0HTCEkBYwSnDQGfpg1IdasjzfVcfLbTzeZ70ro4XfA44d
jJgvXE8OfM34RidVoFZdsgKSu99x54rib2vS/mVZCLnD6kdMghiZga1TKACV7QwtKhJ3vaBi7zhX
1YUIyvv3fm7sbxSmZZNBR+8Y/VfUicHaWHOBL4qbinSPcTUCvqWhhCvJmKEYLP2q1wifleYiZSzk
tSMqmJO4mupN6459VUaa+qpHPn8TRDHOjt/Q7HMvFbaPFq7cDxB5VgTp40GMXdhGNpBVIq2Bzquw
TT6kndtek8hPB49W6OggBs+0zEtBYSvGmV/4GIJ8k9epeKL+VkJTd6Jq7/LUB+R/ZQhXywelHb+A
BQH6cFqjM4SniuF+R9PFL0cg8hM3ioGwa47Nz0SbsiV/cdGSsGbe04YP/zTauR+EEF5AmL6Bqulp
g44+ii6DsOwmD+LBLPjnGM9XLeB0/RNqecGvk6J8Ok2NH5jw0zE02pSMlg3VHg5RVdD0OL3nangc
UHCEi3ldEKoc/ViXibSyUZT5hyVfOz5qZ1TBR7wIgEz/zHYL7rCXmmAGdsHdSOq6Iy5LyZmfRBkz
yX6+Y9rcxqkGGKTNqXim2ZoJC+0BzMJgI+nKG3dlgDSJy0dbuDwXZom03JfqeKqGmnDYfwyJU5so
NAvz/J4K+sFL85huIivVsyR3nGY71H9r9rebQqdavYKXgH1ubGok7h8TsRox9StM6YvXwn6Y22hW
s+XzHi7VH+kmnqGu2QVAeEDkby/aw6EaJY2BklqBDiR5eh31+7hH7JhoAqkiulF6xcU3RrdklAVx
aFa9MxIwXNgsk0OoS7m3lg1noTBgz3KKlXyjv9SRHLZcYJkm4svO5anScD6mZeMoB8Kx23MZ5UIw
9HK7pNKpJU4wK/FwqIfjhuuJMJKrnswg5MO8+Qp0IgAj3IFONSc/UM8EBgNH4noX5W/LicDdPXDa
2a5vd/jdbhocL2Oh2O16z4CI2SgyJJjSwrBs9E4IgWkQ+pSUtWvpSeSDEBBD7qMiShFP7w0I15w1
Y1UEOBBkp2WGFTu7fS+HY7sa51O+QuSVefoTr9+EgGgso5QQOnCRpmv6KXsfIVAnF2bTZtfbALKf
hNcKD+hNBSkttugxWhHdHf2324K7yudHxWmg6DAOkR9fDIiAcGiATeYmREpjgYqVMkQfT9AcYYHx
nSAOdBl1fpQJWocvbIMh7cN6DPB30Zr9BHyKmRTvnbcUaXA2rvy9HXEKJjyH3Qyt7k11DmJ3RPY6
/6iQJhnGmIZy5VkIz5+Ici9PahzpwWvsoRXhQJP0sTP816tmWz6myyqp9zxflNSe7mfRj5DCZ02p
qf//vfc0ndNAv84Eg3d/qkQFCbJHT2jv9eP4lI/EnA20qzpV02JKknw0B8ElyWTuffM72QUbzUSZ
KImUoNOwLs6Q8w9UT+OgqvybqnTWhxK+GsM4U2wfOSsQHtX8fQp0qFLKD/Rj7Mey8ynFcPY9vUZk
0zavS5NZ2ltjFqrywylcFwDX2mEvctWLZe3uDQWqP5g8JjJdh/3JsyHTuv4LbX+EjwL6g5UDUVbh
EcZ8/vThA81cvl2XLoT/bGOqzLUgKDkMb9d15C/rS3RUjsq+NGKMeS8Ji7qBsDKTlQXuLicaXLq8
RlD9fXvBwnV1WJHg90+8w5LHC27Wi9D+bHUnNBoLRLPPWzcvp8kBUdncmeR3Ork/XUWUDeWGR05n
BUxUANctLfb0yWwlwlTYH7aeVmOwxq9npOgrh6T+mvCnsPdacCujzW+q4jWtzPeo4zF8frnjLFdR
soQY04P48JmuI5adtDY+stEuYD0B4rLw4/9ILq6GDK50GsqS64b/6CZJaEavJ8tr0xDxQva/ewHn
sF+Ax7cvOZL47ZdZHhF3N8chvlB+IgKMY5jrcoH5dIVQCJPhsB2K5X7nW0Wcbb4FpOO50E+IHEqc
Vdb+xIZI9h8rMg285OoYvnWFvitQG+2cf/LHmbne3BRd2XnPqbJ061RtXaDHDvzG0lLjQvUgbYeT
1aRoCVI5V8w/gQOjS/v/kNKGNW1BXl/QBf14dicG1kXNOHTHir9kCva3RBoa/Z6Q4bre5tsJEIcB
liGuceRZSyU0t/gN1F9FOMGDh6i/sDtymSttKbGf0cPSp6tmNYCl4dKlAz/6ww3239ESdS6z4/hA
Z476d/FHoj1ruez4UBql2n80caJdbtoOtCvfJk3z9WwdgymwyJWWA0HhT2G50vsPxM8Mmqr14AMJ
SzTa7sa3ZFU7d/KvMs7b+BC1SfsoXthUFRjT3LDOcWuG7b45Zb1IuIyEZrkPw1pS+0OalZ2uGwom
I92AJgQZO15Oo3XjNew07FlUlluJzNu5YcgFTk2eDAfboeiGcgXphIrwXSwih59SkNAE0PwNAoN9
7RRcG+jurdv/hiFTNiKtLkQxanzVI2qq7g/Gijvv7zhjJKt1qtQfcgAn+NBYOsUoHNm7SoyEWm5v
OblHrbdsvg44MG+TjFQ9HZd4opYaLnB4cfWtpYVEWPmMDMLtY3kppcaCAxZQ90Z4QZITXwhrPAa+
klAzz2GE0DTn37+1FRL8zeV/g4fqiHEOVc7C2+7WAzkJs9G+0zwtQgxDzQ98kBhUYokfamVrO2Ik
4ezaDyRq6FCbKZcNSvDqMJRws/rqfm04nao7Sp7drRc3mxQPRf7iy5yLZnrHASU47CPcr/ujwQ+h
1p7RuLAaIWcEF1HzUuVkcwyyp7yiIDhfgtN6qHh46bb+DhOYlsi993r46tr7kFEbKc23+4Ec19al
peQB+fL8CSuFWLKgj7j4eUkXPDJaS018vvzgHvr79S94GY2zqSSd57Pjpfj5riQ91wGAgxHczioB
LtFLISDza++C5cpjrijmiAu33zeWCeOOyEUEXpLqG7qNKPvqYWvr0oQ2249Hra+hg8OEXadp9Akj
q1FvrfSnwDLOfWwBWqXVdOyYiBisHrMdnyg5aznR2/ZjIUXhyvpgzoZkFQqkaSP8PvBTY9IQU/NN
bwW3UF9fvRX9gD9sxTzHunH86B+jooD6iRDVtb1zz58Xu3GShnuLWXUo+nLspbBYw4889fcVIge4
PIgjNTxBm4wsTU/Pr5IOhl5jBdPQ3soHtkyOkIq+8GxOVd2B5qZcSsSVUOUcEyf9NMY23VZRRPCq
elq4t32hIob0ar3gQOEAisP5p7iZSiRLdAdmeHS0z6Pg9FyLEQN0i569cInCkuBtEZS/25Ch/9MT
44ZSSxcvXWSwj/eNFZPiHOF12HeF6wi4h33q51VoseibiHYzWfWi8RND7T0WEq2ZT4er/HSeWrfm
5OkEopVRAhzN8kJzVPlpN3cXK4noSVK85ZGxX3vRWiMtlIgCiJSMBzOQ2Xnvgt0k2C9O7GS1MdW+
lkCaZZxlNzaZpf7zb57hJ5GQzEkZ5NVQpv3f9ltU/qEOmbrwUCs4TrJhkoi4IgdoGWMZubuMLh1+
iQIzqrtcR7rRs4ksARdQeXfaxwNt/8P/Xg+67wIF6KMDGNJp/WiQDt0QcuXbSdg6UnYvDA65BpN+
8xkGYSiWLkTrFdaGFdnH75oxlFbFsIHlL4jimlnEYqSdvYBj+3bBth7iVHIsoPCOf5dr742wgc6D
ANA6C/QLD7xt5BVbcDu6IF2BioJsGEuSSmsFmLxjcRg0syAeSXxNlK+YITKndaAzTGYdbomxU4SG
Pmsn8XsXtuyyL5ThP1Ix5iZKZqZCaND8X4TaIzsK1KEScIEH1eQ6bObzEJX8cvsJQmcswkS/SWmI
e7WcQfIzv+/FVMyCGiuVolJsSyxJAn99+uagyymoMahFUOAZhpOlTZb8tMdtTxtXnC1LtqXdSlc2
8GqTWSrzZPBcr8mnkOSRL7Ujd1Ck+pQc7dg7r/ixfDBvJdiRm688DzOmqK4645YI1fz/Q7kPPv/I
Wt268Kq1gg61wAR0aYtnhvDGN0ozD68Hl575CZ5wdbcG5SXUNjZ6a7CSBJjScmNssXWkua+g9jh4
1iow5nf8VJynQb525Q7HVhgspZHXRLSjsc+nA3/AjE2m4nJDj2CdgE8L3u01kV1FHfoJGjuD6kj5
dznqBffwXDDpA3UKaP5qudoDdDrM8fALe8T3M9sE6U5WSgrpbOBiNYXgpi+jo/xTRhdNHJHwbpRd
MdHCcdtLEKhqa/bSDxv1uSOdffjjUwl+Z1+//1bSBz8fQi76lhnYUe0ue2O9FKHSqRbVnU10Meh9
FElKAmGpQDFlc7NroRTV3qa/eigONeKcofcGLtyKX4RB74X6KV6EXQir9bVVcn/UkfJdSDVO4RYK
ww7MK573AeOBjVZCtAByx/yTPOaerfDQZxOXXQcy4klvsG6TYFAqYlbydOMTA347slFL46UNho6+
ZgYUwVSnHMA5kQS7mUSEwWY90GnA+3iAfw+xTQ6CFMpOehdbEgz6nR6Sq91XoOQAWcHuQeGOzTxT
oMn3LPG2zJjhG5qegOGpNZNAbVrdNrU4r+G39I7CEq/nknGqAQ0/tg2kVmkx5wgZVjM82rk6ygkg
AJLDln+QE4XKnKoMVeGZ0YBAhDX16f85OnDKjovYu+As6ok8klg9JMBk+oIwXJ2siocx3qCb6B8J
/VnmjKkcLMGtb/xaRJ825jHYDrzNsaE5iLGwEyiWedQlC9Pjixw5Inj663LVxJNO+tHOpWYhIhHd
7sOLE/gOZHpvHYE8UCjzRgnlCuv/jepc8b70Z0TvRhrzVZ1RikDwsctK8Klesw6PSpU1lbKyYimF
NFHZjCiKRy0u33JdlG8SG7FonA52yTnJH+pJnoNdE4uBL7VwB1wdcjkLA+YXpZP3t5qq769hNnil
D6FQM1hPEMU2MzuXVa7qRALH+Gfja6JgQGets0zxjH89IiGkp6zrro9/7xuY+CxW28L8anOi6iKI
qIN1GjoAYVcX2ayz7gjcAcC75yetmVqA2Tkf6xrajdc6gMbaKr/HJmymXPRFSMCbDvHJgpanUyEz
hpiNy8ZvOhVTNtLR0xvUtPYmp+jh76bZ401epM3xmI7t07i9we0AhdHhFqB9b1dvdbF1rDrGn3/s
KnIgs5ySaWp7GGQgsgGj6BtD7+Xuqnk3sHhiJWZFH+X5PkXuX+B634IkKBVvUrSRku0gttGHNHMc
AY9g7Bzqw+118JyotEKmVIVjn9H+ExtsnmSusJbw3H/xlaqimfddUBiU9Ghch8Xt9moj8vSQvZjG
7yk67TBwwX+cBYwLFfYbzc4ldYYlHzT8fR9TKqwFX87mmKNV9mn7jD4UXiWVioAKnqqalme/DLmf
SmmFCqn/tLQVKvXwgeCZSUvyx4ReSkrSlR4uJfRv6Z1JA/G49I2BKoOYV/bBu06gOZ4ub5tPe8Z1
mkmyzF7vmKqXqs0bsg3yzJao9i471LhhI77F7wWumHLRtlMr1CfEe3N0S1Gj7QW0krVtW+wU3umP
1zrXXPxVL2H06LSVWTkDIxVpc96fu2iHks9GPthf2ojhHhNlsrG9Ln8FzY2WSHmBd2dTLQNmbzt8
q4IFrbRtYjn36beGSZ8QqilRPfAGSzc3qHsGsOJRmym6tJaP8Knwt9YMtnLeNN8mzYWE1VEedgtx
ffw0IX9EJ9R+08HqlJtj89FuEIT6+CIgbLvmGbwD4O0D6OvNvebGJaB1NdVQIoqGJKvN1snKqXH0
kGjjn5KRzou6zNW+dyx5PzIhcAa0SvVRWbm/lYxBuKNDm9rX6ujMuOr6xPGQYlj4Jzv7tZVAXHqN
P9XUu63tWsIZ8OHD6Ow4nB50wBd6rt1u/nmPflbbE1Yr7Qd2kGTC0LxaiwsEKqT3PJ84Qv45HN7N
VVh3AlDSrO7dT94qgE5lLLqgiikZthjLjuu9YSVbPqvS/aaQJ/GxnPkK6vOklzDbEj++wsEXw2vw
g4sQB/aEoto0wCKgKqsg7dYwqcmgqudZNTi75rQYdU3dYf+TuZsrOOjHPk0vCuKcpyTwIQ881PXp
bCMdUMqGD3aFr2vnxZSzQrY7umf6mkGiAH6ZIL6L3Nrn6OANVaTEwRrcMzizXjaXNWOGtZhHZfb0
V+vvBG3LaDKefdyxPK7Rie6r2q8oy/wjelBv2OjV7nL+5MLjsWeFHhPl9OQ7U4de9Zm7T8HbAS1g
/e70yMv7PEVYOtI/3NqKKhUQ5++y4aYBdg80FIgH6MBmxBj9CuoeGh+Z/AsVuyD4GdsIS9m6TqFQ
L5dgZGStHDup6/lZbhtBwjUA1Q7KHJiRdQMETSRbpUPtlFjQUW0JlDTssQIUFZyh827+a6zVdw7U
RyT8kxPFGCr05kZVzTwv1S0oWnN9SYpZpO8S0XjBAwBuuVVfYKIPNE9/PwNyabLZhDicim2mfyp/
KO12j8drTBNmc6oK+OSyIJkT8ezbEBfuQH5YNcvGbGJTiZi4KOMgn3NUVeTqpyY5Y0hS9RhP5G/m
9hO9XYzlWYYArJcXWjZEDjl6DWioHc/KA45ICxAuHUEHvmvQdqnTyeDMQUFpEhjoRzd12Z7lE+dA
+DDaCU9NArvaxepJfzGe6mTDtDkWw0krHCOrRBvFFP3hHTWqhlZvE0b2ir67ppsGO6nA92O1MVCw
fyaf8Eu9LTqyQ042XOiv/RdTrPley/4WrgmcIO2zjynj9rFKdCfv85bfmTn3IgGVz4YeFcmlsGWl
e+/YAx2irDNS0ZJFWi5kawJLfVtoibAMfw1SW9C0a9gLFcBmh3S2m+OjBqblSLgcAEUrq4RR1kvZ
7PuZG8mR4l4j2Fdys5NPdGou7S+veiVmkxT1XuhOtzPpcUmB63mSZDN9EcXG4HaY0/702RQ7k/y1
MF2nVk1nE7OYwhDyDhzferrfBvKL7ThdmhYHJ81hiCJc90s/lITp+QztiDHWrYqtU7L/V4FkLSS1
TYbZM3xhlltsc2LOJsWMh/aBsZbENGSsRZpReNMyc5QSbUB7J+JqP/hMtpXi49t4rq7Rx46Ysc7H
fUpJx3ZS5y5qadHsWfafYsPyfzhTA731YkzWvjPX9kDgrVwxocrQpOS5gkKSqNWvGecAq9ordcim
+28EqPm6ntWseS4df5Dgmk4tVhl+0cIJ2I57FID+e8Zo3vWt66LUclo6NX39N1tlKEt3ZKZvkcJB
wKyN1GykN9nKwA3G8I1PHRHZlcGIcAYPo2xQhI+0zly47yKSQ5gIft8an3oOJ1MbQq9jNHeddzVf
u58Rk5TKn0FWwgluaIfEwZptDHnzUtZcUDe4Sf2WsvVJiTX+V/u1S++MGXJrJJyPephk3Mz2hF5G
Q3Enihvet5q4xLty317Ue6JqyphJDjcGo/8ro1SyTZ9bCBlo4SnyKiSXNpe7y3QYkho4qrahA5xv
FSLoFtGKnRxQO7DhKP917PXySyFGw8nlBrprzdXEZYXTauDyjlYkINshRcrOVN/lU/BXOyC4ve4x
Hp2qKtFqApxbXbV7SHXKppH6duqScMFUJOnSIV6M7wIR2hmBAoX9Tqr79CO4iZxdQILnGcBt/sLa
y7gTyLuswaKbt1HlYFpYuQG/2dttnYya3P/01OUrc6NrPpTaJ+O+u7isrSghZe9cTcOaR/7DcYJQ
d5QAbcc+AiDPRW2wwadC9U+kWR01MdyvGcem6nbs5yrlscn1B3L44EivsGxUrm/4X6Qo9SB8Byk8
3cfWSmbmMk8oe3/sGtyfESEgZgtIVO5M8TbVfmL8N/pW5lMO2oV0pCRCzkitbv+hRvTcnixilth9
PoP4fyD56KpNCh+8RSe2OUe4/XP1KR8CPGaI/1wEWq/1lSU480KfSmQgYh/a4XKamYAlpWBw0RtZ
FOLyvozPSywhFeH09Dy68wDdHG3DoKguxD8+q1mRtERw41+Av3p3YF6735AOq9kWdrn8BpMpVXPX
kUiul5Ve4NjVXbNlQRTdEbQgCoJLhu27duoM8rfyGtMU7OKBPewY8FMRn6VjeXhtMTndCA3IwZCU
ECcSCZBAIQ13mZCZnjGhQNZCkZwZp5wtVnU12eltbUn6qtiERARkebHg4bj97bXrGh0kC6bLgmc8
/RapT7w3djQ5fxK6a09raC/7Ho6zWZ6UfuwLyi4Ovx0JRQ0S7mpJnHUZKGGrXyti9pNrSM2XfWjs
9lo5tx/vWPuy/zYtI9cbj+aIOSGW7UAWYbH9d0oJtJzolqF5gv6BgvaFVZ83Sr4/MK8X2dLnUGLo
kw5HTlQQiVoyZ2amKXBLhSePExKGa130YumAVDU31ok3SIZ/u4O/+wo+gO0Mhtau0IgE+cBEFOmb
r0rzB2ApggkRp5Kazy7j3gdA/j6kLiWSrsMOfe/CU3tKP9jRP1agJocOP8/OPiMjqDznAtFYF+W0
0gIyRsc2BW/6xcK0KT4f4oFLOtw+aIN+JZ3wvuVkVK1JMA/l+VOHWnDWwDH0jCpyw8YzJ3/J1sjG
jMQf39CQ3SDaLDiQTQ3rqrKLTjywgGD9Z7J8pJGRgtNtFqYh0snTu/rS7KzYxb1Woh9Y4EPZMlbM
yUE7NQIXJJoSGYugM3oeC/Our6QWBcVcc2U4H7mLPpgfQHVdOvfSwelov5CuXCgqjEzqt3a6aFxY
GI4yjAJbN59sHO4UMR+uo1/JAs29yNUK7Exx3XV4uffvNfKpMcpvCUF3o1t4V2z7U+KkOop6q6Om
nM/jOecE6rqRd+Twq5TfKk1dCuI/4mQJSxN7dvUheA/y+U9ATATwQ2jSZqH2Vh3vnqsMD8AsOSm6
b2FvB9DCqVsHL1GpU/d8ICBMJcijIKTuFmOYlvPe8qwgETM2efBsPwhqMbxDG33hTMQPGQF/p9D8
H5atLPIgZo4o+eDuNo3GuF3j8gHQLBOL78pcjkJZS1ptnygMKmNbGckC9zNPZ/rgiiuUqFbhM9eU
kIeUjPHcw6faoWneL/AQHoVdkxWGVVedz4SpIttJLYgpruXO/H/wbpPl0/p+xGUXwEP4/jxLiEwS
xz68s6etVO93xFeg8SXRXknuXPwSRyIxZJ5x03P2BoJcG7z1nmVk6a3SNrf9/QcUBomF+qgN8CtE
9u2tP5j6u7pnpjk/J/eJzWA4BavxNV9bY++l5XnzU6rakqpQnjoMXci8hSHCPnLTSsSMkHDgsb2i
FZg7WLWL1HZEH9tuYe9VJgVQFsaGFn7ZWjIR1Goz+SfsC47GjDZtuMm3g7/MVni7RStZr+qsvXrQ
QAJA6aCio0Bqnbac3nTAHHxO9zKtUHVOO49YOM1U3k7Gqn1CkjtHpfzN5hPCD6bbtmyed2OrMNU3
eEUSMEjHDv/D9IQQBrKOtoIf7QVOpACQN7t/ozgoQiW3SBAv4tOl8WZhEvJddDG3mnrXQxaJNShK
KMSaSZK5hi6mpnZcCBGaqrpp2jUEvJCvvyntDXkn8U4ZnpA0jNcHbawUSUMgHwrW4zLYN1V41LdV
sRkuj6rmSuRwM/YUqUq/nvHshGLt1yWaePn6r8shotlQaq2NXN4AFDZYQ1FrOyO4LfimYV0jVdg1
MHY6vwtSUpJUj5tL7eqXeQMwLYS/4XnLnRMDSCjamyNig+QDLSMvqP177isUELBlECh6VQDYSI/S
tQwFHaoDbjOS1dneH6d6AQrZMx+yWNDdinyaAJVgm8TZqWe91g1YRgp8KG1eylqZHuMsa4N72awb
9YYK7lpzVdovi2foEluKhCmG/xMz5clYKYyxKUGXkE7qB54WONuKDbpDTGOjCfjfPyUKwJ43JfKY
Dl8rhYKa1Boz1aHk2OJ5d4OhpgHsPw702OaH4FYBFqO3bU8s9NbQFIq9NDHicAAGbyzmjvM6JGUa
jsqOe2nC35EdzoZW0BbQahb5bjfDMXmeAKYKUuIZOdoLRowRyxij67T1wkItI9pAmWq5SqE6RC9+
AZOA3z4uUSzvwPpe/PsjrqIYhVjl8EDKdLswa95tAlKFeHFUA6DHX0JMFU7TG+gYCwfY18RVIzfE
XoeFgLEK5Uafqw4ttcFY495qTmgGUGYDFGh8LIsJE0UmAXbPx/zYcOFEYeaAzBd85qkUBhexjjbG
M/GHZLfC0qpDgv5S6GqL920u2srhqHXSBu9nEX9gW7luH0fj/BUp7CzxxsFcfveKq0myJ1eghZcj
fjsSnF7hOuLJG1recl62nXl34CxNfVsetFt58AhNP7WaYgyKDmQ9GwrTF88zmFJYZ5FU6/9U7gtA
++zqI+2AXQ2Nt+xWmEGnvKgCtO/WfGRWRnz0G1OpE222wzJUwLnNVFz6oJjtThgfQLZRj+Jo1hfU
eG3SbZ2c4c5AlOG5JssqfWn9SkN/bitiNzinHqEAbaApOvsuzpbXGtxpuMC+9iwfo4eO5+DDD51r
GQP/TMEHAToOZJ32HXcVoENzJu7pbV2HW8W3mhsCLw90/uH06HQenkHORajrEiKqgT3VhJL3PvqW
mi3Yb60rEwgrRCSgDoimhLuNDvsJhNxWUcKf64vhSRLfnptYDrC/zOHG1Sso0QIlkum0exuDTSp9
yFUQmzJmEOVjnB0k21VfFOQc2VfbowRE0/5W3+Kv9tZlO09GWilQAKLmJtQqXqTH+l37Zrjuz0vK
JG74S8qmRlA3C4aDUy4PAscSPH30HDbJK9dy78zCa9D/wQ2MlvLp4FdTuC1RivctaD+MbHN6s122
R0ujyP8S1PRFwmgN4pvjtRPfvSv8CIEFjAlLaUGZMdD8ElA1tBX3oOYqrh8QxdG+UjLITfdU/DsY
rK0ToqZSoo7SRupQimzfIFiUjGIpkyyU0onX0aGMDWG8fdKkjA/AoO9pmVA+umBJ1RZ6SYrVMtY1
8IPdZytsae1ivQOIXcIORcZaBnSOOMIyXR/CvQIBLxkP+fS/Aqm8Sl0UE1AZmCSOSScHH6fCB2xz
6XExmE2EPXZkpPqhbk/2y64KxgxCiy+WdfX9Be7k1hQKWKqKGaCY9SpIb7JAa7pE+FOm3Yd2Uxe6
sFPjqUGXVocYD4TjrF/1p0LVIcTa+vtQboP+UBXR2q4pjpAI/lhRuPnHwhwQmbrX2NqzQEg+1n7j
4tKaPcPgmAy4OrAHWIpwHJsr/bTZ4V8nnBjstSHBmM4CJb6DQqCfba9gJDxIMoT9gDl2k6yopYT3
/R3PG0TgAHcjC01OWBasPP+CIqAWM2ET0P+LN5SJ4z8jtvam3zrCUvCaIcXmbRn1qcMt6+GJpS+O
LeBAMWphyl1HGP8juy+AxGkxRhx+goN3B7OIHK2Q84BaSDqnPyOW3O6+L9+nSHmuzJ6p8vv4OhO1
Bc73uY1A2CHtcsS4dxndVRaxsrJ1Dx589uaf8gF6tNbNebiG3sdpDcoQOQ+kgPPTHPIaOlfOhER9
WMCm9dtcXiweIi4644uX6rHhULle7jEyAx4Xdas1Gp6Qzib7BtCU2HepxF3sVxPyIDEm63bGaNLr
OmHou0Q8y6h4o4XnLLnpsZ0jisRlS8x+/d3bPbyjuu0vm0rGlXHMRqdE7Zp0+Ngih1ZOp6O4YPQ9
4RGY+lWX3EDew0r8cbZ/tOKJY6xVs0Up+Lc721AiVHH2fKQFXvyki0XGTGh9JRfKCt2aR0U8QWJ3
xYASvwQJIzDgTKXmJl3J7rjyfvdb1DVy+FdDgYYKilu2cxTQ8Xe5HJ61H6PKPd0rda1xPOr5q8jk
IrDiN+MTfcNaqVC0YshXDtveG07Cc6lcNelShxXR7uMlDkX/Dm49AQV73S3AJTF2GyxQFem27kHW
6Gj9wRzhuyJmBtqLUoMcuSYAAbKJV60gclD4Kn7MDRyWjsw1vXwUR+bl9jYCpZ2qRtlKudZKYyPh
EMPSqtAu+o9CZg/0lNH74t2MchzDJR+25OBw0N+2USXxJsbrDMbnpB9a4Vsur1cpjfU4t8G03l6i
NQGSMLaVUZ+4h7ecD8lm1OSRixvdRguGq8sKpAqM5IQgSDQNNpr3nEF5IF3yO7mpGO15zfCVfE4G
djhhjjhHN543eUmuLcKwIvvf/zSf9qGE6eEwUD4sz2PjTqAuete6u71Id3HEy3mapiE9gVnvf3Nd
ehKIa+Z7hKoriIoZrd1EHQ16W42f82oEGvkYbk0d1RecpV9QW4njZ1LX8kT7IRLdtfk3iDWK7rdT
sWSke7+TxDqtaaNQoyU9fiaQAyXrCR6Vg5EY4BserFe0OZQCSB/x3wFHTIchodatNxTHcN9N/wMq
FS1YF784cTKQirsRajNIke75CpD3tB8Cq5pg7DwgQ7ECHYcs8rOBSsq5eFjcTKzdcevEpLdG7J1W
cEzRduQoZN9FIGWIUhE3ZDYk5qwFU9xoRVt7P7ff4BI/L4qXXlb+ptcBoo2+KVje3MM6AfZUXCG9
lVP+eR5k3pm96/33Y58dcHluUKa+XWYX5oqlUInG6xaDNz3551OG72O2sxpxsXj0UHNpHKFaKXv4
wTkMGn+m4zlEVwcQ/HYoKs0NVFaq32yTUVfvYooQHY8cT6J7PtMHmd9k2QQmYElSBb6TYnDmtLf5
aXZ3ayT+fEFYkHOyHSblgIH7Q2Lqvnz/6O80+F4dcw24B8fRzCNpW0G7Eych/pnvVBrAWsR7Kvwd
NcOeIdaGd9pjQYchnOXm/DhmT5FKLcZf6ledGZi8e3cyz78CxYa1vDLZdPNmNv5s1CZxq7lGarTw
VuXG9j3DczNFfZ/rjpDGyYBGNXQZq59lG5dEvfEDfDiq74SaStCN6xMRLq1nnjxG0xx3RW/d44v9
qs3vwxvyUUB5zwQcKaweXpOC2o08zovbGMRkOkhwYux+F1PXWIBCEuoNLLHo8pIXZNiwTfuRily+
nipy6V11DLrjLJlD1tvENuUpEc5NXWSJ49S+qd70gVD4jpCPdJnIYoaZtDswIGKf2W2XeC4fsR3L
rJ8ArZ57mu6Ng/XdBoLPRvQ7TqdhktkD4u08E6mrJvacu1bQyCOOK/8cfzS1tJTZxEGM13QNVS5S
nA5ewlOf/YQROJnYTFtnTXwuzQCB7KyiJtkV4OI6zMOGCR08ZDZ4SpeYy22medfbXThxApNXeRn4
1/EUnRuS7ywbNqpQNVVs/XulTRePz3+ZagxfXl/TzVSOt1SLY8EOvcFn1RDgH9QpXDHxA51Zjuai
hqqLJU9Ug4S+qkdnDYUYSlXHRTZCbl+3XkJSInFKY7EFecepd9DhUub2HohiooGFT2JhO/igbDT9
vzUFNLPlxewO5pAYSTudWbYXnqFBOL0QcKzUMk66ykcfD7uspJXUHviH0031s4o9clNrZjT/M7K3
2MegvGtFhSfWKhFqaHxSJubkucV5KKDhIwBcgmdFqhzIziPRCpECsnIi/7CCSqI+f1wqP/42j4Td
3qa7YdF1yDFvVXoca+4TsFocfuoHZHzliwurD5u2+UyB2bU/rsTjfz3HfKhxpWoWrW4m0RxWQJqW
YMDuLmaJcVQA94S2+HV07f/2LxMaS/MqY6rZBU688ZI5jSGxuZWGsvhpW5sz8ZOiPKP1CqFAwY9P
ZjXiiUSTXrK+auvZ66Y1WulvNpssiuvBuawc3l+pSvg71c7ZJWrI87eI9nlDeqX022d2bhVIlCwf
OC7S6EV4imsfHZoo8ZZ4NoCchTNf5rzLRWrZ2ez+3969/UiW7uy3pVdf4RKaTG2F2K2zlbfO1KgQ
nbsXJ83a9anZADxWD1wyw9UORQf9uLTpizO/VOxIiw2Yyth/9ifWrMh4/2kHocjNzWYIr6wV4oSf
b2J6/sduDTa31Rwg2WrRd3pt9DtMRA66I/a/dzIHi/xavMIMwaSzsyTz5Jrah1WxVxSZ492MNxF2
Bt+cA9Ywxw3Yyi+DstsRbbdHOKzql4QSPIjRILbWdw2jv3Txs3v+M5uAvhkwVl50NYtz4SDIqA3G
C5XvAnBmpRXOmWnp2JExNFqnK/LhY5ITRXKe3kTS28OJiEdyawYoyglCc8kUw0/fs5VhQgExe/sv
EMyPvrjH/VjUUJnIdSsjJltNIKIowUHJn33AeAIMoOaPxPBKHS2jLvJ7VobSPF8Fcjh0kp17RTdF
R+XOEmgpBU7nvJeJ0StpuwUbWyMIf/0juxBFg8oJbxw1F1yiTK/HSUSLs83rrkAeaF15kMe+ZRt/
bJCNVJP0QflXpaovR+6+Dlgi6dJXr0CgOsrlcWt3lHYsIvP3oxESHqM8kiJzuZF0v/ngeL5zxGlJ
1FwsOy2x+ki0Cxn+A8vgwC3dY0TM9UEopsW1CbklV5i0PO46cGSfG8cy+7lCP805luoRkJsmR5bL
e9vqsmuspI1ApCe0SstjXnMS3H+CUQTwIX/rM+DCP5cCYEVewTA9gSRYVO/UnMEVWjFFjFaQiWIb
hFXoqhuHjEMf0tv3E3pDYcsUjhGJNcRY3o1ak8x5Ze3rEPIq3HF8IYrCP2UokG41/Q/Dduhertxl
SKNlDkkgfbX2nJ0Sy5NuIFumc8cBnBweGQSo8GenD7GrqF2ZWYfDErjkN1JZqwUKrgHOfYNaszJt
yIjDsXcNjM7Ff/yhwsuhvEhfN5+0h1bvWMxfp+XfynXseGmIEr4mmK+514Bj8qa9gxFLFyvqdQDv
ToL9+Onpvbz8aGiSiUYc2WAFiidg92VDCszS777pRsKNTbb5RUP3xovLZfs3jV6zKExdRLga/UmZ
bKgfWHM4b46XgkmuY/rBZ0ujaB+wFn/eOd/MTGOc2XoiSCzc2q1zLKPAheHgup+dIH75oKVdlB9P
r/ah9shBc/BKO0ZmJeSgIPnAVd0uta2t9LfLOlq8P0J/AnLBRAsgPeIC6nu27f5ox+TCpNpxm0Ys
+y975przpB8+AxaSoebhnyTVh7Uh8q3o/6bbvA0NCiqGEZyILcVIEjK5Kki0TiDDWdMGPBIMgqMa
LtdV14FUH5pjs7ysH0c0/KWrcqIsm+z8ujmEKwZ16GySe3BKmSRbqfnohcJhFn0uvI3+jR3a/6wc
h1ikMKoIDVZRuNKTs/gMce2U47Rx9q8Fy3cY9In/GgDvKWUUDF/eL8/DlQrvyCpobAgPyRXmx5qq
/2Il4bFFiSUnvYf74+++bJu4u9uXX0n8OuTpIOii7j2/7KR40LHcXDbETYn7Dfbl88kVesXNaNPI
0AMyFTTrIXoyIWwxfz9BFcgBkkTMNtegcJVsUyyaTbekLIBbv7HgHp/8gvLQeigGEyt6bopT40vy
RByQNHofGetsCOpFKTZ+nzEIcBGyLfk4xlH1p7kSJEQv9HAGCri+ePMf8RNP2Lw5UcuBQfUEpn3W
+nRY+fWJu+is/+tP0fm7BGUv5zlRM8n+JkHyVDOBZfgkIo5BBl6h7fyqaB29tjxDnlDEAKAJzBI7
ZJfm0GskgCQ3h6Ax1fTbhHm8EIqddq4qvDZKDdPXmH2Efth9XjAw3HeLycRXvOGCkerDu0AbBW3A
cvaQQwwGL5bZgSy/MOwIWCmsQfB93clWvr/4JyhrqgEJ5oG2asosDkqyDmW2/h8XAc0Xi9WxVFZN
hapku7uqSy57PjetYqqTXw6UZ/CH8Ve8ldXjiCNsQOlpv7uk7DyKD1ax6SjA/wNekbiuCifT1c/n
B69YP+pah4yHvp+9T9JPaHIE/Y/i/UoKixRaK+zOSqOOd+WE4iJIL9db9ZCmuwC+tzS0Jaqxdsig
L0nkSWCBghe0GL7KH6BMTTTRSGoGsxHszX6FZ2XqT3tlE02a9lQ4rlKp6ciIT9BZYs6U2YF1nvwu
gTq+WVOMmAhVSxopNq4hOhkKAiGNOHQXHTHcassoOhcDQqX2mQ6FKIVK/itSBA6bN+VUYpB6dqfv
rS3KCDPEN0ZR0kjkUGpamTCyf4cpAUkDU3j7vI3E/XLmzSXz3bz5ewG/OitpsBGacHxjoen7cULN
PwBxGki4QPpSTIochoa4harpiJeZzuffrFUlemDsB2SWYJFTJEKq49TqhePJnqT6PLFedB0ENHOX
lbFJa3YFo1XIRjJIrTdk8D33VnSSU3urK2vD8n770+BalGazn6MNW6uyvsJlnOZxXI8JMu9vdwEz
xWIjTDhfRRrXeoqz0/t2NdvgrG4BCLXOYYTw/dn0VTpIdyszZQRFQOg2pb2N8bNYoF1KhJDqhFg+
Vq5sk0ROqkPRMw4B6v8PrX52gRRthoLtnSK9iRvAt04HabD/9iC0GJrMrgSR5Yy6Cqm7RczD8aBW
JAV51LNoByM73KCM5MwhdJFeZJRE0UYz1KUQnr2BPoE5T4gw/NEfPh0vL8Y2fkFj6epSGMC+TP9j
n3F44/mdBJrxRLsYbpYnpUBl2hcrl7P0vL8ym9u22gYazVn9jyMyq2kwiipGhv00G49+/DoAN1aY
DiawaJpxv+uT7KIScXNfJRJGakCFkdxNsBOhTrOn3RzhSFB1bblaMqeXGe0Qa0dAdyfLgzhcszZc
5MXiXhbm/fW9bax1Z6z9O7KP8O2CCss5n85HxiBlk/gBy1KkkrrYX5i9xBuL6dZ9H+jluKe3eDG3
TV5Mx2/IFw77l9YFkUOcChCEJwAKHXNIaP6PmNFsK+T4kjJ+ah+N6yqPNYXccLbAMI7ysXztR5TM
LNyORZ4chcEKn75/QSmDvq9ZV650PRfjPNfnjsBZit5TEUUlImnTalNyqFf3LbdQQT0vyth/H8ue
mpbSgB+DwCwH23ekBWN29HcBpt0e3OQXuz9MLbfjLycELjvEJwwQH93mILsfG6ccqulfFY48w/3t
B1jkK4/iKN4xz2Vf2FkPMdglJbuL5R6QzGeQ8Tqlcny/U/QLzKCQ896WLsAaQxIHGluO2LtSuvF3
oPUbhqZLS1A8NLBZYIWNSgQ0n0/ZA8gglv1m0zvkCFXjRWN/Qa6d+c+oQp0u309rcL+4boTcD82Z
0ZgFgDU68MRMM2un/4987Fvdi3a7ypDo7W6iI8fE9OAfhiHyAjzCqAQKKUQsgaAOmjdf0HpBYthV
rHP6tCdihhMF1GNoZEwFZOlREIt5mPYBQBl/vWWPKWUS3uWpberDg6WbmBj6xNFRp7+Piv0d8XGD
i5BnE5Xkb3cmXXUpPBvYz6oJPE/dtlo9yJkmgtcuDe68yfZ2P5IRNbD8pfF53IBUrCNhIc5hWSHG
cmURPzlDffciqohPAQG/wMetn+RL344wsZsfHka+XjgYCGZtYnnsPnRK2SI5cQWjjUA4lQFWnjBh
5NxXkiTZgP+Jst0S8vphcSkxKHrOWl3rUkzTKpYVdR+3o6Z0tO6ENW/LEi9h4xulsuxOC9x4pAI/
qv7BUPwncMfzYWLpEKyvkEZnzDkkdC6zzAVg8SVGTOqWZOFY8EJnpTHo8URxXE+RbPKoKoRZDo2V
Wvrx8G3DlW+QEMKu7ev1tKQHb3J/S8HDvtcEWBq9Kg/ndxZAIGImbmHLKvXKSDTGWWeO0Ld3VUvE
35QqPALFWF0V10dHCPeGRyPU5khRbMy0vMaQFvNxPTHEeAEiPEQY+QVdhCM6gVIBvWM+sntItoAq
Z8CFLtAhQOV+J/z7Ea7Yr5FVOm64PHDIz8tqtcsY7z7m7kigvBZT9Hqb8b2gTqZ5e/oZde6NSCZC
6b3r/qS6L7TVErCq9PkFhpM90q0+Xv2yCGfvwf0Lz7rhjRrC//se217/KOjmrK0pGc7m9qPYEpvY
X/HAWCfaVWW40P3tOknuIkg1kMYHg1muR+GzrZWTaWMTo7HlsNplsQ/zeqzZeYBmzhtx0AiOVxsX
KBVB3vmDYdVpizCwr9ZjQhWk2+UtIpDHBqi9JVB1U1f2u+pGPOjgcN6nS02SiXVUkjEBbnS1txZY
/kSAHYLEwu6e7HblJkR3WnozX7Ar8RROVwtaO20C9/7vfsb7/58p8OibSzNowlA1CG334e4FRHim
plNGBXtSipfi3Voce9vawp5dX7KupayiSgS7gQapuKRFfbCs9S7qZ5OQ5CUyTtMRmE5fwOq4y0lO
weNn9uKTGkx35YfITs/XPVGiSJmZRk0bZQ3O/YzE5bidSN0DK2QrACefqTNYGg6mE6RIa71MbyKY
aiTF3HlwVwm5uoq+cEHz95y/n5rLjgUWVvdpjJ+27w6+heywrKSYJehwqe0kDT9h+LlSlNhT4yVO
2904GrD7lVAiDb4m61xCcYGZcKxR5ol3dTa+M77RROSTEklQne6zZujc38w+Dcco+HsFDFHz3IRL
rQJ+Q9QHzTTwZ0gaeZdSZjfH6y7IxoA/oWKIZG/OqhMVxZZMYJdZP+q6zA8HvbE0wMg8oDweUiDT
ajwvtVG4jGwM+KKO7yfUb9350uh6sgVLSaB5bnvJPLOdOXXKUlwXFQN5BiN9KQGUfema5SQ7KLy2
z28VPKZf+fJszKsfC44D+7Y+O/vVlCVFMtypPpMoHY7AWF/zT5DhyjHJo2W1V+j835QP848mtCXV
fJaU2GgOpKtYzlwtaGiDMMrafPIRGghfPl4disDOzhlBMIvq5s4vyA0NHeluwWR8L0ao9aGVz497
PS0YvcMiCMgZ0wSMSfFpmfwkJCniK25+aUmTae5UsV3+4BWnzOzYhmLZVYJiTqXNliIuEifyHrqA
g6FeNPWzdHz0p+zYBW990PIhw204ltPCXViBHkS+uk6Uu5ePzVWu1lyBoZCgJUdDJ19lxbCY09EV
nAocmhfEAsVsD+bOY0Qhy8A1hyhbhcyEClgDVZtPZvA8DA29ftSq8llGMBFAhDWoq5HgwxZpSfvm
RKkpcd8GSg/YM64bPO3vUVGQWjtbGmAABKaJ5o42E0fQccSKnMhw7Ceg31ievvcy3QUFWOOx5x3N
55eJ8aAySm0Q2rWNTxqJXBRB4Ql4KJAogx3T/UVTXCsm5QL83uU1PqNVmnpEdYZHRHOAX9h/XZTk
X8q/f1S8O0hqnAZl8PuFtSVaOMAs4Y+dwYjuYgmw7L85yxlD4STyXqtoKcmioc41I4p98ZHJUXcZ
k0seoEkUvi+tZrnSb1Pr0K1f0hdmVpPxMxH9z8dn3hz1pA2SdjgpODIN0lhj24wFKc/yBy2nMq+S
DCYLNL9JcEbKo6fOFWm8T4pZ/my+g3hihf2oUzS8CFe6IACA6O4WXoHV0lZ1LGbwIWuW1ol0Dc2U
AhpKBwAWYJUJQxt8bBThMcrRlEmP4+YxcCquKRN5hA+E7P1ShmDH5QKSzwIMTG6eH9Qzs/zG6lkO
/LK3houJi5T4app/OOe2rDJb1DlkDFdOO3ah/2XFuragBU1o/de8dxrVivUV0t/le3mCUo7fH/9y
pqjzO7hNF/af3LwRshKc/Z5dlL8O0b+3k14ZugIp6AWlv8sp2CxcfdvU/jP/TruR0A55uH4PYc3F
NRWhMRd5V5eF6+MzxVsWFRk9BHtgchXinwqxPw/Y2wpcjTNxCt35j36WWrwKcJ9NwVle6qzUli/9
uM0uQIcV2Y8NoNIbmfq1+D4QCQc6pcXy3mizNnARN3WEm8rMVKk0LlYZkEWfWt/ALwp8xPcB34eb
dZfbL+FcpuiVEdOsFWHjmkd8OgInk0tMF6XUXvqzLq6dPfpH+WcwqjDxBr+sad+1NiAd9OCcPh8Y
JMLPYH0rhXNyAbuwo0AeIt/lUr7/mZq8qx8go6Pd1FxdviJQ5/s1SMZB6BdU/KJsPA1F1e5AWzGO
7mKV7p3UNTzGazznsXsdSl0zVmS2Mr5u8ZTGQqPcGxhksdLWe8W0eJnNGf8CPbm8OWeBjbY6mhKv
3UMSznwH2XUsCcjyb5PAe1Tc2TMAKYKpxtbbSfs3cUhYnVUG5Rc5nNgr+BzYi2kdjYyEflAet6Bk
Zx84s7tSDMmnWlDIp2qVUfZl/bHLK3s4ftMRMHwfvEOYdUJvbhNaleyLt/iGAYDNh5NGVXLkfc/y
g6ad2JwGvjjaJ6Rt8mJm9UEDRuz0Fl6AXIp3Z8XNnNCj8DuAJM22dohy4HE72K+3iQDW5BGSOJLd
m1g+5tZ51J0aG945uQk3gaLbpqR594Vih6k9GOWoXl7TAjimhvQBYpV/203DLSq4YehcfteeYQkR
m3DKpXx3iv8mvUX04vIsDlnMY/RbAPg3+KH7sCmkfo8NzSKcbQxqFFLfZRUY+VPEvIwjtxiJXvEt
/Y0o/doQ8NguLT4dNlGkM91uV7sBxVsu2hOGmwNRucpNGePGpsLD+tILc+tlnpYnBAak1nnfzHZY
KDYT149p77Qp8OO7Gc6m53PQzX5CIi4zdfj+eh7oF21iAkWek5sZIdbwjvPPJJ6jaGX5HXWQlpbz
kC1dmIQwwyR5z15Ypn5F1KH2kIwxZvlhSgCkiHzu1Zhst6CTKKFwxwi4d/crnHHoNIvi+EUqO52Z
KyimQrvptNjVgu/kaUz35odUyLn7WLYWMcPz+KsmKJPYiMrwKqTHPI6MH1nQGPCF55chKs2tJQ4i
SSuHevMHlphSHWQBbYBFreIsFjqAvXu8BU90qOvCyzFeQWnMeu3NtJxIUJLi9cHIaAs5M7wXwumY
wXCSz0nF9iOQjVyYTdxZXgCmSxckCcTJNjdJtebZ7ih9sLfU4VPEYA8GixFvSfwX7OqFpqQvqByo
jjH+bay57brgNDZ6rTSUzHhpXg+EYTQCN1oU623KeT5R49W4pLXsJT/6Fve+rRHTAvw8Mp/eTAD6
DzFMKkIVIihH+wGxTXUYGxpQ03W5KrNTVxqYOchN8meB9+9lMCqHsIvy1hvZketowNv+z5W19p2/
uKvDyK/3YNlMM0FGywDuK8MBAQqlAI4sEZnsyjz9Y7i26pza9wwEpWgmKOQ/g/wUqM/R49bPHBwn
XobpUwyMeOxCrKpyvNiOXQd/bF/Hf+TlUIl04cmARLysPv4g1ytmTSudEMX+8HW2uoKwNSGdv2Ym
4wCxlP7D4j+6kKItlNpUdBHMNhzKvwiMk+g2XZttDuOGyiakt4c/MSHQZ4yhfZbwPz5OZLj6y7T/
4O8yfvAiMLLPRsALe1ALxKa+lYb5YCsYck6RJohD7bVnt77dwtdUO2fTn47LHOLcbQszqK92Edwt
6iK3M3XIQkJsr1JpHJAVI2by4LwSDgbc/zZGR8RX6TFgcNqr/DXqUsgfTu/IsMDA5zLYsUdsxTB/
JGZ2QKRabk1vBTZfvGI4Kk96e6vpUd24SPO3SnR5Wmjy5G2c0Rw6Y2+Xfz+MNZjDnhM6M1MaGYZ2
KF5fZi/12VCXt9tXZZuiYZ3Ik88kYwLEU3f6HNtE3Qkg8NnC0B4sHnkX2kuujuRBb4RjjVz/2mQI
ItfI3HUY2PoMTqWC+XQxyr2A6tRbGN/Ja+45j/tl9QiJBPs66+d7DUV/u+ZV3z/JtKS2WecxqMcs
dBvrxs4sEv+QomJ2OVgr11vSSWeKY+1E5RGgPpXpX43vWl61EHgMtb7wKijNO4uk1E7/Z2QKb/UP
42kcP9NCd8QiX3m1x4FRpXxyh4c5r48k1z291arl9AkTH2G4vmBn2ztONmMWknOUpfifxwsXMdeM
qrPKRHJ/SchKTycKOs1eRyRbPpkYSQViiBkiU7Zuy8QeZTwzMouC5t9LZImJyMuwk27VCsv48btI
af95WV5NRHiLnK0GXFXxbQpbohszswiPCwNoqB5H+pBGS2QFaOLBnJZVa5mxXk7okBQZaMWjcrjl
/YBciqUGTPdTRhsC8LsgeuORxX6cLHgBaUqf0UyLs2pPywx5cUQH0CBouMqaE0nugitVVcLyakf3
hyLtQZvg98LTuXWDPQrH3bN3CXVoAmsThOH4RBc8qQatvReVBlYvNO1IWPh4lKa+9l8UM+BScCtr
s6Mzj3RLjjGk7kti61t00+B3kSHFPUzYyEL8WOLuMSoANKr6uZaKbY54kWjge25nUqsqo4POT+oK
jZ1m7FL7scpMd0Rnlby97oNNUQQ5iLx/n4VKBPiH4FOgrKelWKmcdtZG0nbRqwW2tJN5iSJ6aaUl
i0mEJzu7OhFZd+yxcjXYJmLhJFAnQED7cVv0mylAMbU5Ev6evw/vgTMWzV33AyFuOur6wgAdbPZ7
rMBfQVkMwu3YQzMfXq3JjFE7vLRl4sfbLhNuyAM4T25KiNE4EKwnY1zM+EQf6Woy5aMPqOcPk1bu
ag60kkmEetwHKv1VyvkT9KgvMUY/aTratzTSulOPyZpQ9VWGuOBDug2BP5JRCqurC97PKCj0O+TQ
Moy3gbR1hqTnxbzU6zm90Ase58JdRU7pTpBgTTW/ibpwu97pvXJVvUrleqtdLXszu+iAweqHkg7o
MVRsdCVjVywRSfJgPhNwq6XFDnWnbPrcfU6abXN710Kn7eaD6w0kf+fiE0x83hzLX/vrrbJBqShX
BtBt5LH/f5Po+Y3OuL6R3C9EB42TduH2o+t835s2sZOdAp7f3nOY9YL+EkroiaXR0DrdFw0Uv1ci
NZP2qbIgKZeeHbZXPj2vYwr90+yitnsllObfQGuI4RFCPxG991NqHu5QiQGnQ+7np7M+yLNqv7ZX
uiPNwEkmVFkSJqkjhBDpX+2K4FRE8h7mpGloYs3XyKDlJoEx1pNR40s9vvhM8quUg+tI2bh8c+OT
Qr9gus2E76CBIYehYJ74p2jY9FawbYjWxEx1j8u+7Hyf0f95Hf+CWeqfGNBchwoXkJFQkSXKC8D5
2/HEFoVvVYe0jsTVlDpNc68/iVzDqw4RpjgYGTgu965ampEjeGP/+9gJYa3RYUSuL+Xl1FX7EDw3
jVWGdgHaCJKu6p0BqgXElRZbeHDA5gOuaqYwP3hegKS8c0U28l5EfkC5R4EvfoLDIA7BC6JJU7Bp
AlgTTx7fWFiscivLUTqoC1YkNXEUXbrbrXwWcKY0ne+8ouKuXtnhidq5CuiU3UwbdAIzPhRCwi+v
WUwvARtRCT+CbFyA7m9/1sLnYlT9SJhRlA+jTpoViwFLwDQzEwGckIehKuBn9T+Wu4CWSZ1PBMXe
RWZcq6iaxFFc+rNYE5MCo+tBMW7qVxN7wxO/MZ3ia9OvZZg7fjUWfiveYhuGGoYKWTbS7SEerkRc
Itz/CSfXJeRtz+5k5JDKpw8EJSkmSNWwMOmUnmlQPYriWGPRi2VjUBN/il2Ng7+06My7y0EMaY8n
OliYZ9VW6mxT7hm1yyhINXlQdZ3l7ZNK7bxuH9REDKMaYQrDIPNjLxe763CDbY7n2+/j8CZ7yNIh
Jh1nPjp0ZIoPJcqOcvYKOfcvP4Of0oPt0cm0+OEBIDLapenZogE3ekLUyZJ9f/a9MiFCuNWVFsUf
rFeaBvozfAbmoqjmh9hLjzZNSxlWBXntMIDzwV0j+UMxU+HfTSE24ig8SGqvT3+8DtZcByGCLprs
T8nLzZTS5fnMux6V+FZHAXb48yLhqeYpZXfm6zO63pM5/SYWOgM8kNKWx2MElnhx/Aa5JGZx/FY8
qVxHlGddNx3OIyYwQKfcXfr7B3Bd7AOAdBk+zJtCRJvvoOA/oMPTVtHseyMIPD98cGN+43MWSkHw
W/w9hLoy9A64motBjeZ+3OGXltAUsDmNwiNQJ0Bc5+2+beEJKfT2GLD3ETVT++Z3DvNaSWW281vl
uh3vgljvfJIEfAsroQTdPqtr7xRw2CUx71OI2fR5EcZWh0N3YR4xdUbF9DxoX0YWzGvFnMfyr/VU
PlbX8bxe2Mn//4ZuIGvhKwSN0tgBdt385hyRONpNML616yn29waG57FTLqmCG+5NN72GTquhWY3u
1ftZSjz8tti3TL4XwkZDqhy2xh8RpcxJRr+0UwphAyolXnRIeq5+mWa7Mpx0mFIAzxuNEuo6Drne
CBMPTedzrINU2LvjtDl4rvJDUXAI4gCTbyC0+m+ZK1UQLvWCWDhYmd5CWWL64442cVrslQP6LNSS
d02qz+sAcJW7jKW4+mlO3yP/ph7HlesV6O3ISwbCliaYEoOjqJvUljsRp3k/wJmAAp9IkzgF0cD8
HToErgvCWzLeXpoTJ0uMFgc1XoCe2hNrIYfYZtLOE/WIYcari+yNgrm55LeuP5aVvbT7JzeSWVrk
fOX1e/Yu0cZ+R+uZkYKkM0bkTiHuVZOWSqTK52fy576Hy8LzJ3nqVxxo6Bu+RuJnlgv5iuKWwjpy
uvw4+km4nf/tB8ydlOCXV6Cjp+Dw7Y+TM3Ib9czF9g5Q2VJhXVxz15VJlaIxEBeaw0CsM5W3mDMI
W6ACbu93VFV53Fpf/BxDTPLQ4Oe566gHWGJjUZ+2vrdrE5XEYpew3Xc1Ay+AmIRaoK2PtdXLVV7M
OywO5zb2rczpBdJtB+RZsHJ2DyfZ9cT/FMqJbtnFz2FKQKhDq2+Bm5UWJNm+TcPnNZBiXf57EAdF
IKlQqnTF5JDFr7hpIOs+S3tYUZW0mS7lpK0cjxycSTnDT/C6Ec91LDxvWRTpwr+Ng6dThM38sYDA
wD9tYz0bPufbM214iD85cb4idf3eZSOnBuhQlXbt/92ufWQLzd0/wY0jSdV1YVovxXJdGhLtMC3v
leGH3Shu3jwyrImXgjJWXh6ozMcSYCEznzPe/syVw9yokFdZo4t0KU6iXmNFxo3TeUXbnswlfpek
hU62Ug3MM+cTpAQARj8Xzw2ZMztAj1tEMwa+JoVN5H+l6TsbLJXT1hUmt9hnXFvxNCKhgmjH4/KQ
eAUxCLF1OAHBOm5Uqjcy9l5BBUU0d8jwt3lUJZpoaDaWIZYZAtJZwXxIXVMV3eAcyjdBlX3vDYzc
wRuEtNJjpnCDBH5mto1BCT/FTlqtpf2cJRWQi4yjJ7O+c4SeMgq0j8khYhfU3DmmRuKSPzXSmWCX
avRfAt/J5g5jB95MHCpQgaLvdAsKpyV6jcV55jhNzZVW+ZZtrknJCgulcAFMtoGyitNis8XDFvMY
WkN4WKg+ePNsNM3JaJLSeJr4iqJhrpJQXxrABEiqVyUG7xb6O+at9I7Ne1FZcqKUHpRZmpcgVMCK
tPAUxOteOLtQLQcY9YzWZxsp2bxw/UShrLeEV4y7MQ7ydkiij1erdkiPKke9iQNZW3QDPFT19yCH
cnP/bNkGqQJZFkwnH3UKH2KueOAbOG3v210WlLl5pN95hVi0sxX4PRgSYqnH6pW34fplTGP4uYKE
EX+mS1wYdWAYRqx/Cq7yIAlPsmz7EetTByDwLywxyX40wiCrZa+x+6Ltn0PF8ElHkIjhTD+llYCE
VmEqVixNIPyYCf1lQ6yhlWOIakF7frPYIJcFn4RLXjnOBwe1RJX6Ytti6qrF7OF28m6jaQCVutGc
WdSp7mCyGbsq5XFGYBFD5y82BfDwR3QgxW0Gdd3yiW2jce6kn5mm+qavZNf3WSuaoy6vRvliGm/i
1Zzc3DjHdl5Vcf0ouvApdNlBepwFC4eUmNulPafqV+y3K/uDuiyB4TwT0P6lE22RSw/kC1ozb37V
aiKF/Vj6C05XHK5+7XcvhSi9OoU0f3MTgHDDu1hl2APzgvYc72bEMjaK/HTwv6rkPS5ZbNmNxy1r
hkK2n4mlmiU6msCWsBnml83yE7La3S8Ny15ZCpcGFvKj7yulGDIph7DkEpY+WlPrIC2JHrLNUZbt
s/s4nB490WplJb/VfhBrTJFQWZmyYaxver+TPA2Zf6kkShqnsiY78TlVttyBqjoCjkmSSZkmU0a1
Rgt8+k1Uu9iw8Wult7iFrnVp35HGBCLBTpyfwQN7sTqIJNavnyxXXI08UxFm8vLgvXnBxBstk1H3
znpldDEG9JxRTsQYd6tg4ZZN/2ky1sBb/H19y/+3JR5oFbT8awTVaEjfLRxyxDVnOz3AT2HYmKl/
qYmsSuYVXVESdbWWP9YlwMkpOYvlWzOkyk+lVR7FHQHHG1z+8FmT+HKdVjPOVMh19o6uu3B35UIg
U0Uc0SmCiQMAvO/7DA5xoK+SjUkx6FpCB7xEHtwsDL8SCvqSq58hqJMPYs56ZkyTfbjM8SVMKVBI
j+pfjUjB0ATBl0MvDJSdspCd4rN/+4ss0oM66IlXw0u0118+CVdFLefeU3LwXGPzSVmHKqsI8Hh/
qj5ZVywZlryb243vs5aLmA9YYdaCmGoxnm5Raz+WpFaMrtz4fmLHLS7ZhLWd+2+Vk5BjJeznSUXv
vL/2Hn6yGmcQ0GVKtzyVvRU63kPoXct5cua5oGHDb+YVld4Cfsiq7kUsng9yVNQgs7ILtbVZie9/
TQPWyTLOR2qQcUthkni4sYNs3G+ZR/VutfPUc9Nw1whjcdUhY4tlQVHIcree+a3xGNNrY1Gcpf7c
KaJrldS8zEFq/ULOagel91mjNCGANvKqYD/eGu8B7cJIK0zgOzoJJ6ma98Z98d+wE6Vk77AvcDXm
fN00oJvN8bkDDbA3HQXwq1QWLvuiiyk5n1/kRWQpxEpKO5gckYl9T7cZJBQWEFbKnAgHu3LHJLmy
8hTTRsrN0HNYvsGK/ZZv8K0A0vGTwKB+YPUIhxJhG8OkKwnUXdBTjEXtmkvFeb4y1akT1KjLg1U7
fVO7XaqB8NY82SYB2JNR/lThplt2W3CgapnKg8n2PhQfJSR4NZUi6kyYdfAIxr1i2d4QZUcdEQFC
bmtC7Ul1xJj41BCxPXyV9kmb3/estJxdYkAOQyHEz7FzrBOF8ROY1WQjJufT80a65+QnFTD3Ks05
diA/kaun0ByYLwAaLauFL/Ex12QRaEemqo/V2DQSLGhoOTea13q8zkDQciFlB0NHVFKWgD4Nek/F
45Vd4myqcbZ9DSGaIqcWbt50fLv+Xeqk1cBtANmOaFcTnTzVbg+SUYibuX65qJ8tH2FjD5BDlNNA
YmhFtajWnJOK7z0mc4FeLCPN7Q6cZ+lOumFaOrtqgzLB6S/bDlcbd88SGRdMA/AHR/bwUnIWtwWm
zq825EYjfIEmQVa5A34ArIbKVo0Ox0i58oWhdyAjCOF/BNJzCb4Fol3b9V/+fs5cCBsXTKfq2TTU
o6ZforFlm2MfqeMYiL9oif4zvzmKx90caKEnKadOsO7esi/wttKpes9DxXAUvbPKl+yUUxm5nfO6
j2ojyEnHBXPaDRV2KoXQGp31506TB9QhbLTa6gPLmteqDOXNe4uuHzzS+y2k/AQgbq/ALRkZCifE
oWUSAjnzBoqeWSLAF5WTcKUS8c/W23ydJgw2wGIlnivehaQSKyM4+d4S6dEHSSTLmfw2HODuX5aI
aubBb8BsyJJz/oJj4R2i4lbNweIhCvP7cPP+dqCVU1oC9NsyJN6ohTYCnnQV1eTJlJDA2OXrmC8m
HBm4vdYgVnf5ZD6QoX53xJpR13nhuldqsV9HyV+mu0rlwtXeFo715pnQrujNppiPYTDQSQWex/NK
DQyXcauZ4uJHTzvuPuGeqQpThB0vLB1X+/O41Kf7nA6pJaKuxoYpzPd82IxaVcfiEeO5bDoYGtkt
jXDi9+qKnD9n7HO+BMvjNlxMWI8Twn3KuCXwgFjxMMnidHMRad+oqzmxlISmOFIh8BOdDM/327+J
omREhJ8DTOibEG5P5bDooP8f8HdnBu2Wy+JX88tXhmqGFM6KVT+7tGZDsf9OKIBvLZL0z4b27jp+
oCQj6KWPs9iO6qm2Z0tdS/bELhHkFMEHopTBsjy19jBlIzdvTImSQAkeUDbMH42h8Vj172I5OVVe
XEIGZ7qqdoPzINGlv0rzY3SVXRTQxUeYZUlC4EtIhpNTZzDh3wMDFnN9tCc1HsCSaqA6j8k8DE9S
dlshLsFz6cabL/RVmPIE5SCnw8cdjN++sfh9IZPNHQt9u/g3v/8CHuZfJXU0LHqJCN1VDH3IPZy7
5nSzUvPV6TZvbmmG3jkV5pqE5n54LJdEQpgqnuLEN4ELjEj84calGA8qDxeOLXBT3b7cgg398YEF
yTgwrKr6aZf6MjOQBMuBq3KTk7pOSYpnavvbCj0B0g1iB1sOwMGmZyl8W+Ws3fIuVTdyEgHJBsB2
iqTi16Ng7nOlVRQzRLqHShGLBY5mUjGbocNCLTkN+KbvzQSGoq73NrOADaHEx4NKJOqVlUu3TlP3
hBQOqs3FlWDww3ItUbOxv0pZgaDbpeLuqxDP5Ito1vXGnJHYgwochSdZPVl8PuSpvivmKHOu1F7o
w2CeKT39L7flj9BgfJM5+lIJUKMIdsaVR2Sic8NwTS1rvpBZ3ARvmtQnZulBaXkVc0VkweHlIBKq
pdpq3o72EgIv3jKphf4v2nInxIc7E6ae2AkiUOy1Fnn5EdlhF0gRFJL9FEQM0aRYNdMvtx0LwtyR
KO0oVUOu5qTWz/0AHNUhVo92USN9QLveyU2poyzpylOe/BZSg/C0kXB/WGUQ9a6iXBWrGlP+Hr0F
QtomDGwMS3tz75btgXEMQDxYTAm4QNoEZ1muAAlTaci6/+CQ+64RNzBpvRm34eJaWg6AnUXy/bFC
K+90i2EflXkIsP5blYifacsA3IXPev8JSYUSv9xeSbuhymVSa3oWXGhQ9LfuGz3fFSoDnHf7qTiu
jePTVyYJ0dm/pI5XcZsa41tIKx3XhIQvfMN1tICQQstPLH/bJMZ2G8aV2I2CUs+P5bBtr1TkCb5I
FPl06DUTPZSTZGSfjonapMvYeeA/TF0WVCbENc5G5yH7u7lF8WyZr11AMUtLq2acL4/2C/jPuNtk
dj6fL+iU2OyK8xW5h3tvYXKuQo7ZHfq6WUMt7e5KWp3g/Yp6lYq37yhYZtg64aGaiZgCB2o+deb+
NMFbK109mAsrtNPZ6/JKC0BsQWOAFPstC3dQguCnfAVUvcbU5Vx7o8+04KjfG3r/ib37VplGS+nQ
OkPVCCfozJT0HgAP+gTilSBz/5xIKySkSvmhLZ9s5BqGvgeCrqYStzzBk4mPLsRDdd/HVZJj9Q9X
Qh91IXEAsL3Rk1IpqjIy8h7Zu5XKRfQGenuFFbHJ1K/Za8TWw41IJaD8xDaXAr8gxDXBSQjSZ+0K
KqmEtVhx19YUvpc8kntaVT28k8DACR+FFAQqwAm943FcEY9kGqMt86awAV8diwIsWIzSjqeDqWnH
piq0JVBmfBkr+pEjHZ90WCGGds/vy1HhOpPL6sieODUkQj7fTa+WK7mFZ6ZR6W8JMoLFyFl4u7Ss
WLdO0LLdQVGYGhJPv91SejIXrgg/keFXIvcgIwMIswU7ivBj4yGgHOE8J6uZUv/rHyl8aeXA6tvp
IZao2ZEPdGgthrd2p0OOxulpFrCPT+pgi+zkRnhYfDA71zwmyGWJK6t5kY50pGZWkb7Q3M6Eh4a5
6FU5hictSpEj+i3shnoqp5jTQx/NjX0buecquOpWvoQAPZ/wcXg1v3Rc7x5RY1kU/AMVk9DuONYu
tylBk1ruzL9GuZWmsKBPOaiO4ca5iJhGWbMh69mffdUKscFI1PlCpHGXuDzGf3EYLqr18LU3igAY
BEgnK+lrOp0hafbd3ihjObWsAHRTBuKfJDyF83pPu6DFrXix8G+CPLqiaRUoWxTHJxu//9MClIju
f4Ruc9dmfVAVEsvOo9GJaMuDP5jaJMZqSAMJk7TdTPRwO5q7mTOIX37UyJrJM1lXSGEGP+5/Pgu8
6OK4iTRpKy/Xu0tEUdJimev1XhuVCCTXIFIPcrOH5iRj9Dnwn3i2z+IWRT18w9XdMiaDwR9stdfs
L2IS4VuPD28jeZbVFHuz/u+fChLBKAnYRWAYpDN1q/pq8PWUr1peE22K9Bt6I2iuTxhNFVmGZ0Ed
bkPw2PJ+HNp3WE5R9ZYB9nBWcKTZ306IAXFnfWyH5BkoU/0dwvQx+I2ekuQFqbtHy+figsRAZnR+
YVUnL2wBL0EPzMYBYtp2O6Na/8jT0jH/8auNCEK1xS7w64R+fP6GVcW3lnVU34ANrG5YJn54wLQV
H+5FeB+wn/I9wfpU6PWtULvnMMSZSKXEqpQVuQwH+VfFQcsofCTGIcdi+N3DcZHl3JGhmN9NU0uy
xzAyuVWMCRI+t2alPopfFV7MV1G9JQIamdbXTBgVd0Ysz66D4ApsDjwDrdQ1V4GG50lcRr1VgECz
u4kKv15KL7UHWoOIZmHImd2jTxj6XDPpw3/buLoao/fo1fs078lkXaAlDjbJl3rmImmeuu1pBOfl
clJLQvLluTgtuM/0qUIgKCcfysJowwrhLI3SZ0AuQY+rrlIVgc9LIPK2A0uBrZxW1CwxDdReUSyA
zxdtWhgEhFZN40iuWR3T6JN0fZ65HR9HziB/nVXtnqD/pn/NvYax4YKjmEpM0SUAGvj7XkMd3Mdb
N4FVmyXw2OZju/zwRe3fIc4kgcIm7IPiy+/PNG54nXjIv3DdG/a6kgVoUNvF/D4fr82dNyasAHN4
VQqmIethKi17VW5u+aFU2xNaD84IpPJflC3j7dbqFx89HOOnbpBfe8lI//F9Kr0lpfvgegawQ7Ud
e4rXgSsTlWe/+PSlI9nyjLM2jfxGYfK6eClWPafJBzJuyewu8yn/Mr68CCHgO4IECZiwzIzTrqah
9zcTorHADJBvuA65liE+1ciiCceJUT3Bm1CFILbJdS2nq4Al1CO7oxyJUEOvNIb8lY8oTEIQY0n4
ptX/spZJTKez7aZN7CypM++RY4qicWZzYK6MvxpQxrLTQ7UTbA0HgXMVFK3fAF1BFXQIXgsckTgf
QFkEcB4O1hRBw7u1yu/eMFAGeS8sWk4oZiCf370Yz90+CmKxz9jra1kLGjaMTbUzF+kna8wD2l07
5dJ9VAemeGDU/bPZWvkDRz9QPgkZuScY83KWA/YgFthPV9/6OmVeWsLNbWqQ/P9c2vKxQzcZ7mum
bYlPpTTSM07Dz0NPXkzY+QGDNkpdtVjwJRGI+CKtvFLZCprn65ifPCG2PSZ6/aSSZC7F8nyt4P6O
VVfQgjKaF3U2MENvXb28/6JV70yIkExWn5efVWNngqSyPIsBcbo2E8UZJsno+upDr/IAAfoKkru1
BYX46RV6XZ32O64ytdVWwnkJ2alpFgNKCup7VhXP0+SWRFfmEY13RNI6gDPSG3M1s1QHdNKJhOvb
gEqD0yLv5oxWZ5+LRYDp9jrkyVTMjcydnlLYV0XO54CuIMpZ4zHwUQdpa9gbMMsRZJE2RZt3sgDR
/xcs5VLWxw2JeiRJVxkhVjI5uzwApy/wXdzg2Rk8QqvMqxJQlaz1u71lZeZlZk2t6Xdn4b/bbTEZ
iymFG/PuyopIJ8doKRwXKAo6uJZw14dpAwAN87GNEKBM7fQb2kPTu0Pkpo8bkpQybMHPVw/iXPiA
nBSRHS8ZJ9JIbPFC2NkyKFNjnwAmT2whKupF5Cf/q6zZQzGV9bdP92Ugz/T8jPkHRNuxuvzhHgAx
oGWoegOCPOYBVCB+6+NTyX02b7rQLpgMxzYzz6+f8Lo4ygY9R28+k9eCKUvLKdAkm5JVAzw0KRvr
tsMj8p3Re0/AVU03/CopVdCnjxXny9ifdAYsVF8DNf8baFFXp8OfJOdQKaRwZ3Ymk2aY/17Uwauc
S/6zC9+w/heZJdLfdWmPke/Zjo/Mf19sVswZWrtp5CVlc1s4CDU7NVlgymeA3gv3WoYDvli5eZkP
wmh2CLA8e+VkI36LZF1BM/DOkH5BdFY5/MbNSLAmudxwZxE/CRKnaX15c/KgSuEne/kp/AafglA6
9YH+OCEfZiXyR/sIJkIhgQ4Y704IPNtcwY4cOnwNVhyYAEaHZ69KKTi0N2Mz6zbWw0/K6TLv0tCp
2+mH1L08RuBRRxqLIWgYo2ncSEFbgwDLAhkuU3ux+Y4cEIf5qWWPaFN6ihM0ey8DAsVzVlUul0N+
TBQE+6KOQWY7dxUjKdvL3EVByavEmsN6pnPi+aFM8MUhqyysNcgntY3TAkTiCnnL9XmVdLCdzDgb
XcajXmBCTJcdoc5pzvV9oHoi7kmXeBkV2w4/vcNveWaGU5Kk+GvlhspGmMTUbbu5fhEUQrbJEXtn
E5am8JKIxSEqsQH3G7neqive/kOdHpAj6mKbcVobD0U7+1zpDbwYYZp6vyL+MP27AAKzZwrJy2AZ
JpmAEIyyPgEGqLlnOJeAFuksz/YV1BkIwKxZkt2/yu9tvA16aUr4xA2JW62vssCP2hjXvPpan0Gq
3wu2XDAensoUdZxYOF5HSQOlh2k8iRtuEXRDlNRhGtIXs3i2PTqUqfyFOhW+yrHn7JAqWVPOW8UM
PDGbghRt7VhuVDdzpzc0ZFZlD40yh19wgUUF6dy93+xSYsp/4b8T6pUiAsMiXLRzu4/OhPhMTCBN
AjHvPheoKPopU8psLo3R95RicgtepUM9foDOBwmx6m04YVizCIZji4keqZ6yzN93Z1FN77TBH/1g
FJYUR03cGfylKqLncGx/N8DhYTbDNUBMWmZAXyb+c2+NeVhg3c3CCgVKy+KW1jp+BuqPptQHE3YH
McQlvLbkWI1B8Cu9UlNbG3pWlCwNWSkLbuIz/QHmHLCNR36DHw2BdI/tW9J4NqrNyDDee8m6lMFk
mzbxft9rn6RmTfNpAgrVcxAQ97YJSnBTn+dTnx/XzhpRsfUKczqwUCJdj3Yf0nKXyyHRbfxOr4yc
z8KOG1uzoJl2hKUFhyfNrQZQ0rK55yQsL90N6LO55g+s+cGAdYhY/3HmLhZyW9UGK9JBIm508Frs
WtsA6mTL/W/+sD4KTNsQLpZzyoLaPeYhd/VoKVw7eOwVvzOZIzsQJ+46CGEITPUw9c5d3SUwGaAN
1d5l16DCa2aLR2oFtI/crHxZhuuLnyE+XAIBiA3OSGU54qkh8WHAATlt4r3JQ2RxEh/QFf4T7066
XSfYKLDx8LAWaUZurarEdKKcuTbDxtuN11+fF3LRDmoSTpuERqyy5xrwFMGgrz5spNlpMA9boEnW
w6aQPk5c+NocnczTFwF/jS9Yz1tQnTZzLYyLnUxVAs2RNvMQlatbbMAKpR2++nRrV5jjliNiaWJl
gPsvOtAgUgzDLKNh74423UOLNjKQHRqZnBHOfyxEj0nje9S8EpPheWIoCaa4pp7CuCIJyt1fv6Rp
6juXAWQcGNmYG90fGNewurgjYpmcltIkm4Le89pnda48CBPvt+EEXfNd/QIvPTIRB+ejP0eZSemH
S9pi5lwMxLHnCqLZOL3n2CsYvs/KJWh0h0agqqvnUNozGhMTx/d77hm5vNW9tMyU4uNGCk5m6B15
QvKKIz35cAjgMeQrjUaF0VBQpsGqW6A5f33elKbFIgPQe3krqNOY6KdL+iN/GvO0PO9GedMtK3bY
I4YUFrATxBumqxjlL+DiP/j78OCp2qXoDnZ9Ruy260dLp9abv08PjkijHXRHNvPizg1fajaFze+1
OYqdIDfUxAK03KQUNk2wyLnB7+iUbwyxD7zr1l6q8X20ToL05bJIRxTL/jfuyrlwuS6+A/+SNJU+
G0Z/l5kKyYTbmCnRgo0GkaJvhKgHjX+cvbIYn0cUzKw8DDv/i0ntjmo2wfPXAMiALRhMmzhkTxhG
ti+T0l1l9AL9HWkdOnvuIBSRma1C4t/h+3pq64rmoRFFU2DSfZFSzPR3Qdd2m2XjmY/7W5Wg4rf5
zYn+3i9PmSumnmxofiY/gPtqGhB/9wwpkTdUZP/44GebxsI/eR8bjFl0KspUjK60d45R4YwdnOSf
GxmG/a+keg004xxGfpm16SEzqRS1Z9ZIJyRiMNmWiD6f/972HkqoUZRQIOewncIG2zE27nZEKFRJ
R8NYRm3KfUJaW7evOBA5pnLjhHhduFRtWsw44rDiSYUB0eIx+0oZILYtRoUvOpIx9Bc+VQdhytV4
h8TqBuwuC8HZw868FB1n4D1N6dlSCmDSzq9+vU5haCvovh/yfDS6e5n9KcUreRyZ10Gr9m2o+Huc
jHeiZJkbJ+X8eOFjOkQ2cncCmOIxH0JCG2Hjaczjrxtq70ZjHQSi9dyVYOCDg9u/Je5oLkEa1+DN
HEd79DdJnoJsxDyH8agOhGmDD+dBppasvGsFMQSwcX8WqOlMlGjgPd+7eroWGl2pvfYnNEkZAB+v
PVM0WURNUZmlIV15MMov/rzQf7KIWlEzf+J82/CJZe9YDQr5DBnuFawRlqh7YURVCScyaLfKfqmE
Ke3+TZFJPFIG4BpU9k+xyUmTGeQT81nrguzrIdiyjw+knpWQyiNCGVQjLCSBeOmT23FDnXDzp622
KUJWO5zgptycYwNCDTPlOkS2ReaHOgbPY6OI/jur0lFa5k+uBMKyEV8SDA6oMHzRn+cWA9BiE6Hx
IkRXXSVgnu3KMQ2SHimooryWOSIRBSA2UIg3evwFqG3F/3742RRy9Pr7QdyBfp7YKbnU8RdIkwcM
IhWIhrg3Hfl9dksnX5flTyewY61eHVfBC7+Ue1DmN3NyzxMB1C0+4XEZSEjUgGRvtySyrhAdG7FU
AJhk2D+RMh8bzinvLiQq5r9fzeZ/OlnRaQHfhgfVevE7hXxHAPF4CG3Fu34bcgAgHvWu/FZNuxBq
+Wml/F4DXwXRHSeh7bhlVaowv6b/vTncCSiOu1HuAXCy3prKbYkdDmOFJ24Syw4vOn3p6vgnFc7C
1iZs9A5lQTLDrg4nm5lp8n/DZEonriJjS+vFEVANc8HRT8ed3grOVhKBOXaaqZNwMT35sG1dIIxH
WHXk+tVJwmFLqEXQkqKsxh9rOMP5tOY3L7PzmzMj4WNM1GjqvbMJPOh0fxsAw4ZmP5yZYVA8rYc7
O5UC6MODn7XUM1RyucHCeuY5cj0vNLia3ZXWY/KlLYDv19w4MlDJqdDdY7JHSmeWCL/TKCv+vaMq
eL9+57Bl+eZkPdbiyUuCNe2m9g4Q4DsyP4lJcSGRBUT4BMGnlV8pMWfEd6TNs1x9RXsRhzcxvXLY
gg7SCy3lBZmmR704Gtjod8+x7zcl9qKkog/6u58T2NwD2Td6mySOQTuFXxQP69lL78XToQQetn87
uxB3BFFVVNfF95G9Yy+2RCTgqE4X3Lkx1naUj+9GnkzhhWF3xfc+MmN0IKtFCb52Dzn0Xmj9OAry
ysHAmv3+1sQ1pBCPmYyuEnFAeMNwUD/D45jZQbsE0ikedeEzj68h7+R2LZwYeJEwrB7SEy17yDnU
KRyjjJRxUuz0E5OX/eJW9H310tQrrIchLHd2C1Z2EhzUCGHTAkZ6qy3UphFFDDzm3eA/VDw82c0Y
czgEwNxZZx55hSfjeBimkcAChnaC42x+8wQ6cJolmat1wzxyGvKauxkFlOVSSaZ1cEIzHED+bnng
FryKviWeoVwVqbhrxINOPGDSwxS/RSA6uJsUze9eLV5NKmvigDGMii/MHjMA7exDNynkOJWRXdWt
HZQc0DlyQScpoTVukE6ZNAzvxlxPLrhXXPc/q/TjPz+grw0NvDOi7z2OW4Pvp9JvIDYdLCyO6Qm6
d8UuY0Jc/6sY7i6m7YEGKPMPT+2nKBJh2Or+uqc5azRzJMJNlHGZ2J2M4mNsJgr1drhlMuyWzQey
nOIPnrUR7hNICvhxtV30zCUfq6+n8MBO3xpFEn+TRdIHCDH1iFDua4W1L07P6E7O8z2x6DVDSEpI
vuMBleIhln5ULDAl5DFo0mYwVmNyGtUXXljsMZg4iy4NcezYzLH2kpo+ctAonPyUytABd7kYJjB7
GrTnVWE79aqpSfUvyNO2KICCZb57gswt/RNKBam+hiuS9J7l98bYCgogSGzh45PjmqUL2y28/KJV
krXD+G2qScKf41cI2GrvLOn6xrlL0hIrx2PCT4FvS99txexP6/kO6DpjZTWHYT/qqfCNxinuRs6B
YgIBz/eJz9WRihl8Uph1VwcJ0xCXbPSDMHhoDnz/hKb6OWVGLjSyhHGXJA9G+OlBlTc/cDbcVq8E
Nvr/j1zkIHp1dG/7pzqR6G4gReJ4HcWx4c1jJtGOKkMmRPkJvh90PM8ol4dBS/WYhwD+r1/lFiMw
5D8VlN8ud4xcqlIgfK6/30HkpO/yIhe5Sd1Br20yCkZhCLGcr8rbgLFyIPY65iiCTfviRw6iEu77
GMXrHt/bha5QYky0SDy3F8tsFlmgC1O93/jb/c8+8DmqIlcndJvvMWEtyY+hKrTQkygytNn9XD0u
yCZmCUjS0uIJEoiPJ4JPw0R0b8mYlBTiBE58SDORzRMy4oJkD83Z+YF2nIkyjtgdUHXY4GFD09D4
LCDf5yJG1EmcENfJrc6FxNt73aPa5atB4/fBBynjKlvXwMLlp5gEq02Tp30pfDq14ec6cW+DtqLJ
kYI6TAq0te9x/YrdjVGOfE8ceMV0MpBLsdIqyYgFQO747gEDTnYXkNvF4ppGO4MJKZLcBIgzcw3D
051GeXRCPK9iEoTk2JH3R24jJTvcuO/dMf4zid0ivTlAlCh0YBCVMtokwtTA+GIB8T6/EWuJxsVT
2x/xaFbO6Lm45PAGoSqWqpxXNIOhrCscz4zJuLaqsg3bWcoE5fDH9Fy4WppTuwiq1o3EBABv46Ag
EfFqaqqizzDmePS/ECtJQGxH1ukmB81ZmWu2HQD2IB7rD7CuEmJH9Z8ISM3Ao15mv+AzeO8FGikC
ZPCmz5VZLD19qp69/ycw/sj7vPGV75L7vESXcovnGUqrML2CKsIObOxiaJwhGy9LLYXAtOZnOnMG
T8Ipz+VmYugV21MRKGYsKaK9CrqB/g5iAfDyV3FoyyT7fQ4t82SsT7vLsWSUK9bEi/MIsyBoWkae
+ZfgKN9glaAkycBjYieoXZIW/GywpSget+r4J6RrQkvnngkcT4lOTbo64W7yyKX5Z+T2eakd1Zfz
1wDpabctPD5VNeMA/Hwe8bsk8HCWap0ppLni/Exmr1pEPK2tB0qYQ6lFdwT6kVwUEOTvW7ERFMx3
Qzo1hIBjkmNBFK1bEsdyItCwti+obLhqR9Im3UnXXlCCu/C4LI2q3C/lsDMI7R9PgWrL4vhztHfD
gPIICx6Ll4qZ2fj6KK23e9KEfMovAqa5mcL3+u/eWcGvRNcNkM1bM0Tl06xvsMEgz9E9q5CZVRKp
0Roy0LvzntyUSTLjtTEXD9t/j7N0ze7sKrOBT7RE4WRr/eae1sjqPDJT5U7jrgyf7UvZnj+ukwix
QRYO/JgsuvNDx6tc3xhNPlTXJBr1dVYrAuAuu+DJn/pohT0T0KC/6ArRhfQD7sTAM0Oa0/Nj2tVc
fhisCVXTL7ErzmKci1PN6R95oA7SYfBFrVFW0IFmhEEMu9+fBku/rp3tCq4QXwMFm2oK2ZziyuYU
Lb9m0HXyyer0dIg5KYSoyw7kSYYN14V2KGKuw2iQfDTeuG97cJq8Yi/9R8pVW0ogLO1tTx9o4T0H
QGEgu+2Olp+2AKhyrH+A6/jMmtJVAllHY0UjM7U6qKjf7xCg2tJmGxpyPVJt6D6yt9iVEjnva0eK
eGT0kn/EjBNCMJEsR9hlyY4tq1ru1apq6iUZkairXNKkFWDT0xxeQUkhz6sJEdpWSsCY/P1D624V
hpST5NeF02hcOQi6XtCfJpLuyftSzuJHayzo7jMHzBdc/ODPR4ilhxRO8avhGowZspWAfCLyZMcy
J7GT3XNxRBD6zYmvQga0PLFmZzgch1lTGQFm5il61Sdw0IfWxYuF94BVRcIRxyRNfDoi+mqAPk6M
ZTg4njGgT0wI+ENWqGZ3XntuKkNfUpFMejfquWypABwGifNSM/8qYsD4yIwmaZZ4AossY3Roa3eV
Y7Ig/7qUXMpqU+xAA9b/F8waEqR/DxdZnt9NAVmW13YxRVwfawIi4REoo3JIAKytXTyw0eYU3Dc6
ifd6467LI8JmwaMl2AXPYszRwR+2nFIW+SsYD0txuQkXasyVOE2ylsgnuCV++id36GcdikTUvDWK
rrGGjPhcDe06VxFtvebEutbVr1nyuOXTnTriMMvznHQpsr98A8aelMf683fh9iySE1e8rY2++s02
Vcs5EnfBdyaAHZzRmb/DtnSTQqxT7JgsYFh0CA+22+/1CJ3vXfKRl21IQ9QOs5R9+RWsNpDRY/jr
2/H5dRabeJ5D6fQJmbOzrNMxEWKzhhgf3hMQcyjHgoVva3pb1chLNgTKiuNAK0t3tJb9DLwT381H
LBvEzSSg6JdVmCr9l/lHqoPlnkkTF6sL3OrSsIGLxcKjYgWfnX4GXUj5y36t4M1NZpiJKVS2wwzN
1mWJGegrgcrhSBQGUC3JWysCA0S9JCNF3cCHV9mbzB7guHYnfz7iKb+AQc6L921vFJJBvFLewbqh
J9mGpodfskxiLsP5c1o1RiRBEYkJU4aOby+bM0UOZ10GNKp9FVq+ZZfPxWnpThA5Of9Mhxkf/XD4
d0TfBP9itct9U9W51rD7ARxYZOdhr+wlK8NNY8owdOmRx8mMBy9GJSFvqu6Oy0w7/yt9kQQGRkUc
13oOpopC9BY5ZrxXbUG3zUm2on7OUWMTASxOht/coio5AHf+NXDctXhPwPBZ2LNxqeRO6S+5yGjI
UVEDE+m8MP3Y+I/DTQ2D90X/TzRQrgD8Sm9VwVymafxk2rUFhP5RD6f+v0S4YWQgNYP8qz9Bv7I2
NKJY5XhMASmcbG4zF9fIUzoA1+tmW+I+WdvjAP+s7isUd6cD6/1uSXPvDSAuPguCebpw9g4xpHUv
XdhafYE7gwiQ/MledAHwu42Q8kvo/8UF2gD9yz0Pg03c+zreCANpi3+SZwTT254pJ6ojPu/trpnf
XFijRb4aUqTGURPjLFajQyTunabkCUICrdD/myyA6x3L5+WGJjmw5+6zGUd/cWMHFdvtusDoJ+5o
FQeqw69eE79u7yCQquuDnZom/RXYCwTP1bCoaVTX7EYF/Cd1S8ewHCXnDhtxlO8vufMwuWp3TcYo
ZEZUX5pWm/3pIBphZfgeSe9izeDmXH0GB4otqf7qDNlnoC64wCDuds0LyXQxHO3RuYYbFEtp3zoG
uTdQMjRcqnXhCXL90kRKTcNTTnRgqtZiUUFQv6WkgICT1dzk1q2Aum+ruWNU//HnfpEZ6mEzMZj4
galmA5LlbdgVbMG0KVxPhV4Ft5UtHA5Rcm6JRzAxnrMp+APeyFF4EJbxUrY5AJXn+Sqsrhbs7OcN
uLioPpAYsk5A6Qvc2CG5DT/WP4T1wIepyEOpVtHJQfq4idYpFSSYIYOmcrc2RvhpX8TZaOhAaj4u
bRJVqACJL44S+Tu0SC4m5fuODKcDKD87N5cPXfbd7g/MI/lIBfq5Ch+WwOin33bMHdKNIcm4btMo
kTEr6KTSYaov1Mlgif412v2tdO+xaymvZH9fQ0pTguO4zVYITqYeFsJlFM+2JuCrckaH1M9f0zCs
sE4dxgSxQFmVEZ2Slfj5GlLqysl21SfU2dKAz6pG9LglnJaqKPYlnsFgUtRAhAcY6qdfw3KTrtq1
urI8j00tvYvWBJ1gypZR8YEAreyE7iFcz/DlyV4C8jgFqOtyD2LPMX5/CeV50JmFhe6SlWjruYPZ
uR0R8cWx6L1JFjQW/nsYnZFhMWG4OKK/VFAnTteUjbAL+i9Ii/AtyDztOLqW0v+z7PkvSAqAdec2
ofrJUbxtpGn0RZDAebC4tkKNT8z01B7DPz9dSifwmVqh9FDHpTiyLJ8VjOXzU8mDc/qLFj0NKaVO
HX6ITnQeEEOJyDpaQqQxG9XyFiOJS22n+jbBnp0D1Y73/Kx74biL7pybq/cDYkyXW1IAEph6E1dy
2VvZ+9uiK8kBiGPavsTC9QVZ2hC+dQJ7qfmomUVRhyQ3e/zpLJv2T6QEy2AQSB8Rt/szYa1Ppg57
iD+VchHrdLa60HDx9/bN6hVMkrwmN4r3j8zEqTTxLdBo/J69apOKSgScT5kKaL39NjxtTkCgP6eo
DDCvcfsV7akoCKsWnEt5xz4XGoDBS8Lk/HY2nlUYPJoTuvm92zyS0QSK1ZdMAXNQioKip5DLfzgY
iLRp4OXU+kGnpOJ4kf9kcEaFQmblo1t8C1ROgTWfWhh57Hjxk0/MFONVOZtPtBPkT1fC82IQqN2L
6e9q5TuXiIOFpeTkrO2QWfWUrDaQhP+eId3rCGtvasq/QOEhunZTb2qBmqvCxXU52Kb3wEPg3pOw
1+3Cj3Nsdc9N9lQEHLycWQizZzAImIyAbrMdlgcCaiAF1cYkvYEkMBWICft8pUge3wwDO2sDyg2x
4GJFI8wv/V8Yp7ACQMeDtmpgeC0CALTYL39mDe3jFiIgvFoHGUG+nxlaG9/rUGplbaFT0RgoJ2ll
U7YYXE1afPaKznhbs0a3yQKd04zhNqgwRIrQwkBXg9cX7P/KXkd8O4WbW+5r8r4v3RjXj1ruA8GT
j7Vv8CX3CpcrEtnwk517FQi1edJI5jEfBBmxcWx6bvjZWkYhVdynMXblGyB6a4zkuWwGw7zWwVSp
yteHrksKTxLXAoPH2cTqUizb60Ss89TY4fK835dXmBdm9ZnTDuQNwiybItCeFPH9kdBtIG+TVOSa
u0EEDz9vqu1ILpH5EXOzinNyVxGZyOE0Nj0eT+fjoPMe30xohqlnu0wO/4lUsBw8cgXWQC/rPamm
R56ts3EMNcrjYkQZ8st3LXAxsnZ0MoYmZaCh1NXjVrtNu1bUAPtcQDwgGZEDezTYKTIjaEJ4V8BV
RLfI/+vzJoS/Kjvl3/kia680lX2Aghq/KqHM7In35GJaDBvqSBvEbRJKOnXDTLZ3Hujsvo+AbiJc
N3HwJyTlbH0AL3oQS6J6Yu/5Y9q6Pp8PB0ybrN4rPCsJBtbXYUkuqSF9/d/DUa675N+WvLPI5hYd
knghT0um33IyMldtQcgBgO9Gt4IXoScg5oM0QHqXUZzyScsc8ne6RNHeMwa4KBURQwevb0IE8M8W
PZrEA8IkjstIgVAIhLBirj9uCZX2hcqudNCPiFbCOJDBXAu1hpbGtpRVsJB2X+CQ7FV3Rr9xrYsC
jXF4ezywDd9EqEjhzolaeck366xHCwZr0aPox1NU8GOVhdurvy0Rmrz1zHPwPIabg4fccAV08aEH
yR979XBqjUwY/9OWRmj/0DnLnrHGmZtNn4h2egSooOZJHeCNzivUq+qG6YljId6y6U69XA9OoKQj
6CbsG1MBMgFfa+/ctAXo+ekx9qWk9nNtJryo9NDxNEglGTfvoAtrF48EvhfkmCkCEwtCxbF2QX+d
5nHm/45lYLoIyRY7qQ7/9dKpFD9bFn11uIMDdgPV4TAbkv3I+DnWCaesl7ZSIMXF95i+nkDmmXqp
ND2HRJxGChu1lf3SBmJNdLfNbh39ZLPWJufYIar6QaFt1U9HPJWWAXvbHDiE6bxwNg+rQkMBKgjA
iFL8l2Ms2acbn3QE2OE7odVoG4qncEGN2/5T9AjI2rExzQi5P0EkzFa8D7r8nAxXFtn2sUxLbBGZ
b5Kc6QTtpmiicB3VtOcl3ieSJq+LlmdLduNcCQX0h+0HG/7V4gUCwEbinmgTAiO1PINMBK98YGq6
hPMQ5ozMJJZ3K3Eqj4nisSbPjDPMQXqgd8TuZD4uVaC096FMdQkyKk5gA2RJeFRLpGWcuSfXcckK
7P/0vh0JVBR4UtnIzcE8hDrWw4apcrM0ndjAiiYSGDPa90vMro0IdZY2f/Uz9awj6eVQJC4uUM0A
UJYyIhblgRRD76D/fJgZekMwlxVj05oUqdLJZvHhQgn2QYLzyWV1H+SeOa/eX3f+J1Ngsl6Y20w8
MYlPEBXl1XZFfdwxwI9Bdu9Qie4KGvx61544Zk9xUH5d0gfhkr4DxMy5qlDYl40GhycNJswBqI5g
9MRLHv1AySYLiSiijSCo+Q9eZgVPejLPRuc5ez3Nn2ZdD8fKG784njvHZkqLuaeiwQ5jWobtWUh5
sXAaNnrtaKaAr7GcdSOYwzUPQH/m10vDa967D5FRHOl0vpng/WTveJl/3T/i0rlWNiK67yf6LmFH
XFAVRJ/X4Cbh5NO+WeDdFqp/Gial7A9J3y8uq8BgTjhFrYan0hR6FmilebEry/q0JDXYDxPSWOE2
hMYVLvABNbpUUdkbZQYhfpEVom6gX4gY7GzlEw72QZds4TM49St3qDSn7QyEMaxAbPX/cXf3G4sC
KmH0f8oJJTuecMr6r1Nn1RQFUgeUXam4wADzRdmi3Bt7qKnPEirbgHrV01WWOyHQqoiXzKoONgVV
wCgtIH8Y7yq/AgSbVFFcRorr1d5/60JHsDXBTBgwIgIRYj63mAQOKXlB/hdA/wPGUWUUZxuEDl1H
EiIgfLkxSKMeUcPd300rgZ+J+88STkGkSRilJxFyRH/GavHYrqjyHamrfLwT5wxWluEMtXmktPdz
fVAG6TLp2WPWKX/kg31NY17oMlo0+Ao+zTgJcFGO90VQAEtVuoxqayEhKzD9pAvvvQQWP6OcEFOL
2oa/uZZ9VWPZ1ObzzG0Ro2yHDB2pIsQ3bUwy4TOgDpDz834/axKuWQvP1BjuPr14mNaXosZxneQ1
lciDB4JeG5buYrCW5pwKzlM2oyfQ1OLBcb33CtvP2O70OE3K6wiLWkZhc3kPW+MsHpsReg9nDG7o
GQEuNFvr87ZsPinjlBU1SG6QylpkUk6JQ6cz/c0wk8FkblXePm7LYCE4wfKyEbMo8mnTLwywAQSa
pfPpYzMt/3B65ERYTDGDjWkhv8OMkPGShasehFx4r2TclqVabWH3XpurMPq+qSUqTPJEpWe/QemH
+CdDIr7gQGsBzj8gDHF3fCAV9uLIzT5xAIcvFzULyMaGw7T82dMG5sACE/TYqzRtSjSe6RZH7l4q
EtVkrMVWqUIWSvMgQx8KXmegzzPhVsGcOUbsmVZNAMhssQpo47eX3kq4uMhfg+/SuyxOJGLUvcjD
NM2mVDcSS3evGhPfGMKL28wo6uXe78xEEfGNf2MHMT84ejCpI9RUlXlfEhH+TxGsl2UAnqe+VGta
ZY/sQVAXYpd4H2I24RuVldrnR/co77lwSoHCiI9h24wwFaUnSoGhvOKfZMJTaFrN5nyqjPHjwjzh
HskHcSyPNYLNGAXVDtywZi/6bGeYNEVSAiSr7QyVXvpsOcaYY7soriETyIysQ0WgUA37y0ZIyOTE
9/9WzfY+Wrin+FnhN/GquSvhUEB5hY2ILpb58nEQATkn6vHKY6bqMkzt+Fh0rSjp5koINmO3IRYx
qBkw7NX88MmUclH6pPsOpm3emuhVzq6+whuoGHwAk6lIaPlfQG2V2C9GwIdZxMyKHL1ssKHUsnOd
loIaIz7du91U+gQ9+NQ9HPg491RlgwbOdlCUcb7J3hJzCRo8+vlm8PN65vxYAiNGrZRgir8ETXvL
wJuCxwfseZ0KocWKLPIO2/az1hR3PhYXsUNdthLmPtmTKhYaKdlzEYrCKcFxcgS4j3PW80MxHDJo
HKvRzaxAKI5pjhhi/vuN5dEmlw+pljoelE3LU8BO+76DmDW3X507STcTR/I3CYlN5r35P4YwDEO6
YCPUsnRPstPbB8Bo051ZbCeFGGV1RjyBR0UKTLMYT3r+YP59Qutssv2cOJ9TyBgw50lProSGhgTa
Kh5ZBe+zSY7N0lvMt39/0Q4GAy5PcIX+kJ6ZmrZm2oW4C09Hy7hkua4Xr0bbuHDU3tL+VO9v6O7O
VwyL9KR659sdr4WBb6FgomLrbodCbisy75bnWZMKSwcLrkT9at4n7ZVOEgaGehDbYZWfJjjpTXc/
j+tAxkjTuHqLRPUPlfSP2oahUKfMoEn8EAwLE27hYcaEjaHiL8dE3mNXPSxUI6uVAyyVDIZZPNUe
3b8SKrJ+XwBx7VjKWGZp86ORWKMqAf2DpU48AHkfacYBEnLiqeaLZAvOOpt4+HpiFoq8h7qvJ3hx
BPhpFkB+t9alKNrgTx6bk5qgkU6NKmwoZc8EXg1P2RpCKmELESmTLMMJC2tOXQL3Xpz/P+9Ak8VD
64quk1MU7CkyAaHFAAuRNO4WKBhOz3oqwZEQQAxIMft9EKoqRIzLy5jSViMa1yNgLAWL+y8XQ0Wo
+RF/yvgECRftdjE+q9PECsOfwT8gohMxjSF1nJnqvjwAJ73d3eniu/LiMirx7BmobTns5TXm5NNt
G3m4SzN+jdwUsKNozShO/TFTcAfM6V3WxiH27p/acVE1GDQHEUQtAKqYas+uQBh1N4zvfAy7qdwr
w4NEb/uVFLNF4l6uaAnyaSZAi/WEnIMxsblkhccdS7u4VnDIu/6X/XA/7N3px4stKPYkv/iT1U4z
1HJ8b7xZygEwrFHFCrVdbM8k4qy5MgbPhFe5JbUEttUAecrx+lB6oJPcb1Ljn8NdZ0EJvlJp+kmR
FlFCc1hnlwpWWF0LeyacqxZ/Ks5cX7mJ4eqmN7R3MqKXwMUKK1VmFWNHoYMdY3S/KRt9P/b7+Kch
pN5d08MbF0hIiWd4Yrd6otpfDNv1ppubMEJNufErqFToJW2crUlV5+LC6Da6IVlvfvAZes5wqH2N
9IylMramjCve/ZdRDxRFJm+hI0TsPEe9B0OSq5oGUjoQxcRSDiHm34MoDVB0SRuRuwRPYJHV+Dig
fmJM/6nyNc5LA0au6/FafjY7yY0hqb9bdeHYk33AGKrgoXpolekstn+jZQx5B6wbpLZbxFkiRs7L
Z6psLuw0ns05vdWMm0Bwr3dM9mrkaQxSDBanKuPWXwJ7iAGjJQWTpKQpA6G4r+u2aMI0B1pF0p1V
6KGqHMLc6VnqVJD1wNVCeA6k8Khf46SCjRQJ63/pO5GcGEUDLRLnr40JnJ1M/mp5IaHXWjGsV0yP
9uNyEafgsErUU2iejdYjOeAlrRicZp+GPfEw4wt/705ZMifVUHqccSQFTmfBcSeQHtUfi8xCS5dx
uN+PuciBGpZ0C1J05g0bLYOWatxz7fMZn6pv3KV1V3rDGHcqLDWUeIJx1saOfZRBsSdHXyjt8tA+
3Eh2aMkHklGI5QgFn/Ah+zJ10MGQ6B8PQRYJkh8EoxX3r1L8s53jA348vJLTyy5qGrToWArAACkc
irxIDpj+Ve15P8UN+v9/Ovx4mn1lWOWKntBY2mwPXL5jInppr6QGZKx3Ih5vNEGQta5fVdNZt+lr
CH4tcQ2kcjrZCuQc1qpqSG97q7xvXvfQ4IRiQn02J681KA/ZL8SFUebc1WINzstNUz9mgCcg3a8M
EtghMUf8IUQfYYIGoaiViaXG5yFAeEIqHnoXsONGFUlymfD1mnhcmgqbqqF1iqaIMXGYl1xXNN2o
KEyaAMzzm8Qu2+hqsEYNyHKQqY0ZGfZVqleLJ4jS6YwasGLDYAfUWtibrBNFaWFrNnoGzypCRGCv
ZnQIwpYdrzzhU2YWIuzEUcdKymzKfHu6OLzbnzr0PzNzowfkC87mdTwqZtxniXanfpwk5VMRRLdf
mcK4PvbnsgkghCEnjmGqON4zafZeDKbZ8+kmT79W4MCH5E8rkQdeKycDfUrwujwxocgiGBDUEJ6d
aq/PKoFH8INGDa0n0Tk02+8EmtFPDWUeDx3gIyjav5IMJ5D40akx2NPMmA7Fk+s+EkL/O2oChBxH
oyv+PVMxf/EGH9xc6wZOhA1uVk/OfJu3VDgix0bIqf5k7ecelkYDg/Ba7iew/yaNniauQhF9UfR3
QiynK3RLRvR+gyBf2mbGl3Iz6uQtiDJorPcVgSW7zbWLuLTfEn9FiH79YNoS5MnVuQbWqLmHELlu
7SwgPTnrktoyXzFxodnd7mtk5RaH/VbgrRFxt6f764Dgoxu/71Y1k+T/Uou4ntfjbVuqq4BfMyB/
pKNcG2fcmM62dbf2iX97JfQgEBiYh/VgnJCxXr7jkEX3+rsJebRQXfBhqWIaPezZ/HlzlyHmIa3f
etgu28kxB7mEZ7iv3qjcrcBQwa5UGpdiWtE3BFRv881sKQgsrHvN7r5MUY4TyjeKMica8vlxAs16
aY6bXlCJWMQYoHrzAksPF+0c7B1xMRCFWbUmGuw5F2OAwIbu57GD1kjrfH/B767bNidR0PIZskqE
1lGddDTlwvOWZjvLrL1tn/prh4/HY9ll+WG6xYdSfYhBlkhtldHXz1QOcInaXUMHteo5bOzyB1dG
9u4VMmbk+IoLeoD/AtWRHOd16BxeTTT/HCJq1r8Ojrf4588usD/Lfy0vglSE74G/edG3EIOnmYSk
JT3ke+vEqbs7S2pw+zM+orFI+hlR8NSfjsNebhQb8TG8WlNauwC742fxKXShKZkVra2Ac4/IGRnC
U2ZXPfwO57Dbi0aOZCInDDPpC3MRPHCNb2aRSgbxQkVSY/McA8PlCCFjrsCY++KD1PXZUapj8VU1
nt7OGH4EEh57HqAejN98lrgFV+7PDLXquhp8ri2SbKTEV9lgrphMKBVxMeBDM1kj5DuMeuw7VhF1
QIy5Z2FcX+pCOqbML+M+fg9gqP7gHwG59/YFP2IRlK/X9NN1mnMp5YPp75P0nZecB3Dq9nZ1jwvg
U8cihY5LUdUNr0dx6AAfFquHJJgeiVFoWQ369B8X6y/cI9TIuyoTJ8KqOxo5J6szm+XkmUjoROxk
jdCmpcJNjGfBPpW+Mkz6Em80WNqmVN4iVvMUoaWfJmflVOyWCFwS4GS2cJl4zayXJMGOqb/C3PLs
M6WrpGeOmA577mepKLYo3FelCx7JQt09O5fKHoGBMEvvCIYMvMl/bVlITlFHQrCqiiZiVLr4AbvV
fd8LzzDVVizJiRV6RiGMUrMLgwzG259a5oZYwH1zbtBeG3O1loTUkFZ2wFHer4lu3Mn6mPW9xzDR
WH/+WKPaeHBWCL3WZ1Ns23kPTM9MlW2QeF0gO/jc/u1TZLWmza+j6a0ywwVsv8yzlaNcKmWrhQGL
mJ4gdYUZMvfMTOLvqkXKiImpwgO1syrf8+CUCKjEyErMRDjnSCyE5FudhRgQZmFEmB9LaFkb9lnk
EVQ5Opcusfs5+FatvaB4pSvQflFtFT4rrkw+3vgdw/arNzlawHIlcRCeWDy22A+Rg2gpdRGDe0/W
qmaRCOSgSNeyGd9GAyrZl9WFVw5u0ULA+z0i9hyf39IIbxxF1sVfWkACdB76Qd8uq1pdlUfcfiyL
ND35yYVXPjI7bqeoHsNPr0/1DouoNA68vDSBCVhfLzBx53ELyVapZPeOoplAlkhLr4Zkw1lMhghO
6DX4Ugr4vQx/nM/ab4s9+u9J+bvQjgHfPkieGvQQgdPrWVFkQBCosZ5c3JDtYMf3kSvFmXbWnilO
a8hJ52szm9yDjaeMTu/rsMdxEzg3VJgZYbDlmlioPSaTtZw4Bd4VdIfOf01k2lO68D7ZxmUrVJiV
YW87kjuiVzn9UTF5eSJEsgJQTrmN/x7c39irpUGY8llTzMvZ6hce2eIjLN5TeCKzB8f+MW0mMX+v
+V/lfFeUCOP3/tV7VePoJgMihq3XzTWEpqAKzE3QDwGUhjyUKnQyr2jkgPQyFzlqyW5XbsBmEUWa
dxx+eKEX0aYEBvRT4GurMt8+dZli3NpO+dtM4YsoRcMNBxtZoHxh6XzEftHsM/2+490pt0JNRwhU
pgZzD3NURwuTEaST8dQR9K89P5pNqj+24c62CXbJk/u4jPCq1RH3I/Kxyycpx99jAxaOawwdqQGv
w8p1DlnRc3InWxesntkxzLOJlRZRheFOplp0BQO+F+0BVB1Hgxpiuqaos/m4YEE+vQNCRe1AdOKV
pwVFF5Th2sZRHCPBJyX9A8UDxNm5a/O5H3qXFml0AFLBYTZuzaKE84AE4+/+u12h8bjqQjmO4vFL
aXiNIn64ADlM4TYWmVMMpPW0vwBGUcWAkD1ywxZ+Xcpe+omFvWwczOCT/w473cG5HijNUE7EuVvw
k9C+Qyrj9Dii//Yiq8H9fvh8NPS/a1XeL9MTZXNqKMjU+RzWf4BRpJWHQo3kklnpmcTvRiiSJaHp
NYZToPikR2lJgL8juC3jgE4ARSLob0/0AibPfoxQO59wdUfW32LwElmgFv0q7nX9qLjaC3m/C+Gs
a1lNBr65x1jEniQ433/85UH7iwwoDtqnEtDWp9lK85DU11yLpBOFTjIhCFAEYuyjbWWoaEoftU1h
nuwc8xhYilPHzKfxz2FdbEvj9BlrBWBJIbysybVHW8hDsogUJn3XZiVoJBu9Qz7KGkbOIAhDjarc
FyJpY0wZ43/8V/t9k8/26cs5DBMVz730hitbGuSjrI7jzGiN6FdahUj6Urcsv9hC+ivlbsVlEYI4
TdXIDnBkTMnpqUcgNlx3HYsMQuJ9sfGbJWAnAxIOfmiK/A2mny7OHJchn/0RYfF74zzRsPvOLXgR
qn5utAwmgCI9YBdyEVaxBI4Aluix/dXHWX2dp/mdKbBskcWeQZ0OnIoV1wfdluIqRCAfH1XJRpLj
A5wOGBmpSjoOLGAe63cQmBUCfHHuPAVRll7oiklRQ11px9mcozEXsHFOZlpuuUfL75R5hdPvsIIp
wl93KvULpI20Lzwd5lGRNcnGDLOslpHgIbRa6v4Riewghr8AIEGkTGSKGWxeK16DOTA4eUkOJ8FT
7zoIptifD4gbFxrqCL8vEkcaSw9H8OcTBDsgDYAiIUBdPszf13XqzRi6Aip1CcrF+oi13weBe8jP
KutVm/vTukSTU2CYJEg34BA4tDEQCm1YCij6P6ZQDGYrA+O674pyKGV4O22ijRTGp5y4SM/mV5v5
pjY9MFwtuxQqH6mkB6wZc08bHNj6jGuM+LmCu7kNnmaObdK/yLOW93W7rsZCgKSViKBxHFl9NxuG
JE9pELkio2B0/7BuMhaLeLyQ47bJYAmEysOhBua/uQ9vXTZKuRVXLQxINATZCWeLzw7rvclOebmy
AMXw9acDTPybz2xJj3NEPpypYNC+V6y4aRgsFr9BpyjO2ikgrJTP+eQpK6HyA31vRWjn5uLm6Une
3VS08qhlROHNutZK72fHGRcFHh+5eCF7djKS0zB+a/cZ/UTzMbhv2pjDuIP1x3Xbl8+wOWc0jnRq
p8cmvolgXDaNNqMFfNIDCB7cDSD8TC80b+Xal5SnY/vBXhnJH+/iT42+dxVReuGrovGnt+yI2s55
NKfb9z237btFPBgx9agS2QAUhVeiaMhhMLAzTgVH3E3L2//Fa0PYchduUX1uBENZ6z+RHXcRglkn
PduqqssbDkG0tMt0UL0UKSNcN9de+CVJeZQuOCRdakI1yDRQZFd83Oui2sYg5/yohMlxYcQ2e/5G
h9EOqIRK9MacD4DK6jGnOLaXk8ZxbdqGHewCXdCk7yq2H3VVWWI6yNA8bQ99Jq0YuqVaq1yuaYdD
Y9AKLa3LIKwddpFZgdM24ed13RIyjAn8XMNFkTF9aU6EtMgAzFwmPQj+CrasK2PQL+LpO0Kci80U
LhjdX89bwYfAuczucBKYzZtgXXoUO7O8xLAkpiUdEQl2WC9S3AjqFrF6ofV3SmISAaJ42yHV3J2p
36eNtWDjsFmPfCOnXML1Jqo4PvpKeuS3vP+vSsv3BydmCE2H6hi8UydcoFSFnYxq6HUV+tCWbbjQ
g5ymv9kRMnCYvl/ytQqLs4DBVgV5ftrAgguFwkIRgl8xJln8+xfgllMqVu6JStkwX6O8MhGcPcKJ
cPx0GISLDR3bhRq13yEcDA3UOrZQ3Slt4wBIUkvOLAJ2XyQr76egAN2MhPfqXaPs9nRyskjaY2+v
4kZZClyhAvF30fy5190/5a/yxvyJCXJ67vAauvCK5yOJp+gRWDvxe3hjdQMcFg2Ru6Otp7fjKbrG
tyvliCOu8JpYoluI+BABMaOJHQ2j1nYEv+67PQ8wTaUf+pCRsGjVKzd+CyEQc6AaNxFuHJDH8mWU
J1jW9w+iyReJdvoR4pCQ6vd8dsLFhHGYzLCUzUy36RUuCNfIBdo66TaBOcJM3+o8QTYa2XaQ+qNl
xaUd9g7uBn0HT8/z3Q/IxoxX2gu3Az1CQkssjIpZcZMJWvCeidJfGNaTeIXYJINHrkptJW38V0ba
tKRo3kJTrtd7xRBEcLkyotrUBCikNQ5AUoH8k+F225Ji+ybUGw8874mq5decWjtBlsmfmHCjKyCH
NKFkmptpI6GwDkJ4UgYN31mQakSQxE2xZSBBTlFvb42VRBrMWZAKBbGJ8DB59nFc4AmELWrc3OLo
31L3R4Q3rjZrBiA/O+AR/+AigFQ4fp1jB68xq7hMEniLK3YvMSTWcmmfXeHlrdxVoY++1kzt8a5T
7uUOPMzt6iWMnnEupkRA44LjV4wf2bHtGN2WXbEAH0w2cHoEAdXb1F3x9PhwpDltx7Tl0uws9DJa
ZKM1apgOFaBRgkPd+H4l+jdBClQqcNAhZY5jOyu4AM/Nx4WoMt0TZeZ1o8S31otg9L6yqrijT5NB
saGd2tnTUKjE6kOCT9NIDnEfoBYwF+cgZ9i0kXWSYIfY8AVOvK/drMxARJnNGT/Na5RmWGpts2g+
Nr07ppRcUlBy61jfB04e1ayp2t3zJC7zJXgUdeOm7KAN+2jGdsb7AYxPjGCU3/IgvXM3CEWjkQh5
XIXuBv2JALX/tERki4H1W7ASoNjtRRLDBcXhE+cICl45Ryzk1miWkh0HtN19oM+4p3DqisKx20ku
N/gPNLrV+7blW0GmMb1RDphEkIFknY9ndSMZuDn8oEOmxa0bZ5cq/c34gC3KdCqvDT0oy3tPFRu6
SNHaQWgTqbGD1XDtX4ii6w2b4fao8ATQyosRiAEQsInJ6yJ889ujf3RWrX6xF2kXuChySSG+Sn9F
/fRA2je5gt8BJmzGtyAfEHueR1X9rhZKY1W0G51rCkcmMNxLmjwaESnEpqKOAXRk32tjv+itq+Ik
t1HjJZPb7+926MyNXNvYcosnZu0Ksv5G5pwXquzfUtU/M4AHofFrPFILaDXucJyp5dAzRp1r33tu
y7D7fzyv0iZDFp8EUEXI28WYHhLlt2A3AhwX07coWSifyL1k2Yx5a/ZDpZWdq4GO3sPM0/tifH2o
VLwyo+OR42zI6BSA5RUKsYh+ZGOBUbFCMLaR8V8ixRrw3Cw1500ioV8kwIUbCgR/vVuPVVUOV7CU
vhiyVyeJLu4frEJNsvVOD/94TDNg1G46gapjLIN3jGl1N4YVAPp8JFODSGrESJEuaXI7KQrj14lq
d+fddKM0BMhL8fWB+EiHx84doN9Gaj8bbMwUkynrBdhNZOFkEvRoYS4LigolABLzFd0xnP5RAzka
1O/qPCtC9tlYPNYffK6HVOJQBtKT80ZU5EFFEmM5t5GoHWk4CemKjGrg4i+9tFmuH8sEJ3MvLCDl
pAMjxfQpfz3ItYexYTYOutvtjdD7X0LuSUSCpccYcO8l13X9zn4T6Qli3FaZvRO+a62lzrZSfNmM
z3x/UycUEZcUuF+3xHtx6NoMqMrbOzXzuEZBsUz4tlOa5c2ngU7nD0KoPxtIYV2m6JyDdHRr6gF7
VCkmrR4sQgsE6tX3/6m3qYWWWJZSK6q+4IhpNq6iKPx5vjgI9nnVtug5cTA1f5MsbbXqKMWm12jc
C8YwwSM8fo4bBhFnNkR22jx1WVpfEzI8L/ClJQet1Hui1UayIR0JHa3cl2Mi7S7140YeCHxUo92n
asTiqpySWFjiTK8jXTlJ2+8Oj2bZROmDnR9bbWwmbSqSZZ2nTMaq1d8Kq52sJ0bIqMG0qYc2VuZG
d1MdGcFQqu4Ff1ODyhP5pDQn1wxclJhCyLzYltb/Shvgfry74Qm6D8SFdMVEsO+npSOLmOOtXd/H
R+Wrd29OTaYM32vs1CcuD56cvwck6K7Vld/KPLXfGWvWgq5rVGJwEZjZ9MU3FXzfAwOLzTnEEbeY
qZicF5WgZtzaK2QJzjlWY5g29ICq8tI0VGwyfrxtWDyagVR86rWaJs7dMXCldEppU5yafdkowmFJ
Upxl8RFTjPzuvB9UTMUT3enQ51IN3j4TNcVfj1tMfGVSdN5BV7lsUlJs64rZfHXGa9hdL0MwnRR/
Brw1ZUKlyFankAX/7Af4gpdS+FfV6EmDYH90XEICQeug7qxsO0axGstxsSxrk0jHP/41fGsUmmYY
MKK0daiQbabBR4/ymAbkWnCIoGvobcVzQNk9NeJo/YsEjlAsNW95xyxEOFFHKzkHwN1YPwsBDq11
ksK6L73GvdHRV834BjdPy/jJynLHxClKrUyFNTLxS/p1afC65T8/Epgp/z45pScG4BJyruRKLWy4
AuokELSpWzBsZOCASLnxB+jyRMOThYt/BMeRjhUivzd9TsequFwPbUcMBjhbrMfNnu49NvTEW8V8
LJdcKlUBSIsMaQjrQRForXifpfLWDGsRNj8zxZ1CYh6Mbl7yV0QlU/BysaX+6eFdlk5QtjHU7HrD
2a7Xguy82S9iVAFjxEgQBG3hhyAEz6E3skBbDnALJBbAfts/ZWKz4LjOBJFc2p4mFxIiPhI2nDps
74O9FNZTbWsHtCm5a5DG55jMpQOuPhIQNVr6IY1uBFcgATdNYnDeQPHdDIh4q7MSzUfXe8K5wtf6
e3xeHOwf8a14gEEYPvd+n0CRD2uwvvoQdz5rIQkRJ+kmFeSS0Q5WNaQIdQFlGGgjwTbs2gmzxkWc
q5tYfFoYOwjRdCmj43ulQXVp3bM24CUUllJJYFQlHM+t3t+beacv3Ma2EAVZjm66Y/qwb8lrasDs
fS0YxqR7CVWFFlwDAJO9pecZghtMREt/kNh+7daZdyjmh0g1jePH8hNWNWu9QNHYwFPe2Pfr+Azd
v8QqkdIsr1sMbB6//CjlcAkBBG8ECGEaGyAmdS/HpGspviTtXmXhF3+o3cOom0VLChtfYmA9iLw+
cmAlAZIOpABNbXrRmmV3Zp37LfXfgbeYz9UMO5JSaWha/UdEPwUx2GUIDP0wBBSdSpQkw6Np1W6A
MrzwMX72dtURXGgesgldEPf/teISjEJfvKiTb9VWjSCruLoOAe0fuler8Xw8iZLa3S7dMNvLBBUF
c1gX9GvD3rzWKO/N4ePBZ8vJa1xYd60bZJ1fmrR9MjJ8djFSdZQjX6OkCuXMTox6VUA6pJSvYaFW
b8oaLzRv5a5KEEuyTbe3p8fO6Jx7+87gbyMRVfo612/AyxUovppYlu4zaOT349UBtj9C0gq9bg92
L6auPlHMeSvvEKoV0pGBzsxqswZk8qip26rbm9NvOjSo1crc2oHwnVbpZ5PJhSv8sXLdmr/5icDY
xgLPPD5+qZU7R7jQV4zqWcEHHpkwq0dhIupQ53knsjfpe5W9rX6vTJ2t4+mVwSxqI86ghvw5jcTo
U9WsrQwK9U4ZxK0Ufq+vK0Cz+v1bi+n+9tTrtXQOwpF48Y1hFdgJ0xCXFomQoneHjL+T9OEYiAiZ
34qfeb/BdB2DqqcxsTmJZG/1ux+mXtwzHz2mqjIGEVY4kotD26979TMapPA2tUzJTQjx+tsSIBkZ
K11afxqcqxJzckLYgzP+qd8BSF8iTG4K7fZuNWP6InmmJA5vUP8J9rX6ek6Z/aoyJ4C/pk95jwJB
5BGiEd+Cingg3ErrNWEu6vtO18RzrsVYWiDMZyHnd1LTP1cPqCSLBi7ksjpCC+3yBkzL04RVDADC
QPTmFWxxGrcVh0QtHGjsOjFFi0qA+jMQNNyo31UTU/pIs/czQ4XE47e89PgI5e5r7TEyFd2D7/FP
7Sf3AvTqunq9rr0Y9eIBleNigVPFHQAXXaBX6K7BPrgG/B3LcRuqCnQS2CQ5HIMwCTa+isBQnMTr
eh+HgX0LoOkPN/mVQwlVnlx17ghYyy6aQ0GFez9E7cNclWzZOARwmJnL2Z0B0Ysoey/GLTJ7fBHn
LnnIXEofCWH8VUP8/VZv3NpzRSsiMULRyedZOkfziMfKey+5b4EKzHNeqUEBsQZ1S04cQi3T2li6
jzl2dBM8bz8aCUf/V7pDq8JNWywvg8otN6zqXOJKLO8id1yWXiTMZf3AvumLwq8TLRZl3xazfJUi
NB5n6L5B0vwA1EY+r06lIm2ovsTQkroGDqzsz9YIspfaBZ9zQaTubJkp7KgZBVNQvnNDtXF+3eWo
RTwR/C4x0va4IlQx7WZ8wPyP/r2j7fia5iZK3rGHn56+cE65Vww4k15LxLwTmgCBLfLOS3itmJIq
GbY7LLzrVYMlB7U2PwqUb4jqACjdbIwieotIBkTWOh+YaNMB0IAXGa6aKVZZ9kL1zEHSay2hkgsm
K4jAqHhxwV0aOsufEn+wpMeD4iZzzn5HR+jBvYFvlcz0a+6Kb+MZODbhJnB0vYaiW/nACMyxu+Sw
RNlIQXoPwC6DQvgNOwfU0yO0vtSaeUgzdwHSCyVjkNkJXw+wgvk1LkwfaaSANxOKkPeF6zSEuCCf
E9DGdurxrhIQ44wW6XmcwPQn8lq8ezjoSQ0KZxghsX1Fqo8KzbYgmAsL+um18wCan7k1NWDxy5pu
6S1UJtNjwEjBwMsuvqHErj5iT6CkX86x5NrMKKPv8C5Wy0DCPP2Cb2sDmYjyeUaoY18X456fhUqm
wu47oh3pSRYoWhegvo2WvowdZLxT261skc4QAZnXta1hU/GSdYivlxmwiMNFXyxEMBnQUTp9SYSf
Rrb2Vx8k5ax5+PUw8y6/Y0lIF0uNtGL6PTI1TPSgwXx864ZhW6I1ci/iCdJh8OGhOjsb+3VzcXQ9
KWoJJxkSq+0r8b4Oo/aE63TtBrrkDPpKVRLtgwzj1P632DVAvIe9VWVlfG0rgYxGe3xnmwxLGJVE
axVmz9VIaXNnvum4kt9J1Xy9PkNWU7hzRg+ii6KbTg1IMY2y+BySxWVQXAGpV3C9Y0X1wZbkY1PK
0AYngYDti0VC+FsH5VMY0swT0kEPJ7CWW5Y3xJRFopn3hcLseYuWFy3orvaiOwqRaD5UNdEqXQOS
YZjHgYSmNsCvXaWJSBXVerW4tJt3ozu39IqjCmmlGQ7iNBBc5WimZMZrhFKYTYW0rXJ7BgHB3BNI
kOFUgot8PWMAC9sCEzCjnWr3gh0tI9wysqoCnflpPNwGNZf+i3mJibI9Umky1IiKXuT+B5JNHpbu
R4IJY00YRBQbbpoN4BjyE8/ZxuAfgMvFxggn02BUhiputNNhKHtvE4R94WRfNoEJNcNd6zJbXyD+
t7jrPZMPvHfNRsz+9VoC9Kl5muGPbMhr3j1zA4a88uf6/kbFtxWly7t6ANhSSsiPey3bnAOZg+da
zwDPAQW+UGluciuiWzWPhYPH3w/HUma5IiO4c8dZ//HWgWsQQeHxWEOpKKZAJXYyi5TUdATyX8Vq
+mderzmfNPnVzcZG4vQZ+1s7d1w+JX6/c81anL7QByVg/kdKVQKqbujIw/ZAtW2J7/bo3W90D3RI
lYY7zQOk+9HPcODYkXya9Nu8YxQHwzZ/HfkZZC2OD3HUlAXYEvuPadbT0TYLe/6aMKUEQqkw+U1R
i1rbxHKNC78rirI8h+i/HBVuwc5/X5bAxN7vACjbv2RxFQS57J7twPkuj8ho4TbQshbA0Ahl+oVK
ZcTKj/DfX+VYDKZMixCvOBhky+IkT+2+39+cPrck4NUfzQsB8RkxZgyvWflcB345NLOiEc264GK8
IoF/sfoPOFZX+vXqU18cqa0Zpi0VCc928QATos+ltlprONlao2WavlX6FNpEotmkPGITxLvP3AKS
OJ/9bo8Poq6gnST/BXAYQVCkSXteZ//MST9q3qwQxGJNbYF3DAs2G014hI2sn/9hGD2042eyoLzQ
/KEfXIP5HrjOG3XFtUfFJTAYH4Z6FZr1ZNGaT+QDkRYHJqj+38El81hvVnSG+AVnADKcmgCVQUiZ
kGRxdPa2yOTgWyk9Puv4FfIQoaXIndPgcr3x5KoTFn2qo6lXM4do83jRaXf2zlXeEi04/fFO+Fs9
DU2Vb3Y+Jkr1zDPEAGJq44//Bif2Zpgfx+1+exnEXjIApPqU3ovItY5mJntcWVkdkKNOD3sf4kkc
TAWELT/7lz4sRWKe8401mB8mASxSbtKAPbt1TsEiv/D33oFsuyxMbyRnDulolQbqDa/85RHKIP+d
aRBaXWLPAEmXP9vjt6Jf/hg2MSvJepkMB12LDO5zrY9Tqhdwm7fk7ltGgg2zI+meMQ5QqDtJ/1n/
zqlHt5UDmZ8P3KipxcmuZ4Q2ui+J8u7+XTHpHuWd9D0oDMlUWJJw+BdN2L1EyOIAC+RUk9SqxJHW
qwKAD/uWcF2ptWYAev38XAY3ntIHeYGIL3dE4a1T5Y8l6uzuIFMKPCSjlb5Rx8Cv0C5h4aniYA5n
wm70OgrYmJB7B+xzJ3q0715JK7ArAvUI56PFD/Jg0RDhgPthumSR7BHICLa0s/dOPb8UX5K5q1iG
y7ZN2k3zIm7b7AVTs/zVqKQqGyv4CtJtiGWAenoA39Y2dJc9ZKeAEQJINEvNIAv9EnsV6pNUnfXN
U/i1uGUb7yA0XgI8bcMOx+PkNwGEXeo0Cx6G6tdgL5TLk9/AojhQlIddo1SdkAYIWAW8sNTESzFg
wu1CU2zBYAgpfovvdu3uFRgpCS2rwcnsWK+uC27HX1L22syr+Y4tI9rEJZZYrNBYVTPi/Ksux5RM
LtVpy54737YhF69QqaHigHj682ALeXXKIWV6PkjhKRXSEjjwks37WliExsnMzykxhj2AKlH811AD
WOU1TttiGCDGtCEe2av0RNBB2w8kZeUx4DvbLH/7D8BXRADknDzys7302PdV6Jd9RlCLSH4RREet
xlr+50vswx2Tbk5h+b4KkV7oWaLSuX6cpYOgEWVA9zO6ZOuwQA4aR32TeiqRWjP2hlQfsEZq+g1n
aG39nH6Ll18kinWKiiEwwKbtM8OCJho7o1lXOMhtV6n2mPrhMlD9oWRHE7+ZU3s2L+LfemfZkh6+
CyfnxZzGEP6VgH4Az1vO7778/7Q+w4lJdi2NywhkTY4vr2amoZx6RAddelKyy0/6T5ZrWHJhMKeB
4JQkxrWQ0TfCjdj8SK7RY2jD941MgLJeCrx5Mb0B9WVf+AXvnQq3P+QdU353RgTA5NL0o4XhwrvE
P98D3069t6VA+e/xvyW6BwK+jqVY7o90fh/sqeowM93EoYIYFOGWg1TOpkz8/YdXvBFa8jbhlv1H
DS9m1JYtME44SpLmFZDnat9tuUD5RdbFoVj0B5iBh+XFmb2gs+9CjNJqdXyqdc3o6IH41F63coay
cedeusG0BR6OjSS7+WpjdcpFKlTDfw1LEXXWzTQxB9YAAnizfPIKJCw9o70YYUEX6s011MVDzBPi
eMHePgW2fGjdmtwhMN0qJXqAeQr7JfUsqyuTF0elkep7OQk7svFDIkjW1pmk08IqhgMpggf0gZb8
ZIWvbk54lhQcX88i/W0wUxkATkSVlj+D08yFH2xYIx44DMeGJ7426KLjknNnlvNmJtWFItrDQ0eH
KnzN6XB7ChhnKtSLIEYwDTHEEGpx3o9ogelH+UvL0V5fKCpyG7D/uLDaH7R81mggoWDC/aL1GSos
sT0kO/eW8GZownUK/yi2Gpq/LttTeLSidShgTfIdMtTJfwObMEE4USUE4A7s2rutOQvPAQpTsTPy
9tHYkCff6i2Ye0TQOSWmcNjInAPBYBq0qtuiQbTeD0VfWiROyUy/0sHE7fm1kwaRy7DN5ohB5K6x
PTizQ/fDJIZt+e5QDcuVU6rvpNG9vwNv7l8yhXUwnFn7L0UGVRzGyqlf2s63LdCAhrnXitZ8B8xS
UsVSG72l+XWJnL8AWksBL1RiO3J1rWYzcXEkMtrPWptLeGvoflk89AGKwGFOcXNN+TkAbUiElzcY
x49QO0rcEHTfNVA5TDVc8HE8vB+eOtMZVxklK1A8/vCdYIPGVdAQ8jWhMige2qlFHsPkDIebO5cR
ZCWODvc4o0+ZjvKbSvvdtsk891VpPKMixRZx6NeGyteBZ6kBdftmdyff2Y8jLt1Q40DZN5Uaph68
RPqiCr1pML7+CPOxsHBj8C3dZ3oj5rA0Z+e2MR2Xibyme3KG0fsUiV2sbfz+j5uUaguU6IrQUAMM
4GwZSxCxfeM/90MjhCq+mdLcUSdouw74hfYYCizIFKEcjneEqM/KNXW5vCG5tOlft7l23Sgric9g
IDTqQDUWDcwFqZIl8v7nsJQRxwBLkXnLS6iT9efnKgbIaqeiA070uZCuGa+m6O4YMM3lSh6dZ2DG
yyR1DO6w+rcj8EZJYBO7YI1EkrG13hfhfhwoVKeuacjyNfXh+jS3KxSYENMm1O+Pu4/WPEFKSpHJ
8NkxxSaVgPlAOi+inzLVJMXLqNx2qFOun50ytZVmUMfTsPB2CrJ4c+iMIx6Ewu8+tLJYxiirabYX
MZBTrBMYqEMll0CedKkPXoXsqKPaqnBu/LCmyGFHHOV720RgY/0AQzhZZjcGA0RZnSyUBjr/sbfN
jAr1fPATgr4mU+74addnJRSXlyfs157ka7CNYaRA267hdnSh/zPr0tRS/5p1ZxKGdrcb2oJPDT+6
TGudqcauZdb++AJUNJWhrUssXWb5aCiOABVfpXNvPAmkd3H0JVY1R97DunH728wnZbZUi3nV5gyf
+KMoNEBBJkfRj8qitPCunJIGG0z6bMFnTC7sKEozZxkFgWKQm1tGa0ZrODobGUuOe9NrFpgr3sED
Kz39KdKm6K+KwdT6Cuqdn68RNuG7XKznHk8wglr4iTzxuyJGxD3EhUMQKM98gep0FjxkgjrcrCI4
xjVPXXGlIWDEnnrrTgoLxSVg4uyRW51e3JXJ57a6RPHr6LnBsLbybUi511SKJv0KSYLPrRKKH7Rh
H6dyuuorVGhSjU8h5NS5VF71MPX9PDbGnH5J/yhw/7xHpnwf+0d2s3RmRCwZ67ndMe8/KWQEQhDO
HeBSnz0QxSVV7q1924xh3cCJUARt3VNgMDcx9ouf6j1OqSdrCk9JAjJ5hFeUKnOw61pU/jR+TmtG
OVL1W86VmCUTxB8kUjIj7SgERhFn12aL3xe1s+BvmgIJ6UhsZWV6vEDNsJiqZlvgKWingu/CowHj
UxE7ASWLkewElUcvEMQpPSVgFnUS9+xWYWyuoR7KE5Oxy1iVYDv+uLQSi+32wOHXWn6Tx5wCTNHp
EFRADoJZ/iFuqBKvMJLM3WR0zsQ3AI+Uk7Vopu4LvDzY4nuzkREbkoXqIUZQDjtFy07XpsuxUGCH
okSs+7J5cRJSNUSMMIYs2GVDx4em67TQ5d79dzeA+W1CjLuvvkW+24owwcND7Uv3tHz6xVfkxakl
bwsoQmPNmAZnWodbIYTff4ltkcXaYTE5tVohrjU/DiJ9vPQDDwR+IK1wQDCjtaAiGc4ii8bInNkr
YbnNqRExDJowRd0pk5jY7NLSvCzNWsuCiV8gXA/8UFtnA/arcw+73WTQJ6zClhMMVR/zt6Ay3x/r
ZJWGS4UutiqEEubHURWAYMZLip3i3cXPuBP9e/EK8cYzEWXvvU7B/rarUZwjB/zCyllIDU18kLXC
+gK4SQug4dh6jxIhuBM8wbXDF2w1W6z+kML8nUmXB1MSMpe47f7BdVdssuJFaqF3k2ycpM3EWN17
dPuwAZK/BACFkiK84t5L6QHneLRcas3Rxvc1YVXgH6VRxFvtwXs5QBlCTaHPrLtuvTSzWwFsFYVh
AxDCP6RAg4/+Go8iRpCl+O9UN6dbDKs0ZhcNOuokMnwXw+bwyyyvmQzb9A9EOPQbSYtVtXPuBZJF
WeUTn04ZxRNPivpMr4JIZWgsdGLiSlJJEVIKUni4UEiJEApXmTRw1zI4/pqZiqV7aKXb+yVK7qQl
DBl9IRN2j6DBBq5m918PvzQQDSGWumqg6RDvH7EL+OZNWVBuyTiHXMJwygvSvZaK3L8Ch9H/qrwA
1+rB7m/GN60E53WbdASB1nFu30ss2Hjgzgv6dHeaDUJCQzLW0u3R+1SKhsupK4T4WeQhJcmKFhL+
04cKD+7dpUiKlmrCQFpUpvuTXmrNgJlb7y0BrfxI9xcLCvbDXwfnpucCsleWWGIqp+Z0dXZ8FnHd
FayAwAF2LLwkeQQQvqlrwOHPepDn1tJQ10S/jLgGrxqxyuVmgQ3LBy8ldfxR1xXLNPpqfxGqm9ZT
+OceNUyfoqeu+xzS6RazpBU6RvX2Fq9tGwJ1JOkfQhFTjS7402aQoB2tCbWV/r0bAUoZhY7nVAX0
cMdyf6cfuuZ8ec06IyoIna0s0uIRkgdE1hGrxxqNgUjF5DFULUr8dh9+NgyFvjrzEaXralRDyShP
pZgwX9mxyiFvKL89SV0+KBH+p9smbYYvbhn4Bjl8SZGg7Az4Wr0xkX6xltbJjvOB+C4LpkchEKxs
lztJLXMLkJ0DpSmGEy6iDFZu9LBW8mkpXIWq/B2O/hlAcgmmOBZPgn4UPxGEmmBB3mdLehhYGXer
sUwO7yBHVPlqhruyHg/i7qkkhMMo7E9fSlTj9Fei0RtUD7bGN9ITundiPoEJOnFkSUSByc+xIBch
69lihdwyDXf30+Mj3Q07qNdLhOveC6FXZxCBtF7vpydoHCEsDi7ut1Nr7Vm/ukrRXYaoZr7DIDpl
KdpfV05DQBvGKDeCYy/kwyxxoSRkD00bbUv83HJteV4uc8I7TluvsIaNw4wZrAXQMvxBeIDgSkOH
tyPtQiSFKCUW5l1EmvRWk7gdbk1YjwPoKnvQRFV5avbBB41iemVX5Y4Qee+q5T1tRT2rA8nbqFH0
hWIU7fjWOt/6qhRkx/jpiyY1Rg5AclH4OMkGmoItFtQe4mfgf8K7Xtn80YYbb98FhSGBAKRs9b9k
EjxM/QWmzS0d+OTmaEZ/ghC/EJEJcz/zpHKNGjRYs/+fEutjhU9ScnwH8QWcMYAreW6jmm55aP0r
oeG0UYkeaWT2axfl7fbLcuPbABLqDQZrTecavcG0WvazNKU7jHOHOVNkfaTgCvqpCzaQ0hSCUasY
pXFsa692fLmOQJbOy0Xr+GHoZYP9p6kZfmCqeXgeWestt3JqKWGAzmv9+EejTm4HZWa4eEEh8H0C
McXB/7xOTbIeD8IbJSaTDRS3+YnA+YMSdntSa/3WtseHrRTASS3MpYsCocf/PoyKpFTGG8DdikrS
uLThuFPcDtU49tahp0M8eBcnQuZEkDTS7uohlMzKebqGXQjHiyZ3Eh3KNCoAIJLRJ5oMcDFcdM+w
Ex5UsU2+K1raPZfPjwsvr/gp+C76KctRo4vfcSWdkGZRve9culo97DifabzkDy9bo0micDgBfhjZ
YunH0ENH+oJ9oWDuovQDg3LKcAHdPrhVx4Ap8LzxYKZRw0sCPcHChKK0u/utozQ4q9li4vX1uOSo
S/sh6n0WPiktUhGlVwmciPPKbIX1IYj50VcqeTxXXoyubDH76JSrWAFOQIFmWnXt10lv3fWh9K1p
tCB3fTqaftu78fvVJTKpv9oBsBIb0qOpks5ZVLL51zHWB/DpydIcCR7O2WTr+qGmedOGgByxsoY5
nvQkPFBPOi3hDF/F7pUNZYdUHp70pCq7U+qz9jXV0X8aIsDwo4invNQIN+Y6v6rqoEbzDiKiNKaN
jr3mcb7p6y4GbpnL8N//8bkJZL3VPR/lO30n3HcBdnvQ3Q431AhJIRlbEa+fe7iUvHs8WgkuW8dQ
1hwLO8PrMaxhsAIxbShemOYP+aCTiDfer2md2J4WlikSbIybDs22+f3El3XlKYZHtAsaUSvMqHlQ
VNIsJKXRkfh6n1RQUae1fq1P9OdI4uIAe7l14JXeSdz9D3bqRmfWZmL1Leqwcgr3bZOb8d8PAY0B
PjsokWbnZSEqGG2KiZadverey7LE+u51dpE0x/GJhslNi227TC4s6ps4ZE/787UMb2xa8ZtFlYxI
YelYIEh0qpCXq5CVKBTn20Vpm/HZOGjKACRTtXCmSALD3VkSMZNo6QGGH7GgRLzc4TtAhI+4YOY7
7Y+Y/InHNDYgtrj7ZwEvGCCdAKNiQTqqwG+RDL3r+8jK+8Krwd4wm+duzFwdBMjtaP+iuPd9zTfY
Bp74OGxPklnNAbYbLu0QYmcSQJU/qbLSVpuRxzj92q26i6KNguC25Mv7yN/u1aas/COYfNK8dqnh
mIpnHdw6lLQiDnR3tfhXRk4p9CqPIZ5om3nBz25rUlmcK0ZBLAH6Uv9cWNLAWvWxagmN/S0/oLwV
ZirhbkH2wnXIdFJdIbJlh9ByKPeeRhvm/NlLyYqtTlYbjzAsck2qXjqMbk+WlFibwMy8vvywIDBt
B/UHhdPAB+1hGXgytgmeZJ0L16ZoJHx/HyWQNabCMQy2/9G5UjgAqpR9/vkQLTxhzhJRMuQdJcgj
KQ72e6GSNL4gmJ1J2WhgwVd7ulaCIC5Jf5dv/7SKXZ5eJmEyi6Dl0SkC729My6w+v696pP1lEA39
/1/s9yWbi4/BpBgutR2mYOFE0VkLdpXVB+hTvzs6rq9YzlRXKjTkV39KzjDy/1YeEwbMTBYoKa28
8lFkUbEazLy1AckhR4Rb+qhWU/3FcYUu12Oor43caZd1cMEIokhqbHb67yUBpnyq26Qjrj1DDzUR
OmBPgpcoopvHbwu+c3pUqK0l/meoC9jLkYGZXnImkfa0drxj/PYh6cxSs3mUbAZR+4qxEeO5/mVw
sjiULRNkoq4ZYT8xEemxmbZZ4aEsCWoCfKN6UOyJtg9lfti7duktK0/sZ5tiDx60o1Yl0lyMKEl+
BidMv/GjmuDrPUXI8Dt77QZPgAhWn+bdhREd9zX59rHiucmVVab5H5E2IGd6N/J5xOnq4phg0OlQ
O3wxeggMzEwKQnR0igTRF/VX1bY0GOmaM5Rub4c1+z+Et/HUAxwk1nloF+fYLQyPfCRIHeyBd9Zq
OIiu7accIKFc/INO19oDr1mmnaFNtDndLRfEkge6VasTkwqN0aqcZGxYdfoUOB7TzVJjqYF15Iwf
oaZYlXYoZ+sd7pS4rOvrCwz9nB+Psq7lqhfIOff3Vxxwz8fjC+65zjLJKIdGpp41A0zn1qvHoueH
b6pbK/oN0CbVLPO2FMeVcpHxeB5rua5xCC0sayNneE2bYgkhXat7RoJLZz+7VNKMbdV28CJh707P
meZboF2o40ZBTDgutwUOVVGd+HU6Ab6ZpYeMU5tgn/fYI+GgvdbSOtzscqGoIZQI12CBix62vpn/
kv3nt65FKRvlCg9p1FbqYoA2N8dDLiZ4iKvII5L77XGBEBwQs0kqKRojotLiNui64OHymaBMtUn4
S17eGBUgEls8SnIJ70A+l/+l4KdU12swE11EXp6JGjBicIuGIUgr8viQk95aMaPzRF8WqENVMvLx
c/mORokOkag9PSC1UAkO+JzocxeNquLkEmiESEc58KXEEWmPL72wq5PF6zQZHmlOIdvOBCI48oTC
1mWLRtqovD1pJLTuzvtfDF5v15gbPUHD6OEOs92EBo9I1HIS48ZSJnxoEQLu0l/Y7ogp/nCZ7hDb
d5/UXD4ymdnX+qo8FLCnRpritf1TI2OP+0td2yKqS6eoP/iqmg5OK1MpzSkAgCSQGLjUgBDRKtIG
Y1KDDutBTOQMeTrty+PMZlyMXemr34OR2qiXd7WIbw5sIQO7BE7Kl35bZRYuC4YwD1JIfEi8A7Rq
PlmwRMznfR46qevGJ2qmI4COTSd+m8Mr0uo2XwsLiY4DplSFiy5hyivjg1X/RMTXhxC1w0J7IbKE
eosHviaMXu631XgJc4ii23sVFTKHzMFz6+VjK3fRxA7mqbRoPy/2i7jes7S2x4DY/O3rURIdqM9v
o2cA3gKGRmjdpdjemxnyjzQLvJtDE3aZqhc3SZL1wkdZ7jCMBRtuHqaF3W/3eXQ3Eb81kHCKq7nT
Q48manHkH9M0kCWYVim220h76F3NQOOiED3DbWWJfbT5qP1TZ4EH6NF9bhqd49biv1Em5T6z1ouJ
B1n42JMYk9EplSRTc4orFHtoLyqIweOipL5zWQPNCde+s+7Z+HyjeikirwEgpkfaCoxDGYXz9CaW
1lihElYL6Yjj7MDfSeztgG+XwSGs2W+7l5dWYoLaMJfou/fMJ7MNvHt1fS3KUkcYVajBwUiS2di2
VOm18z9ZgEVC7Sg8q03mci2TBUtc8pNoI9+swcHB1iYD5PBfW4c4MRFGKIgKscqv3JAyKdLDIjry
2B99BlmGq+tmJgw9u1GtZo15sDN03a/eW4znDxYka9j4f6MCsVW/G8su5gEGG+Ox8yNfsoCuKXxN
Q/KYT/jmCQ1o1+qkJLcbzptYarwlribU2QF7GoYedeuP44OjdJaVcILKE8/tQm0Q5DxeOPDZ9yzp
lpDvKyYz7r1cuagg7KY/ytrzrVrzsDh/i0nhvIJhU0gmUGz7DKWjoyl0pECOz9afLPTnyGusW0UJ
JIKqbwez1UJMz/6xGunLvSk4mmv0k32PWuj8d4SxQm9h7iH8g7Fa+WukYhs9T3C7ub59LIFl+uTg
xxWYoXVUvnQto88G2vgGR/j9t65OiuOrVQuRanef4m2tRb3l9iAEG2fNz5H16h9AYMb5WDASysEY
tuLUO+MwYQMHMPDdGdWepW3P5Sr4MwLtZkKlXY0Pza1ZoTH/iwa6Y5S1uVvYKNJyegvougC0OyIE
FtBG+U+yQy/cn+9hA1h6ESGv+TkVY5NTakEHjijz5MEdvGDmFYf1diy2+VzdO3Rz5C/MI0COysZ1
QEk+99JPJHtbyt2+ijKf744WQT09Xb3Vzxv4TnfeTl4AsqkQeV+1Slmdr2W3KiDMJptn44YIpxiS
s9grck3GwonEsb+LZ3GFYjfQarldss2HNuwluoE/qIiA3aYnTfU4+LCsjqtP7ybjZN2s82s2+P0/
GywRp7jAESh766yhPX2MM/WebGhjUHLKSwg3cbwLOg5X097nflVPGrttwpsVTxnopswaOwXrOM3i
A1vwx4Kp0TEyCTnN+otfiTK+IL9/Ux98Y1fBT0n5fOr9kgBhO9j3i8oA3wp1QedtouTBiZaVQVD/
e7oRpVB8Hu1+edRqyYs/LrDn6PKul0peY0Mfc68sTv6AQztnO/+S7crWT/MwY/AmzrfdIyh9Kulv
MLAbopgzFiW3qDUyCHxLaGrckYTmY6NiWr/7+rgi+84H+ED7Y1RgceVjrKzz2X6Q3uYdxoBErgOt
kpIvvVltfQqd3aLKbbzXs75e5H344S+2wGzNeNQiW/Oj0BSBMH5LgKOxsL337v2sxpfpfUgArUgd
McHOAlBdJB3YrbyTaAkXBfTMTxtRO7OSBiHjomaqqzC2+dKKa22W2uNNXI0WMLd1XNIkmBdxhG3g
qTc8b6MpcLBS2deHorpLDCVuTCci6Szz0/p1tFwFsTURQAQAV29Gyrq63XI0oPAR2M8Qm/TuVjvb
/FfinOzDOxwNb1uTkuRTjaL3jIkiBFy3DwH9s2piaeyCsy+oN87LcyiQj1IDfJFD/HaoBqhFOkTz
m8N02Wg9STy1aD17hSBlWRQkb0yNeQV9Dg93bl39e57/UORhE3C4ijlBkcEXJUKSpDQ6JKMGv5dT
BLZ1eqzMbOKdWUuTAZFNGkO9iSSTcJgE6XX0noYs9jNBHzuCRoEhIZzV8Jssr7M5LJTEpbn7t0OU
3XEZSexw9QZyoW1PiBBjDBMoGmTlqik/rqUd7G+KhLIKo+a3TkD2BiQA+eJmxfiF1s2BejdE5Xyv
k0kKpx2hFoNuBJPlgotSZ3ShexMZEOZ5WfUcZ7WG5FOX+NhPtJ2Tg+9ACn5XxlvGENyBUm7FWVu2
qI+WauH/fU3qV7CfCINgPJ4r6oZkr3VZk+Ju2W5hk1y91n0Qvu0J3Y3awLpHTPBgB/XxZJKx5xil
SQGwqEFQGaaZziNrN4LYrMCd0csrKmYs7Cjy2sd7I6twGCDt7lt9BF8DzVRYIkhDxgu4f7QLE32A
lyHo4vZoRTGIx0gpFOcr91Wn8EBng1RofT73YkntbLEnk/4z/nLNLYE/FZ22ZvGNLk7xfGC/r8Hi
iN7SDdj89gvakvRzma7I4amlrSe+r39m97HBCOjiVoS/KmpQLesUMF5rHSUyRtpPfwRE2o4jkWzZ
y5i7mTvrELy0s7dmm+HaCcKfBfO8k1Y9CX9Hd4m3S/t2Bjou1eDa7z0sagSUHOzS5RTJeRNW+4xW
33kvHfX/YmkTHkToQoChBNFdSZ7Lpn/fatPPtuJ9UYnkHdk9v01GM9uSV+jwoeeAIHJeuvcnSopY
cIMOj0gd/6wcYZw1H9ZpXdp1h+Vvls2vJdjy1O64xbsRaz9oS5elYnvF1a95p7r/bES1a+6D8ps1
XoNkD8cyHo3EbwoDFH8jOHgdY4Pbqb4OgUVVaCMiaZIRsofzWIxe1MC/P8fkbz+SinfJijItiOxz
PL2wJU8qRjMvTIG8C4FaadSQWIw+olCjkV1UjUufQcIevnR61vkv/7ISjltGZ2vV9PEVVbKkmWg9
+lEelntl2lyX/Hb7OMH608UTvvqUbtaJrV5jZeQaSlk2kvUpy674Wb670lJCnjCq3ZKVqXMZIy5V
UEGIX14UdNrUDzvbZloOXOTBLZiTJrXXqVV7NOSW0b5/W6kUvR0dnuIk145MdvxfnoqHWa1BlpKv
lcW/Bkvfq1c/SCkesGdi/Qk46eEnyPDFcl9Y7N1tbwTkxAR1AdgOX+t9LsjjaN3aRePYniJH32qY
XTWIPvB4UdWsMKYPz/PCuysXeAAwa6/2cLvqYiPKKsOH0WWFi+JVgIHgnQ5LAW5isuPohYvrH5It
T2DGsO+Gm6BAU4bW7PGLUbUolrpr6iJ0NHRyzS4ve4TCoVnr79z/LvxkYpimjHRgFExdsPo4z3Aa
sk8O0cVlbuLvyJs8LHJJ4AJGr4xnG74buvMb71rpRTP0murGANoCFV5uY0PBaleCeT3VAq4kD7W4
MRlHvD3pZgc3EsonhFjNqZ2mBqG+IznYZ7C527QRttbsM7vFB3kPvXZSqQpsrnTslToPwSeVRRwv
WOVN7utaa0QTqwlI7RdJxUpF2zfKXgtpCrTVyP9f7oHT0O0qZ/4+WTp0JTmY9HoUMruEWXo/AgsQ
uf91ynefTQChKTsBEwGfE9QxB44R8xvBbZs8QCDvahvwvlkjKEGfTrelz6RFPJtyJ5llrDc7qnao
x2Ua7l5w0yavLr41GmBaHCspor6iWcu0kM7v3xDtgvHY4FoIimqtTcZfRh0e1jM3GHUBOVAaafg4
HtDsZgWgcQULeQXdrJxgh8Ahmls3lrfFGTTiElyYZsoSZrajS8XvlKpHLW6qiWwB9i3jywNleIhG
286fetmjlqiuVHNXmyNGNxVEzwrHxzGRiridP7uas8aeAsYe8VEHNElIhyi30RfyX565bP6UV2Dx
zlHZUS5MtTbXC/Dgiy6spbDpP4Y99aJZhc7ZqQy3KzYMMgEoqIlVjMFgu4iYecZ5fIALYQkzwS5x
KMGOD1r07H4yrur3DGE8ON55przGyjRjAXwgJ12yhd0dDwcAUuTP7cgB+nBRMArcTRmHuDVMYC2B
fx4HqCrVIkNpIieUI4d5/fl+dcZE+7INCFR/7rGe2N/94BsHNIJ5ps5ELYFWSUjTRG1EjAHT4wl4
WQspv4Fvq65HaKA1RQRHnRcH3dZpRzAT7vzwMFfY12x1CTXTCgh1NzT7smgD30ojET87t7eLm7/l
H+ih3bg1i37ghdPMib88F+XdiB2ywDMDgmUyPAZICjKrlG9Z1C3gAcUDnlk2KGacHt4+G6fvXwYA
VGIOaqgYx1+5rchP0dRc+jJ86NYZVDBAz39r/So1f7pVhMlLVJUVjBhFsquWBwsGlPosZAN1qpRa
9r4TjMhqd8rOxErUaxCUoTITLb/nNXWeO0iX36sYT/lnxtWIs+UxWkYztS1ZpT4q3afNct/Bat/H
5Zi44v9oTGZ9uU4DgE3MdShgTpq/9WBkvaY5hBw5Rxegknjq1bvCZYCm1biFqJ8rZWGP204KVWLD
fM6MkNNyAmjuBm6+RveL0VVELMMmTFqQeCz/w1fgwi2fJvF/41A79ysA4bB+DWgdfYR8mhUFteVu
FOswJ6hQbHKLnU6SP0foxUgCISVIO7nk7FUA9eCNY2J6aS7Z3o8hJgzlMD4nbsxwaNsfZ2+0qAvz
2WF5SK5U4N6hiazAqsNLn1vrUN0pNCr7aAOv94VofPLsN6MBaOGHAdyL6ccg1xBtrtLsEtDEFpFp
QOxLc0f2OASx8JjJeIFhzYgUCXw8w3urUzAonbqrTrPrnhByKsRUHAlmE1aZApY+5B/Zr/LoQShd
+aoOGwWB5Jh/iNFVaWhLK/mkk4jK/y6Bn4s4wqwlkJAlKL4u9J17ZfCNKHF37P9izgD9KKaX7LL0
oFqq0aPAIT1JAZ85PTSnMi4rg1zV1n+5mJlpNNZCZ9JaZNrsaV4Jim2Rt0ctshDrDpC60QBG1fbB
FgczttU2HhKLhWGUgiD/XR9Akp5eQCXxPA2hCENNLEsKG/Wyn6z11f+o4/Aeo9Yk2pfQ8O+B7ezv
QHF55+QQLylTsqEm+xfZZzlpYYOq6/fIH8l/AUc8qsRb6Qe0zKj7XBq5MhviIupx+v8jamhY03H/
eSIYS/wzz0DPKd2IXx0ELqzEwyir9VQaVqwuPfLYLgrB11etO0bb6EZdSwmag153Dr0LWwa9Lr/J
VVvTkGvuyMdHCaUL6mD4pWfefXabluapYkT/UZd+Onvtgwjw8pMveLkSDBVKmBgbr+gRwxc4OwV5
OwMWqoUXVTtcxHJLmI1UqVxr+aZiTp8EqjRJw05sq3HoFV9uhN9NXMgtsQJKU6se99YxkoexLEas
s9hTw5VRDCU5ThxDMRAf58hEEOb/AUADPTc8iqNbHDa8nDSKXvjvlfKZu9lTog4z1H73Hd3Y98W9
n4PeSBILBrg9JSxXyocdcPn8O+pcGmfc4dXY64Dwhp9cX3gF5fsq9vFbY2PE4ppRKfclPmXYFFIZ
bg5R01K73NMEJzf9c5KWwNcsjb2xPxXPW/c+dIaPkC2hdBUL7JtqBFJolttD5myEjpjQtIhiY80g
V1S18B6vonIeGZfkErgkWSuJBIHK59rIJ+GmT/0oZL8h9n8xnfwC19ZOuHLCan0wQvcjHxqlsDov
kIk9ct88LBnFKfCO54GUSLxvp0Ojg6Jf7ZABz0t0hynevijeaLylp9pjSu471DR08ht5BHoC3Doo
MSmDBtfOfEKyn4cwJSG0GYePmlxxkoV2tKD74LjS5PVFSAxQIfSV4j+ZIJIvM6jpjv1Lxzgq9MER
Er+sv04GpkMRvCuBdx8LiZLjTKhCW+pb1CnwOVGFGH6m6zkOTb1arCzCVpm48cdQKd/+e4wwp0cp
baEwzDBCRGH859+YEMPkq2hjLHLivNP55Tph2nYa8cZGMtG80yXBJWjl+PlYqUFEMuUh40yUERYy
TcqvXO/tR+qqPHNvr1SC4uFkALo5fdqEacEKhg10/Z9uJY5j5Vk5+EGAxDT7w9KVy4uJNOMOGG7I
rQANIVes1g0bBbg3Px8dmstBOuZy+DNfzAKn/0xiYy9qiiLWUjrvVPGlDWejFTvFp5NAVm452pwI
41QZZtLN6LJZtZfTVXe2MqQA0xD+0ucOJ9PhB558Nd7fUrPxhfLIZFUlDQ/zlindv8PzkTaOgGQU
kj3+YhjU822EBMeDQeZ02VZn7mjaCyIYkxbFb97tStHE/+EKYRPG6kLT0iJ5GrzbP5gj3K4FFfOq
AaZSqMnkMNnfXLJezkh9BfxEEwQ6YHgQl9jIiLDddrS+rwesXfOdBKGXjwvTXMDsb9LeQiiAyzTD
hCp3DCwtfJwuX/nx2lnrEw72uhmvGCST8AFEYTMUsa9QBY0E1ryZ9CedSGhl1nPJ1g8GhGyzfajS
EEM43Vxjane2DPFrClX/nc07Ap+RioS92RYR4hVILWaHwrJVYowdSqzm/N/GRy0AgsZa+uDImpM7
HwmErRILup2R2Pqm7RYRyoxUeRCxhhszwQCox1gW/B/K22r+JwCOcI6YIt9URdjwZ0YL4keo4Ef9
7wQ/RJB42zJrjza/7aLtdsAB9W/Cpsgb8SUw1De5Du23M+Xso6iqe/oNq+e21ZZuOLi3cxLAjpZ+
HoQF/y+3RAf7TnL5qkCUJUBd6Kohxe4qxnLpQfm2bux/fduFA7YxpOO+lKlop09vlhN7NbJ1EwWO
71IDshEC22tiBXf3L2Ak64THEXL80HM4ZfrX2udp+FfvEocPH0NiaRuD+trdMAoYuUxTml5fBOYj
6jcxvnHHp5wJgGOM3ZFktW4vE5xEbYNucu2ENfhkz0DZdrqv/9W1p/iDx5ZwYXav6d0C1UN3/oJX
IMZmeZrUoqyTRU5B3QewONIC8QK27GsbJv1A6Lcxkf7CapQKGd+kfucW627jwnGm8W64r9lMADVw
yY8vvlOneuh+4RHYcr/2jRsEpcYCJHw9HjQjlmXS22GOQ9qYzuU4P16WfJoAOVBnJ1Eb5DG4Fft+
wm+b2DP+jbF3vXNSXLdqh2YcxqsJuZ/8ogbrHd2LkpwCMoQDYeJw/kBxSPIx5pdkJH9iXs11nCb4
GgOzfI6b4Zq3AKvtYtL4czWYD0ouEOFTrUjxPv8mNWP0kLvRxDwNk/z7TTe+JL6q30WptAzWhR+f
zz36Ww0qcnijBaXTspP/aQrnW7ZR6bA3aWGzM1UkEgEZ1cvC/lahOQ8lanagkeWvl9KcMJ9tA84X
/FNZDyy7Nz0Fco/kez0ADluetBXZeFJe3FktadpByOExkecPqvYaiJi/ivPPJWHrxWiOaxQr/kM8
YO2t/+eOYiMxzIybwwHEzPZgyA8IaZmT1JmaEy3AHKn4JUaajFGCSnmG/945kW9H/2bDXXBTjLaL
ypzGTqDYgr3ctoB37ln7BJp+KBpkhKimRRjv8CgMCFgW8YJoeHX3aD88RkF+qPJaz9TSRQCn2nEs
OEEbFP8FhFBJa34EjUMv07n/oEuIkksPfQdNstzRkLzvqswk6dR+ukMwFeMK/AhbqKq3zqGPHCNg
21oZgAMatRJiiI/dDEVLpqHUZrElALqW59ir0mgpoKk6giG0Spq0A3yxN4uXH4uxQpvesN/0Zq3H
JPqVNRiCnFKjtcGjcmzY6ayyDkGpoJno4g1IW+ScsH58ncqse+8dS60Urvtijyzx1d7oKu9BNuwb
nq2GHyfQw/sWcJYb1cmP4wGMp9Pr4XI/UdKcBgmAlg+O5xf3oakVfOgKbFzzvBf6n/j1faQ+4eRB
d7LA+eAW9VmUxt1RMdSTvOaH7XKA6Wa7uVRBOtD4EtOeO59CcvAdjlPjtQB4fsJT8eAzEIdD4knV
j0CB4XBLZgdlEaXS60m4uZmpXsRuOGio5d22xkvBKgAr3FWE3frMyoDqpE9hQi6avvgXEfjplXVt
nDaoSomfgQuQ/PECdf9inejRlg0md8RZsWVJt70HRgdDwoVjqfSyiY6wX8CuDPogWcGQLZICKQ9k
bxnuHcCM8loqQ4tS9RKD35tG0CP4YTd+u7gRuepZHXYIbBwemRGzf7awaeLu+owfvD+mdOHFW2e/
WCkzRjedB4F7J2s+7zNTDUoteauepJfmrF1HoAZKshKgpt/3LUMqvVLOMuyY2GsqD/CIguejA1ND
ZoJTleSiFvFEfpGh+ahQgRZnsFJXv27sbd7IWl0Eu3npmtV60PwWfVC1ZZLjPpSe7XnBj1zWKAyw
krGIwsbrX7j3kTNGMlI919yFqDhP0cKKRD8BPo1hl7t6zAbiFAURb5V8rfbe4t39YCIeytK9MXwV
Ouf2zVQEl1iR04Ge9ZGTff6Wt8dA2wznVsCe0wLrEqQRy9aN4U2g6fMRfjBZbasBkrdRKuULbj5V
D+r8PecLp+Un5BOHQBs2akKLvY4mE1uwm2q/ys/fBAOWlEn/U8p8Dvmyx7n8rkMI10gNq0VI2pUd
5OLVmMuJIHAWEGliVdsXQeKuCfuIjJ2tFDaEBp39XdM1BdL1eH387lPmE9kzqNr/SgO/o6x0KhES
nQQzr9eNpRhRZCLwK0BmfG/BI5C05Hhl1Ok+vJu7+pMItO+JNLeKaHdZNk5fodQj+4Z4KrvYiXVq
AX0zI3NijbLNz1wIxk0cQ08YYWE/JyOk2o8Ta9zuA+LkBYtF/N7sC1V413xqIwnY81Bs4bsRBPP1
kwBZ7aJBTv5/UcL6DXGYlDPzvUdWYjVyczquw06nTEY2ifNwekFXSJf9OxgeuxSeZYH240j4dQc6
qwvwQ0m5J/Yoj1aOKRKCEFDRYywedXuvc+SPtHAAZq19fkcgZU0fE+D38a4Py+n5+GMSYpFA9HlZ
+/bmzK9bOMoVgF3Vx9SruZWgqLgF2hPWpunZ17Q/b7Is2HtJSvKHOuzlaStdvcDmiFigLRZ6ob5n
u1w7ometAQBb+WEMSOlATwrqgEQLZJxzX1Q0aZfR4d+8mCRuBJHN0qFoiZ1z8WcczU3rxzlqR2Jp
oC6QuvUQRNMxBcsMm7cwaHDLZe3TpZH1TnADh1O57h9mzdzmmFHbuYi8jNV+7UvtizeIQwo62dnQ
IBEy3WiCC/RWbHr4t0lHD9qYixo4LT8+0kiV413Y/GJiDA2zD5TVbGhxLq+lH7LG/NTD8HBsHzwk
3WRj7CuluA6tv+6L1zKzCQdoIrFNSCW+NHaInNodGkTuyEiqYlnRqN6B8t0Az0X4SP1UMW+4ugc7
XusMFPWjbciPSXiGpvCIckWeGWGoG0w6/pss83A6atIq0fQq2NZvEBW5+bJJkJVkRdw3NIa2cOPu
xz64Zzu15EZBEwOuh5jsOupVDkduwubCohmAfRVnnarTdcpm9AX01j7C74jAZruFve5muWJXF/Zf
VLHbMMp9R4SZB9gVJPyZIXDGWGIUOyrZ4NV3XT9dpp3VU0FZC0R+dOTfsiHGpGMNuGSlYVXl7kIY
XcMHEIY3l1bNjuKaOGDrr9frCjeuVFYmOS78AMuZ77+ppMvdN05MKYxEXJmdtBqYHn6zoaBh9Mrj
yy6mx1vvzP8vUcgdiuUaKrFxcK/vIP1ow8NK1kcozhkYxqQLhsN0Pwb9VxjORxKER3WP2uKEbqCl
wwdb9SJpKUY5TCjvj+eeXed8RjXLMvk6oRCpRLasILBbR6KNdO2uNqA2Js7BrOLCvS1EOjfNyXNw
BCjiZ54J4XruT/EZfhvF3hnoW0ZldjBGijEWlKybwFzctQ7q+SpOtidneJdJwi1hm4hKIP3KdOuy
qgQAmjXn2EGlBCJgyZ7QzwCt6Eespcz1vTOCc7K0tN9qTHxjTcgf4IUh8CEi6PqMrLMfDOoFOjPR
0K+KN4TZxDH8uj75wG8Tl1DhYqPuNI0wDatA5twiYA6AAaKf2TKvHUSUHBvBOJ1/CqWnAMbYyb8H
AQWxj168yzzEd+MjdFmbVBjb1tNhAn5BjhykcYLdxtRLAh1Zvm+7N9nw58dU7zB+1sP6GESDJT6W
u8oLq6xMyB7K5X1mnHqFBKubFNQAC+ePcU9Ki0MY65R8uy5ceoYangQC1CDVa79wj00GCzPhKe0P
a2GMzOd+SPp/OOqfxmBcx4t8B7+teliJf3hxQ4ijuLHye63jME04iS7LbX+mlt/qGQDZay/w89SP
Ic3gGVr/iTO1XU/sPF+TVBktHOzL4Tvq02AANw38bzztcu+hQZbi0sU3R7nUQ/FZbdwjZIxuENWt
Um2aH3f6MtCcPkB0gpRxF8P27Dp4ikq0QX2KfchsOROnGYBj0KSzs2D1uxwVLFg/c5Q4kuIrm0oc
86SVRRptZMg96ONlkACPLivz4WSXztbVC76/qsgtudYHXjpmWphB7GX3196eWP6dMJx6z/21WPGM
rDfIhewod7+zurVheLQdPSJM/Ll1MdewWLVZHqUHWq5Ce1ZRAPz/c+vHxzo7hItOimGb/E74o4nq
q4hfNoUSE0iB/27QQYoUM8uYmbQI1DOMEtWsoQFxs5SpxxyCbq9Ri33hvW4IYrSvJ8znseRxTbgr
W04xQguvOX36EwmnUCne/hIudTjfaVk871VnAerxgokT/UapLWIoQ2GMOyKzGlutJbN2aezSHQMb
TfKZgpzaRjnABq1/7QEjpdImMuGkP0F6hMnU/fOxqrTINoupeDvW1yDZ+x1EXiNqNuMkyNMaGU3g
Z4KyS/C5mweefeOKfKiTRknvqcZ1+TeW9BhdiuDMtedTmK8ZPkfFMmz+RShf8oSNo7zIKD7ZEh9t
igkFObqkBFIwJQtupfD91KLzbQg1RdPMLMOYROKNekZaJf9jWwH3HOnd3uCkfZj0ZOXTmljP1Xgl
uExNtKQm4jj2K4kij+dnYQrDGo92k1P3VewqRMU1TmHwhu8uf85IlKoqEAq5J8kNr2zKonn9ITC4
yoFMnOWTuBKrLKbbqco7/f1XuMiAEkbg9i2dAEREsyQlT+EgGNvQ2USZ7hyUAOoWMjjond9z/mo7
ihy73L/vAYhgF+ni28fdzq49rkeH7mg4p5a7xt1Eg/edRXaBxrdRtxzT3G/wExRDakCkVF/6mYFn
o4vDLM4ly/woo9zpVvN72xLTz1G2YY8RlNI4VkxUWl/BO8BAAn46G3uUo3wWd5IWrqCQEXPeypbN
j+XKjIlr4KYw7d+JiN6yF51f5npDJy4Rj1Ib5kHgrq+NX11FuTDD7W1zr5yeWR8yMNxSeLnjWaSP
ThdgJ8SlCoZYMt8XGG7iDvRMWcSMZF9UQT9UwTxe1B3MhcNdllb/KWKfHc33GhnjywewNSNBcuHy
zX4UXEBkjqwRrLK+Fg9pIw8qBDycPlwv8PC8KuEoC/k16i20xcEKRacJYA7d051lBnA+kHQR85BE
StSXWN5AakWuy6dzQ677htOu+xs/0ydzRFZl61hpp6YtXQZ0mKDgopXHfLN58mILch+U14/9Yyfg
AdT3IeRvqd0O0yBBhw1D+eA6fN2konSDCrph5W+SmmizcvgRnzB003UAP+Kyhlj6UFHKgu9NZNYX
a0hcti2TnJNTq4OHsqXJRktv5aewVVnJqEUR0QOmjPCeh3XoJkRDHAH97g0h/0flMD2ZnFvsqheJ
jh+2ERND4gM3QHbg+NvT4OvaoRXGbNkGxwUzGcvqX4f8ybJe1cNjX69GYi17fO6omaoeuktYZxJR
IsGVrFtROelVdfxaTIPPspI+1T7jqQjr5Fk7+YKm81LeMOXHMosB2uSlFx/ABqRb9Gr45/iKH9Kv
GNKaSftSbkveUEcaMJAJh+LNYk7RwFwmS2xMJNxp0vBC8vOLAYmY9nwmvKmvtgtZq9q0rGM1m4/c
oB1BYqiE2ks0srJcJkdnjU7ftP+OcFMka8dD4doLIgyiB3WGGsz+aHT9Enwhpam8nS3hFUc7ykqn
XffcvheT3QDbnYxP20wGWdBK8esjaBA72q/NBMv0JI7f3m0jsM+P5WKpFp5a5iRlDDMwdiRg6we3
+8uiVpWgZ+hilS876WbdUACWbN5sJouLLcqMk+sxc3urcvCVHsK41jEkk3aO0VJVggw7W717mhjr
2rHc951KSf0bPSt+q+sppBEOKu+CIqInUbEyQ5Y1HRI8XMMGYfe6BBkhvUU0RSLJasiyZc0ccYCK
ahMsMYD6tqEGh5HxtUp35Dc2ogtjwxJ9VCVEt6H/2AJHVkCB56nZKwUrRveGnNYHIeFVKSHC/SLR
1iAW5eU6OTTFaOzRtwE3D5/cFjstpV0kwIm6GR1Ra4tVRREjo2ORgF+p8szcXfrLGYiviS+u8Odn
Kt/z1B5yvqYVncJUyg0MZUMplHq6ow+Bes6IhcCSSuptLAFM0ONVxVoGiEjAHuAzsmBnz/DTzMge
xo9QYQmLaKJ5a4WaIfdUkqyJ9FnGmhPwPrhNbSpUbZ1pcVBLxKAUiCD1WP4MXgAPlrY7bqafjAxa
FCvF35rdbpCJahG9GjA9yVeQjvFyTzicC6Y9x/nzuRT84aTMir6Gwsmnv1RGib+nsZzI0M9Tq+tw
tfJccCBQQFbD0StFhcUkF592ZQi005UJ8FU4mRxXSr324WX+Wq5L0fKnjvghkCy79S7I3Cj1mj3c
G/he69yImss519G2dYcnimovvI51pHy1fSfhq/rg56AKyFa5FJwoHtVjcfVj1JSbRNFHWswePOfr
a+jwU8PJ8XgflHSPInBPJWkKOdm7MFjYmARj2mjcNO3/7MmeFiRiILfB2D0eLoSlUsXBKapXIPJQ
BhSAKfXjo8KTUQt5flBkYNkAhjegLTJjibkVfs4wcEAPv4hPODEyHrrgeB34G5sUtvQOt6m21/7Q
m5NvsULgr508PVCJhvxc6QgYeX2Qz5Q55q5FOl81+xPYiG1+ghD/k3u0s3cH3h1mpwAwIiyHwIkC
2SwxdxcJYZ8GdCdii6eSuWlUBiRc19ipOrhEvCPGiPwPh6fhj44t4qAGyP5GURbfH8srpOT7tP/T
gu4fNWiCp4Q8/upR7wEtnLI95Xh5oRF3qT17X/wEfpFLERKc74X7YBN9I4E2K5hk1QOzr/90m8A0
CQQD7gdH/sQ0pUR/VKfVZpRpMwnIikbQJ2Yet+GtyhZMnhnrtwarseKR5Vp0G2Del6AB6y/XYRMo
XAuQ8N5PFbWBT4pAjPeiTVhKZmdc5hJLCyz9cESgUKgWnWfTIQXVRGT4UeMZAod9pVXRTJ+uOE6k
syXYx+JJsPgD27C3pBXirEpYjiYzZxAw1rSysnZQTS1b8/mlpggjxmjH5xLI+3oEZt5X09L/p6Ah
DS6np6OmR368Ht/ZzhyTl9kvWFWONQgXqNy+n91pKsaR2C/0Tpn5GkBX9M9mNj14DdGZG3VGBAME
PG6DUf9ABTesHjcR0xzc5LZcM4Hsmy5L4JMAh/8scwqFY1qMEhc9CXd6CMOpXeqh8HuKiKGwZpCM
HUPZ+2qswVg88ig9CxecJNMWEmQBupcEiaDCYFMJOVc85s1rpAjQw8TLAtbia98LQWIPoL2QOAuJ
He9d4UilNuyT/bIuXOJ/gnDuQLLWiGOHZcOcLSrIMzyFC+fJwIAmaT45Tk3Io4SMnZDUb5lSMO46
EnfqT7NMdsw/8aZI6bi/Ru56d43dH9qZMkXp2aMhTn7W05JZLHTA0axA7ku+dVsQJtIuKQbJJ7jg
P+Z6lMrf+FoPppMG+sK9R33AEVijn+zjzmBoPYMhu9AcA8A4s1RHr9ud5JQoo4Nx8PhvoabzZ/wv
G51ovR7N5XIhmwncZl1XZBtctqlX9UIOBqXG57+TFa/4cFAwHR7lOqAFd+YbVRSByqVZ4u0bxD+w
aSXzhXt2YLL4NKDMj/CvD3qCk1oLhcdd1mNMgSz4VWkc80dMMP8bYAf3mhqX/Ge/6pKWIV4Yvukw
fheRQz0H/G7IGEf2/DxJixxb7gFHTLv4BMXFULzdVxHP+RaJqwTia3l7UFG3VOfsxbmdsIMPTChZ
wLIWBrmP885TbvUYOurWOKUZleI0+pBaOGsCc+eao9gBQJJaEcYu8kNg0ozMBKKvnPaaxm8iUA01
OhsTpCJt9wiDITWA9Uj+P3vHa/eb0N+zdRF1PmTL+sJtolD6hbWLGSXFu0kU1l3l7quzE8B5eD02
+b8YzOfm/ccr30zDRuy0ePK6fc45MJpICTQGzkROwZOj4UR3DQ46TNAWWvZC0iTujTNOkKXGXUeZ
SDhpe/4p1qEafMjJiEINkKpSxTIiniWbBQh16cmVly90cBXbyVCMASlgzn+9taDwOuxEh1LZfho9
9MIGqgtZY+cyEmaVH6UTNadB4lJLXJm40LjInkjqYyHE8ag7MQxKbKrnO8OXl8JLFy0cJFI3v6L5
bTbIGTrMPZMfgsmSxqQjm4eynHMe9R+viebiLuFw+888N/l7rZrmCixnfxyJnHxg2+THRJwpDJjw
0Q4QB0yVnyw2AJdGuXlKZVPLwPY4pPRsUM4a1WwOvn9fzGgBYBD3oTg9pODKAzQNe/8JCyftAmQA
u37poeJxGIKPm0UXJFJ3aE2+GrCwFs8fViKuts9QkXCk89JEqfNwSxCgcJ/oumxPsRJoqrO4omGP
MHMBw0hlxZlsYgJX7KVlJhMhJElqD/zywvbys8D0aGXzGiTjlMsMUKKmFPUukvBn6COaXxDyKM6g
Cx/uPcXNm7NEBpjdaLZdkAxrMXSYRZpkbgp1t8qffWWbfeXw82fwqWEHwHoDRlqSDEEmORaniuAZ
34CcAUYkIV7JcdnIcZ2UtTZMFAQZ0ryO99PJAiaKltWaAoHHQPJzoXIz3LwSGEusbF/Xnm47j1+0
DJN3aIZuWePAbTVH8JXQ1OCcegRQIMfCWyaDTZSgNUoPKc0n48BJuhCVqzDVwyIo9uj8EeEVbJnb
cBcH/0X17jQNVd1X9N42wp3eZHd0WeSo8XzhXTByDpFizaIfV0ZXiqn3XvUYpS8w93zY/nN6yyz4
USdEXNLcO3UfVhzoWx4Iy0hnR77S/ByBDwFZmvVb76XbR8+a+ukV18uISaSXrnEw9JNoJY/rucTN
cugtf6kdMIJu0mGFuQlZ1lvEyQX8QuYGWmO2j/G2QFFa1VtvQe2DILFJpbl+f5r5UnycCyQ56Irr
jY0PDxmdHYJil0PCR73aqm7geucqtwMhQ5ogW71mNEZc5ADEwe67bKeIIbCemm4+FnvfYrhZuzOy
owvApls3xCtgJY6LJFOUd0Rm+fq+0ad5k9EfGqyxBDKnFl9yiiECuTPbxI+h85zQUifXlN0qBA95
T6GfFWOSAkNexMbwle4kna2LzZvgNdo1VePJ5ouX6WYBk1g9HBdYd5LndTfXugsHblTZ6C7C1tEt
VWoyGs4qBMUtosERw0Ifj6jgiBrHYOYDOCKdCCf+wOt4dn9awPETGSFM6wy0tlqGLzWMAItDEjln
/YqFHYilP9vcQVDxfF6xc3a1RSLYiKLdkiAm2AHHdH8BnFn3aoF8rMwZj+R91/7Yt8p7fqfXBfI4
aRI93k30xvIpNs3hY7pAFPmj9qIYcybfeJRVqeqCZnPZ/hc9BrGJyxs5gt07eFVziBa9JbM3kk25
ar01OHr/wiwbIp6RDMBjHumC71fbg3HH38qqu0t6JGS0h86uNdv2232FPEanUAAKWXry3pBRP4OG
biPaHYqlY3bKE9Rf3qKosIUk8MKf+khlQxL9qBrW+7XvzPy3uw2RHIwBknAxsrdwWNWKk6Nx9/ac
Yh/ZHOKSYI+04pa3JRVzQWsQmazXeWi06KKOOJSUYyqU7w7jivBNi/2zxlgX21PUKc6u+4GHtLc8
RhT5+AUrXIbk6tEevBzwVjlSKLO9nZNhmTkJz49drf7PXq4BeQrj+Y8jG+P9gUqs21/RpT9iNHyJ
ov+Uo/9ZmrYLywyXZ2J6GbKlNw/L6k4w3SFDiBfuPq0fLXVPMCAYwdQDno/Rsmo7Ds0WXjx3ta47
VqPvbIlqr0WA1a9F3fBI5x4cbublNto+0eSteKu1VdzqiBF7PALJTgTYQGUkCndSrIR+TmMBFDGs
hJ2IjQtKOKOnPiZuiXkw99v4N/NOYjaePn12VhGwTWqPQXOaqpx9D6g1bpkMWRCpaZnzVOXWUdMs
VovAcXXdTL8ICLyEiLHhFLeOwxfzyywyDgamLV/GEeq6hnxIriI8F3qijtv95L2jWiJIME+EzIBq
FhxRdU/2UX+vqTzaGaw2JyTU3WZOEjypno58O3SVSO4C1zeLt4mWKheChFfIBvbVfp7Rg8rCefxe
wHqovvWWL8dLbJf7qf/3hX3cJxbgqBGRiArFI369wIt9WKmuZUT6+JA2O5+0LVK9NzSLtWXA73+D
2T+BXltdwM9xsuLBiAiKJK6OsEZx9xY5bp/peAL1omidI1drCVsyAijXp052vfRU33Kk3/XOKEDS
hRAv3Q35SUxYhxCgGzJpzujyvqbl2PvTnfX9dafyhfNsxhKso7mo30Dt+EH+KJpR4cVPazmJ/06h
Tg4wTLRUEJp75Nev2XyzUGt+3N8OIIWyOZUiHb/LVwx9lusEaKuzbQYILAkYc8VoiKXQqS6kOEvP
ZYuZEIfiVArSq+NwrMAHqKAjfDYzVnwsUj8Jr+mKgHZVM33/kldYfIeGcvWkBkR5oVUJOVn2mf9D
hfbRJ/V15E0Zg4OpQtSYy+Wl6y9FCF6K2EYdeezM/Psupgwryg0e6Wh5IHPgjXlAB/nEXlm+Dri0
iu7RpRyN3ijFQMwYuHa637C6cBLJnR3DPMMiOm1LrHd15DXkGP+ZyAGN8xNcrqN+PNl9qLAL6t5G
mn3cXd34JlUxrs//NJxg9iixsyh+62WWqsGVJI0nY4FDUMWaViIgEfN7W/QV/hQCtyHmrx5Xm0A1
LPrRphHBX3weXuWQXcnWMNGuL/Xt7frJ8HiuC0EQwpKO2sWXq/UK+dN7bMYb3xlcy5VPlDubljeL
ELwYIqOYwV0NlbjwKRoySm7aWtE+VnAX9Bo+VR/BqP9cAMShm+lTSbhcW9+CYwthFm+Fy63PxNgR
TawFZecjiYTO2/5bY7ORoJF6aucAVJa4h6jb3xYvwlRngQbhx/dw9NbFFY9CPFar8H+6AvQNVYH7
CBRzMs0uahK4chte0pxQTGeWBHecsxAFhWWp+CKzBpfKI6bh9WLTZ7v7arcw08DkogldS/RbSvSz
6i0vjiF6ZQjcSXmt1LO3g6gyIUFSYfREPnZx4+qFhpg3YlDtIfMPHvjMOFODTJ2IxwpjLGUzn7ye
BOrMBi69Ovn397UUrUBF5/pLsQCekCe3FxNqaFeRNCJxnMgiNpn+RHGxm19AE0FkMJ4UTuJHjS1G
gZ06MJJjosaEvofWGkOmMecu1+UdmaZ7WV4tbpnCjFf+YHiYHu3nc0dQk67OSrREPB+sixl4v0M8
fdwHsZaZ97yovzgxwC4b7MNqDFFDIEMRxHGIkL8nxT1Pb2BwYrsBy+NWMxNEx3UsRNEX32YbAaPo
mndJE+NuH9iKvc0R2wytAUlVc3leoAdaRn5B9v2RPl9wynYi7LeCQ6DYC3BPR1zyAG+TNc1r+JJS
1eeWZhb9mZ6FdKXC5pWm5NoH0OXib/dx9Vwifctc8jqlMn0Y+DA51Br/BNZf2T/4VU8l2Alceo/0
UWMSuKeqWi7V+XTdXp66Eyh/T6J8mp1yd0ts4d8W60TtJu4WnbS16D08owH1+06ph408Y3ATyCmW
kyj8N6CfDx3u6G5DJMf0RZcwVK9aUaM3HtM71DK790b9Ug8ALLealkYfatP/Rv39VgN702UsGEsF
DurQXbBNFzCpLht8CtjesijDsB4HZBad+wb51M1qnV5fue0hXYX+M2uu2TisAM9mSmgOaOt+BJ0Y
w9lhQD8CwJSdlu960QrcBxkdtEgUM69npNa8N7AP2c1Qy0rMeo14HFdFohqA/LsI0UhilX0jH+iR
xoJhxxpjl7+7YHoAIbQ2YhsloEXQcFiE2BCchFHfghigLde0ta0lM642ijaBAwCi3k2ofY6Aumcj
Da4JptDcoExI7qDnlcaKxEROlDWzEQsdrFyikjAdTjocdnMNDB1+0UyqqLcv5/invGeiR+cRBNOJ
924NHjAdD0yzzv4ugvo57UtTeTMbB6COqJWlX6ciOlWVZtSM3Yyr4BWcNjgegheBsNHJdEuSWqhU
8/cR+cmRtTEp7cHDQ4wD4Vx8Oo7ddFcjZgqlg92nbxp4qEqXjEyiH9rELtScBUje3UnXMjv//XTA
0bpFdTWrgpPcUWE32AqEnebfQMTUlqlNi+k6cak/683LUeAEFUj43RwaGdrrDQ53uDqZDtlo1LLv
DO3UFFRWsfxaKkEUmom1rXzLMBB0kY0M0xLm6hNU0kjko8XgjO1NiNk+mfpCTFHvtHu7FlKS6US6
BDWEMp1xIA4PX2YU30mAXx5DcqV7QRCdBzihNY8WIUnkWIB1xkXlqsch4iM//TmJAiVo6O5bk55q
h3rplROVM1lisziWkEWz963EyRfXfXRBAUpNTa393XLktLoWDPVxuvp4Y5D/jHeRdPuMcJtiNSb0
sSIhTXW75HeW0DeWQHb9WFmcVSDO5eEsDPslI6+Wphsdp2YvKO7pbNo2rjwiUB/88b7DORyiCqpM
JOc6d2kelYP8pBWKQ/sprbxxGkhbewUDE/TxNLjXV43Lv8tadJoyX9CFkEFgi9/jnme9uuhLC+0S
nT/nVFvDeSR349jYQxtxSiWY3rmgtUXD2xkHsDFRKJv6rI2PVxgx3dRLRkV8H7DfKouvkKR5RNir
ZIwkn/TEiEZXoTYzQFgutisjUgS9I5v3CiI93Gb/z5D19lBxp0v6jxijDj8CCCaT4LATXWLgM3jX
2pMlXraqIqs/AhZycsTBbs1tTmgCzcQWy5FXZ2YBJvE8x/jEBps2owUfuIIcw2oTJvqVGgl5P3W3
gchJCuZqzrxLVyI2c6qDGIlppT5mwTEk69KO8LRYLp8r0/E8qGnc+oLzbHnxik1czLx5YMyTqhKB
1grp7sW96SBrJFiuh0TF+Hm6drgJ1AMUUCnqcSAmcdMlZlFRVxA1RhodliMO2HlAZkz/o2Ji0t94
AkPGytXSQYuzf+ysQTPZHSeVrhYzgwE//lrKqMdAPpTZf3bU2Pn41tOooV1LpEruGk1WlCbc3ViM
wMR40DxqqYUchQJxk4psY7hUaMP4TQwJY8abaiXVKB5aPf67nNezPAeQYXUwv64g3EVK7JyEIXjz
GrhnU/3w7qClpD00Dv8QZ96QnAQqMICr+ndxIQwAyEuszzhjmUNBjHljD/LlZWYHI41zCexMkmJc
E7XWkJcmcbvXiOCb09cKHkUMk/jn7FU+kvPqlLu7OQzKHU25QWgWoMQUk/uEboQ6107wN2o6fsax
0/q5DSG+i+ildsFQUbbVHz2reVdP0Lb2nUXnjdOfw70iD6GEKlF8ywa3KJcseI+hmnfbGzPDFNl0
IZSYzXOn/Hr/KihuQzsueQTmNnV4mBnpo8NB7wMg0zsGZUbzkvxPzTdL3E1xsdrLGfP8IOkV166c
sMbBKru71qzrESq4hPCMMw/eIhDriRw2L+j//XiyqGtbBdtViZR/B+0x+O4Mguw5sRLskzpnNd7U
R+0ziSkHEojkoPdD+4AJ6528U5CmgESwqqKHZESuL8Ft+uveCAvoh6pHQiPxgWiDiJsO2grvgS7g
ujrA4HyLMlFx4GIwkyD2OM3HnHVpeP9/lTkiaXytpwxAQtqp1vIR5WAGecpgvVFTXX2kJDqbdn7w
YBrzgdjUQXKQIDgHZCyNVGVidZOiA21NJ62PuOn5dPSoGeFr+t1eo/n8pCiMh0K3lFg9qpUPcDKQ
Ju0dKXGYQbW2ZvO6K20W6SQPEHfS/jDS8NxuwRC6K6cEV9lc7skhyr34YseQD3LtNVdSmhAVkaIv
YUCmz2goP5OW5EHYQKV+kTVTSH4eedC1eIgZRMfqExmu6yKqxvKJVNQrewIcFGBNfZoBtxRAJBMF
3EdTQY2aoOx1p3miDhrX3/a++zVFxlh7UrkU9lE1y64bY6oLtbX+yhZ/ENjq0kAKwt5SE0GBxKyK
+9mbZyF2YjPvm93LmSq7FAIb5515P+f4dEMSGwba1EArWACI7aD4WqIbTkLsVCThZqMsKPbohV3X
QWSDqfMdQjDOfhNZVjOw20/y3uO0vxW/Sw1v6KgcpdGftunIlFCGfMooZSjleKpa81ZKXvhMutw8
WIQsJfX+DiMalMd1cVvpZLloSjXa2ReugiSC+4KRAzqoAZx8nshg2nNIPithDPqb/3aUMeRpQO6o
HANEeTcjgB9NZO1JzPiZ8SehDJoMCyu+ybuxKUd1fy+y5gGWyyVvg+dqfeLVYgca+ASycyxbm2ee
C/0eCSFk31WMAKiNp+Lk0LN5UnxE0QDYd2gDHZdrhoMbEi+pOwtBtnMxVVqQ0yF+4PLDWVwcyPeE
crQEVhuV7KSbW7ByJiFIyzIgxT05HVNBMdY4h91FDx/s5CI7t1Y01pZvgNEYeVoS/3PQ1FEiH6qB
IId2J0Som2JcS6ZDpFAEiVmNIRzX1qyGNTszADJpwSjYJDHCXEf8ii5K3wyMSdoO+dRgIcWDYL0D
p9Sbr138AzwGxiBAkfVCCgPaGo+ICT6BHcWGK207IFij98HgYlO9jHSY4onJhUzIjU0zpAtp+odT
VzTVEbGh6zYmbspBDMm2hTDZZnNkujjb8dc+SByW5qiF1UKsafmszpinq79B6KcFAGF0r9Ffaz3T
PgAGArPDY9kGr79iB6SwgaBH0rWDEHrL64ZRTAM0nFQ2YhBai1CLeB2gpCuMOmbf76m0vGiyrqTD
SjnTw9kd4q0+TYphTpjBu1dH/PYWY3U6ZAAx6xn8r3oAcsu9Dwa/qgWXSgEbnVH7uik987VL7paj
dAoLPEFWM5KOp15iL1iFN0v2B7mB38zVg9UR0bLcFWznH5AzuK8krSNttVLIxSFn0fBmIMojkZu1
3nwCc5Jf4JC8YF6fAhRGn5Os6ydX+ji3USZK9rrEC2qwtehcuRRE0FZ5633Ka2UTrgylMvL5pjVw
t/3ayAtfMvHNf7EPBoNdz0IiEGcnlFlrOjTKNkdvctcxKHTtP5txEMAJ9yUdoUxkaZ9+YXeihBf6
z62xRiETyiYN+a6iN8ILcfUJXGD/VcGTbzpEG4z0idC/Xsd9bBAj7rIxE724Vo3gbCTkjeSPtZdh
OPD+zQUfgnhp64EgB+8wg9PeZWKbHWFPM/19792S01tokXd/O3klapd97Lainh5WYSl3ijaAUxy4
GZwktcwSAZ7xd8KKBZOt2GZHah3SuO+I/ZkWTm7tCzI0vexe7DAMYro02DVXDCncwWiLniQhhH+D
VzAm+9s8hzqj26t96ipTYEywfp3LqLSBYneoVSVZ7uMxFfAQFkLx7ldSW6pPYQG8c2CRQDH3QLav
aGvB4Kvgfc6QygcHQ73uFjqN+5yCE66PQ4M6yDjgXznQA6ZkruoFkc6HQlhhLYUAKp9tfP3r4EW4
cdHKoGoiCU+7AntIj7PJnnO4xXijm5uqt5BSsgFPpBJ2KZbF0ix1RfHQd8kiuUeDKE2iAbsEQvbv
x6n/jeQJUzp6YJ0+bbEHc2eKtfiYkAvj53ni6YuUrEUOOz5MN7kgq7nYsSu05BJOffF6pavQe4uG
hZXbKEadh56O1XcxdmtBaejnCtkc0e4w44kjZ4BdJb6EG2Vi07ShzABGaCiX+MaW/jVrWGlbATJG
wwgBiUWykKRn4cIQbrQ9z+Ve7aSnlySpRLSFfiBlJk2HU/SbTRaWYp2zxB8yuPbKkuaMjQqxKc/t
hNQVwK7b2tpe8lq4a+TWFxS2C2QjLwdSqTUk8NBR7DCjwEcKzlINBFg8QpyaxLafk1Ub7mvqBgzr
BtNEKK+WBi5qLQK1/SRwtkFd0xJ1BhWq20BJnVIfpwRiia+UQTqKtAYc1UJnQa/FAH3tL+qHiRiX
wlnHJH1zilO0BcHj1zzhNVCIlI7g1zAcAlzZDHPdNdAEw+xaKqMCUMchMvbLQIj5QqfL/7+bjaW+
tDwyqpKjAa6WpmlGWlypy9hdxNT11fvtL5s2DCodiBel6TsdGXM3fzdQSc+cHnvcheBjBl1rZeyu
pt2cOBZLlx7wRcGSKYbUJrb01bZNhSO5/hWFVf273G0mYNqaUonYMXcS2crxKfCPXGJtPiXyVOC2
+abb+Qcr8QfpNQUZFO9htfUH+SaDbC+EPrJyUFzysiedS5r8D+r/iL/smtCzSkTu6r6Jw8NLHfmS
tH+MYlQ2i6qZl1L90ZP5u/VnWAA+F7KQ9gN1CegWDbnnEd2lODDbLz0lee2oKWXtj6F59LNk827O
azmQ9/6BPresjoLmCTXzssk5d9alXA45VoX13I3062yD2DYnnpE9IfuOh5fWpovvupCC8vyeGIZH
Bnina88tQ5aB4HwbniKAFKlA+hqN7iOqX8CDypU72BNOAHZuOmiwABtUjNrtC3KnB+xc1HZNWmk+
EV+IYQ6S82OtQZYuk3HSW+cmzd+g9cnPiUjclAsFsQNwS8vvOHBJrXw44ddrQ3ueyXNA4a2ABTCf
H2PCpXGIL+63xMeKwZbWlRcWO4Jc678JR8K8T5qI0FVjsOsoQUvAK4p4FjSID+JKoNJGIEJBYpvY
1ZNCGi/kRZ4pQ+ZupmsQvwIupCIQ7FKjPRiaT0NcsKxCMaXTRn+dH4kCTS60adfyX87rjsIrT47r
BhI1MPCjGuSejEENijdra6LVjHc6iIAdHP21eU9D1b7EsNhDe/EA5w3xhjBRZRfqT/Wl6hDrkB/w
K4nk6LKOvCPoXfc96rf6crzox6BhTsl93iUP5XLlY0Pu53Er719VcCpcQwbBuRgMyJyHl3R8t+kn
SP43gMAqY8saXhd9CayM8QrN2iYJgUXu/H4EvCxzQFcT1pn9v4zDsFtu+Ylzfiv/8JUlHDP1YJy0
6RQOh6RmwffOYFV6qHKfSXWr5pFLsexswZ63PkbPmX6NJQ54SpPKLub9fusqPKRQmUHXT83N3/0D
/lg31UK9il+tkXG4KhfCvHd55rk4f9sXGH9EiWsSTlvIGT0NoTMnzzB+k0VUqH5H9b7iPxAttobA
dWGRCNwH65SaRn7B3p4gnMxRtr8kyyHkS1veNQKzFt4AMcoD6qipm0ctQCCRckA57dGY8xAJITv8
+SQH/mShdG6tZKag8jcUtqtA8PugAsgm1DGzIqX0Vmf+2X+Q3OEOg6RnDGCibDWlYR6f+K3du3a1
Flvxx2u7mHP4l67IQognW+fzT0p9fryztLvgSzZkBS9h2gNg21CewcQk/Tpsy2GNVI01Xq3qGmhM
LQNV6Jl0uw8eKWfVMo8+5X3+9zmlQ3g7LZ53+4zLIuNqXTwovIYh74/1bxauGvDUkgd1cbHNsen0
NCfBZ75beyPpuffGmX5uPXZG1Y5KGGdn9RwQs3+vcYXp/lrixBN/qRoB7Krc6BEY3GOLHvovxMsK
zWBseIDXcQ/PSiAjfU/F3Lv8E4vgwS6xVtifly6lhc3kB770zItTiKxgZSkKrwW+Gw5CXbGkxN26
r+f2OIP8IEPifLGp6NWoJUchFEBZBnoOqBdDJz61xPChphKwLo7pXX74pt0gvMfV/YSYrGOJcYsE
jMzWKyAgwMUpmfI1UIi9IfROveuRCie/PpriKa2Wut1q4yG/oFrQb7p1EeJAoBptYFiEq85avolB
kh5xw21HQMPFgwbOytjyIKF5Kwi/QNYxO+SbNmdP0ma1mYnu83HKMtriIvb3Fc1TZnYikYZWxA2v
+mSGHBbfurKY9rdFPcmOZl1jaYI38CXo5DDOMiVaOLIodZFuzbBHftNHDzAwzZ5WtywqO3VFxYkP
miSpzqya/TZv2L0kP85bEFQIVBz8U5yVWQsPpquWRXp8cOmlI5b5YQW5xkXuiLR3/b3u/K5ETcE/
a2CgEMMARS8kIK/zc2/iIESctcTrA4cNcbmgpYdaVn2OnVqHbpQiPeT2mLMaimPFTifzx8xbucqv
EJn2jI+2BTZPKoziSseiYbjzZ6djg+R/lzeqeNtMnIQZqKV9XW/KDbFojWPvEZTaPUjR8nH2g5df
9pVjjQmkvJdeYft27UQjslSurI3dFBIoqwR4Mpyn9incGbokqO7AVJFfrOg3j/HhnlIYbHH+CQ9M
m5ShY6MvtDY/IbGH37suFEnDHTmv+1cdUKIRgRzrEI1rFXgXHnu9aTmSFrKPgLWFpUNTGfAOaq92
Zj8iCNMRbmXD2uBTVe2+kB3vs2GGv4fe3fxgNMK/vpvxi4h6Ir+kwPWwG8W/Up2QnF2xTwJZsRnT
4K6tRhMLadl3VKIw2JKPRCyGlaaC/QcFIO4BpRJi7/ddZtXAjKVsIf3hToUtFUgYvOtfQz78GpcC
bICYToRXIR2/xEcA2Ie3DLuXo+g6XrEENSP0VkMBj1DH4EF3+B3tFUYunkSUGpI2diYwVIC1XuaO
C//UMLYZwFyqENdaQvGYVgif0cu/GSnxt17Li6NKxe44hfjsOSxfvWRG68GDigw6fD+GGwmZ4iSA
7ny0rBCEl7pXx/R8P8JSETaMha1uDWvyYa0bG+d6/PkJFXmcBh3dvYfwOvt6FGvB0gJgAT+nX5fz
ac87MeTMBAQblFxdIuF+mob9qqT3UROFWowNghxbyr4IzHXKq4wiwVfuKHLp77I7DCrCjF0XA4At
H9eXZhJNJcIPVR/2gjCDKLtHnq9fvoDtXVnmOu8GsJDESYEsvvuJUTMv0+U0Bu9u8jEM7rXaXU+0
tEQgMhWHb9Qp7ntI/j0G5ucdMdp1ObleQLlLzd6MCs0r7CuIRdRx0pMAJG8fUQIhDOYm9DbMDA1t
AqOKxOpKRJqCnj8Ul0r1LYwcVJvvuuCiccp6A3552y3+IjiC5QXoOPzlH3PdUx4gFDUE3e27HrK+
4yINQ8qsfQ2Nkx2z17kcw8CzwDwJtH5FAtbICCNtQ5iiVmMIDazuJT58hhwb+8Gmo/7MNyQfJlmk
yhSs5ea0pXK8Q/tE3S7nBquGTXber+yRtXSKd+RvCX/UJdnu4Jnp12G4Eh713rfi1P5c9G7acwQa
aL5bYyN2/XyLI3vkNNs42MTF9Z54BMyouvwLjJ2On/bTeAmwh1iebwdK9PSsXoHxLXwXQ3wFR7Sv
wK0FIsFkkb1xDeGAuYnDxunYjkPnE90xt9/43oMjI4UCasgg7KVMfnrYZ7MjjQvt+beUqu45Rqvx
ak4UMq5RdlPaZtRRdGy7OUq7+Ww6fhtvBV/fUop3uypmU+UYLTz4pgqT9ak8IqW1CyZ6q0Qnm3lF
bM39RacN5p+JkhxDAeBrqRavQ9+zpXN1os9sGBJtFv0aQDhjoiXjZebmpO0KchU9C38KuT1WLanE
URdIqjHEUcb8ms+rQT/GiGp0q5Bwcf1RIdYIs+CC+q+CrQ5TlksNMh7DWPc6heKkPxKvKilVN1Yn
irjL9PJP64ZWbomrqgrdfwMasoEaK0EXF26LK/ZH9RbJytnqOFXpAJm6tGfjJfcKNy1diuy2YrkW
SB4Do48JAbGy7M4C8yOTBKS5C5oN9ZgADtwSuUHXQ88fcWOEtb324lxKk9KGj56wI4esJhYfy0ZZ
p3gx44zthFUrSQphnhQDwXdRn7DqAdZmkSOJUZwhSHRMZgLFdW4+KQhdLL6L1qWwewzzZE9FTx4o
ab+lyIfdX+ZU+GaHEYiWFGWq36hZChtlnBkS6lQMzSdZUmgbv3spYJNsI0o6QSswRc7YxrlI8bL6
z6CecB1qcG8p1PVqEI5Qlqs98EB4eixPcGDFAUhfWQhNvPH67IptGwxhgmJMQJYeDngQCzLupxDd
8yR7yFgPW+rl8qVp3sOWXPaRfT3zWUJVTuv+MNVu2pBMBmr2GcAqsmcFq/xULwmexeXUqcUVStLr
lunU6r4dwjPaPOokbi6qD0WECQIB/nhnRbt61McH0X6hckQJHo4jQZrURQ2aZZ+DoKeQ36L8Ywts
GutHI4wtxeg147+jLM8EaTbrFD9/Gq5UqEH4/4PXuRW4MkN0xMfrl2bUBr/uNYWPfnBQf4SfUT03
RZVfIBz+goNZNU6Jiw7vzl8xa3kNnn8ZMVmOq4Ee+loY553nV/AFbvNnBn6GwjO2S94Epc5SSIh/
XrDjVaTZTxKRNM5+4mK7C6hn/83Ek3A+B424RK1EtSrNuOCpuaD+AG9zgdg9lR6EQNcsuf3xftul
SGZlmaB/UPTu1xjYt4UX0g8o2PMtmJvFcs5mL7WmRtEIN7sXXWX+B9nnb6IjnZXWBLx1yolDx1VI
Dd/tKB8h2RpK8b+R3yxFu4o8TnsVlgM0W3vIgbKFMrAO3VGAy/VyqL0SB7jhYwC7qwUUh8GxKX/6
7smM6Qd0X0Uuh4qM80iWrZWipp14QKTARHQOV9ntyc5I2cawXvY4V+3dP9UVI8XjDum7EyyCFpCR
hCkJc+kEZNWjMbF3XBaBy7G3rw8ynqj6fFsDMc8nwGgDDS1ah7YCIOxr7ryFT4/iAiAvBPNzOQBY
qfecDi8TyuvjLjHGmdc74j9WCDA7wBu4Z2cfc+HJ8GuhKPNGjWmxgtnCkJ5+5iy/NmVZuPHFqFql
T3bxfz8j6RfpOLIW+bagqqiYw/LCMgzhUeL1hlZSHRHMOJRaSePdlqcv/rotdHq0j48LRuuruBsw
n9JNzEe2uOoeRXzPgH1g7m4m79NnTkYOf89AnZj1mnHLSEbLc+LlctWg2CqBO6vo+Sw6aC7myv/8
ooENKCL3OoehuMM8FxewNSb9oWCAL2AN3zKmLYnoNQoYgfQm4DzDT9HCUz8tMIxfLLoeJxy+idiZ
1nS1hJN4p2YdW9/ilNnWxpJlccWK7PzcxUGK9GvW50m1Zew5HFillr5ogC6BuRe7o7/GYBUbuAkc
FsqgxI3Ji139lrHwp6HsK2vSjz/n3TXI5xGy80K2YN/8iWOss08e1NWHlo6AhtTiOmEmeQDdcyJj
rjDxECqq+CtxJtfvVAJU67VosDRaEkeZiZrdlZX1IactTgfps4i0960kj8YAZeggJck7FDXDtaQ7
RM5YplQzMX4JrWZ4NsyhGIi3BjBC0cctfDZ/2hsmIaQSsB7JLkC33x5Xu6zWpLOl7oBEWGG0JYp4
zvCBLGaSnDsVdrp4IrQ9ldhtRfWLsHFv254OOIeKQuB8SYDSBcB1WK11gpNT74FHrm1NPlhN9wRj
zdhVjcSYLrVEecrvOoQ2Gr+BDTuUwWm06wFJLqmoc7S8nyPBRh0nPFfsRo31OybZ7XmQnawuTsb7
EphTRPRZJIDGzPRromcdNeu9oatJRb+I0DfR2ksNjQ+SkxMw/e03cqYymnZmWEsEEmpUpSWjfB9F
ErKZd2yxHWYtN8g8iOJvAUevRUqULTBltUpqSoIguLc7Bk3OsASbPwo8I5AWrfLivIcBcA3NmTNL
uBlhNQ3Gk4TmqkeK1Skj8h4WhBPAl3K0Lc7//uEpCzEAod+WXsavAocwkYNPrYbeL/mU1DwPD85t
GXtS1d1oeFdSkXAp+wtTHu22CoMiBjiYwR0Qqn9lVqSsKGmAWEQcxpA86AD7PoyL4c0zYEiB6xvX
iaVZKHFVaStOoo7s7RbOet4VlgRuqopOiwcuKc77N4VQhvexXCDt/TM4kTDdQDoNcYpohsfJ7DTl
LE1qbieU1oiYcJ4Thiv9KwZvDRc/Ky48exQF35lcUPLBQRYjgp4ypvYmb+vwY6Vq9TdZu/M13uVY
spBP5jH505hlLNFdaHLPIGzGR01xPkz+0nWcDqzpKagNZr61dfRdGHs36zvbrE77HvCsKGrL5uxw
aaqAi0Bna45j33ki0XoEdnRS0iExkA47Bzhuo7NH+ZEb5rrsWfPOBcKolJsBtTwOSnqtNLg6pavK
D8KAsaLH3eZpfK3W4s8mi0fH84GcmJnyHbe5CUHXHNWmldZcCNLU+5cJPlVluYDtD/k7HAKzHlcH
TGA16j8rnGeIjJBzcXey2z3FUT+No70KwSo3E+iZICLwxrwu6/Q+qQGqpB2bfoCLVVekuGBwtc/r
dMoXqztjc/DUaHMNMZh6DUpGNaAxtCINKkWDOVR3sDP8kZUdsgDVBFu2C1k+G6Sv5JtG/dE3N+sC
LvB9lbYpVHF7pNUNd0LE5tr7dHGMsnXumBF33eh/IIKcr2dMAmO8+yPZa5oJKwJDTRnvRVaiqE4Y
rB/2h4VUwhmVOzJBCQMfMFfvZahb7MX114w9t8jEVlEqi5GUR699NBor/ZriGI1BTwlT76u/X0zu
PBdDJdOV/Q8shHgQf2QWaD0ZDYrk2h3Ccsr81r7nkOmSJJN4IgxhPFPHGnVRv6Oz83i5O8ywFVKx
79ECzj9jIGyfrD50uJal4FD15aeLAhWph9bqnSdsgcVinncKK4y8GubJmdq6kzVpuLSmiI8Era7G
uF1AnXM+s3M8OQ6/hWqbFXixo/ltaZGaHcNCxjzQ9aZc0IjtuUfZkeilLjwn9YRDUrzFH4HBVWy3
W/ii4lWk1SyuaV07lKz+6YrgKMuzRBmbzoTUIuf9YApZfNtoTIdUH4myIaKuDw3l/G/wE/4fifho
qpu05NjdRgvBV4cWT6RVpdxLJTdqAqMy/smQef02eTodgEh4EPCD8aKjjqAPM84b46aeelV4VgXd
bSlFzRGCH8ns0x5ieWSO363GeqfcJMUcIHGVoLtsu1ApsRdLzJhQtVloP7urygie+2WvHmpuldFX
I33ToS4MzKsfDg1djb/sj6XDEY/OLd8OpHH+xG289GPQlrUE6Pn+HwELYhG7af4PI9p7EUqreGrP
DHFt89s/wp9NtBXLUZRf6AF/5lvKKSUSD99hKyTQN0qY0vDa7ncMK3GqC3YmAKUcIsV4ZCHkvx+v
8xFH50hRogr5YzWnv6Yum8xgMqgzdFnaD5eoBo9Kn6WMNtNSsf+I+94u5+nUUs6NhV1Ykfe/5yDZ
2nhfH1oolIwlvx+Zyf/ueAvtKfZ3ewYIOcfHOuT8qoqsfyOMsVmlXw9kOLq22uuc9UKV5/lnag4R
K7o5dkD2c2FTi3Ln0OF/BcINAIWeXlmp0rGksW06VeuOmdKNyplehYy6c2plJn1AVv4GHml5Y4Z5
rROe1ZoqKo0hjBRFOmbJdybFSGESH5vPdzfW0SpczBjCHuFQpqDUsgDjkJGy0Lm/ZvM5XvwYyvOw
z8Cv58qc3W0S//sVU2g9MiJ2gQ8i2/vtRh09W7bi+Ytw37vyGY72WrzLtx6VpTkcrzoVh5lppHxd
dOU+0oeQRAPkBRYOOajNsMY6hmo/5fo/i9LUupxYg2t1ecu24mnG7d2l0K7GJN2LjYzMqArWdNCA
OTnomZN5NeLh5yf+A6V8iuvyZm4hHkSw4ee7S8YVULyKAiy/Qr22hDzEXdSsJdArzYU84cyOF8sl
tKqE83YwuN/EmKJCCIMwxCO7rpL2QCOlRW78VS4kYPuWQs6+E0L/GQSMszdgSY1LTVw5kToLyfwk
UxlkSfzqBfCecCrU6Mj+UkijEldg9fPbFOVuCCwJtaDCnInbD7Yg1CNeRUrKEG4szy97kVUp+sea
L4m7bzCt7v4gknNOKVPzgXoF1e8aP7E4YOTOS4Tw4KDtan3rX3Ljl9g1PiP4jw4QQVFHTrW4TdUc
g8uPcYVx7Fr1/Xx6XEx7nC13I/dS50BRzxW2/8p12R6Q4mNUnr7GUOlPoOv/awyi28AHmIRrconq
rJNXep0FoeBB/+tFgsjcCT2V279OzLPCPu1CtYLljpBMakEnU3vhUuv+C4mU4iRt3inUjXdNz6o9
hrqPpCqFgsJUTC55TFC4OvCmfHiDPv1geCwFwfVQgGx1+oMnS17NasYa5fjHCLaYgkX830sq1kQF
o4dRWPQNXpRwOcd9vTnyXrbj7Qshgf3so2kGLaxCquNOTB2Lm3ZzMtSOLpkFA8vrI6WsuDZlcFLw
XMI3eG0EEC/VU2zQr6NbYKB0S5mF26wLczBJsf1KnaaSoYKQz1J+9ZV5f8KoukN9yxG73f4iIdbL
hQ0OwgGevko29n5904KjRMJzJBrxc54j3fRtNBCt6mo461mKsdc/pQ5nfTd39+KYC+u5gBVBXwsl
HA0X+gCueXMVpfqxebxpyndQFqepSzFLLuuP/4Zh73hgis8klQGU7Lqay+yeaayRUJFM2epEdWwB
qOHyPD0EQYWMfKIOAG+VZFGwF34RpbQQQ20LLF3qxay1Z/s3fA0g9036pt89aClD4EJEJgzWSizJ
ORPAuibxnWPQmtx4qX+bkLd6eeuEQNLPMttUNYFE91UCWKNgFx4NfWjOIdy8hvEwd6Ot0+a9sZvD
FEXw9QikeOCC1GM5F2MZF7vVdsKVuakojnT3NKmi91/5LEcQeUpZK2PTZe9RRIZ1UDGVEUfw31X1
9/JFsQLoEBNcbdD6aNrKF6ZxUvBvsX+ITajDz4Bz4zqB9O6gvhEtHZ3xen0wd2aG5D6Hsgr+Cotp
LhUYTuFeblLfFxI6lxvczu0ha7uC3I6e4gw8exoRGQu4vAtruaUlFdAiLCspHS5kLXklfC09CFq9
wzmihdu4jQlEvrTLqI1xY73tPwKapEMSheJkN5LKLt+ve+4n03iT17i336N8FKPYU3c8O9+Y2+fc
RydAy43gsb2FRRkkXH7GR+rBehmjKVgRAHGZoDpAiRHXkrGVXL5InazWV8XCCqx12HaVHsocXKae
PgDiBrEPz0HtUR7xupswuPAbqlS8ZeBhh/sxtZ5bJf1e5WdMdkf/g2WpcFLZx9Ggy7SHBSdtflfJ
V0E2kon9k+3pGUzB4yZpR1G80pE4Ra2p09GyO65mabgA8veeOarHhPji8S1TsS1LyrieIWRX0lEd
LcHroG2Fo3ULqApoBDh2oyE+xDMbR/dBr8N1GQbuzXJy9Z6AzgwealaMhWW9601ijTpWw3f0/o9u
F6jmL/KwPBrHk5aZ55Vrbfp5XNKjtmvRknUOgdRcnB1sjsreDvl5qSua5UifZoATIX6G/oMaJ3dQ
2QHXWoaUoYl0nOPLxEI+Wu1SbaL4531YFjXlnY1rYYGwY78N9eATJTMasqmnjy7JoR4LvM2nvYS1
YfLbNlXxSK4NZplDA2QhJnRRM+VzBt6z59R6scbtTtZ1b3whe5fBH+B6ZMbQ3fh4YoMQRxytGGPH
PNc5M2IvGjAKThJZ7nBQuw9kh0LHZ0F/KAQDK2Mno1DujWT6UWdWggkrSgI5qmE6srnkw5GppbRj
bUih5Qj2mY9njutmnntDGg71Va1eiTKb/WlfmQpen5mGWezdr52bccUVQfVJHVqY1HZYQlbJysNL
XHiCC7usZRTZrH6ClqD2GlE7GE24Atz2qF7U1EmHtPUKMFmSNnmeKVsyvJqtnp9tydZIcKm/PfwH
rrenged+oJ0h8+ClBlaC3Q54ZxldCfDN1lyt4r7Vb0MC73c5JmmhNfW1gKaAVI16Z/TQaBoTBSo3
EcIQU5FLJJBgUuberzTORjn0TNTCDR5D9m+xWfpLU7S2TnCyYrAeNmWBLTPk4uMU46ctqPVLz1OG
LKpk+quIb6oaODOrWlFreYNaeIe8igqRwV+Gb3BYcf54tPj5GgGj3QrvPn5HEs5YsahfOT9ilIqP
TejANaHCPFAJXf0By7Zm7gkWSiHiOKZnNZR+75ydP32d7udhaTQwmCRu1xMbC78VJzOHI0e4pDCK
PJEQwycjH1dblv9/PMacCsMaVDsJ5VT0ZYVOXrm9Wo8xbpK5tLKzvipojigLZby3O6ATZ0LoACrI
ccgkeFbjTc7rmXYWJ13gkIFUq8bMDTSHeujafjkKXa+3XiWH3XYiX12ZVuqDvSyXj5+0OaIlB36Q
eb8XR79ISrXSuGjzcd/UvIifczn4lr5EUI1b4cdJFkAk9CB53xuvpVjuTQwMh38fO4BEIieUKvhB
FljfNv5RYxTE0jZxR2KB6MqE3yGSaCg+ubR0zyh7OLXNt9G4heZrmL+uPKWTE881+yh2eYgD/6ZW
2KK4lQ9rCu4vmH9jw/ZQIOV/w1odDj8Fw5eT5yDUVnkPfjegS6TTm7ucqUolvCEU12LawreSXZIC
u6wPXrFiWpumnKOguH6Sh+b1Mud/SXOPdl9PvhYV0ChiGuCktYHJwLlrCpHxRcbhB32QE7uVLWYP
KbJnAxedstJvL9PId/YfIjrrz/rNR0wJ+3qwwQA7ixap4PXLQiCSpLX4IGTbhIy+ruy3dq9cGDFN
sA0iwRlxg4G3Nm5EpzoSpbwlZ2fA0xtSY2x34bviHWGbQB/kb726ecpXmPRivo6J87ScdbS27W+H
jZLjhWz9tkpHBclJ26voYmSKqbdBFmng/Ca0GlAMuPGVj3yq1hwm2o/VUusik9+FbUUQpuGn77l/
bmPa7RcB2KW4Wq6iceLrXci6N5YvlBTjV01ioBxbOJDk5D2JaTZ4SyFjBZxgGLpo0BDoy8qjP5Ri
rfd2sJ7Ex2lERqapnWijDcAE5SjfxbpPm6skn5JqrOLnruZFU97yvZwgJON0FnuywIanPKMYbzty
XVpNV/6YZTtJ8UG2NS/q/JXExUf7gXWDvdAlkejsX1hWQUN94bMQR4K/YqgwfxJV6VGZ2k7s7Yar
06wB9RZ8hZ7sW/KHTLOZDm8YRaVu/uPdhtBk5gGma/SN+PM82yiNNWI5HWip4qUj1cX7pdLBtpZ6
zX2TOis2uNFFiK99j2mgi/AJKMjixM9Fth5PhkRoVDI/UcmLbntS+LMYzKvv8Wn6iaCOLTAveBbA
DSJPCeNLfHt4LGuNxWKubYJSY/69swNwYJPexT52KAOZPwM+gSlFWRqgynKBCU7APW8WKF75K/vB
U2yl3fhhNoO3wW4taUGjceqE23YLoo9uLZlb+mFNl5xhhQvnSO89YOYFiNygsYymCGOkXTksy0du
yoywlYNFkO8nsohe0easd0MV+co0dGzVVJnfnLnOV0IS7DN1OYTl/gncW5HJDk42E/i8A225Xowi
VR4ZvwcxvIyGzOTmOJJ+YRYaj2dk7JIqcBgEhBYacxHczEHI9W2TblsPDy6ypYlb+h8clD8yinPj
T/D2hSd5DnltkGRDeFyEQ3wCgtYfUlaSBn0+4bOPBSqD3RH8MMJOPWBpdmWT2mCOqT22rAhoBGwK
id70XbZf25mD/jl30a9GnR9e7tUmwkUs8BUX2QoP9+AiuS6UVfbFeHDML+ZtL/Fb5PXd0DhHUkT2
5oqwYZIaKtAKAI2HWetZ3lrIxskc0iEhw30vE0T4/iwsPYBcSUTKbV1SO2wS1rc+RXp7BibJKIrG
jF8r5TyxLZXTFaBM9vMEwRqLdFzelAHmYxg9aJAS9Ck4GshmDe3gJmrej9o4HPNTcpnOCH1ZHtt9
KqyCQvP19KX0N47o/m+OP72pSzsmu2ZiV3+oNlTscPv/Xn4Cd+BOLbBkZsia2L1y3PBgqtMQhuIt
KXP132KXWu+S9v0Z8NgS6/BWJuDD7W/nz4isgWgdz8+2/RloDuSOvORuPd1sKDLWROPJoZm7BL14
3Jp762Q3la4VJ32Fg7ZOxzC2g2rXJHz4sjJ8syM8kmRuJ0BD/3yhjVooLbnsA1eWmJNAQBviPccW
oS22DmEJqOX8u4xPyQcQtF0mtBNMJLS/ME40RR+NAB3f1W3o+XrEMgze7g5xHBzn9aQqu8FHvRm6
0B5m7IMHMzLjIHHC2q02ExGsLrXqnexYOEkwdnn3khQDDmZ1Ujn6SNU6zHVmpUF9hClnoSD6k0wU
pX2ZCgae2w8BXXwMYbET4f78geWyQc4c4KqxEYjVDW8vEh+eUahOJ5gDhUpJmqNvinGZTV7yN4Sj
noNs41B+Vp6INo5qKhkHRHlHEgUODSnvpmh75e3p6tErX086e+dbyGEhcKX5123Rx6wFRM9lxrxS
4/ftaz4aQvm+DvFm82B+SqQsJzIq89lBACIbQs7Qcaur/CqjuZQnmO17/cyBWhPO597FkFn9KMJG
2mYvS7Q2KlKFA6PZzKj0USSFn7SE6dCCkSQ2hP2mLfl/TAeeJvojD1FfrUXCQDmjfimUjQjsz+Lt
oMMifFqXA+Al+WTjeJugQ9o93tE8HM5CUZlWgc1DAYRWa6sL1SJOrCIzZLmxMKLoVhEgU4STaNby
3EKo6RnRctITCr7tufiZO5eLiU54g3TjR0XK9azARBQvrExqj6kXYjeatVfptYbPaHaOT8PcmlCi
+on4nStoJTtqbnaoPwAvJc2T5zciyVH1FxJyzi1F60++B8WhCX0egxXkigs/yvVGwND5FKKRbxFO
fzKHQah/G/MBNTckLpzNhy5i8Ic4JrzNSGzjCVQPRSWs1OjEXcpP/5VOZoqQEp44qtihZM7z5Omt
jJEwoOIK9Y+5cZf0eMtDGoZ+sCRiQElrxUkKW7wuB3ZM3WUW+A27G5e2QkUYwmLuivl/gAIpV4h7
f9+bf9jJubYPkzxybjOpyinNpmgPCSvr8M6lzo6bk5WOmc0txJgclLE9wkgKtD/tnunkiZhQmeuk
9G4ci+KAzEH+gwGUSNFRG+OSx6/WCRo/lOdZEiUTHyXNb1IWHZRzGdR0PNoCfAAr+b+V8zj29dQq
ny/V9OAXmk3V+y6YcMzQ0dNBOuVYFxleQioh3cBFZENkrqte4rX038IGj0OIDD9u2e4NH8+E7DhR
qT/ooCUHPrt9gFRCaHIjB5GSGYNlkekfuKXQ/Op0guyNEodfDneHGZi05Udau/ssSOVxKu5G1vOq
WMKeRb2Bn9xVovgopbOBl6OlKKHxrYmcCOq5ZuinRAkrlHongaN0OY20Rx8tSn1BIlQSxxRs4wqB
smRDAxqFHX8UvYshKmPBOuP5nYiG095iGw+wi29M6jsccwATgOBtpOmTLEg5kviG44ExnRnTpW+2
+ufG+4LLvqT0eO+aylfenDndSwKwj51MRvhlb5n4SZY4xvZHIYpBFZqSJRjAn+13dAvuzKQ0ofE5
P/WncCB6t9xnn6wB8ixOtdsf84GWrX2eyj8fxqPJqFupWzwM3MQSnhmlfz2KYTxxlOQsDTh/TJdn
Ww8LoD+qiYi+DEXIYT3fhmAwYKRGfzY/k/kb2xVvB46y5hApPFdedAgDTZ4dFdVe2jidzK2XO3r4
Bg8zh9qBc69sL65LlhDd4stcj4wCbxKBfmLIILdDhutORuwVGMxxp95/up7fvk9L6iNrxw/DOU8N
yCqPCXXlpsSt4/C2eAta3VRxREzUdjnEu3KyExzLehG0FTje9Q0C0+B4gapK7mr5NhN5vfCdtKE2
C/QncEbv5XJyqoOfToLrthVe4kteM2/4xcsUW5hS2GI44sFtyRRhdAdAG5kytU1kW9MdLjdY+r+R
3lKiaxtzt13gl+lnb56FD/rznKKODzpB2FD1ChHRW4+YYzqAByQ0a3grJsDZaq3TtdCGUkVWgLdE
KKEbN75yVHlQXnczRZpLdWW2weQiYsggNcS2r9ClSAzyW6gnbiUpz3fz964jmIcdAOi8Xdeippk9
kVnl6djziz4h2wMuA/2cr12iuxcFrvXeIoIIKVtgpLZOMUUnpRGjnrCu6y2+0oJH2QRMHz1B88D8
V85YFlCwZRkmtoJtgRjVZVNkEhqTJor5x9+Ctk+P2dEaozrhWSHXhbwLMOopIMp9H5fxgOfYeFc/
cpmPao1iHC6oZd3cWBx8DJY4l8A0hvOiOgxK4N+MhDq55T9CSC80OeHoW0zdiSro6T2g8J04TwWB
TVS9qXewxvJ/a0ylSTii3OqzuZxlhUH3ln+/FqiKS0aLgcUkKCJNoAK5MSnsPAvB42aJHTwhpxr+
G1TBJfszNMWS9poIwbuvs560ksiSUQTSVBmluqb+NfhcGiObVxDu3O7kBooUU4llwTBxPz0PwBUE
O5AYv+vaL/rG33R5o3BkBL/XiJPVzLnhPMScZQawSMwZPKdFgDc1PZooGHj/AFQ5GI7LE1ST01oV
ilIyqXsQfwgW86YekrIiRWUFdjlISX68f87kK6aTn1NlP0etKO97CGIFLJohpsjcMIECTK5bwxyo
WCYUZ7k2Dxa4MZQBa5LDQ7gYm+Tw9Ycawp8oUbKrS3Wwp7BzCpjrFdsYkG7t/HlASAL54dNrPvqd
92mrcstCdxGpJT44qMZFulkmuUdcnD5fmD+ohVPMaUSqtiRcwpHEvTtxzwnMJ6LY5JsQJelcu2xD
iyOVuwUgFi/Ii7I+1fes3O/lmCvs3oFioHy7fFB783LhpBnMPsnTzSg+eZwCx2z2xTw6CIoiJvDU
MAmiPzhOQ1gorBq7+4nhL7/7/kzv79GjC0374jfbbp6zJR/PwLfPB6AN2C1fLeWm4g6ui4Uyr50j
hSjPrT01XGJf+WbEnPaJzbZcqZfY0vG7+NO8sjYB1orQXwejTjY7uI8WbscQvdFYRfxKClIFZHFi
Z1ot+4GBG/L5HK+i8+U5JdokxJBpizdnKfT9XlgPO2bGfXhleryqpdrGu8muCtmDhTQvAoU0ee0U
Ho+lOi8Ij6rStunQ8NDdCwwnoeILD3ND9bzPdVsG04Xm/8cAw9XJBf7we88MU63dTbtPcGlxA/NT
2I+RPgHjsmhMDh60uRRkZKuoqzP92/baW0UF39cvStaYdyr2ASgLHSKgdeHUz7xHTUQibyUy8S+P
YV/ztdCC+nfTEn1wctAu8xDbAcaoA9d1qKrPKrC87IfWm/CdD3w+mq1WBK5DNq0YOG3PgrWKMF/e
I4Y0Wm4sEyKziXxVMjAVqSY9Z3lraqvkgcYKumxpxODmqODbtHbcz8yvbV4v5Yl/HIFOJhB3mNaU
nfLgzwanVevFolJsOwhsOzIj7/Zm0XIa9kG5mQMxuWp9VmgK1opil67xrXg0dQnFl8rcNdRzfk6u
h/5XA0pYZI3/G00RUPHD/ixNkieH8FbtKU60KoJW/Fp8AnXf6eSosoC7OAppDODVKcndi7t4RjiV
05DVUjgkd2Ogd3VW/jpLuRaZgWjwIN5HSd5b2qds/G2EyFeMGuAn5MWZlFqvsYRQ9G3GREUthiYM
M/9WdEHuCsFSFFiR3sfd1z6b8XunxJKjEsNZA7YeeRRLc6k1yQ4lK2HXlz/GpmWrtN3nes/zWR2N
WE7Sv60eDVYmMXC57NriAVIcK3OoEJVpjF2mulYTeaqOVHKzqenYF2ueKecr/I7sEWiNRlEtL/Gr
Zs2GenY6P+ezKC4nhGBE8Aokc+yEDJjpWEJr1FihfJWTgnp5Z9vslMJjl25t+mVYmIWcFICQ0IF+
UtAqHVWW0MQs4GOnHkX3l6mAAh1RqngpCz8G8shTyIKi7PNTYWUw/FC+sZ1WRjN2O7mIbpEVDuya
lFPunge9qXYWUHcomgJAQs5FS6lxMIPqBwrPkXfCnQE0souaxCdikSrPIWHfpzXMVZKUde8+BRBa
KfejGJSzhT3XmIgnEtyXeuKQdtTR6F7KN3eyUIGaDzy6gBHEl5bZYX0QRGIx6utBJzJgdis6PGnL
z2SBQbGDB09Cf/I7zIIrBaCCC1wjFXIwiqiQ/+fBAe/x3BnpOzryuKgc2ik0DU7fzbcI43PsrZ5t
L6l9yoykuHstKLZxMtmnV9K4GU9fE/nGcLbEtmu4wMAJX6FyN0wuSZSLL9txLZo4LWyUZjniGyxv
9BvAYbTHjoZFobHXro4VzZGb35caTHgXx/y6j/SItQ94gY1ppPxOLGCKeIe/9U8RC9ktMNvcAOEl
dpPGMZnLWjZjTqYDWLMs4TuSuoudWbyAvuZ5ik4F/WFXA20EvoNGmy3FiZ9CjePdSptH8eD3QKiY
HHHyexyYOqZ0DTB3oLMfl/UamlIa5Y2T3yuXWIgOY6712ahdcAvgGP9RLuSvrk2AuBby1W2oRyT7
cQ7e4TA1qfzUtON686C6tstPCdOapHKgWkxu04r19WxZMOhZqkO25/eYVkQYIaiWuhzjlC4IE+MD
W2u/3Qc776/XXRZns1B3oSKHK6zf5OVgqeLiW9sAx96kUQtjP7UUC0Hzk8uiO0cETCg6RZgcWdIY
PGjm0QeT9kJjh3NtEisdwGiywC3uMTkXHgsyRGP5iriHaL5FyrTHINst9ae/7SFomK0x424I3FgA
l8U8nXYHzINiOkTsKlQ9M93A2COiDHeT9ZuOk8mcf0OS9kQN0voqgs2X5T9hmpf0hy19lPVip0oi
rLbi0etyzr5KS0io1mAHR1jPEvO95EMiXRO41VPMY78wcwSfEVK7oE7Vnrk371XzzEXvWK4wjMMO
Jz0AgvulZD3odvCKpxyKbQ+O15hx0Hj+s5SVoaZgdioyINMyF9oabK17V6CCYRa9Dh414hPXx7dP
8aSm9gbR61cg7zEVMRmX70YseU8vCa7vawWHjwICkZQHy87hVqfTdyRRcACB+d3O/3FVE8Rp0+gd
rCOHVQxczj+LaI0MhYBhhHkPTFqYl0bX53RkuY6BZKqmj1Pk6HidvsTYxrmJTWiKrrM5GPsGFoHB
0n8e1CYAiYy9IuxAEMOjkivKJz+dKSZUHwuRKP+1ZNpF2R7IkD5sIDVR6ZguQuxqBlK/0dxNVBYj
knzLCAuDobhiKBdcVJyopcVsVRdqviiMQo66gZcQgNqktcDJU5RH1yO4N1jNvJyi9D0JOSgX5gBv
2X/tsmMmQ9j9nITA/P63NiNyWVgCj69UNWoTOT/DsfhxBklNIkY4ZMYcEEbSdrkbCMx5gQHHzzXI
dXZvm0nz3sZbSdSF3MCmXYbY94JR1E+h3Pub9ZLRKE1QeVy2JONpo5kv7zo3coQSzv3pC+wAivbE
3Sj+SSlq7Vp7oOoa5JKjoiIWjok1vjqTVRcaH6LvY49pPDt4MGRSrgOkPeQOxLsUIHdZjtgNevTQ
YINrLkBrFhcM1km66sOxD4zPhMrRiE/jVYHfM3Nk+YONrU/q82ad5za94f2+DBivaqgb43QpUz5B
Q8NNEdK/p0dFYLGOtRQItNnw863yISMAhvK6C5jeYt9slU20h7gb8vPAVLQPUAOJURzrAwn+ucRc
0N3ZyXrN8yQqdSegwG/szz9lIkGQu9HLWcTL4uGEsJD+N/gU+i0s1tEphkRd2GUxASUhat2Pz0jU
MaZgwg3zj33SfbMaBhklds8kq2hXtIQH14s9ceKwpyHUeONXs2MPr9DnMvRDsppcdQg/IfnyQa8A
pOPnywWUkkSINB0O5i63x3Itvw+KmgktzkDZ4apDWPjJkP8kmfZHU7KbGLYudpwqegCh59gGTmSA
pnyd8h67veDHfk34i75j3JmRTW2TFEFkoXKlfyNdeziR8o+KB8yBnzbQsQH1pVenIbqMxGLyCNzd
QAR6cFGxSngZeSWugcity1W/vaXM1rNK8K2zN7rDqtH0wQh30Uw3qw4TxHO/S6h9hCIC4pGKRnI8
qwR8oeHoY8RQz4ZA5YIWpIzs/tuVSgHopiXlNsC7Xq7T/TQTOWx/mgMDPF9ePbv2mm97HVCIqkpC
2mB8v5UiHXsYbFSF9Ug97Zib7ZINgMyt896lGVCLPXwSwirsDQbNuCldu0PypJKt94JygAX4XR8H
dOg5HWeSHHUbKWgMfu2yWXEcNoMhIPRNSoW9uJywwJyJkwiYTuP3jBFtyyUtQQllAsgwDITRGzO7
hfRhbBxB3A7CZIDtXX+Nx5RRFxniynkQ0FrUtdZsDHedPXl99tlxWnQJ6B+ubDx4akCM3M+iUwym
yuSpzt28vWxztCmDxIkmjB8KtWqId9jj0R7Xyc+JxchoTehdJunmMmK6ixhUsrd4zHN9Xt1MCcZw
bwLJSsMfxpMjQJZPELCbkGNoHYK30OWJ7Aiil5nZz4J/o+fsidlSRXT+Pn+xYogSCzc/MOky0zjY
24QR4dcVEOE95fReWw2Rg6D0N0qLNpXQj/TWqx8pN0mY+ob9KHbgJu8Ng581WM6aqwebRHjT0hFo
v7Gjgdfs4My61cyP0LbNtofM1VCoRPUcUDHd3LNIg7WybFpajTB3hRrdB1e81zQOD0g9+yxq8AGP
tC/QVNc5m/HRYBCxIsro8ozPuN/4zu0HEWMUpVHcjBngxsjk6qfWM+20yCXlyg0i3APpzaZNXAaT
fqN7CvMhUl9d4X6yVefIWASrk2kEdPZQK23KcXnxly/ANtypespf0Z4w4uN9gv/MWhvWz17ecKbj
IrkdCTF2ASZQbSYGYeN1WHNrrHm5uRWD+BmGiAzpLIjg4++BCxlqA2TXX7ndNh/LEoenkHOENaDc
c2/DkbPX4FlrnfG+/Q14x0J9Zj/2HME3smOC8falpp7r3YGobj5pWOH6DTUj9YSdiRrS2ufkADIz
uSLap5sMJ5GgLZusEjUhfCWWuKl329xYcnAR7ua1vBHaNbuGcAtdW7jyynfonMfHrDFhgJbU27Wv
buXS3U26qSJAi3GRjAodKSmYia8S8hLgP18RQVXc/6ZTIu/oZ1E9TCDrkwTocXOTPOg1TXlL0lT+
Ie/5v/oT7ZvV7ZINglK7CQwz11d3lp3B6oowNDM9omK/advWjHbFUvHNB+q3Th8Clda9HD7PHbkQ
KNe1gFKjmKOkN8XFNxFkSNvD4z0GYeV4pHkhimNyexoWdM2lU9k8jTFDmvw+95n+zpKD9NLjY8Xx
FB9gVEv8pQNC03wSzyoxByMB/aZM9dQYleY7Pqr0VsscFSv9ZFnWXWd5Qz4MlQVxxkd82IK+ZZ2A
gZDuMlAnYwTTyiB4jDg0R7kLduWSoIZXF3DwXGs77iDHfTxVLhEVzRbY+g+RdTxhVQs/tt0Zo/q+
G/pWYrmOdwtFj6sVsRJ+9YCg+A8wj8JYXrELeXelelb8KwHyhcR/qD/j8y9zxYaegnIbgTUAoj/m
QyF+4s6gQ1s25odRQypX36qb8WEPtJZ34MnaA7xBFtSOWFmrTtyLdCZ4PF8dX08Snwxth81eLxOa
5iiu6UCZ4T+0R6ymrt1hNzYQft+S6pDymnsClRjIFzqGqRkneD9hgknziBWpHx7UwaVM5uKCS28d
zJD3SGlk3+s5KsBG8NzvYFSadX/i4FFv9IzKSqybYfe+th5NPEaBNxuhgxgvWooyAgUi5pTgyCAy
PYLOQ1Kku54lhQFVeh8YiLZQkLpj2tsLjGNPWckVV6Upjnqq0EHjH51Pu8ANSPs1S+V3g0qcfFjK
5OxKKUVNMpiJ1vDiKN8oNORyVxSOqXo2ndC28VGT9vPkxiXtQSeVGNzrKzWLMnbr6H/3KuU/NP+W
aAlbgbphensZXHnTSviLV0/al5utUM3eHWiUmhZDzxS1jT1C737hmjyKsnISrDuYXTZrmIXs+jLf
4eeSKOQg+1YYhUbEhV3I9Vi7sjp7dNAN2jOVhmDSKNTogL6rkf/6h9KonMELCiazpRCpvrmUjzRs
zVKsaWNmV3NPqVVfCb30YtfIKkJFopVAk3kYLF2zF9rXIbbuqYLjfFFa7qRc04rQtZdBAa2Dsfzn
mHRvW0A19kCGusN+3WrFCfSKShS3lJMc79cMXP0buYI+5GK4ehXhNZpSsSaeqB7l76gEvpJLjrUZ
4xuzSMKbNEh4c+tW6iFLpSK/vviIv2b09O8o6cCcWwmzGxBMKwUReE3mNZR322k71k3HctWKf6rb
AtqJGhvd93qiSHDT8MvEF1rV+5oHgmP4etht+JvifhVOnWcG5qS/r0fVKGlSzK/41D9yw7iX4EOa
/JAklPdFnJTBpzHAx3Zsk7R760oDhcR+rQmcuFmSWLsNwBto/HUBle3N4F0TDDC6Hpmx9usg5nhZ
UNW49jjyG6jpct8Oh/Y5tQBldNH99w4HZT29gbX9029xBGG4NcyzGFupQkx9xXmiidGXqESjs8oS
Eb4rR9rVH3kTQoXp1vuemOP3d0Wg2ImB6qdqek36IusGkkauPYNVZ9q5+Ju1gr1nLApizi3kIq4P
VfdAM8ViV2w5s4UZlwPVbKfhsv/NxNyR/Dgidtaheb/c0+HAaT4wjmZn9xckVbCidP0I4np3W1JG
UFu1EWcDBqGX+qfs3t6Xqz2vr5wibV24YtWWg4rmBK9lBUGHmp2958WSokwlXtlDGiULIzC9KdnY
e9Ytsjd8jy4nJj3lCjIVYTJoRRjobXWJ4VFZaV78kJN/Rqcn7VWD2rtTTWOHg8cEUHjZQ1r1RUnR
DNiWAofzE8B4y6Ni0ttXCIjpme5OTl3/wgenrsTMW8XqMuFS2fitygAJEm12hAa5AwLJe5aTiRuZ
8RAxr/sc4rBLRtaUgmvUXdi4qPUvrxcR47PoV/1b0zCqpT3ZTQ2L6U7zbjZEGFtB/7eZw+a7fxFt
Z8Lr4x5lzTvaMG5LrG/X9varHDL7E0/6q78oleNYt1V0oHyn4Lf4Km1scGr7lw5oIB9OUdSIoEGc
t09CTn1six18Lsiv8VCAYHtqdrUz/NMe9A5X/iJIc+8m3cl12VpY5G00KKCQYEim0Q08mQ+sF5CM
vqKrmE8xDle5c7lPf8i0V9F1BxD6U5TWhTNrXAu9npKpxcbYd20c+Ru3bSj+ULVmh3VIhedWHx/w
qFIgy8fAu9Fxc1FTW7Zq1w7b8bwr7p+g5xaMgB5wLXFI8CA+P6uHE2ZZPpmXqtJ6nc1jtO6XUY/Y
7oT27FKmO+7VhT39JOc17fkUNNAFXmMxyAVZNuxiirJnajoVfrBk9s93dDPM1czMKEwQoUgezGXg
zuZH/qnpXPnpEOaocgtaYD/bweNGV+OpIB6S4nY3N+gv4arjuXbaEy1CrY0RcCZcNbiQFq8CBM84
IKKOEbnQUlTFsIkcQjcB9Do2E62y3bIhzjFR1xMj/z67eDwp4I8p690vfhOpncyFqE8Ffdl2bEXe
THdp90pYRHYjekN83dCUesGvBoBbbbkK0aGlf/YqL9PJqj5kbks58zp0Ssdp//qj8LY55aRxhIN9
aiZwZ0c4JS62ENk+qy52HT5Jcuvhqh5n3ZPtqQj332VYEXgv25Q6oafegmJymwA3QcrsM/FVbeti
HjQ/N/Ks05L05mRw6KMu6X0mjLD8PEG9Y6yXxR7+CzV8hHxE0pHYd7TjzrdgUB/ky1IJrEpcjnwS
FJFqTgHme2P3CDNu/nE0zNKxato5CV+z18p0GL59qTlzXlCMMBXeiDGRyxcoFzxfHb1mwmeZ8ldS
34kXH8OzzNug9OrUr/f3YefFOSSs+zaSL6N+jygkFqz+0bZr7Pr7PfaDBNnF9izt7MHAVLk9vn1u
KJc1zSxL0s1yigFy1N1+nRX6DbeC08pdrAM21N1/G0IcHI4/2+5PVyuo1SCD5Wj2OLlv1cmGju1D
oAEF+BltDAj8xLCPplIGmg3yyoU4ElYbsPDgjdhGjkXIiPakS8j+Mhzbd0yUQGIwYUfBeIoY4T1X
wVmkURsQBr2YNYT8j0YZRVZmsmoaxHLWxsjQKNFw2eEwrKkifSJ2+NCBaZJwoPgORVvTWO48tLGV
1RdrYwUjblVzQw3eTCTt3WOx3bGexzv5nmXUtSm8pfqbsRb0tXij3YxMJkwxJYK24CahcGoc9JSG
tAWNmLagDWZ+LTsjHk/k7JlCsOzvWBhx/ls1EEsp+6nky535nWDeQ5aBdeVz3zis8veWciDalL+c
TWBd4lpnY80s/WNmMBWuV/yZHZWQVluB7gKPlc8EGRSslKKpCK3OrIy/+bp2LDiR2pB4Shxk438m
xftcwWHbRxg9MO9RA0u8fRyad8aOUVXEgExV/FQW20piWOhouNxbQ3uSZ/tesPNh/eiSSqTXZiXa
x6FDdwSyS5dJ5lWuDH9DNsNIG9e3m6aikh7ylRWb4nBNsYkai4IrlupdkmAuTaDLOMogdcoJwLG6
n5iX+KLEi4oGqdexuS434qxHC8j1UQwgUTsHhFD6u9txp1TwaSfucDsEPZSb+Esrv2vdqLYHpHDO
7aesOANpE4NeuTXiq6lhRO/0tIBz/YbZyax9CgCdlnfg55sMI9Cr3rTlHNkoqOFtcpGOHCDphcWM
9RRkoSPRdY0x9cv+PdW9UwURaaITe3Ea/c7CRJoM+ypwythLKIK+zPuhFCH+F3EbE/devfcxLElm
tkxlB4XbKThBW4RHgcuZ7fyF2P8+MgFqkx8sFsLCyimHIVAxrWGb9oePE2RKtiYTL0XEZgp6q8D7
Rc1Qm1rMUrVKbsq/nhZx+JraDTfmgiYf2NZu2Y8urd+Lb2Rd5ocXfinIhV2qepLOOU2y7UgVd+N2
JWt1RtKUG7zA+Gb+dN1oHzaQSHVOHsVeuMdQ5FdL+4ZFuDJiDsV2ggyewakL/goHjGb+rsZm/lWn
76CnQL20AzT9zO5dpwgDSkWy9Cac/hTI+bn3e7aDJanqPUF4x2RWaKN3wTEIuLUGN5PpJABd8q1V
8KqLvSXsnP7dSoQlDOg9NjADOjTgTmNMFCmPYcDOaDY3zvJD20d//HmQKAg7LSpVbTH0I5t7uiB7
0QMIuVB+rULi7gN2TEmLVB0k6Kdkd85ZwzsXF/bSNyBAkRRllno/J4M6JbdFu9IbYZ8l1zSzyw1/
Yg5gXRZZXtEvLMLaz2CIaQ3vrk1CbIkfp6WToLTqaZhO2k2h2UICsUqNok7qknIChAO2izHljWi/
HVT+8D/qTqFc7+wJB4PrZoqox0EQS06egeH8zKLAfRzTGwUUI996P2QgF2dApU+f8Dzpsh1KFdgd
wWr0UC3pGVbBr7ozYGOTAvSclNzVG58UmDZiCA8ZhSD/rfQREh/4cWn5itiS11CUjHhGbhREhhZP
BRK/ZQu1YyQlgzaxF7QStUGrcXVbt6yFHKzstVc4Pl9MBOYiFKMC+odzlt1kmDvhpNpzR+dGvvYo
1CIG6by6/pHEd5nVeAryZTyDcUgoRQwf9MUwlRbiRBmMJvqWzN8bMTptmlH5kUficsCUmON0k7EY
9IBNrnE18lcYkBPxN0cAzFsiB6pW6h15GLaHCKu7Mb2ZsdRH3RgL/SXoZWDq4DhgVlhOI9stnN5m
dN3OmFB0DXT+XZaVN9riB4GxfjVmTGoTeJ+Lzvk/qHiufxuAt1klaL4/w0VC6Ea49lB1MC2YYMsJ
DUo33lyIumIarVGcSurGo7yZsg5tYZ3wiDiobULqhw3wK62+Tvb/IHWFYXqygMfTGlCUrYZ47urY
2pMItbn2D90bkNXR8/Fp9waIy1nriGCnux3mZPT7az/WcyDgKeteJkHX1K7Y/uXmZQaHj0bA9axn
T3W40JtvMrb39l4De+qi3guebbf/pVz5CqvIrsQa0ejVIe4ey22Os/clSHe6ZiHdQ8kUvsVkBucV
qMkjZiOGl/dIvs9QnEoOEcjxWdy90nU6veOs5u8qFU6CAZzh0uBlxt8keglCthdpxfQNPjcTUubQ
xoIbQaogBEjqsH66M+emt7+7zBDNMNKYyzZi6MoqGtuVRevo1PEdWp8aIW4zOQTMLjqBPpVOC0Ca
flpHslbphxTrHVdYspdNuTSMnrfrUL+ub3WhSlrUpKhZwInKpqP8JUDx/Jn9yZwdabjMfxNvp2f8
TzQoDxQXS5LOJ4ga9Hvq/tEFILNJcEUrcA4kkvwxt5LAa3ABs1Huc1hordZ2WteCIey0GxcnQKRK
6VugTSaWAISyUr0DSwxouL4Y4Ye5DgPibb3VYV8LDXfHLbD1Ng0dQOz2ap/dOHdLZ0bcLQbjNd3k
LoGkVve0ydJL7xpIxUVBoERT8gc1NoCinJFFfRFajLYzMcUQM4GIJWUlrdJUNw/SkRteU6GVf7eV
/oImrSfY+JPTpXslF3n50lLTiOQvz7dvY1Xxp9Gkq/Sx3Axlmy4kt3VxGvQaMiZ1U9PA23u8XadQ
hQbTonvkWLHrScplFNobtwmePDeBXlrs3JHvRLgxoQtFsKSrPj9d1myWOk90yZ2h/Oc5eYyrLVx4
ADAqfnon6g2PpZcFJDGO4xnpUfls2QHYv2SS6O2N79p3b3bM4EktABhkWSl/ZiZoKy3UZsol7gGe
eEWNd4mqHIWnE6PisKPe3J04GOx1Wu6FQWXjPQR8pypM4uFq8XduosXur0EQHNB38pvq5Wco8m0W
ExH67SmdiCTJXVQeAqzZcBoOfyMk2mixJJ77dobhQsdxZhjqW2dgmvZlfcuqJZHmeSsa5Ga4aOYh
PAnxFFEh6Js2U5rR3ifEMFd7+IWct1d82EHjYJndfeCbM0mG1zkX1nlLvOe9IC4QX8HPzHV8+3oi
WzgXqYVOrwJSxLLGxus02nKdbta/P1gb/DNFXMT8j/oBvY3nrb3eh4ODjFhjeAcr+cmfyB/it1LV
1+AzHLe5PVo1wDhGoK8G35pKbfAFsei9aTcxL7YM9Z+ODARxOk8YCVtrdyOOrSANZp7PQIL51hnd
z49FHmfeiLQLsu0Ihy/x/l3jo8vX8BqERxp8eBvgYl3X6sLMe8+nxtsnjBExUhuRC+CBs7TYOtjn
tp/tz6JEU9QfWbm6DjRAPPkAKCzZciYOrEqoRepJOj5cTzOLMDb0DHIpfATa8s88M9ZLJ/5SBDId
IMa80prZP9pVVjm/ZonNC2Yol6wao22LU0zIYcfAFB0e9T5Dk0mBuJmdSW67hy2yU8TLj1eT3two
chk/EFCUR2QcC2hW9Xo8X+/s3NqiOgTNx9YmpS76k2WLFLA+mREthuwiY1BKvwgBYagNqgPqYdwj
mp7VBUU+AGsFIzc7pEWUWaEce99lllUxQ740saa1ZXQfXvHtLH1SSSRno09fqa/TeqPJcoo3SwYM
eOg1/qktP1pALe1O/pWmlo6o+BenUvK0XVDPLXGsLQje7QWU99djNOkop48ydBZQ8MOYH/dXalHd
foaNh1et83sBOrTxYL/kOAHKjGIjXW8dCdsVczGTsLu3gXxsxZ9bOTcReKgL3Y6uneVq9M+tRUKJ
GgduX501KGLAS78F0gXqDp8N1fACo8rcLPa2S8J0YTbe8D49WSAGFYwUvU9zv4NUpDQPIoPT14yA
45riwIgFfHz4iY7JiiwmitdYxIbRUi73I6+LJX8TdfXcY5pO7LWNLfIjJ2tOGNYg/4h+X7dKf/7i
yFXNrRa0fKuNdVH5+DMEYoN9Ko+AU+PlImTEW4pLSnvg9bBH5smqEFeSwngO5lNm9Ieva1rx/CIR
pszBtf8gZiBGvOLjFCUrog7NKjJhBjniZuf4ua/fxwJEXMZmCjAICZXwkNe0mj+cVbE3ZEeiPOYP
r6mZVhAxYPWh9UY/83S6wwPNV5M6sNCCyb00DmH+77mDE0Lw03t2RYdLSvyBFvOSrLBt05A7a5TE
0ashAUIMrKW6Nl1xCa3XFNRnV8o+ay/o3E5PD4QnH0dIzLNDuz61Nhkkv2yJLAQxlcs/JjsluQ38
iFWmznt+927rxor04AO4PQZtsLIYJqN/WI7Tp1w3QW7xcGXAEsF6Vvf4Nbnfi8zPWuQ79JTAJ5L3
uDs+Y7mjI4TgiaBOuVX6rdxiATzR2a0s+cOvvZem373xg5f6uEL8KfVOwDx249prnkThKkfgEXTO
1nFahENR9zmCondQa4cBjkg4Hw262dEvZ80mUQ/ECfLDLGVgotzKq8uN5Z3oEUOt61hfItFo5G57
Mbhd1wpunKPB6F84313XEejL+NjMyeLVrWlVgbeQUXE0qUlNGzdgnj/e4DBF1Gogk/foT181ouHM
JgDgga+v0B2JEKwJPeHjlLca/Bk6r9A4P4+Xf8UYV8nlS9MH0AmD9Cmh+BiqmobeV4gy1azBjnV5
nV6wztuOduNCqtSBfSFTsXnYGaKkA7TfpNX6qhHCd+/cd/eqiduAFW2jp3kEy1YTOXyYSzXeLdNm
+CF+d1vBo3B7ZS+bt5gVjTODN77IegNigGRyiy9VDM4bPjYQUFGAdv9DBcFHmfrcgACi9/JMHEHg
qwsrbblOrR4aTUagNK4dYK/xXmckhCLoRRQ9E6efr8cvkDZ9v2i+Z0K4a5+ukam+E2rdZkzqxLrO
jX+O2NfU9S8rN7RejH4Jc4n+QtqLejmsZ3JvIVwJbUWbuwXuwE43BwWp/kKO08cENJoH/u/CPUE5
99edzsON5s1Wa3wRNrnQwYiM6hplz5UiaQh3G5cTpBirLLq9LEJndoFOZWMc2UZxprAP7sCClci8
ZQ/1X2plhS8TWzkvw+okbvvPzhcmVuM+FYzyVMxPXuY19CiRHwcCe2puJSP9gosE5Deqk+lU3tdx
eE81JeX7sYyFWvwqDXIrC4ZIqsObHJi2es/pMHTm63b9SQC3LK4NInHAXRY9P3NUCuvHOsmRvlqY
47b++5ErXtxwdAxBJZKY6vsSYVh5aZape6cYY77cXtdDpTc7PY1e5eg61gUYWsxmCEfFtMvC3YbN
xQhK9H2K6ETPAYzEP3+/xFl4CBCi2c9eQDfNzUeG5xv5dM6YjhEZS3caoN8ZIFgM4FXoTXICkWb8
MibIOz2WWDBpV9KNhBMGhQThAtNHiuzCQfdjlel06gvltGHaeXfm2Ov/xrlQe4XRn2e3nji2wevz
EbzbaCqJ6Nya5N/9GKPeOUeN2Bs286xNEwOB+F7KNILj0DL3/qbn02g/pkRliQ8BrOtIpincWrh0
36XJSowaxUVp04lDr3YFjIR5nx1ei9C3cU6zbW2DePCsTwxZHF5KgHYnwii4vjEia7Uk+UPKMccz
6hVV1FTVLDS5Z2I0robV9yxxxJamuGbEfTU3tEAC92o7OrPiEtbnBup/sYqZwTTwfSgBKlYdXt/K
b4vF4Kn0cAYLly7WN0sc3DAugtSlhJltMNlf6z4ioHyue512kiKmX1rUcIDpsWIY6njd9D2h93bo
ng8bqdrLNwXjCF7xAoxSeLnWxki87DgXrRaBbdSqMN/ErXrjdP4xzI7Gp7Wd3mZPVlm8KOiEF9KM
Xi5rbjiPLDfaYnmRA5MMma2V68OwWrPG7+aerR7kPQFEpJFDpLoiTSiPX7RyPNd34slNrwyz2vW7
75XA0TTyXkDtYnOCbSFZ9YsF/JYw94SfEiMZPt3Lnd1GRsByMfo4XAhb4fqP7mjYJLSSuXT86pR6
/usyFI+aedH+RB8CTlT9QgtWWSMGQJy9Wzk2ZDEpCkfTLA8ZEp1Z+tTqV7CFBbtmvayl6aaq5fHk
/PUOqG5XU/E7CNoO591ySAD7lfl7CA9O2qjB3W6O94jNR1PKi8z1wc590Aisy7xCSB4mU3HmIXDs
MYgdtg7hB7bpoAGoX6UZp4tJffJuxBPsUu+J7LwPeGq80WDwQscJoIbUpS1Ox2kXVMRTvNrWhhnq
uEVwSwz7jy3uTIt2AteU99C2E92q+G6BxTAKQxJvsoxwdw7UGk/YteJ3lYlbaXdJdiWGzb8Dipw2
tFcP6+pcSzyuiJq3gywGYP0OCp4tgnDpGGU1mlbiMDCH4MsDS3gPC7F8tF2GrStBEwUtB6T5GxBJ
cVgIaMnm19oyNuCtdjS5mtpuhVvFxLXgqv4XsjCKh8Xond7EjdlyCCrzfCTuHjV76xnm+oo2evmu
zTgkr/0G2U+waGmdDp+pRD0x+b4WIwcgn8PL7qXR8hB2ac5KNQgAoHKIwVzbhQ1vk2tDZiyDKQnz
KRXovHrw20vVsq4PRYmqDjU4ZpGSs9t5Q4u5G8/ggGltt1slNQ02muawI10fODVAfPyu7s0iplzJ
AZf6O+6Iaw3OWif0/BOK91ZMobPgrsw0nvj591MNAWBA0lnW9BQlhsWl//s77ZZenSy3jevS/eiA
Qsq1UKVjhtxeNTH9JOc8TjkcoKsZUws53GFgtfQFkcRT6z4aJPKADHo5TFssGyNKGFlBiqGMi4tk
fVJ15eQVj77wUcxjgvVUyNwjzs44GRnUUocQ3MWkO9eeMqK+Zvct2uvPu+ebqYEhKzDTZm9IkYpT
3Vps6BBErGegsMIpVGuzRLgdybdt08Y+/9jyvpdrizve2rFvBql32WLTGRzIFW7+DKOC+U6/gQv6
zLtpN6b4RGsHjUeO6Y08I95SxZTlXput3Tenu/wsbzGhklhqy7+pGz+0T3J06kJSQ118aMTBGTgg
5yFF/q2NwCKmBDo36ctPTc8wk7jg+bliHOsyA3dZlSI1jf1N0cTwqLyIOfofPSqkVegb2R5yKcKU
p1ZbuSU1BsWI0tt26RLLz7wMHsNspuMrsjLJYYElKCIL0sbZw/v+5YGiPHWmH/AIdgAQ7YmD4oFn
VDX6Sl/0b2NIlnyLqnEQTzxqt+2bwn+wdmpZxe9jSv/qIE+SzjELCgxmwj7OS20My/R/IhM0PBWr
UucUTvjOCeU4biYC1M/h0O0tDbj3UI3v5NzfiVSAZgdAh5PiazkBG9QYgXIsYT69zQxey6SGvlLY
zt3sSzfVlSUvAI7bozxF1Pf/gsAte0T9pRoHTRJRIKvS2EBL8TC2rBUGGfftDas5gKItvY9odKZf
+F54xpkKI01QC07y/nVRsLXsiSLPK9QRKvVpHlwdTx0UlArqNcqFG6zUa70W4i9DhR+uwNky0fXs
q55fid+vI9MF9JY2JwoCisvVwP8RgCVwUV0m5s2dvNW9ZWUWoMjozd/y6DYxSOLUmqXw/Ev4Jyj3
ijioj5lgx4l/s0XEQxidB2Ad9hbdvQtnzgampXBqSjgh2f+zNaaMXVjQ4BokFIJtF+HhYSQ6kR0g
LqdgUoWNMZC2f7cRKavzOK2YDZaMI9rfMvLLrdc2q1IRREC6G79GcG9diW93f0DEIYS1AQ5dBPWA
3GetAqZbMEYrUwettqTPjwSVN3+GbZ0K3gv5YDrx2pWcu+6OIOyev9QppoJgFyJOq7p6D8dl68fq
SDrNUvKaDsCI3pvQAt88wj1d8WMnEzu6R6mE23KcmCVruwl9cT+PHDyI9Uea1q0qTllzPqxAwh2+
25b9Ip4ybbznB/SibimRaOuJG2V11eVPllnAI55+QEKo6bK+P/GU1vsA18O/m5Ry58/JHG/Knrp+
qKioWVjtnF0PH1jJMgCVSJr0jC3rn4JNdlIx00hwyoYpTDdjNXqNfgXKCR/xu72EL0Fr786PWxQV
MTC2RPD523HD6gLZ9AoLXmFplBGIceL9aggyJBk1XkYvVk2tSOapp0t9PizzoSyI9GKZLnUNoZZg
/lOdxvcq/97U3UBqYlyzTV6Wfvxaxfm4cmHlXrgV4SI7cgCr/+8GYUMIDVPy9o/6ppnJF6yfJsdo
62KnYy6wBbFbDCBmpO0BjRvITP2fusG77iwrRbbKMr+zJG7Tt3PbQJfRT+itI7fAoMsbNGfQ98sJ
RgVAmyrJWComQKYlzrEPRvBpm03AS6xFdKOTxstyN/NcjMfku6I4druJC0vcNfyZrxvkd1B0lPpH
k+9SYtmeB+Ntz//rYSM89FMVQb9iPv1RGCxEugj9RHDJ64JpHFB1r48iwY6QnrfLcoOENxSZlo2N
XR4QJtTbzMoihfiJwT0jDQpPBTrb+WMYRNWgrPG5FxEcZ7catED3Wr5fOMIchvgXIySJut1JdrDP
ndV/2biJcUZEs94p+EE97SxgrzlvelWouzGyfQpseY9ArZJtq/OJDuo3ANuT4AJwZVW0b1o48u/8
iv+r9rpvbsrrP36uY/NfJy4l7++r+0jAOPrr/tROEsvcjFe6BH0SicUhNDpbTsLKgAkdYWBSsVV6
SRFetLY9eGeUksvpetkvANQHVL7tpMEhhenksmFNWsw/8sNFmchZxnXSihITZW7uKh5pA3MBq786
sRVc1M4qSXhBvXprdlwkCHyCrr3P/MsHPlNP42VU9Z2G1Y1Hwzjc3nKue5l3FbAfBtsfl/DLNtbh
CPheH1KHCndanokwpXE/NmfDWrAy6a6Uxfqh0S8JXEm0MWSuhJLIw33p27390Dgkk1c8DaR7mAg2
5dWQYuptcdrXqAe0TNG1Mnngnk5SMSuKLfkFtqHSocEV6N5VRkzlU7DAKcMJYkw+2PB+a0k4JrVT
PdMd+P8Pqqsn4duUEbGdbqOILcJF7zzGG4vhPGo07qqnS5k5CMk1uX19VKHlKqPYDq1irQXM2ZG0
hFNxNx51GH6EkyD19K6QrvVFs/mbZ+PWgG6OQDhCESU5BQKa7wu9JYfuyPFO0f0y1dJ4RI9ggeDy
5VbfSbEFXtQUBiIZqpBHm93Aolk/iIsaEZtOwAkY5aq8thVoyBnOfqi48H5Qhbb4+WKsWgrQzRtL
CXzA5nfZ6ojSN329NgbS99Of4xriECWJ3abCl2FVsWeKYxWwZwQ6vigE1V+06nKOLYxrynpOXuJJ
9aostnmhREfL6wDKHP3ygcXA4feZ+qfg5zdsxIpW/Avjfgrx/6F0YwLJ5SCW0EGQamcRAE4+DMTs
p8g0DopxgEhYX1bxPRs4SdDZaZc7fsT9s9oiw1a9coiv122U7OJMPFiiFa2ZiKfbe2y8Oo2BBRlY
lTbS9xBZCqh9xmR2ILWpg+ahX/BrfSW1NTKTSnLTFrUxJP8EmpdsuWDNcFXi1bh90DVDrki6/hDP
jrsB0syaG5d/QL9ogUiwl2E5tBdTUsHrgoFgwnvdvE08vKRE6NTm76UMZ7n9u8x6M0ZU9JDGPY0I
EL6zuCK7HYYsuIvRDVAaFwGZbM/TZEbyop+8JDIVom/t3SQNr1HAk0/VkIOAuhVO2HhO8Huv8l/6
mUK2n18+bjVdNoBEpXGNyMjLVlHFK+bOufvlYMiMgjbUjrm1lQrmY7TiYyQ0Tc642EbSTV+ZpRyx
9+8wNor/9pFiZh6jLY67Ybri3Ugf3tWNaFKhHY23Z6oTcpySmPalb34edTMrZv4QQM3W4MVCVtcj
9UWP3ZgRS1o8vXsQKs/dLY8WDK4RJ/MpVH0iJZrXOnIPy4Vnk53BBDcW0bI3T0WAaBKIzHePmV4J
gHvvXRJ8XYM1tzwm8W/p6BGNG7m5ufDC1oGBKxGutH8z7btpgAziXZ9YKpiSXKWMfaom6SwoTYNJ
5TpfqaQWEP67cjtwDtAvJXRmUBI9dGx6Or8712hVL4EUSOSxpkDaO/yCMjiB/T9XY5kgioEVu/4f
YISHgUOVcpFf0kAceBmx3XCE+QYc7Nxxeu0PHMF9VXOdLfCA4E05IMoGsI+siB7bTeH+WdSiltzC
YHuel48IhwH3WkxQqcgw2cCCmSp7SXPJ32bR4aWrqPqqr+SFBr+EEM5CG0DddxuCttJcDqnQwirl
PJbK69DBGMoAdBmqov4HKxtzFaOdspy+XU0MlAvLo7z/HQ8tRPbSHp1CtjtksMiUj5d9vTdn7CnD
NMKhZ6dN3poiRhXKqpdDk8ZATFKbD7DpaJOPmuKSe27rbPBGMxb0X4BMKsD1EyS8UDqk/K3qLo2Q
VrrDMCphQzSoJofTkjBh62hNSUglrq/li5RV9RsV0nCktYbi/H/4oUOQVH5soIKmMMZUQicGiYYh
epT21FgZcExOSpbst8Fnsguz7HFjjWFPnSo5h29hBlBqZcf4qz4A6AyMEyNIKSdUKwXyl7k2W0Pr
BnSwj7S9CAikHFPa+7EAdm75BZqJFlLHScSnQb2/4zTr/ar+cZho7ooXKrycUX2EHK7Fg+CC6WtU
ba0HoO4Z0SGNT6m91ZfbRdmDTSJW4l0vuSCQXtu7yaSw035iPQU2n9mm++ImwHO+z33G+zYcXFZN
Yt66fEmxIvhXqaqv15DZUSb8KGghlq5TBml391bnEnMUevFlcDkUxtbzmwCmoOkGW4iXbDtHQFP9
1Fa+oPUsls74vSWnXwibA/jzRnYUzNrt4umaAi6C3U/QRb1MUl7K40w0feKHoKl1xhdGKgnXBSDQ
2nqYZjdg/mmT81PYX8U8OjxcQ9CsnPTE+hz4bYz0PkBij8AaxRU7wfSJNmoAZ5xsp6e4mPiS+EZ3
gzwCb2YHgqNT+vEbpSoCEPLoS5kxP+sngAiIbZ97ST2RulNRZJUreXFLMoQHjhYggOrEEyEky5Jf
7sApacIBffRoM0cCmSoe43jZOIq3USiZbTcTCvNGuwG8xkwxTbxLbybjzEq818fckwM/QY6cEHN1
8irmEXKhk/MKCg86yMxbnB//EoHnu1kDIIxFVcWbDTW7jz7FB4sMZKiVmqiNftN4EcZKrIPO8cvK
otubu61QOxUSbWst7dZixmanl+eOxodt3BPxjLIKYRijRWQPro4Cx3kgby7nn6e3iXKGhf/a4MAE
4aui7sKqBS31HdoH3QdJpxe5iyDdBYkkk5sKTQxFgjXpEuqu4JGKAEOoO0GL5JQ+aY2AvVcJ+1ij
vTMBKuSsjdSO7SIHOFa3LAZj6jXR/LPjjkisyqA9EiEvjSlkipcZqnE3GLk/j8zhXoUS8T2tUAgL
XnGs5quX5Dz4W5fGReJFXmrG3o+w+XPOTREUbvtijEIQTyvajkWEqPeb5HzNtb8D59V/MJdVgocF
BYHTWSW7FH+ixaeULVWFSCw4tFtBxhz5WPxsSlsk4bsQxmoPmCX8NpcEGidyPFP+7sClrLEDP+jt
uR56z2af8pMqPiu9cLDPPlV58eXEByMybTUla/kFJ9PGEPWpOLRKGEkRZoXlk15joXqRM6qXVL3z
1yTVv+52bLucq5iS5tg3jXkzxvKEHEjuBFxoJpGToecAKX01BN6DBbAJU3w+rYMf3/LwmkW07Kbw
eNbxV+Szfqml6wFwh5cpAN8YrxvJdrHMS5d0PSEY15GnY6FUq2uRr3Ho8tK/q1Hno4BmPd/5qFGN
mjkX64LtdPSHb3V/hcSmgNZSIbp2mEsZc7qlV3Ri7oBq6l7/m3Y8BhwHXFptLC/3K6y1YZgpbx+c
2DcvI4U0i1Cc7TCgeAiJgGZh5ZeI7rv2IJuXOXEw9wxzaSgFQGmoiSpc8FCoJ7WtOavT2Rs0JX6f
iuGjoieF6pll4AEFXrPptZyHxULbjaEgnSMPjJnysHzbP0IqA1FClkBmRR4Riza69XnYXu7kIj7e
LTG7UroKYg74nAYTzzK0SxcROoiUKCunsa6B1evk4cyBAcwhCheyqIsK0/Fag4HiNFJbYatD2lQx
bLKVwFX/utEFz2B2DchgrhnO1IKSDeMF5T4udU6iDzCmaBmHbR7MiE+Orxvd+p0YVvEoUe2Dn7P0
zHLhtfGtudR5J8uQdnJkS/qxNwKM5+vEO5HIff2RaiLcbqxZ7lAv87eXidhq1zEXw51gIupWuYZ0
+Fpu5IEYpAYLGbzH1ETBCWuu41/Dj/tZMmhlGKxck7NsLDaCW902OCu7wBKhs2zb4/PK+gycm6tg
zSjYKIFmHbx7XM9xBuTqNh0zqJZh0+w6L+lLBseN/tJox4sl4B2oxzi9cwE6Ef+CGvfYDsQsJ+W6
t035HsPwlfEA8wBJAFLRGc8Wnvmk8A7j0FSnYNMUyNkP599E/8vTOXD28ZDKzablIcKrx+4HltF6
i6Tj60VpwPL0/EVlYSEFkJC59Ohk/75aGY8wN4oLr+FgWrrJjrT2ZaSZApbLEdjFC0V4mdp8L0Ro
rKhZztZZKAZeGrvp4RUVl9HchxH7pvKk0rIyO3YyCNqW5ss1iwcETuJqdrkiyApbK8dLVfnY/0j+
5kKXdGpRqo2p/DZTL4GOLOICOsanSNfoIna8o5C+OFN2WqyoFJG/+RZOWYKytHCc+ywqUrLQBzKG
xLnYvuCwlveG/MIslldih+RgWJu+BZU4GRBIYJh0Em3pMEgqAZ7KnQiiG3JOxfRIZiCSAVJvB4KR
EE0oJMs9t4L4ZOJQ9DBcVc9lRlsGY70m3fi0+zwRuD23NFOQ9CJIoPYXe4ncnsIDC6U8dB6QGmBb
lF0+E67Co7sMJhlaxGiQB/qWyGfpHXGyG3GBGj4WMF/6GmagObz89k8mRHaMy6hkU4oYb504bcGU
9oGi93Tvt/ovzXa5ruqm4/ThcQWh23T7BiJqfxp9lFdTGiNkPmsrhzwC3uAPwySiO52v4RIMJZLO
ODjjsFRUVGeXhxg2MAJY/yBk8Rdg+1qYz6hRD3XlfygWe0XoDuicFwl4apJ+/pA1ZzmJLwMrzL0T
vE/srxE1e66blkGljtVWReui1pfS7AWE5wi36QcAkXBa5Hpvt8U4rVtplc2afJAmHOAqD+TTm6ne
Yv0RgKPm5epGCvKcdTJAag85JBvgHU7eVlAvy7DZFW2omrpbRXY4+Li/k73czyCabGNTO8Eg+LJC
YKpUJ6ckc98EU56sbhVrtMAfXXL5lxfqJqzlVUQc6CKkzQsPWILrJpdiUfUFvjHDLbekuJyPcfAl
UAnouC0eBVBfu+sehvro8Qjo3GOdqbfqYmd1kX7slUwF/rv1tj0sybocf54d82mW5RXgPRVh8tnI
SRfravwQF/sleW+fENnhx12syRAtu+EhI0JEnHnWvfh/SxAmYefdIYvr6KOjMlwsxDeOHYqMMH/t
TyMmodL4HIS7yBJ7b0NV5cYLtznGXlaBvU/2L3LfPasRCuHzNyWoMTpT/vufu8HswdnqbIOvohFe
Et5gGoIccB6YbZlMqmhCTPXVecrN7A1p4mq3kK4pw5y6egGXz8nk1VahK4/8j6NtAS2rV595J2lg
HXkEZoMuZrEXqOCEyQRK+As0x+g6DsdVkuRcFtME0cnLOihxhQ/dBw+TxwPvMlRfyZSZNMga1Toc
6BMkz24TeazMXJXsIe/n3IKGC0Nofjik/OJi+ONrXPDTNImCrkjVTnUzyl1P8KAzgEqcsha/xFHK
2kuxTHAs5Wsg51uSQsFvLJt+ZNIsTjRHb7Cd2daZ7zt8VQXzFfC5XVHN2svcsmZZz0UgW5jvcqKW
86x5OYpVMozW6Vqyleugg1hC40E/yQfYYLLXqX7IIntfq3wLTCi2n8XhIHdDYQahWi1KKzbL/7/7
5GWTf2ZT38MY/f2OjEMN6KNDDYPn1dBvxZ2C8o0opq6W4QU11nSTdgHoj3YePeeMeYyhSv9SZZ6D
3P/pV++7BGj8khDOX+FLSNAMmnkeWNHwJP9xJyBukSGgaj/Rqfv4v6hp78nDqtLeyIY0Oac7ltZz
DMt64LBgn/qzqe6qi/0Ts/Smet0fKBPoLoBz1NHCiV3uXxZUxx9QK82+qoHolh3PkVrQBaA2oD4g
MTPsGw2lLT9dXO6bX8hyPO0/KZU2e3Rx2CVAlnfP8FVuq3IoMVsqBWFmHS085Utj+LXoPlCCK0qC
EEcHJBaUEEF8t4Xn6ufHg50H9VtCj7V+UosBC9+Ka94TPCYYIuy9K1w7jpmuova02DC0Dr8tJOC1
XwWbsfrfhPtsHT/veDxRwfBPUSBH6dJv7X8ymFe2YiPJNRD0dO43jqbgYTMBuL8vqHEnkIOgoM/Y
BcSehvtUMLcAUb76wZ/7qo1DyH6n6K8+7b7wfkk17iONcwSOdPIk6/9nbqkDgiLDSj2IoK1hG/WP
KaziXGPn1jpiS21S+4hfwL8XpHUupQwXsSGyliHogDOwLJFPg2xLhf5sbW/J+lCN92lpz/0FJkt6
866c9ZOGjUWf1wCzye1DrDSGx3XZhWuYwtLx/7a9sTIYY03abOqgkcJPgAzHnCgCeKfGAIAmJv5V
2d9BbecrmIMznVGyf4ycGDk18Dv/rkLyf2A3LIrXU40fMcZRpIlIKCr8AERVHfLPxvNTYiU8CTID
LaBjGexgPsEx4xZPOF8ofEWVw0A3SxWcOW4zyig6gwWkUufUi/i7oXzEc5BV5e4irHX2ey+p3Liv
SHOl0Bq/3O4a21XLShSizqRHkqdXAH61Y2jfbNeYa9WZl0xLN8YfI9KPNC06hl+0vWm5HQZBjPfj
GuaLRMaqiAW1hHqXshOdeoaRLWz4lucm+Q22k2mrjaFrVyHNI/rmno7T0J+jzOg/+l0qWq7JvrJH
Tab/VZqhW7R2ZulKZcrZp9aeBSM8E+z8Ewg4nen9Z+9GYZyNbAR7R9KDMP8PKzXNVR1AblQKitLP
OyZ4FLmMJJ3qUaanppNbHSnCVELr87urT2A+9Hbz3ibD2dR+rjD/rWdu31HCObxUC5XJq4s8o4hS
d/5PzEtwwsh3rAIBisEebJfwfpsQYg4RE+UDR8b48nCw5sMy/hlf+huxfYWiMpW1p68BNu11n340
LB3NzvKOhsi7Z7ai6PjeGr9r6GT25BzFrNTJifSJnd+0446owzsTEtQClP6HpU67BWxPj6Jvc6je
QdG6JSoblsJOEAt24YH/uvo8b0R2RqAomghcWW/wKimR8VnNpQF8DyKX1LsSeYU5qGSRrF7X18Iq
lxzwMz9+2Wl2vkxujf90F10bg2WzbgA4LEVDDfR1G6dX0iHOd9UUT8b/bBuest3uWEAvkEq6wY5H
Kev+eoVy8vHZVvWyJ4elVWMePMzwtQYpe6VkMGGfoyJalUyIbgz5poIADYKtOZbg5Y3fExYAapo0
YMrjHTQghVxZCS0bLrYSi9sJhPH2wNSrs26PuLBjEdeFslVqX4Vk+19d7jYalHeE6TXuVuJwmIjH
liPUvb3+YiQ93Wzl6GQE7P9FF+HAzAFUCPJvrz2QbrwKNuoEZHP6YHz/XKCjaulMHi67YgT/iMiP
tSYDvaw2DqMoJUyrQewcnAzosKzAqgVXv20Z++dBXAGE/nWJZMckHEiZiRep8VKmEweJGay9VlL5
LOVDUBpXSevFm+2OC2djMAHkSr2y8dRgmx2IQHg+8oq4LtT3UgkDMflwlLYCXevQ6Mn6RSnV3+2M
BxUKlqJ2RSDhc90eIaodbfzEwubkqDkXSmsKHtYXtrJ9rQJ+sHU54RHClFOIOP2+c2Jz9Y3QcgQe
5LAICo2GK/IbgRy2MgbAf0ndT/U8OUHOXeMGoZdHm176VHYk1CVu848oOju6JbYoyeIPXFziHl2b
vtqsCcHTHExk+/xAONRoN7IrRRRaPeD2G2xKhKBU+L1/MWtL2RBIJzXz0cAx8m0RDVEtI1NXM89O
4a0mWUfX/ItYWK+QNCcGad3Zq8OyaW8VhBz5tJOBlq+6Utx18huBn0/houUvUDcsOBh5tJG1kdWL
H0b/jCxLkXxDSfBPZ9cLp2fj75BjE/VEYa9g4BTYcaTXvdrKeveK0dGcMDUrLUDqlbDVI8ap1UEL
6e0RzR3X5QMG+ERhe62i/URErK0p1a0++++RI26sccTAzMr4bKU5OaVMnAEsGZsgG9Jra43ySnex
TGi6Ara+H4o3lnrtKjdsj615C/v8vg3ylGLHoW2qoG9b9MKp3TZdf+frYlDvj9EKcJZKIbp+LTQw
9MmdHQoX7jlSu5mZhdYj24wRO/mmAUrL7937gxXL3ximRz8GlUZjLzBeNjehaYVDoCnMcgObbJI0
2j4Q93q20dOFOPoaFS1B84Rvx5ftGv/Ahgfe++NBTDMM6YWe+0Dr5epm0AGAIzCfvHc46G2MOqS/
PCNYpp7m64nRDQms9oECSqMGPlkudCEOBJUOU5eFOxdNpEpwQNrz4MW3H4BGldZ5LbmyNJ+4430Z
ywOW3XCWObloIg71PWnT88xXs4p0qpTxdddIMmrydY5e4fvlKP/TdFsmw+/RFQRVSBb/OaME82lp
fytE+wpeJ3h/BX/3F6MuweshDMIMJkvcgJUjctLQ01KVPns8NbQisTicQfGMS8wUnomFkYFhFt/d
KhZ1N/zHRgCSuxK7G8TT8tDYJELPlggr5W5fWk26UtehhtJyzTMYTZUQpqk8aJ332jkV/iofXzFv
WnJLaovsjm4L0ZMHvHr2M6us5bLiUtYflnmrCCynYGZkY3b8WdsPvKPj7G8Zttp8Z+B8L8xPiO/1
UU1bTi98fMkP+m+8QgeX6q+77RC8yRv9rI9huWRjxMkH2TPjIZTAXVdyGn5yjS/rijWColnkMn04
/Hr5R5B+nURVWogc1ag6pfq9sGDY9xmWAWSIWB522f9lkGSwTiltZwLVmTp/RXDS3H13+vnkbhXq
6kejvNM3xPLuLltNBXfbyQIJ2dlIrLEDKWqSn1S7UgpFJmttrrJJ3yIg0K7I6G7fEo8DjBigSa85
VMqBDz3jIgfWgSKkE08+H2DextAR13oQ5rHAu3mbIKeEVQN6HCVXPpcGsGVp/5GWJ4z2YZi1DuxK
u2tKBBLBox41kk3NZDCm8oGM7ffmQyLYArwr2K1X7QNSl2ypGjxceahdEs+QYWUCbYOXpA7hiEkl
cZcJfQ4AaI0qLx7fclt/WqH9f0TwDzVqfdceDJoRsr/5XxHeOYWwtspehoD8q8DAZFQGuu0ajFqE
2dCB/nAG3RPMZuN5ihY839RiyTe5lwIUzsEoNX4u1Y+HBDJLrSqJzFphZkafBcWewDTGtB+WiB6L
5i91M806PNhQ7ivez/jSEVS9LceJlfb/VMQHPQW4Ak61zq6UYhBd6TAdGGhggqw0LExK8BbZ3bJi
qq4BDUaYBwdxgCms6VBwglvMohhcbbB1q0fbH7I2H0yO44HXGlfO6rMKaXw7RqC8V8Drtc2ijlVO
h/I2sghDHZCAye2rzO3zdEPi4XulzhZIqCzPQnynWYgtjKy1iY9m6koFVb89AMLQU9ZJgKafrg5u
4GNnntSRqBVwMS6xkDkD2lF8rIqM4iGH57KH5hl8uIAyr9pCXOoX21Yo6Y/ZRk0pAuYf0vETUBkA
tbq9b8P8yOilbBtZqg0VuVSJVZ+bYcEP7JNK9EYwpOaOPsKKcVDRme5KMBOrdt45scheu3aaRS/U
D0A3vbsPlbss/GjRQgZwhD4X/k1KKYALPR6ZdOYZu5Zq9IyqDwns1gvHCGHs3j/0u1ubjALGEvkX
HuQD5MxtnElZJbG4XM4QXKCXeFyDkqHGaiYFoDwoK2nb3IdrSFUCgG7Ld3fJ5jbH5o5Lf9WFiB95
hwu/K2Rds6VBsk/PixwdNCf9s5M6Q6Zd46EgoGz39q5J3ogq/ZTPHw2/lSy7NX5L1zF5brvkwnhO
5MarVGkknHMRf2bqHCEsfhY1bSYa1gajRavYwDHbAmhHE5eVal9RDLh39dtxaNXlKKTVPVVBBJBA
6T0JiikS5KdTL9iDucEud9b6J/EqlzdCEsQNYa5uAxpo2w8XO9QCsfUU+cosM9ZqNewePl+1vqR1
QgydqJPq2xu+wvWU1DZyYM9CU4YpQ81PGEX+AgcSA9Si0rZFeMzMHEPMawnWA5rz4TkXYaDwdSBZ
UcNfMr7BRWaZ4aELgdP/PRwZedmuDr1f21zKw0aqQ4+peZmNFmLRaCTRwuPUB86oqamQw6YXX6ba
0eO/x5t0nF7AebDYD1YFpc9kSOnal46BxxQ9cwG/NVg+0FHDcDKA3TYqEMPZIst1JV49Wzc3f1Y3
RHyjRNec0zKIYzBVFeVx5sHkRj3oQVkcxy5mD+4HAOIzlil4En26j6d0DL8E5HPcwISRsMi3JZO+
Cr1DVRaTkNZFUUGw5GF1py+D5YpCY3Rt640zghTusD2B/vshrU8ZZLQCmMQNMCnyPUwdD60f+D9e
kscKur7LWurcKcYrIiM8Rkb9X4cYSFAXCZ+yh4djHHk3rZ3D33K7mZ1OiLEpHH1aQrtp9N7uTg7W
C6YnCvGeDL4if1vOQxSmYv5HOzFPEsYTZVHM2kwLv4wqVsChkYdoIlDV8OJNTKIMXvsvIyNmo8Kz
/6bAN0maXoLI74LqFINIO9b6A4Z69J6DaRmkeWquM7w9ftqQpF4f7jY5fNPwBKF+LyZ6Lc4ccOTS
SQoUNUIt9qPNviNh6bxrnes75W2TOxfeIkT1lcKl19NX8UIwLf5EBODCDqR6YA4YNz078EmHQ7wR
Ssy7IRQTdTbSy/20cn473uwnUYnqYlv8UIckiNfD5P3J7Tq814xwDt9WYZPqd+cjNuCnAEkii8iK
plNN2oNjsusMRI3cABBL6jxxbyWhAf+pm5X9RSontXchgK9ibd13Vgkv7pSjFCamheHl2fBIuGCp
3f4ai7Oydv4Grl4ThLnKIydJkEU02SK4J6MzAi9ngqkc/WS4gK00fO0PVQPpoii7NkrsnMfrXCtJ
6eC1zt3mZ5AFqZJXhJlf2KMGoKgOTGHxtdbp9LitIriEHMy1AszAd/u2vMmjyZz8ovEax8V/Lcjh
qKEL9e1VVgMlOvNdcOHwzWMcmOuM8MTSoQK3faOCoH9i24y98fMk3nU5apiaaAgf8wAwpWVkVymV
HP+qb9I6OCrI54mOCsIkkDuQKb4FriXzpUBEqQ07sth6cBQZklLLavkF0g2HJUPAhcHy8tUP8O8K
sR6kItyqEXHcrO7sBdJn00AxoqNKZFSRUUnPKZBI0VpSy7aWY6UEcxCZyzI2PZ8RJYkTtf79fQa5
AYJhSEAWD/kg4Nno3WylzRzEcunm6zm+THcFrH6/Wu0mkoduABflLkS8oqlL55/+PJcKL9XLFSKw
tRRs8NXro/Zpv5C/093QgzZX4tFEz/LXNCIg/QeMeC5wH7re1rLDn5v20zrF7RtlqpYwZu5ysgTv
rINBBeWMdi2bjvDTZZoaI1zIJNkOr0PjDuxoU3zlbrV+AFaVmIz9UEFp2Qz8vcnU+nYH+zKJdwcu
VsqPeaQKZDjH1KL8ojpfLrKvcYK17muk9uD/vWrd6xPTuEOEPWTmdTZIwtUHvpdRI4OzKIw7KivA
B6GZqX93Y9fVJOreOoyLtAfnWiNQ4G+totvHId8AWRda7bm0EFkQXTeeSF4bas4HaEukOxj1KV3r
KB3TYiA1WVyTxsDw+UDKoT2h3ykFt/hov/g8On2NQIFm7zy1VWwYH0b+fwDhpFQcUkzAGHN7gczH
gvVIP8kjsPAuAKUfg3Ko3VK1/I9oGDsXbYekXLWMy9f5Ic4DNBNZ8ONYpoZ1pLaSHEqvHPuqxfaE
+q66kbNcvp3XI8pSjbdnwv/f/P9tAI05AnqVvolaXmKJO0uNJGg0EGmUHWZ0LnqWVlnVLk+NHPOb
peON57PW77+ZJIhcuCWUdxKFvVp6XJNDPP8eeFRFevwZWvIuGq37fvaWyU7eMLdv3TN1vEBKlfPg
8PUDBXYOQKiAIfLmLy2RjrQ5RDWKLchjsbqTRd5PuR5q70EVHMH3ljcrNCmVyB3bVpfUnbhh3WIW
3IJknC0b2Ns+EIQpQnWjNLhQ3gjV8GRMUnO4cvFebx29hmnD1CR0qp6XR8CbmONUe3fRPMI8rFh2
f/0pRMnH7dCGH4dMY3MU2uJP2rjD3oTn1V7NE7OVz7tDXR+AMJj6k/BPRL2ZRvS47yiVEG0JIkhy
dmALzd/sWEUG2H725RGNTVmd4CCzsWfYGaSbnjKy46OZdKNySlLGgUA23j55F2TPeZAk3P8Eyx7j
AHgN4NGvZUOWoPZ67DQAXHECqDm8kPU1cfWBFHu+eir+w57yMlO7lT8aqgGOPdq7B30XovpQPG99
hpfisrofdxq7ZBO+Qw0ChHB3Xh+NxXOxpo9r7m+zPer4bPrDLbdDOJqpQYpClXGkl/zNYoQiVkNX
ItVOp/7M31AEnl94Ac+Xg/nT6I5/+r9tsNleW1V2yqNmFxFbZd37BtwVy6CQo4hnbt+6cH02Tq9j
iEblseTD4lM9u+wmbD/KLdOzyOdKqVGi8NM2GW40nFXL+KTyfjSFgjxuXxHIy0qSjSyt0+MhwvBJ
Bx5XdvBmSsgXEQ7Su38mYRR8tzd4+zHZ8m1TeKx5jdnf93xLI2UbKDSDJabxut8eRdhBm92ygdu2
a2esdmDq3/4HjxlJeKMt6OQTqwuXhBK73BGyDO22PIwUQ2PTR3WOW4rMS386aMROTq7K9agdXdRR
/ZZVLWPIUf+8shCQsatQpB6uo3i958gmMhs9xxuCXVuRgJQu3gP1i+XMtroHqWGAwa4M5IoEF7LJ
g/+uBRO7/9mjIAfmiY8iWzfiICPtdxt2qEzxxaArWQbftLkXkaEttfSWL2XGLBrFghCQISaX767x
UnMyRrSWsLSWA0Cto1pkb3ti5+edzHN5blIhb6KQHp6V4AwS0/+4NFD72pVbrjhdwixQpL+HFH3M
bzcMFA15UST6MJKBtIAt1BAE6dMLiPKXL6/0++EIRs/m7OlqTACWvdbKPU74Wu5jpMf7XHqXwb5x
ZLNXCKLjTHNafTwlzVSiz2oYB9vGSMjaxYLwcvIQLOmlXdfxSN5OoKWB+EuAA01l1JEdcxxP+JvI
HrSjnWsDSzi/Yn9A1CFDCsE7wt/GsCO/aYgz9LEw2+PYF6LpX/bznnyYTQRJBRLrB1qHNutEq8Cw
hlQOZlse7xmaUxdrCmu5ZYTAwSKKUINVkXf3cE3Dc2gCrkVQxki/+/N2dfnpfF6Bejq3q1TytXwx
eIOc+vtuIvjp4g/IwkyyJnEUm7TZnnzYE87qP7rNpmmEuHIm6bO5FdRH6Mo/UYmmb9ZXOXAt5aDJ
g/x7f5vRT3PhXBV6PmDs1enOIofdZeG4gkXmbDNA3z5U/JS1rGBkSeK0ICOYcYDqeUujJtENW5JC
VdwI7NgfIzqfvegyr/oJvqIdU8p4dWKsaF78v8VP6ajpxnSH+Y0HD+jAuVE7LU8cpemWX8mAtl7J
hEyidOPPsWcnxJ8PRZb2Y2HI8B5gLMAhdZFzTKhu/IfeUa7tJKgtD22dXfgFm/rZbfMlgp5MmMzS
Ar/8MzyCy0EDEJLOdVu6F28klWpg3ACWuNjhD0daGMK1FIMMIghZjWbKv+2OSktEHffbaLErW1t+
ihKN+i2yd5TgXx6u/jFeCLSAQHMMC4C8xedNnyaH0fSQj3fRs+T4pCG/ivnF2809fEkyIjAsL7S6
JGm6dD1/tMJy4aPVV5czXBZ6PV37zoDNveNypmY7AWlNzoQj1pP/4n3KrKfIBUsYlckTg6rkrmI2
E/FTr+YlkqKmAZutsWn9hlhiUBPYVGRAUMVZauYS0cbwYeNN/qT/+eV8tSaelyM8bPNY+2p+HymP
WaUhZyH/3TZX1tTvtzKdWj/6hBDqUbmTaaOMTVY7BWTBMq5UrnpiOna4YcZVuQADiHYdunlbh7n/
Pseh6Tsz8BCTilhxwmFgTcp0HYjfDnQ7f8ifZ0h5IXWOPflEOQUPrUJR0dKjQMq2sRxGb1r1igGk
IuUXnGbPT9VJEU1EbDEJdw9D9zDGs9acfx02uUgN4VhzbOjhT6aN4pB+UT390/nh2WDuNG42ekps
oSgo4GRBF7TFIeVDTqPdi6Z0nrwBd1rd0TM+xPGnPt90D/uM6OeD7NgilGANU7GrC2s2Tqpp4sQX
mFYmzw3XDqngBoGv1ZbE/cuwGcQZLVpsbe6gjzyuw84PtR1ss56DN5g+3C1dQlnrL+s4u7PSkMSf
NG1qmAR3mULsyKUQ7FibUAsnbRybk2EZdMSse9HoRGTJ3P9rWHdxT5tp0X5/eQkLMzK4ZJKmH0bh
Pt5bU0amNI0T4gbpnhpkypdmFjOvvBLaj1WlODFiid58BreeN01Uq66srJivK3jYyrWImrvyOw1Q
xgfBSvcJc7Xzs0epWrUammBnAHiQdPrQkvauOt2zhwxgShngS/bX5DvKSzElrGwugkIF6okKTVkj
ZpJsY/Lo1nce5Ssogdkmz0B87W//Y440n7iNCFAhnyxMklT+W7tPFWk9Ndg0/dGw8Y42inwTTvRA
90OTbx/6Yla1N9HGu2/7Z0iK1O2c7xQtww8uPXa1GFUxObNGSosxnHearOc8XLW2JKUGDy9d02FT
gvmpc6p84BdWLOKknpXUfkYxbr3PXCuC4T4H/OWFdqyDIua45wIftUHhO8nW3TBGJNQG0M5xOjc/
2LT5PyDsw/1x6IcQrP+SWHuPf/C5rcEjQM1uEREkrSdYtpMUK9rk2hQ2NAkrd5FNvlC/kpDHoNlM
2qcLNNQga4JV73Th9y7q/jhLZrdA9e0WDbJDppKjDuWfsdhIzriwmbF26X6pswRL9LZ9CQBnSOUC
Z9KBfw3fRhgDoVW91YgUwqSdHXgU86z6Vb1jrX66Vy50WZdz+YbwYg/4TrxwBUyPrJaqnJrDHZcx
oq5bWwPIZtyb041g0Oc6ZLSBmUDvK5jO9wAO4kKGaFEe4weYMz3LWt2d3oCISYvC3chXQIer4qZS
3bQ+yJTruhieopPgGWyholsXBHNscttNYrbIWAg3ZqtLY16RzyklhMgkAaG+z2OXx3KaQFUxjfki
2uV2ihojOesj3VBJ6wwNZSSByZ1ekVQPNOgdbJu8oEGLTyHXs5us+JGiQb/LSJYQEAadra8jTvCq
mwZRUioCPce2TB22gRikK5TnjzmLhafM+8Xxv94fhx+sO0s/6oLDksoOMwIyU/Qw5YuXn7jeo5BL
gdtuFCwnp1uMOsmj+KJmxPlRUYkzpxL+vJN/4cWImELQXEypcTA3hRRteJjlHqsnZm6395Ap2e6V
faqLUzfVaqA6OFSJIPuw1tcyALbBbQukEf/Y3nla9hgBvDd+sJVkB3gYKOh+i/qejzWsi0g/Ny1D
TUihUI9pUHKPJImq5Arn+IloPNQsFg3mQARsjbmzHpPixMI0499qzozHSHAG8zSdbuURIOl3jB72
OqSIidPpwTcHqvCf16/0IefIawYR/XS6NR/BMkPPIbSZLRsM7zAD1Q6m02nKtS/0UFudGW1aESzk
bJMReM/WjH0CzZ4PBh1C3qaJnhOaRV5BL5ERJcLnoRS5sPFPTn/9HWJGGxezmnxzplmnA2BhIjQX
aYveLij1ejyvwcNkgyVwddOu8I0eiL3BbTcrmBlAj0n0KZ6qqa/E0svQup+vu158b9d7m8meHEOG
x/OaO8jKK+m+MmcOPVW33714vOjTBIxFVX0NGzmduV24p5Jg5RglTPLxgncc5We1JP0eSXHQOtqH
N1TvB76HCYEp9eNnom7eEdMj4+oJ27m+MFLxDcb++BXI7cRTQwZHJF/WHRKVZp+C7zF4DdmJdYxQ
s5nnoj1hJ/RCplDYYyJnR6HwgyMTS0tkAmIlvB79MDXToqbe5I0WP3Pse6oj2RKt/GRLyLKlY05g
efSw5JSaqv+QJJ9j5kJN0d67egsbmF86TVV0ttSJb7D/U1ucehbI8aa2cFY3gNt2t94kcqXzY0yI
eYaNszylZ3E9uXgQTo3F6k5pxZZm9lrNgd8sVtXhCAKjjG4PIvOo2jQBVz7JVDNqnX7op6pPS6Vr
BENhUDp3gYGBZakW5H3ZeEj9gjNxZVjE6KjXdSBwwK9jX67Tw/gB1TUhTxtdzkC3rTsu2oqz3UN0
76oUp4jCTGX8xkxXXUSIKrk9RbfmVPf5AvVlS8/0KGOer3hR6zmkW2EyWr1Zra62A12Cxqn43Yoa
6E6dmCp2/WSO2gMbN5cgtQOBq5R/nCIKuVEjuoQsfHV4fTiY/PWDe9iO1eSXqMXCjnPCwQY/KKiP
I5agztFEX6trtIBCbwljsU/bXQbhO8FpGl7y/PqiWpdzC6PM5AsHgRmopg9has25AtQaR64jDOiV
jnbGOGQMOHOYg0DfksDne33fK8HMmMS4Ed7DJ1OklcuoNYc+TNvttArJ88FSej4nvKlmnJeEiv2g
LalYcqzkW5ZIlymxL4lbnf9RsceZDQaFBKVmLiUjQyeWOFVVLVBYyZ9plA24FtotJ7+McSefotVv
nRQitZLY9QBhCozPd89YWxyN0S2uywCGQZvbyVkxxDpPzFHCAsXqQHOGFy9oNt4v672SMjktbGik
Z4PNLC2PCLva9fVDLjk8ODLuYBxjtdxAOvnauKkKnJw+nH14r87iQZmBxKKvNo8wVl3qnpCJ5IOG
n1sCswL7dEBmtNZNe269aPNQNqzBvBRKPnJRGzh7a7BIzX6+fZly2S+PqiYFpSwzzTNnhxbbOE1G
tk1WZSDeY8ZR0SJl3xi0Vlv5GHFwmhQ4UyZ6yP5QUO6Tz9Xol4Tqz3q31wENCoDMGh6eKAt7ysRt
E9wMURcHv2ofYy27PDJlgUqzVF9RFEAVdzApa83SfLXsGOIBBbe8GqSwKZNHFvPffBgB60WpPWqD
/ZzqlZ7rBFbjSaTxxpcXlAZs0UtgT02XSTGW5ocHMJ4V5c6/CFkyQIftlSkKcdxDQ8OtdpFnZ6Ca
531bwiMGY939C8Om4wiKnucVjPhp6BjklypNgx30ucwqSts7nLS8I0+8g2QQ5Bo+Gu6V57OH42yt
CkA8QAKIAUrhetKYf3U2PB9BrF879RE5e0MtiMwyoHEVksd+5nOdtvyPH8TH5MgHzZORiQKWaLGY
dJN0eJCs4BodfZnWkyjSgwL6lrxAbl6Utb+GQ1qOkdiUyLPoQeBMmlLqRIjxKn6GRaUWb9bfq7Gn
UVzsiwZnhYcQHB4Dd7k3whN1SDuwFX1d2ONPfU5EFBMAhw8UAjzonYdpwfngyOvDQUfdEPx2IXDk
kvLcM53U5fKiZnc5j8fu1uLmxzdQsmveHTT5TMs5k9GYPhdwXuSUQV6Z8KIExe9xCAeUVzF2XmaD
pyPV4XlxROw+jR1dscKgP2Ar1jf7AirMcPofunBTHaj/Psdn488+sK1clQYFAu3tTXbk6WVEFeyJ
FHW5Y9tmkH+DVcWd7tHT7z8n2B9vZrvk7c8WXbv09HlQjo4FpXq+au4RXtCk9Wd4mmjkHyHa2QiB
mHM4gWOXxCOsdC8DlQt02dewQwpaHQhiYjnUsQoQkcSuUHQUZrgPBar1zRco97vkubaT9dfEWM9z
B+8SazAP0PMVHhNu92tjZ9ujL2Ol2gY1Ghp85Woe5NZ75CheRtPr6Cgz7JN3dLOL5xXLFL3KZN81
8kcMldZgARnq1vMd1ZbRPTatMY0wY81sgJHwts+MGrIUU76X2xbBm2pS848mY46eOMH3CBd8YzpM
FogHZ54r4e138evhD85gTdcC4C/bFNzCjP2TXqll+6YSSy0DDAMmHUms8fkUjvSjv7AycPdhDV6d
AT71GZqDZC0C+JXltLAhfkfTkNbLoYMdEePjPgbvGw3UB0zOtYG4udXQxh6I9iMJIY5Zs2IVx87u
t29U/oE9xz3NgsOJyVhUURWnIm1bF62qkxg274uoJ/4UPlgBeajHoKQNE6rysgZ9S7sK0AVNk1SE
5Pr67r2GdNrTmVYsvufkqalbMniQ+6wm+squvATEyeZ3IdgOHaMA6Ph4PodACE4gwq/UurOZ3g+z
+1XTkWzaxtvRH0GmdI88lvVcZdOVyHrB38/xDQY8kPsHnNZCrQIkpNApDN8VSXomUESVTch+H+lQ
inEOPWFzKUPNs/bYvKSW6lhYYlb7HLauWLQGPBjTSsahZdLwV2wkQxRpv4utiNfWlMKqmiDjlZFX
D6vwkLKJQlL2HZBGJS6rC0K13SQ5xa1UA6AefThF3l835OCDkEUyB95NUN/eZfNJZiJ9bECp9+u1
5RfPbYwc39AYvm5CpFRwKxH5hLiCSw0IR1to70dG66HkoI17mufP9Aapqf1+7glzds2pQMV/XlRE
ExIMNBPClE4KScfwHFB8b7sOHi793ySgidso2NIMC/s/4lNnhnS+8VCzpgvQuzUfV+kw8IEdNFWp
QiiDhie6gs+vRUqMDKo2DCcKnAuSyyQE2Pep6D91LFJ3DEXCUNAIfgf6SqfoDreEK51vyIFFylxO
FKASKxMXtgpKEJxzQioHYazwPNxm2Z/+h+R9XEJV9U4m3vPa5YdbP5zITvU/MsisNKIy9ggArxlh
nk2Blim+5JPXZ3BT0KZTqIohRBAAmxMuHiP+LdMGSor/invpqb/x9qSJX2z/Fagl6ZiqZ9yKqOSl
Zdj0EnMzQCE+uL9vLxe24VkjSJbwlv4ocHZZgWk+T9hc6ZE1aL4+UxPaEhC0dm08avqcFbhWhaxr
kNCn/nD2uqME1b3FNP0+4GnerpsYZF+Bgv2wPaimLjL63ioXCDEVxmUSBEkWz4oZZQ3B5Yrscaez
WLIKrvpSWmViFcrG6zFmD5GpLOgYfAQLEC4QITx7UzR8bSHGv/aTnMhMftxm95nkQoYjUc+F8LNH
z7E8naLxfs8vBhXX9LsB0rXjS8BcJ/pMSo94cQHPo62hfcc5XjO18O+1vZxsGoqOM1Eli/fvESq8
mrvf/Cs6baCzJ15Z2Eb6gc4UMO/ns0cApTc+cfKoK+LYerFm8E4UCPnlv8ptSFTgMJprROFAyQLe
dzvH0mxf8yTzBesQCMt03aZV4CNfSY0fHidyFPt6goDobyUQ6u86OWv2cbmweVSs7NnDfiucwJ17
vBI6INieccYklig55epYn0+2IzvB273B/oANT2jVTGyhTiYEnfGzeQ9uKoPHkHg2JVzKG9HxIboF
vR0TXz6F/l6Pvprr66I0VdCRM2nQcbjOisuaJ90NPGQCZkXl2D2LEixwgXquL5CwQrFJ4HDuLy8e
tWm62NKWAtkJUvpbq8MRdQp699K3eAkiiDpYyFEO+pxsPlqCpBQssjPB9ATCyXmW2dxNhutJ7k/a
pLoAQT/xjBs3IQru5WQJ+iKpZgl3PeQGNAkzmlN4AEB34WGcQIlR57jFoF2QLWKV+0x9GNxslQFS
ZF4MeC+0KGsBeOTfDBYJNt2ScfJOcwGmo9KzYl0iFvskhJBY0peAAwUR3e1yulKOBeC9jiKl+Hny
M/zbvWz0O7Kv1/XiIiacO+Q+ximNVaaGrXKgkoj7dc0YCLczvqKGeheABkV62CLScLVnjaE9w4Zh
YkAegt7omfqsI0KpvwMaBls1Y3xwVvBXiGjYTS4Sm2/tiNgpdzl9GVmaDquvvrr/PFoeLdFd1QOw
Kz3Pl/9YGEN+ruYT/jTxbGwTopQxDA4jXwzaQ3FscUShp5sEVkUCb8Xpu4QlTizMw+fLPtLnhpsA
AVuEtXt31ckMF5gS1ch+oOuooaHD0Dbz7hvskLuSU3JcywqtsEvmMLigmzGGFvQIVV2ETD9+Qy/U
xgRhRFg/P4lEXxzWxK3rONYah1UEriwh4ikWZbrLuBIWcVRZuLMGNSLq/FD8toEAC4LcktHV/Jgq
Nnwmhuy4sJzRsKSEuPkajUhjd0V6Yy8LKausrqjvVzZ7Dqg09EwOR5J7z8WUbncqrva1m3Ssaaws
SDFWZ4pM+fI2HLfs9CGZq8TyVeKDa4UiJPLutZ6jf7v0YjXC2wZmg8SeEWd9QyIhvIqolJLgTjbr
qI6WtFTvA45tK3QfExPEeFE3uUKoR4yJ4dIhmHmjIpF+fGxW6soaDp/YhsI0idOv7yKm+3VemMsB
oiL/a1f5wXV5OPOgfTK7S5R+p+wk0ASMjpRMcuL+edfRRgT3Ldx7j9Vc/iOugLp6jIW67RixvjqC
lCncw0xYSK8ckvz0cZajweRYPnJT7IU3QeBSdBQq/PisSr5wSocGO/06omfyJ52UknBqr6Kvrwtb
sECb1GCSBKu92MahYnG+lYaQ8qWo68d/YFN6KL3kZ9l16lsFAg09tbqPu/cbBvwy0O/aEwhX34X4
4cHeIUeYpWaA75hUcbzsqqFjEcxFpmWYe5dxMb3cyg9l4BoE7iEDOn/qlUWSPcIsBAi63OUZpYu9
FqrZT++DitFSsxmlC8kFdZsl+asdpjc5HuZ7KGs64Y2M5haUsUnzxN+kNbXYuJEfMDUJ75hMgakC
ay1+4SFQv+uDVLm4FM6P/WVXh940qMumR+pEeQfkhWkVBYj1XbXpEpFjBKA7L96/zhuUdicRx0qV
Xrty9o7cFfgrhJlGTrUV081nXzMzhYjJ7gcAmA/wHnqDZmR0s9HcmCIhx/Qs/dgmsU/2HdCx54uy
PVRC6OMjxjB+xdSYRcMX7cnVRELGPGDe6Gk+1XH06vUeYf5XjCZDiubhBGrGTjUBsbou5sD6d4+s
4W5qQktNAp4Rhci91gn9aMKbPk8M2MhNoiUF4zWTnmhJ2TVd2FlNy8no/ypsKaDwbtRpzqH/T/Fa
xXHgYE04i+HDpeTDaoeNZgwlVZmy/ZnbKIkskrd9iL8t4s7hsq+7Z+MHxsWjUnGMJPS1W9hkkBBU
BrzYa27gCsXAwCBH07/5Kd7SGd193GhPIjLrMFPOa9x3fL14bMACyLExeuCx5vAFdcxzbFCvMIo6
KQ7uh5OFUYBSUzFb676uHqGvgrzGnJVm+6FHMe66LbjsZS8yq/hKquo7WAHT5RkMoimFqDgG5xcM
B5io/hNrBUwjgAcDqTPeulTa1gq/0n+XidPHXo4Lf/EGImXzpU3MV3EPShoNGgT90G5msxMaqD2W
mksAmcJsihuZJDepFFQWzH8bsGRgihzO6NtIQygOVfWYwAcW9WvB8cLa7qCTY623r/ftfuz4Wo1k
LHqn46J5Mf+vIvAgCrbfEDO1RBp54RMAIlJNO+Ql9nWA0G8UkqdHQWpls9wstbqiCMpKNeF8l8Mh
f5zjSSUgUUcZnofgHrES2+l8sSz4qaCDXc79d5odtLX/soWIsdeW/WvFXTqmAGLA9m/lVAyIftEx
Vc+q/+djXBRbOVRfUaZzlPEJvTfr+0Egmtmf4G7vaV3F+DiUoeqayfd2or3llf4mQdK+d5f+GTRa
n1G8NMcfP2NiikLBjsAyrVsuZTy1AH8ZyRU4eeCD3xa8uALqnLeJ6IhNww2SoXYTi80HoWTc6WnO
JwCF/bCbzAflCRGedfZYwhaYw5MUd+OjyovKJG7s5iTZdgq5sAzqEk8HHX5iVXSwKivA6M9cGCIH
Th2zJD3cywmzjqwC9pH4I05IM5uYWzAj4umvERB9o2IAFueVTBSQ9J6B0ukhmdbYmUZdwcRXOJjd
UVV1M2qsCLcma2q44U7D7SVXjxzS//vJnoh5NY1EXgYy8a6PArs5SNI5eYSbzMiheUdQITF08RaN
WniIlv8qFfH98ETD+u1xFIyB+0fZUpRYtHUJmqv29Q2sTVVRngE5INEJeZ85fXJwDNROtT77gUHU
ln6V+bvSkR9h4BrT8mkZBUSyf5E5pXkqrDktzQYufi0cnxx18f6Off29MAOVw8WbMtDiOi2ysikN
+KER29HyuJbXog9vry5neInNi+vuQv0wOgGGF97hfGCCK1sUDayuZ6v7iZSjwecTg/1cvhTrQS+R
jJW6deI8nlqJjyzKuemL3xxHxocMefPz2NBiREG69sJOkELFDIt2SkClaUfskRtpjWK8Pe2FWmua
zUKl/ETPdsn9GMb0gxxQ9TwfD2i6IO3evKPVvMfQ0xGuXFeg6gN+cm2GYIjj8HlVjoHQEPw47gld
4/Yv696LVpRemRJNji5PcHYtYzNsJr3xjFj78l1kyn9kZPh3LB2Px1YzkIFZDPxQESQd4APu19pP
/9Y9n7VYxaxq2JqrLBofb2VNYo2kJnMPjUhJakpqrX/87kDiRYAVgGXFMineSJMZsV5JGy3/J1T/
/D/WpjY7B7es9FAWPWvErpveYq8SekbGIsfWnVPQ+X4prVX2QGdx4fkp3aqcPjDqDeM47zlqcp6a
rpmCTXaQJJwWz9cqDbzYvYrVRYTwtcHKEfDR6RlTL18tK9Gj/v8Lt38wwdnmnk/1kiCiFBQ1efhz
vzJ9bAlauPTJjXphmF0LKOjEw+13Kll9WED/z4A0YsnLFieOOoAaxPlUzW2LGnbY/Gvvf6KgY+E4
N2R8TfmcNQb54bklwC6w1nIA2UFD5ZLLaoiJedFeUcMS/f2IOw3+1pG8WZtgKz9fqiWTh7v9ekXh
EpE7JHkG/KZuXrurLXhLYj2RAi5mKoR++RopkG6Hmja5PlUD35hs45lTaVx1ska4kMtgusaXMb1p
lXSqaQf+sEofHUFv6ODA6IbPFe4I0XwfK63LYf21VvKDG8oOLDA2aD8NWNT0cxzT1f4j7V/EW9DL
/4U87HPzPtsUtmUdb2nXEBJdU16/6AQyNB0t18fg86lMMi/VZIuzRXHULAVQEsZWHv2e8Ou8/E1M
KDHX7/2WAQTnLgbqf3RfW6PtlF1qrLWQLBcdOl7D/iFd3UIIXNZtbXLX/iJ78MeuaXcZmuyl+QdV
/H0DAdhdJ6B8dAvOQlUtOOsjYIvpUWYWFyRL1xf/ASAKL1+Zp+qwL/0DgPcTLrlIgASCAKnagOB9
MEx3T3b+8l6kt5aDgRtzIuzL9gCL1oLBziIQ9rYzVrQWH7Gu/VI+vlnMLSsuufCOcbDsN1Ncvv4a
A/d67htm06WkGPg59BMgFKtJXvOl9328CDSx2nMghtXOi83+ay8v39bROq2fwDH7ykoEK8Ylpfhd
pOTD7Xngg2JdfwJmcxSoSTGW0dxv0tCu6kC8YmWaXxnGVSZJmGvngtVUy63E3AITUho25sP8Hlpw
RSqAec3iW9dtW6wpeUj6DhZtpn8LYQ3JZky1MGLc2gzLIRYdZIa8avXIeUpfjr/nxEIiDGr8B4fz
LmdQrSzNrsvkt2tTEnsN36aWTPwYMas1koc3DjTNosWyxNnPS7rRYspTv7t8clW57VbQiHlQKOLJ
ws0bBcj+/t0Gr2US61JXErnLQEMK9UXXCJ2nJ3jApXd2vgup6UxhIgNsnj55ZKsllj+Sg0vZ3fzt
n+MIf/lvcbtXHQpNbroeWtzm7Ybd4o/ZHB8P2lOSk5lmTmar72riM+ZActnWG98K2lr0frEfi6wc
Zo7lqv23UeQsuPKVYWbNfkfOyl0tpkI4jjAQxaNeHw0yqFBVSUbq76op2EklSAKRwEwt2vMj+f4V
HH3vQdIVgRWe1qfjq+94EBIgk4na9OXLVgg30r9U3KIzCMda7w8h9XlcLb6ceHwQ+KnUEbzGGWiW
XRLNusWnJMr3GJlz/e5TfNR6zLh9sy2pNt96CwPBZqkyr5VJRd/VBslu19CbAaFFn8cqZPXUhi1l
hbre0mWX0f/0gLbMU1booPh1/H6mcNdNaNhdxEtcPUt33OSnsP7LycMMbtArH+v5aolHrOd+mDEg
TmkHJYnvgw3+9AS1mU3h+MIIDivQD8bi79IFD0iQ88G+7GhhAbrUEDVBv/KwhuWQJK7fEQhTw0Wn
CHWJmoZXOBh0JQl3RynYdUnpA6ZJiCj/0CX7Fos5ejHAMHxySw6KVtdpB8Xa9LOHglvHdwi/crvb
gFVunITi/waj8/VOMSsxJhct4sC7t3jAus2rNXu4WH59ChegHHppd0fRgnwr/xWCh+WdDboEtvZc
kU5o0BFgQJ6b/L9p9PestxnAD/YMww5b2+iTsA+i3rbNcILypVfgVX9E/PZWoKlYoWmgZpDZ6DHC
rUhIS5bMRT11UCAOsqkbuBBLIqsD1m6FTt9hBbwgK5WUCopK4M0Lo+XhR+pcdJEo/34yutEhr6X2
VcgYciTOS04FKrF2939XOCq03RbnlH+YRE4SIxa0pCsP6vq5b3TTP7PsT7bmHLfTboAfUht/uZAV
ywpRV5JoP91YL3vUpy8dgSV5Z4YYfz5fG/eQVx4oxSEkD1Z5U6g7PiwKg9/Ppa5ZYDZZNcCehAOI
Eto06ilAUw+5mNQIGeCL5U4jX3enuVzmP+yrVJqsjBZ6AsNJV8rp7RehhlXGfQF23xbAMP6OzMDz
LQahkpRA0UXKi3bVLLNyRor4mbOPwCi4o1ZqkSBQcumbHHMl+o8K6x8M7w9zrSvkdtM0neXfZ6en
hZdNRCdGAJ5/TdBtwFOi2gR1woylHURTkxzwcXiG2WmOILlFy2xMKnxQCnEv8rpdOucRetI6oUt/
lpdM71FiLjfAOVfB7bhO6qBM4/0vgAq/b8Kk3LbpfVinRXHgAxl+wXIJP3m/+xe+fzqzJ2mezcPF
XqJZz/Pdd0p5JROJ85qcHk44bD+9ATJRDIs9CBUCnuQvWC2b8KW/qP4DXq2WUfLtRDxQ9Sn1iFaS
kLA7VJHQT5qVqwa8KjVzsoa+Y3QVL2XxsrsAeJwbcNz5mlko1Ztjq+cBSeh9aJSQyTghTrrm829z
Sfhz5V3aqsOIKJLCe+ohwOJbieckwydD+ZAvBurgGjZS3F6ALX6y+6YcmTacfxoPs/xAAN0F8fEU
yoOnx8iCsbVpWfHAU6sANtayvEqd0Po3ZU8hoQoO/S29gG/t7C4YfSU+pD4Rb1YcfdUCecHolxC+
RWKwc/+grM9q5RDkjuUeGzrMLCT4VhnmfLslIjAFennkOUpsw5Luq9Js1ajI/m719dYmVEFo0baB
UWFkDRzs/NiAilUg1Xpl/X2ZxUcCRv+LpytqrESSvhQqd9/Eb4k9KexjnBUd8Kcm5TfccMTdmcQA
ndKzsjUUZZcHgF3pxyJ10SOpIlhwgUvtAWfhllL4Cu6Be0LLkJYbUHnLMuGQQFpvl0SYB14nwn8J
4ZGKlAlV3RGbyrvdP9axb+B5U7eHtSFF65xlpxW7k7U+ropAUPrUj5aROjolEj7sneIdKVwwvhPz
nHLXfx+Sc0DOLUZTK2gy1Ep8GifKtv/JAXPCb7LqyIW8UU40D5TQsx2gqf/FR4rJpVzEYslbkZNF
EkPChgH5/0oRZR4xqcifSs6yxU8120645nPsOF9d48vBayKjsCnKfkl3w6VABy12XzVerVpFcoxS
qMVs0uv2p2yM2CxnGNt8AWN81sMjmI4/v4RLlwOGZ3bGME2H4yUNp/Io3sXog6LV99lTArwNvcrE
aK3C+O6Q0NK2b81N5MLP+1V/IAjts/Cave8OU+bB5H8TcalCzeC/Ltcd+i42wXRiGEEgy8R8iPrD
uibW7JvMUe+yJF1qJRARk0UUroVro1uNjBMddYEiSNJ4jpktD1Gh3uEYOwoKnCLQdDlI6D5hTV/7
f6pXKdXQUDw+Gfq7U75qu7VYihU2ToIyML8+x5SP/ZmAACsLkdZi4RHSaS4vOU7aRRzLgWwN0Lqq
/FaepJjDl3AfRDME77cjn0LMVamvaCJXMsiounVtwU4yab428uL4tUYIgEWk6qlvUyHESyhzmKMK
fJyfZHckLT7ChhnND4ce1dglt9KBuYb5nUbbja+xzXo29zhdDe+gSUYgQhPCxLEiEnpRdSf2fYrp
OvlutwBh5M5834HXhFmRObF5tW/PZeSM/Pr2Ak5jhyiQqBNRMqiIIVj/+yPqKyZCncxqfAsUnzCB
EwCMdpOcTPosd9cC+ZKUtoxpPG0fPFvATlXH1xGRusTtzMok52iY4IeljELd62adLAJ44WDEtnWe
sHBU00190ndcpZ/xSs7lOLuqrRWHl9+285/pHooPpGy80GQyQgYNsiaON29Nj/0FZhHznxfluuSv
711JEE8yrcCRN2GoBkDm6fZWtRoy7yhNR8chRM5Ysd3kia9nu9lAbAJ9NJaNWXi+Mxwihu47N5qA
zTBtf5XhE/OKEyfeeQt0+qjb0Yigv56oSJeQ79TT1NjfB+7Y2SiRpWXJ6qGyK3B6uv8I2hjCfppl
GQL0wvD262EUDem6U+uMkClWEsJaoGh/3ETbV29RNqEXuJRguj7Nr/Dkq5k7a3soAjhxNSxOKalV
qJM9NbWyKwRz2hC0TuHB0BufISwuiMm/i/tGelaiD0HZQ6j9J0nSS2e7OqI2vSBNQO+m5wAFFLc6
QvnnQBUOuLh8LBioWZIUwI+rLL9CvBvyiaxAXs9cZXx4CPe7tVv9KrE8HMsp92CxYsRmLLqDcq5e
Z9xHgmsFH/I935V07hntcbq1Wpo7NHgcYs253RlFGATNngrrf3a8i31rtpgOPdubcpGgjZ+Q+Vl1
2iZTKlzVjolLym7zYvGgPkOOdJyiNqT72oH24lDcd/NWP6tKOYHOIMXr1JKfG0asadx0Zk94hQeg
iXBEmdaZSBQRIt3QJpazY3l3V2+jjAe7ZOpHfQXNTjqzsL5owGZzQdnBdB/dEslhlFr2VPc2rQR2
GgyZ0jgfQ/BYlswE+nDKDfF0Zmo0YXFlyboKC80aiF6izNsq3BfCF4JUxtqpNkauyWtkgW4IS7N5
K2EOJi0u7EU6Sv0z8RUYT7kbY+nqso3hYjIMkudhNOEXO4aFFcwx08+dvhxe0fCcbfgoPGp/YB7C
ZYaiwEQSulcHDcGIPjTSN/j/iXKnfCROES6m7Xbn+T/bUvu9Pyw5tl+TuoPiaVa8o+jJKRR7LDw3
oBqJ43C98Hz7HSwCeU0/Bp+b6HuumFtGhf1do9+EIBYyUtyXSrguOzaheqSM0cqAqi1H95IjsyfL
+yysGieqRJfnss5z/cQnbXVlcQeBdj3nNSMVn12Eo7a7P+jUyjW99A/5jlkZsVRyYKQN20ABkW85
OvxieyyFKRAxQayThrSERwjrLeXkg4eNCEyKUMx3FMsER6BpdPv2rKDa5GU57M/bjLaJmezoWs4h
94DjcHtBHIheO68V3SfARLCS2t3e4hoEN+f+CKuFTvAwciihjNw8C6CdAZdqK2DzRuNilV/WQW+Z
FiwhhVe/BU612e5hIJo34U+P9GxZAqfmsLTPm3MbSnSVcGOJ6DJZC1MbO85769WO5LZi6UhXliHI
fkg5VNj+BTc2eWawWS9QstbeOv2O2d/m5wpHFhc8IwOJ3P2NG92plrTibIy95Cc5PvhJvqUpwEGl
mRB9N0rPSzEPLg4sTVv2VRo426ePq4AXEiVrBEaCfZ7jxFtlrcdVR6Xrz3uIG96AMW+DnpVG9neI
ey1/75L/EnHUqogE8iKwavGTzPkhP/dNCMoVOxQPS/fHqFySV0U/hjsAuzDDSsD18+VQUCYbggKq
4MeWfxtCTQ5riW95KP6x2Muhw8mVq7guY9q0nWqFEFrvpluwzbydnoBfIL7ndefGzQqKAmm/J1L3
LJvjg55JMjMlKjY5PXVxFCXYDEkwqb9KnnK5c6SjOViya/ozwtd8ibLPLM0Uks7wdDpUzY+geXNd
glqRceMZPT5Ge8dU/jLw5B84MQq74Ww+0i3cZqvglMhKMn0NgbqEQqvjVSwtIhO2oPlHX7ByG7ii
FTbZg1iMdpWLYgqzmkFRcgEmBYY2G5ZLjy5hNa0rN+n24JQd48bD+HTRknRX5ns+2HmvZOrydVtx
o6eunMAsDqAVcRFjwjkSMyKjNLnicQ2MsulPVLlIBgTnD0C7y0w7WKrORKZSFjg4keupmc2obFfo
mpMD95YhSkpOOoKEkXzN0vA7OJZ/ZCDQbp0NYY5Ir9z7lMBemJ8HN60QAKLrEq7r/FFDvfCOQhTa
Ob5GOOldrAZKLy7dBlc+tfbvPW6E1+aS9I0uN5pRGLNQakJYsbAlNkvIDdWX5pKcIkbreXfT0ijI
4+szkoSlh/qQA0i75SRE/FoHnSjaCVHHIPH5L9lw+zgsodZrZnrT86Z5BEECT1VOyYPlK7RHZsvM
EGdJVXfp9K1a/T9atVMIHXIPPICGi+IoEXRz5wZqTa+KB1Sv4AMeWihlgsIohy7UBXQb+nxhre+9
KCjNWUJ3bgY0z7SaLSV4mKXceBgxaWEggGTO/WYNyFAtgbyld4lZIbi8X7xgxTQey3OT5ObQTYEi
xpNsEn51J2xYQblFhepc4GJfVovDv1Pt9MNXqwv3/0xdgh6E1F2xT/H7kJmv7oWl2LrC4dl/dIZv
MY9Eh7zlikBdqQRPBRkjTrbT61JfaZm3HSjkaeCl1gszMAB7oAoSCx4zXORfLwI+7edEssOMsOY7
CLELl2CVRP1F5YwuSB9SW7pIdsngel6T02aZ48PvUA8WpMfWbcNrT5+ufxZm8/lXaCvJpcb3MGJ7
UtR4j8S/xRBAc4cg0dGZVBnqj0LwpBEWNxFKPOXFGESDnpi7SE4wFLlUjCjlEwqbmjZgi+VTcP9L
EKrpTsIoTNCb7MqQjYV68/80s8SlpRFKXG61FcF3DtOhcaxjCZomdDIpt46JdM+7dXKPUs85NTxP
1mgekq9F2FZ6a3njrKCC0Zu2P+wvt8Ytw9DlNajCOslkPRzKzlq2ZG7E6TX+KU5xXV5N8/OUoppq
huiWjESG0mwo+qB4ci44PDTJbknJ1V2e5mi3gFmf7RjULzReQ24LIm9eYZgE6Ibw8diH32ffKPrS
TQA+C8FeJFaa1ihK83fcwIa1COi0LDfUC9qOYni+7nvICsLCnWU3DSCLcJwla3gOIH7UuHHgWezP
8dMgIB0u0mUWIOUrMxfEvK4mHofbpbBcaC1rSPWRep1sIacJ6AuuMmTnPbI2CzmCFdyaFYf46liG
TP+oEwG54EcPFykOAfgNDiyxi5lbmGQFf6Zj5MBFYHfKfeUEnx9rb4sEs013Wyc7grj2ZKsHO5eZ
adl76Jznz2oD/EezGmWcFBrDgCTEeBR4zmrFNzQr168EvdyzoUFpv1PpyaoE3OIgVpn7E8guucZc
BQcu9kNh/yg+Y/7Qa/cquQ1b2XP5KIC9J0nkP5LllV1zdigf6fz6y4MWShBy9SgEbBub6lKNWDKM
VdteTHiukWQBqhvCPTN3vJ5Xw3xQo0SFDFfr9JSMfWrzZqFSLOedwh3jnC1T0wOX4ync1cJdWfPZ
vwPMFwhwjBrOou9CjZcRp+tfDGKlPhl/phOgH67A6dgAUAL2HRAZGaOfeFJoZkZeToJiaHwmBgA4
9SNia7XgDU1Q4AABaHS1VCzaEFyK/PhYxO34juJp0VwE6/B4MME6xsJ8Ql3xJenGArbMIS5+l2Zd
YI9+ZiFe286yexM46l5JTBo0T7FAO3tNDDn7666BiupxdraM8QgWUUDRl+oJ6p1nB2eqatuGzjJD
CPxoW7WZ8IPOQQmYYNGmUKWmixY81aIq8tEo/vj7dIOIs/dMTH4s95xjSRAB+w9fUUAqINHOWN8n
bbq5Pto/NKMYmUwCnOBB86+3w+9ZYBNkjUxyG305gXVGeMeSzJwWfSmq3dk4hhi8b6kU2oy/lSZH
0gDyR6118r4PGxP3HYc4bOSxTl269wXU1BuUpmSF+iz03ifKMNv4QlhzDiw8ePJ8rpHDk8sglvIF
KAYc9cfw8w3PmWxbJzbdml6eW0b4IcxvOX1WjRVelfwhxeqKJoufXbpQEcaZOmEfTr8sm8G6CELF
ZCI6AnXgvnEPeEW2UpzNtKvJDz7KGy90I/4liU9BUax+e1AR2N1net3vBj5SwEqbmtCBtwKVE/3Y
bUeFTnvGghKGJAtVS77w6IkyLT9mn1lIlqUvl12OnXpoEnOAtRjs0Zt0OrTUAGDIDn+s0+aIx92Z
c8k/ohf/vR5pltMKQyS8mGuqKf4QoPZz54AbMc/cDME4bIEsFcOeIUVnNmwDBwhnikOA7K9z0pur
jBWXrKDI8NEjpUwg5aK2n4bqKp5izZfiXtY80YVOBtJhSiu9VqCnPKd/CAlwUHEXw60NBG686OKm
j+ZfP+NM6NO4hcwglgPPMkmK/ZBhS3+MQL0hEK4sfCU4MKmiF+KfV8JeqUinszWL6fVEH5Tb19nr
qa5DnCQbELiGkbkS2J90rU8Lsd8sHORcojaL32/C0h+MEPopw/Gi4ix2ybkN1L4BLJlEu5Tux7Xp
/s1iy+adWah/OkKFeIVEcIj9Cgf1xQGCW3Eza6VUa97wq2fDGUoTiiIPCuxvyiFMkAZYHTcGao2/
1nAUhrRpkjb4WfrLR0NHuD75oqLsKhdtJkLQS9OeZXOMps8UiQa9IcwEpsgs3JhfQ7pDEJ67GbaV
O9Ln7yKMlZ+h76mEQKoyqmbplGO5yer9unC6hVsCi7q+uvmsZ/LojsIAvbTR3/L4zR8L7teBGPeN
AdFS9bdYbuk5yIC1l2kGFxELeaZew3Enr0DPV7z0fdXYR5hPLiIL5J+bNXQhN15oJJ/JjqXG3uxq
pHt66SeR/jVrhuF4tBs7UVUlMBTrTDyhnCqm0eUpz+T2PWveiP2z/Vxxqrz2zbakCgE6gws4r8vH
34+Xs0+egubfpXTYVOlAnEiKg3yjWG6/g0LE0DPR2/TZSjO8ABNb7ztNmEACyL6pLdLhgWZfpvl8
635aGDuZ/FlVJBubN3gzq12nV94uf7TXZQVHHIf+IVjMwkFFsZ7rFEGnvGJjmUbpaVVVFBddc1wn
BpemSjg9e/JZxk/BqlZHlKzQxG3wVB78KURzi5xzliN3/qRpSgWSsHZo0QuEnd6unhbR/QVoWI9f
pFXnevt+ET6Cy9eIQhrHBJhDfnmq8uv0xTHIQx2tkQ9dzmy+N3zBXhtBrn7LfNdcGE7oTQCWIfnz
NL7GYkwOL99qQwjT5MueRj94KmeKYN9ra1u1OIN990hcS1lKRoeDEIgX9WhKUHKbGiPVfbI+bGia
fssGWZGEiACa2K4FTWZ1l8ljFK54fYWK6RchKij4OsA3zVcnXm6UuoMlbmK8lalsE+dlJkQXhwLO
NooUQ5DaibhhiqFQ26kC9vVCyW1kizudrTuuVFam3ZvMulp5u65RjzB5Z2jlJEhGQTxwaUkK/wRu
6J7dQ1n16JwyemqUYEOu+pcEYkVxa/E8ZAavVvZodOS+TwjCJDgVdR88bTIDH/V37MnSw7oOun8e
pX+I+PH5AB7MrTBbgie7Jb2Xc5CtMoTqK4P+TQoZjS7h4F13hZRd8+9HbFkqcxw8n4HM4wJUvV+2
uHaqv+ZXx//3cGKa6NXVrH4yAJ5SVJheYZL9D3Kr07hmZujiMgMwpkpkGfzx/izFziIFalorLqkq
eKw2JAom6hF/x1g5wU6tNKDczsPvPD/Izfpn5KAJ1PvAcpfDoSMN+A5dbkH6fn57/m+C+aqfZMsm
9/4xdogRjvogT2nSfoVKqYB1UTeYgXg1ClAaSqSZkZOQCxAsaVlMv2G6K9VeGsGCrNNmeUzJN0l8
IeybMTKD5uXV4lo2VNwJkLVjeFZFc17s4KVtkeLuvKrdKA0YuI0Gg/SvFduEsurrkpZjb6xGIS5U
1gb3oSWdW03QarI5s0bMqKbIkfuC5x/vO2eI2cnzE8gtAuxqVbuH+TNM2Is3VauJVhVeNvVi1igk
ha6FfB7eTlTgDe6MnwVxBq8XQJ0tgaBIvUWj+ULbl6mlxfUDzsz1Q21Ifo66V4XVEEb9UirALsew
BHaMky6H0k0uv3QU6b1L/u9sjPruxaMFTOvhLO7terXGN2Gk4fS57/+pkCNQ5J4YwHEhsloxIl9c
pjCidDwyXcAepBoenZYmLtH4T9CaxGi2wPNW6RydzFkDGOx6adWIxsQW897qKt/UXimVHwXgROyL
xzG8U1hz1vC/WXx7ezHxaD4LV4BcohKPhDhOQV2OAB9inXlbS3ySuQQwc0aEkoH9Gcsjk0bofjfm
75BTRoNnByKxxnep9ZveKwIQDKlLVqcwAPH+ZPWsR6AfIxQq75uCkL2/l4tpeA9BsmsbZZo9kWtY
zK+aWpuZUlgCR2ZV/LGpktPc5IXhpCo6oPXg5N2DyDHu8l7fO9ld/wOOIO1JOINviZ7hAyZmYeZA
9hZcvVOOo8mafktp30p8nimPNAmvMo2KijyMdtwR66sBvZi1Xh+3oj2e6iH2cSJPdCVE08fM+sd8
EAVFjxQnW3uRfW1u1m0J0BMv53R1ONyrNP/QLtiHlql+7GbwriwhBTw6Zuh6jGa/9N+E1bqYULvO
7HOjq1oiGkIhMqSU8DSxSf4I7LXjrVxhnDGHaRE7TSvRSWodIAZMHg9bFMFeQxLCGx/Nvpebv9sl
1LDp0uulcooXIEtnzP+n5CXHS8JN4SSlcNKHv0H9rOQZ3sIICZ9meZA3viOBHSN+BITlsT46z5cW
ILNEhMbikQbYWLtAN3+4HmT3bHCoGE2KgCYpJdg8sDr9KIOcaWF/BG8sTs1GoLx3PZppvwxJ3JDt
sx5a75t2Z+6gazh6QnI0Brx5oBJvmdz/SbunXm05VBjP3HXX9z8xI7X8yHmU0teRHu1yY0XqGCEZ
HsErgwBVVA/plztUfykt36PtkhgnG9mjw+Ew32u5UJPVgNxYLwOc0or/LUl54wirTxShqbagmBVF
cOCAWp+FUcp3KRZJuPdLHa4ppaMQeoiRURHZQ+dTQd0XJ/GSaU76ZLPSHUD/S/yHRJH+Lh6gv8kf
E9HEhh8QNHkUD9EA1sbumtw6HwSL2i7w0BEsIhNJrNSStI6SEeL3MhTeOUTy5Qn12faJlC3iK0S1
IcG71ebWjXJuSjaVEwwPlpoTXbAdfW90ADdvkT8qxQJ4552R2ox2p/OlHKOSQ2NmKR+6hvGMjvk4
l8HQjEZJpEFSdWS0rUektmS+lI46Y3+wzZPfqUy90+qPBCb++WqszRzNVQqHOu7lXE3nxM2aRRaZ
p41yXwh0VpDGP8Z9yRI1bpqhPAw0oMj8rOedYpkGAHZe2jwLTHPmoQTkFuO/yWFhHN0E/2QmSdr7
qO7g5dgNaJHfq0+rmIy6SuMQARfDWcYFF4fmgkIkFJrGdO6tqDAmgJWoFaoiEKM9bR61hym8F8Pb
Z0QgCPevMJMYrf3PaTpQxi/6bLy9ReNkQnQgEHhnF3eJq+tyEssnR9Hj5lyd3PrAAUccss2I1xxO
3z2j32nAeK5RQIVOxDrXdrOykQMWJcdr7/VA6YuWc7Fcp6/muB1fCQ+sK/AJ/GGG9QTaBnNCDa8/
gqfw4jWI9dNLWXCTEaa2TYzAl6kFULZOcunmzdXyq5H1q2qREVCrrmckudmoAHMujeBvTzvKuHjs
HU9Kh/Th2aNZZX5Pg0ZSh9Vfpolas+VKX52+nQWK6Dc6Sft+Y/rQXzCkJp1R6Vkk/C+NGb5nFziK
2FRzO+u5VDJJHi+EwciKDTrJwPMj8FXQNBq8hbuBmt7P+Q1N+YnJ7r5Qiu0t69PxdfO3pjBw1sBl
SQh4NCZUXOuJtMFs92r0KknS3Wg0frp1gqkMaBS/b1eShEiqfwRuFAw1ZO+vxtX1LAxRu/ZRt40Q
1vQxLfRvB4QOkGp/GWryGBB2tGPWrXS1maR2iZPfkXZBr3toXWveZbWlOIrCDR8nWkS5hazaLpi+
u8RaneEWq2WQ5G4raaG+ygfB0bjxQydRc/foTh9xaSs6CuQhmScfma+BPmHOpDIdIQWSfzfPs5bd
F6iap1ut9pP8hNbxN5bms165hVQ8AtAe73KhQGjp31b2VlETFwKLJzo/IU0FIEYJx5PRjo5Uekuf
obLZkMKUqCK38LIoFxIbfGVFw0Veu74MT7ETNLC+duDnpuZyISJyma2rkZXTlQtQaIsU3+yC8QAX
ywT6JfXe5JFevih4PJydboDRc5ZfSUly4oHvViNTOPfzGI//Je8XK4mrRMFVvkErKtO/54AjwWM8
vEHmalt+ID/l+F4Ges2btB4PB2AGMMrIuGrepcqT3BJwPYQTu1kEIp3EceJus+lJJO+VROWpzbwQ
/zZJj6ibuC8qmMfVwTn4A09faL93mVnWxNPxZ0XoA/OAWa/ETQTAvHf5i9vekxuVAa4emm+vodtn
7r1B0I3dANhZOLBau8gdSXQOt2Q8sOE1fdwSKr6I+s/PeFpFWdb3oRI+hQ8ChAZIdV312ngD+Uzx
8wxZCev9yy3VU2ACFTguF8KeUzUKYv6jydTd0lkWrWugmzGl6Qphn9jruVlEnkgMpb38JrABlyXk
lPqBFsrAn1GGk1t2kcC3BOzvW/CgEFDxCOfXHEqaJPt71NVCVqJUvjVT2zwo1tfziTfbd1c0dACa
KK0wDCvz7FOP1quC9noUzSW53zykHsjR1vJYvjJo0IV0Fz+qonKLbyKRZqpi0ghsVZkuOxvRzhS+
9NpoD++Y6WWv/SrLIQ+h2s4xXzC0/U1lu6CgKLVVYHv3g/2T/CQhBDBEUuLTyb0WipDHa7jzMj+G
yY3qndShxHeKERyzvoLcftuyO+TkNBd5zs59Q+oIyuP8rYVqXW6yowB6HAFx77V0iDWQT1Cz1sQO
bBhBAd5Dpq0qgyL/CsU1bSksn/Urr5sDMVa34usqW1mgCo8l8h4/BNZ3aKmixWc9yC7Hgb8+iVj6
R0xWWCf9UzFjLlgHRUzw2DchucaqNsGJ5aMraHHhq+iyYujLQtyH5MDBGWe+H/vMz4DKKNdD4s0P
vMrZPn+0ueAnbxGyNiXXQZmm164Wcl6MZ0Xn0q3vc1L36bzodvNB41B3NjtMMXdp1DOt2h9NJDHl
F//sSVtFLaeZX8p2LjD7qfl/hJo8bwreDjup9KJTL0qSfrBDcrKNtlA2j2mwf45ubdKh3D3eXlJk
taiu2nyFXnKJSqK2snrB9Hb8+o9JRHEuttLJbyTuGETwjC2yAiyPM9WavO4ToA8Ftmaiz24txnbV
burRRhafK5iXD1bqPNsJ2yEonE1mZ6e/k0Dg4YJyhJnz+XpnjO0all7Vo38oRl3BaTah7Xx1G9l5
YUCirgaUddqe257e9kl8EKhivy9S7HkDoKBWgXp6DaZx8cp5GABnySiEZ33b6WYwAYlXGRc6NGFo
Z9/BVrAo23mGsM3k4gbPaIxfIlC8ioHIINCfreZQyy3XHgVrJLyQsIC0iCjQCEB9xG6ubx8UvktM
jMqZ0zD05TDYWWRHkH9M6SfTMpVewKOmfr1q4K8t8iKjxoL3oKYxc+827jO8IM3AiSPQKEeMoLCa
Skffo0NqZ/Vmym0qIa8meJtfuIrdRdANPD0TV84nWQ58Kr4GavpdxxjuVf61ocjnEJ30s9f+krXl
ZBqZXw3EF4a1fgKHldnsk6gNCw1ZOy2tIhfYjk5/d9dBn27mQ+OIt26hy4fI/xnl2wsiUZCnyAdL
lH3fc4zuj7gRFcUHLsQlMUCcK89jVbZmNYuyk8KF9E80lwvOvy9OMSvdHDLns/6t6mRE+EzcelVp
DcFxsXocU2e8RN9O8LsrLQGr0LpP3cpfAC3qMDfWCpFKhs1FHIFTIlP4guGR0FI+FXnTuPLk8MPl
jups2XzpkjcFZDuS0T9fN2LUn+pgxwIXVcvIPMIkDmX92EsiIIxsaUlcL5uNnih/Pt7iOgXrorwI
XDdH2frcOLjGz0kNX9rU2V96xJc2QEui4q3IVgG0WohdKjXcweH85jCVvXq0EjGJy+3h0ja99ykE
K6zYxkaKYDdndmx/jfTHnT8hz+LPA0Sz7D8kcctQ/+KuyqXL60fGim6cOanZCV0r5iCGb2qDrJgh
gfvJGa+r4v155JIdiGmAU5OPD815398n/99e4lFq6uc0tHuVr6u9ycYPZRTbO4zvP79tDl7If1eA
F7UJ7XZ/4/ut8Uw+Lh2Mzo3B/i3N8ikdmhwvUk8pJMgj2KV3vKDE3g6haAWr9oUwOfe7LG/LSrVM
TOR5A7QWypm1y6oRTY6GgzFO9ZLd/tUE9cPUuj2sVX7QZk/rfBKJLRtW4pRoxs780Fmmtyp5lG+C
7OmYCIZpcKXHQlB1lKJAi2STcCNghQOG87yv4c3otXCAvdbf4/NEQTGavhnjdtuV4WAViTnNR8GT
hEYVr7i2ZcA98xQYVVwAkWMum5NigFxLzCxixIw0P5tQUsbzv5OGF7Fbt526qc5uvdWjwAbD2yiP
dD9ijiIz1CIBTuxVu7X829E4ngSHOJAMOUJddxBbfS//9G05WW/bRVyrvrXbedXYUgx55taFDIVU
b1l8toRkr0Nziw+ycBTr4sxh+aX6km5AIEVWpJsahb0BifQ/WJSkyZuO9s26TRAG2SUzb21X48nT
upztXIIZHmM7cQLGweCqZ5pPUgyhPrSWu6cMLZ48aPC6T31+ydR8irpBHRxfB0C7oTFQexqP5isb
HWi2NQVjEEswOaoo/s2zn7Psybzeri0fxMJcHSri0koaSNNTZKPnq1mPpQ+fscgqkGUMbiOubG3i
ePQqyeq9rW7QYeqzkBym/Fmm6ux3sqL1jnDXFIpq0ZLh2p8Ght/Gb/4h0s6WAeqWtLq+ZHGtwfBG
nv05twbASuhQfiW+G9f99DsscUHhNaP08+9mQoG11kuL4ZnoFcDthVxKrMp7ESFE0Aavsnz/BQZL
WulgBzxnab5hya3q3zZkw2+Bn6/eMlJ/5wTXyn/puL/j5O+pXONSpvL+R7lpo7majJYH3pJsXttE
zG899iWnUM8QBVLDwqqBsR8h7Bc0O11BWd2ja3rlABbI9KUdr3BPUWNo20D3wEI3G38+34mF4XAs
VJLLJw+yc/Vp1d7/6gVxfNZLnivYgkzN69FeEtI46xSZJlbYaYHyBp8zFf5J8Cuic843j2HeyA+P
hFFD+Sw6XV1Zk2rVz6F/AEn0HrXP4HF+CwWgGQRxK0J7nYAW4j1UsnPaCh59Y2lHkWcUZQSGIUps
hW3cxfbNX1RTWnbtbJAs4DZJio+e2QcTE4hGttM98xcvAkraV1RMHTVP8GpGxR0LTmJORBdikYV8
r+Wm7THX/7fIW99/rl36ccImomBX6KENhwdLPpvY8H8XXU99SxWsvfAx2A5QDg78929OzYHtue9S
OXZa1PDKqpHMC6yltYE6o/YSkUckUVoPUlLE1d1zmUdQkjk4n4YgglAnTJuZjRVnwCVz1osf0CGQ
6gDtkex4AUNJedVHdj4YbFtwBjcJLCOGBBEI3tYQXNSzgZFpH2Y79jfRFlGN51yH5KKF9ZZioa7a
fACndbZnG7aZzBOyKCcHE79/hKD1zRMusIG2nrYxk0/R+aGJMmuzH2AsxqZbp1cQd1RE3RPb35LD
bQT0PXd3kYpzz+JVnPUvkqwv9IH7aOnxVTc66sGCrHHSfoYotIwQiVZ2AihvUz1CfYug+J6Nx/de
pZi5izYxPJTfVH5EzlvRIAMymT/B3kFlMLSMFb3YEfdyxqH7uZQQ3QIpTOV+2lfrBL5rrz1Y2XW7
11AEoiH/z6tBJp83K4L2X4qGC9AE7KATaFWzzlOHWyeUUTTk9QCl1oZ69MKJQmjJ8ntu1wfKBURP
eBFPW/cmOkwuBlRyM7Fkm+oAwE4qf2MVHWNEXXhukE/Iy/UoVMFggrPohHTMfNuMG2jjhLf3G9Mh
nISYkR1QyyJTpuG0CCJXEz27Aqt0E7QumC2qIFQbSeMP/jh59VK9rgVVt64/xr+3DDzifU1q3nT9
HppfI4F3TW9uOH29anNK8JntlUeEZVFSd1QyzQ9r2aA53ZOeleSo1CFsw7vR24H6HcABLkKZXeQf
+GI0MvhhXD/RkT8jmiCcGXgzCS3rvDEdLuYRRbinuOyyOKzIYYJnAkkh3VCh+TxcvMpLRTEOiiOs
hk2RK25t5vAu+cyIlrw+NJy9+Fz/nyeSnyaXkBUun4pvK8M1ez1ZzpRxdEV+ylAloOB7Htc+Z5GZ
JxqS0RJsSHhuY9RrYA4qtEnuUBvrUHwi/eOlEw6Z+Kdqr9vrEY+dOnUM9+w4MgoZRfkzWHpaRhkY
StNwtIT1MhkyObjQ/CuIzZiknQCYsE+vaiGOHiMyedI+LpKebd1Giq0T8z5WlcGERIYfDUFkVm4u
Jt2K9zvP0GBrauNV8d6yZX/QQWDq6Jc4yfAidNO36TVBZiQbYOJHLJ5+5vtiGu5pRGSN9JZf0pZ5
xqseUqUXRvJGIIosrNcW7jj3PIJMX0vuefpDWQXFPMPnViN9wHl3fib8flL/GdsuusQTzd69jeLh
n8SGwYZmoklG77Hw00nQwB1hNJ0kF1+12haEPh1IzF8xKFHx21734ygMpkJk0kqvJXMYRH6y2SpI
gyE/fPankjoiQAVr8ZIpjkzU/ZBoxYJmsF6e3c9igyoKEdOPh5v5O/KXyEEeBT9hW7/Hz0MW29RE
q5ewLkQC6yJOQ/WR+4TE0KgUuAuyjFZ0KrZ4VgtTgY9DP8R/S4PQ5AstA70uVD2FbmoFeXRFmxA5
yaIqe0igIILcua8rReImtZtvBPSg3kyg8wgtDNvL53qY1VD20wPvyiigmH3mY+C4IZ3nJ1slU7eR
8n5yun9YBjbwTP7ZowL1h5HfkoARYZsS9r+Sqt95D2uoTY+x6evwJXGuAsJMf/TwSkYEvXf2JKKk
hJPSYp40H6+djYFXy50SX1AhgKTQwJ4/dtqfTVi1T+lKUVb91n6MoOh/v+jdTkn531XCMciVpfl3
Equj1JOTduHNapMqD6f0o4e+fGlHyrdDafY/PdtxYmM7ajpMb7FQY/7VEpO2ZOjwtADg7eMXMhMG
DoNR/4iqDvgXR+KsTwr8sCkDBu1JMaPEcRfaqW5NRj4AMCnakcRbTW8et5tIPMrP9f6FjOa/MqI6
1vzshiIIDGWbCUWK2SUfF/qAV99lDTVl0OMS1iW2eWBHQgBVH7ivAL7lmKd+yJcmLlMyFFW/5wvr
MEeQbtxB09+6Ehqf7MbOIWLHRrd3zjuXlmKiYZGB1Qp/XfNHiOILUTKQywyim1qfMbbiYU4TJb/r
TC7lHwhMXEj7K1sAz0hu8CroY4g7aVFswicr7HGyBKCJ/MM61Y4oOlsHpJi4C7HH41IAqN/rCaH4
nExFwY4wJqb+POJiU6d9BHUD1sJhiA8egvFgBAEzGqIjsLaFyUHW5q2xdpzGlr5OfsztUkWYqauF
eFxTCl1e+fwy9KAaFayVbcoacqlX4rJ1aDjuiQcgyUAdqNHq15zEQdWWhuTfCB9+5XHx/pL1/lMG
uuS5DF5cswuxSFp6lDAP1n6pQBZWef/E7dPoOcrdw/IIYV9RlAgyN0QPWS4k9QAOvuBfC/ecYB0H
lHZ0Y2Ssjp3OHGYb7aVY8+a5dkb3kPn/RPpqKBtQt5NrH5JxiQ00kxYF5gWO+mtQIQHE4HmGtH+4
NOYdvJ2AkISrQXB/qghBf0lgkDTor4GAJVHaJ2ceF5RZ0pU5ISmq+LmZjdUf9JF9E2eIJQhw8T0h
Ljz7vIeNwo+VocR/a6W+pQFKWWZurEm+vthW34LlqSjU5HuP1A9ns8egNd0ZuyVFEp8CPfg43s2L
WWdTsDD5gqY/aQAZKmO69gix4SHPowQEVj/JYl1ctcnZE8SGLS3GhgruxQPRQtSW1VDQcccyOkqc
AYjDN9cup2d8dl3U9ddQ3qBn7vXMSqVPQsMt/N7StiBeXTdNX2OphTIy+ZvgOCmDC45KR02MKDgB
WTXm3G0nYoUsug8egieX/j5E/h4YufJxelSk9oTL/upIGhGoo38oiZxI1t1kaJ3Fak1woFvSo5KE
XqIZ4+IdLex8TLtS55rzoitgRH0vsfYGhlEhnFZPd1+wxQa7IYWDo9dSMOjI+tLGDlsySJ4bRAgD
geVDLvRwCHCk0+7CLZSkjRVwPGHlyIeHBo5ALORviQYlqPDcBLNNc9pu7DC9XlTfSAxjwFt6qfLU
6CF1+Jtil+6w4kdD7wOqAlo+Qx7juNu1hMpCx9fGG3wS7/3NZyqNPqy/HqG8J8xQ5r4mvGcz/quW
F+ndrHwb596S8dB8Weo9tr9PY4u8A4Vvhj+K5f6eHHKqCm9qWm6Hn3rLn+MGy63xkNFh3EZuXbcv
6y09XwXbpAKW8lUaL2m/C9kVtxe/2959aIr7Qr6CE3na8qLDdH9PDFlAbNu3nN/gptgjY2h+FjjZ
+vpnFMU6VP77sGERmKzGdoduR5j8imyBQOj+M8MnE0u/R+FXGzjQHILiKGgQTmMqgshPKQ6MDf+I
XC0Usj5XTReUbLJLhcRyhA3OWL2cGYeBAoD+3jXAfLHweMUPexW6j7sgdEzhTQt6uqDSJm4/xX94
8FmAF02DaaVsxEgiJpyC+xKxUiq2m7N+1+mMN+SCNjr1LU5NJdvfA74CPoVZGg70cP/ZLqtIpqLk
BuQZvjBCAIss8v/mZbEbi/ZeIh/zXLWM0qV1akViWf9O1YVvO5SisdZKip3M/Rw/HHVk7/iWn8TJ
BRM78xGrVoFgr0nZUSnMS7wE9mnnYHtScDlX20QRkStF/4XI6G8L9OhhicNSuwAeDHNUodLgNmlb
R0Jfrkgn5lGJTs8BvCbat+yFILnTb3KtHJ1bs+rrQH+grdrigd6RVONDF7K4LASAI9KUl28Am58c
23inU/NCF69+MxQl776Nm4wT1Rs4iPPwBanl7BIjtgRBnmi4Bc8Dt2ftzGwlt1Nnawyq0Qt9zFi9
ab2dDlk972A0e/EdQ7Vgt5vRaP5FQN2j5tV9zN/QbFnumBuLb6tjjhme2slWh46uS7gnjigpM/CF
dDKHH33afL6bf4vAQsk/8aMiCoBZTC7AFZgIp4eNuC4QUqmbNsF64W7EpXBsTLTe07Jeo3ZPFba1
fO2ss7RbVxU8oDtRrpDLbB0cdQYn8cMuVxPIXscfEdFaAV/uUTkW8rc+dLPmYPCezqT4U0EuDKtd
5XSIO++5oE2bk3Hn+WdbglpkyKWpQUJhcbbf2SFm5F+HK47jbr37GzpzCvaCCU7duXFsSEqViOEF
41/qGNU2/zvU4VhY6qXjGlZpbfwjJn54uk8ssdotN7LDgBNdRkf5AfqMD6EKr2MOB0GLnkYdtuIF
FZIghai73QXzQj0/tYqgM26+xa6xffhauKSzRTHRrDIFQ/EEWtBjsj9F5O+OzssTRgJdxir5/fRc
3kXGCP3mwjH44b/kdN70dITetYFdVx6l/JEv0vmExFLpw0GuDplUw+0pjYpvrBn3MfaiYKR3psoY
Cz8ngq0Wia+HrEATxx7XBXqXgfpzrh8Da/AU9H3HIJMaB72k3Bc+gm/KD+344foJHRn+JimQaY76
vjxk6iJ3CObSq0PybgAH9Nso1sENA9LZxF7owNZ3BQNEh3TNAfahq9maSgNHHahqCUWi+ePIjC8N
nzUMIQ5+EU/a1rp3bRVQwokILS3nTkjuG6OF6Jm3RtZe73wjlCxT54rxGK3SFFmigD4NkA+rKQrl
mU5UJXwTTsZEI+47YkfKTf+i/hFwkKNcvKlsc9IMGOuSxCZSgJYs/N+8LQwcRmgmfpHTzxPsRzjB
o/kLlcn4t4XlPWkNZMWZ4TCYiXjgPab9yF/F3sUQ42uuxKJYEMPrWkY9IfpYzlmxSpZIQTICiY8C
BS2qBye5tkZi3nwfQoZI99w5/xNPmDckC2nsKt6/sog0mWgdDFWbU9RfhSSVX1emUpu0K2i7UASs
tkGDQzwBuBfcm0jRS2yM99OvX99y30golwnD9OFqJw/Q3eBbPFV5Ivolcad+CFveLqXjJpko15+7
IZl3kDJ671fU2MrhoIBy1hAY2HBk7a2wLH1UaOJIxl7wOjQe8g8hk2vlcytZ4gqgG9DS0RW8LDGO
b5DkTgjlGbteZti6pTuXsLDDGeWnzo+mFjFxDFA+PRTLydNcqGPMiBbSDcqEFWfr51mGbzmlrahp
U8nftFlBfYWY+vc0+bCJ86Wj4CdnI7W1/Cp5jc0j6e/zQxm1jpXJ5OZMMljcibLBy5PzY8FSn2SD
aK25Kb/QZ+EHYphTe1py8livBjrNspdg7kmaSJL3xLyAfwBgu66o6wAe68uHfW7jd3RDRGsAA5vN
iWXm9TP5iGUgCG26hxV+q90EfCbZqtPlkq/eSwTvt1rm2wEWeqobVlT1emLUswLptF7fpVMYkhzQ
Aql9wrkF2pjj3NokpVpZIR0q4JieL+osQB1gvoyp8gUN4Pf2/5gMWMzhIqdLiinWvP5Krpx+0FPh
5GLSuGXfhmOD8lbajqDnZL6GoK+TU18fCdkiC2HebQb65JsmA5DWP9FtXkRKp1WcKt8ylty71OTH
xLgXEUBFDy5HHOJu4f29b8gyB1AaG2n85pjVonDy97JxvKtBqQt/+Pgog6eHs4VLJ8wzZikr9pic
ubRY8OyOzi7MDcH/yR7YIKm2tKlhFh2gNmrkFOEanHK5L1gWt2Pem0HoYJoqgrlSG0DpfdKS6cIA
ooLgwwLSl3HkZPALoWj33OpcJHv4VcpLTrhBCQh/sVDADe1aEoLgeJp7g+6R+DURveQhqw9aM1Zy
bkl6GmeGvisEV860Kei4OucuerhZoDF7QNBZ9GYhNs2jW9lLjR0pUhLMtAOGFlk3XbbvVDUcyJIQ
4DZFeX48GeXYWpkRKpaEBklg+FHJai9hu/BszKKWhb1EjA8XFYpmN2eMKCcs7lotU9m/egRBHPIq
yZEeiQvA2ojQWBTH22ISmtq88vuZgDNDvDLihCtGtEOfFVthTWvOz5w8pFmANaJkzxMhqQ73jEAW
4ZxsMVKWSxmAK1MujJLISsz6mad60JwIhRnZM9LM7w6t0Ac1/gIbQVQzQ0bNl2bnIw9rGvMQWJ/j
SLrNjPSL92WpTZTK5jnKu3pV7N96amvdnuINXXfUbcqoxGizeUXaC/6RoJEbuLsmQ3j3PaMwVGVU
cu83GlmhPEFHKenjFLGIELVpvyIdTXFZpV49cJzW/QtB7FEjvesFjHqndenC5xO7va3JbaqEIXYN
UHjo08liLUmmz7behedthAs3meVpOVmK674uLX99Qv3fcmFVyyEhTKwlWEEP/tZkLkACd1docIHp
GAfC7zLlyidNTF/Gnpg0/JyBaGvtAgikR2vTpOAm1TfFq2ufE8366y5UJ88eUT1ANju0M2927mS0
InwBte07HcF2VhNjuYv+34wz6I0dcQl6rh4p6uPW3cUuVarTfOS9JoCOCDTxIHu9+3isdNLCxCp9
fozaYLYrmQIJmukB2Ih05B9pR5jQdVDXuLfCfdhVU5CV2YQ4UdeTyTl6n2UbjoFcHfYmxdbJAhjf
gZorCSxuVhTg6Jx8F55O7pVp5Zf2OMEsIg1EWdX/21uh98hwJg8/Ci5EBdUAVVT6CSD33SXpaBZv
ghk5iH8ADmvqZs+aaPbySU6wxNz68Peq876RhUgX54FIHxIGZAhK5US7uEdd5sR3NbFPY2gx7VGV
37cYazKxVkFOfQh3zWyfefLgkb8dAFviZkNnFdt201Xe8uShKeu6ypV2uH+SSe4MPe6VLRqKKUVA
7e7jdldzZ4JkGCyfLy+QHhlxaNh7U3rnilCj4xq6ax3HWJ3c3EreKCrcMZN4JSayRYh5LXAVNRKA
MZPW913rCWgoBEIhfQsdKVyJ4ExmAOKnrlMg2yYcoICWBsS+XlHuXviowa9/NdvZvto1hHz+GIq+
8588Ru6h5wEic+Jh1rN4gVE9Y0hcGVLkOusbctIZI5SWOmNhigpVybKukQaryD0Gp1nh6atlycUn
81PMXETdHd9rzQ/ZyMQr7ugevr9PXXSx81kVNIIkNFMZ4+OKctnNpu785AZSSbwwgJe5wjOs+nf6
5k/nyuZFoFjbGfwZwmnlDiAW2ijlL9PXhiBNMSFqFAvQu5AWMq3oj+XPc2uD+NctBYcZGX/PBRGS
TzvzWeNO/9rLj0x7iFRGlXb7JtPUxQvDJoux6Snp0PJjNjRWUUuyNiZV9QJpA5gR+PTQV6xX0L40
lkO7HzJNA90FrYQDnIeGu05e2yD4G/iPZ2oanXhwDKQiDc4FbMz7w7oSjmJvfI1asqf9QoJZVN7v
jvu/DOHBXOIQYIHM3UfTW9JSjQwBOyAe0K7rtPV4N/gpfQ+T+WzWuNArJ5Rfs7Em9z2DO4E4VDBw
TD6v6P1YlYSKp9QdP9GX3A+GDXbM5SRpPFxhVIX1upVVXCeBItzSB8K005+kP6lJFbP9g7b87cT3
Y1eM1+TyUXLuRuh5kXHGGyPe2D9ZAxzR/zrMXyMm/1libRYe/iSqSmTFalBDHznUIpKu5b+71tr2
GrIPElZKwiTX/JYd5YUmFDImyI/OinH5TomVT4L1fgjlA4EKTJo+fmxblnfexDG53OUu7fz0QAOT
M3zUdHDA+lH7fsn5VsHKlI6eH++8yElHrW7PVhd3FXAGaD/LvpGe+XkTiGz/2Tm6S+k56JN341Ti
C90pvksyKtkthbnaSUirsgRcKsTBA+XIwXWwqtaN7FSCfSWMRg+mNhxrorE5CWwXfSsqmwvGg2RG
zg39p7toGSLIg/0FZBXZvnelo9uRXlZu+njXMERvMeE4MNMcPeRCuFCp4ItvC4jy+CNo6vYX7uSb
qIDaVFvpoTSWtbSKlbLvJqHLe0Me6/gGFo3RQKPilijhai/fPtlCzopqalLgaa+VeuqTtl1RYZh4
HZ614Vg7d3xwRPqM8OMhpJ5GVk8+oir18pbXLIBPqWCtULSoOlZK73OICrop2+0ozVUg52k+CMc3
Tc/41hmkSXPJMTaYyuoBoWjDxzrdsdlnifEIWzo0o2hZaoASHgG+QuymYaI7kd/wnD0hEFjBpFWq
6cKwKmhmjEjXv/ILfZsNUWBfCYNtSE9G6UF7rvxCl7tqqfSFeGs+DO79bTJuRy5zQcn09T7tE6kM
/XTLMMKhY5Wy6LMZeRjcUERBSD3yNl87/giR9T0+0wB0ED5ZTnKWm9+jbKZxQEbZ1Q3ducWL9nEk
TYWrLxVZEwS8Bm0BAvFyBz7TdSGAkzhzPqPcqs9m390A086k1KJrsioxp8ZKPSQCbyTWDyM/c4T/
4AH9/nE0PVq5OPr2CkJaM7zhGpxbDB7zwoa28CuyVLKDgtAA+z4nfyjnbciqENiV9/Vpdhh7gf9j
ubZe1ZBbaD/BUUknEhUuBGR9TV04adWwn7cu85S1K2lAX+IV3UL9xLVNOLjGjmK7xM5etc9OG0I9
bL9l2FqJx7FKYrpZwllAxa1pmreyYICFVPbJIIdZC20Ewm8MFv8LimQdqziOaUkYz5zUMkFd7yYl
aUOPxQdyknhGb1d02R5HCcHtkYL/dydo4j8LrS26Uqmz+Eg1B73Ovu8i16C1/qV3qlC8EEuaE7Z2
xK++bdxO1nUwxbgrQb0HLUHzoDIIUZ4mtDRghR4bGLfJZmoc+OZ6/Kjxah3ATWybTpL2yWgou5SK
Ahpzk/gz8X5r0CTh/N0Q4Q0tTBWirEcUfkOffU6ofOFSXNlrP5pLvw7U55Qd43cliou772oMQj94
FdELrlplxOT+YzOT4Ebu6lGM9oyiBl3ioaVLZ93iL/yaTqRKoqLy6eq2jz2HdB7ZUrP77M82XKlb
t0WEYz7dSYB7QjTRRt0nMam/ibljzrmshROrMZz10fgXbJ9ubKgclLJsGGanThonQoCPOGJPIYmp
YaNNKV2SGkL40j49T8U/QWthh/VG6UbbkgrEvyiv0H0D8iPLjNM5y7k+N4yme6FNhA+5EY+hZm/g
6ejll6t7DhygEHtLpX98bWqp19zWF0XxjTzE+ct2cYEm63c55sKzH2v4pefHnmLH0krYglaRuWBC
fT8I7x5u8bqJnEVHa+m0uI55//4oX3CPt/yHOje2SG6IY8Ig6v9UC0YFSqtm2AMTAbRzY3674iYI
cyvHd6PO9ljE7+DAcq2XG4qCY4LXVg4PBKluOy6T0HpBz6KXMOvylcZKfJKQXguqFqTAMyDB3DjO
DXnAObQbbJ9TYWPIhDjMZ/1H2gGbpVQPIHqqv4Hn05MuPQlTs7WCeYmLsdS89AraR6DJf9gRcYGg
X+9XrEWCoJZ2RrtY3JyeBnrDlsVn/+5IRuRIsWH55Rm8+Y2oGRnThC74xXiPdvRCOoM2C0IBxLlA
Rkn7P1FmbPDT/01aNW2hncCk0UKEnfVB1uSsEgyCmVvdFdhFU2g3oji5jL8ZDavuhrYuCuQDUpaS
IqYn+82ajQjI+a5Hy60JxNXtWxR/EppPH1Qzop2i6J+Of2Mt2q5U30HKBlzuYsxI9y4emcGRoJDD
ud7M9tHMCi3uqB+ttsgiAc3IizwW6NAFbdZedbGOYH8LXWJTRIyv1UqBbmnIPluyDaVgiaQeyna0
k8sc4uGWP3v5MD7kuY3KS/chbPkMRLb2kNWlKV7xSrm9FQhMkcaa9Rj4ujElhtdZBhI8f5ZgTBM+
ITz54NHRw0jx/755wpNMmwPMVFCu456fcIRNgJFwZhCofdBZnnS1RYh/fZ4gRv8KaD0M33x67UeU
RgIEJcOCLdER+rfN6kzp7w0V8lKft3WAwLlPY55qs0SJZ58VEqqnSrHl65ZKj4lOVj7CA9S5JXd5
Gm0P52c7bPQsJUvvlAkND42ywoTAfwOotdMUIYNoDyLuFRNl+royRK3mp0TO34IJbipptDrPd9aW
tOrVyHpzPWxlbFhyHtGYCydwori5fxyBwrWWYm02gDnR3dEvjSoXn4f1uU1mfSsdUXn2zBL7fKnF
P2+eq8YQlZ0H5KrJ2c02qOdn9xEfmlrjbaTO4a7P7P/WMe28VdmbL0rG7ZH3BoK9blbx8f0ddutJ
lPXgSTYRczJ7Mmphgx6eUngpJ1RTP71ZYwWVlKba1BU4Ta93cijxyR4dMDbFVIaicNTPx7SFEWqV
pUlYlO7PBIcdJFuFcyUU1rSZukJD9gG/BCWoPhk6Qh0VGYnCnECzXb0QgGJ8PIQW/XuUjafebrxM
GbdcFUtezRG6LrPPyAP+4loZFknpNlmLecvCkc7wQrxejud7p84MZwlCujdgEKgLdGg4YH3yP739
1seWx7/mA/RIMHgpXCcfteglynzMZ4JRwr45wo5jRydxh4WqPL1Z3tHD2ajK7eagh99UWmTxCV1+
4Yr1h2eL0F83qSA48OzZxlDGVoUgg5EKRrjFs5PQQT/e4rJ6nJVCh0vpFQjoVF/y3vDPHDgSCmJv
jertxqmzVQ7zqTHf6yNZlVxOU1IysEk+GeUu/abti8ApeX/kASdnBMlgyKpLf+INoFjn5I4NLEKh
vh2P5jSlZ8+f2eg3PwZGDtPeMQi/ozHbGBMx2OefG1rKJZB3Qg5vom89NPE3A7PhhGqclRqDbxoT
R5wY405A+F3znm77MvLOd7KlojdHYNm/ZneJEa/f/Yl3V9us539SH+zJGR4gNRdvTil3jHwHGSB/
vtT47icXHbQE2OlUqnhCsMjnsSSrYl3jyKil7HBvhe69DJplFwq5YyTdS8LvcMYsN7YNWMwyKRcl
FgZZoYbQ7Zwts54SX54caLdhdfV++CfTQRYDxlhmUyL2W0XrFzA17S/TNE7SnreGcD4ah8Lb8DC9
OKUo/s4XkYwAtNUD4UzMkwa1gkr7WcSMt71w8G0lQQhMu9fvvPHUWgli7eg9DPXRPqwwqtUp74xO
f1rW7VNtybvHrNNnELg1CkRkjjMvJyO9b3RGLWp1snXXMDFcnkR924eLZ7H7WaImvDIKys2gHEXU
ioRtg8cBiKLnurn0vukwqWBeiWP4LYr/hXyh2lKzsvHdDecKAIUiDw2UJhGcN8knB30OjJwjWd8J
BNYSuMHXLqF9M7X7tX6+9iOSPoqdTXKKKy7VKY5AqztZa31BvfS9uJBpK83npYGUcp3UY4CYmqmT
xAst1iz1Jf9Z5RNdePu8iQ5G3YeBKtmQnq3Q2jEl01R4DuEo89ydUzORh0t9HeGHpWn7kp6XgcpO
rKMxJSzOPjafx+23yWceAitWMSaogWdmRwGzDL92cib8BNZ2pnFIWmu4uD6GljwKCXZQPBPRANgE
f0gnlewIGWSoPLEsEau7e5bKyOs31sUAIA5zQRF7ALETvIMf3pLklp1QfusC2OEl0WC96zXMB9+F
dd3Jf/luU32PtoHF/JLWWPIXV5KbJA7rGbLLVjwTy3ni5yVb+utJwktKn7ds/XfIdJNLWLyoEPGF
aBva26DLkqFO2ASYwgxzkVa4Pk/rE1ZShPOve6n3Q0B592RIZAIJtkVYnsIDEEHubE8CMwhjiydq
CCs8AN1wCiCDOklUAMwSD1joLLdB4oNntNKtlnkkg7vJ+z7AsIK+A5LsMGIpY4lJaGDSvVOTBHi3
zi328LC2vDN3wlHc2723p/8o126Dklj2GRj1BgYHFG17XktnTna/V0NRqCP7pw1y4+FDIfGpaxYh
IUpw4Nu6w0BmPHzfGqnF6o2ibnwlcUKEb1m+utEf2DHE0CFiwLOkzueVU6FPRxQ9TBtAmvvHWuWK
Yprpomsq5JclmmWLkOb5gzxcIIljQeVWmK69VKZyaMW1MbBW0+ttLAZgSwNB7ccGewkHkjo+L+dQ
jSTrg67581FiulslqLUwzrfbrMpaVCrDZIc7Ew92klMQ0p9XfwqlFHvVIW81evR2Jm8JDrT48Cd8
fv503n5a1xmxtoAMmkq0yDzdrNLfgtlWPEz9kLNzWiNkZG8GsBt6z4CZ1ADd17iCJCzir4aJvxH3
ZCsEtwm/03kIFRs5e+MfXij+L1EY3a+0eygQlDQrDQT+/RiOw095+2vrXEtqxS9D86o79ZC5qBlB
NENmXl9dPcIE3LCe5kJ1YiEAhmns6D+nQzDTDEToe9Ne8NHRaaLyUpsBbHO7jX1Hym+NLUufNbrr
X+54a0Pu6bIfPpP3NWRGaadhXDmdj6VSGA9lxqUKF5xRYtjCpduLVpZpx/+BCOeQ/mu4wOjG6aMr
iRTch632BngnQUD3a01+CRJECK5rJ+s5uMHc8h+xYUzStwEA/9QgIF3goWhTWsHNFqC2Yem4De7y
myBFzls8MdfwwfVy+YHEDR6xrPJkYUPtJt3Afw+ZEtfPmmNDYcuxIFIjz4ZSYCEb4I8ZBNIC4qhL
n/aVfLjMHPOugYe3V6/wVUQg0740MI2uGIy+i6IjUK1LWAkMNS1ClyvZZAqMQkJE5UMh+wfmRHl5
3wJ6QG1Qx3K+CiEWQke0Xfzf+2IFGfnr4NBceW65X5Jt/Xhe5WYTPax/e/5NgvGe5fnNbhy2HNsH
aaPagfylCjK8LH5rINA5ynEXmUDV4wgZ+Wzq2bVL7ZECjreiXa1RxF4tHbg6aQ4EHwx2kJ/aag+S
ZrhYjUFhGkoKBGbp1OxRlPT5hLgVs/jiamay/76MnxQsFG+tB/kUE4MVdWByJLsEYw1PYMX/8rV7
+5u4IdO9VA3i2Ei3sL+0ltUew0jYTGrL1BirxSFe15Vs/7gb+GvLEbAZMS185wjGaFzOZh7+pMwV
kzT542LnXPRA3+qQFMp1R9zma5thSSBYfOLNfGNchFwGyYWHE60Ja6p+ZDcxpI2QhoD51q1vdMX3
JF2dbh+2ydsnlZCCf7FFHtI9BwbMktPDdh68TW3rZTu7IWiDW1Z5Bps+Hp5MVPFqh+HttH15vP1E
8hzRmcH2a6yZaRJ2krXxeJ/P21Wl/pPCrBMEYl6STky1aVi7xBhwTsssmysIy1OQCdBFSvP3YIH1
lYaWyH+Q/LGHDI6LvHKUnp/tnyJgL9sBYEEUJ2C4PbpJNbyOEh9OF++V3vz8+6ZWxSusyEo9/3MK
9HDMwXyz4zp2Xcwgz8Mm/VTShzdaIdJiO5NSoSsU6UPqPz4WbVONsUPTpL+TZucsKl5cRvXsA96I
XQcYragmfPuJvXqFLSVGh/ocQuOq2kPNnNXzG5TY/6sIiRCgAwZDGnJtfkqlHDKUMFEDXyNfiyAh
IKY4SLi33ei+vSIu1Ad8XcNmEHhC8pmii0K/mzTpmny10B4+e1ANe/YuakTt0mi+3pT829ykEMjn
N3erkOOQUIilKMsTgReKwGWK/loA2gJL7/WOYdaySxQmdAjWXC5i7EKm9hKI215GmiFVVR52AWny
ruzxpds1HGDCpIQxc4FBzlyT3xEUPXntB7PPT11ovvOBbzaurmZM5OscGByyuuWw4aTlnoi5mswA
c1uqMDd7BmZLddQJLTGrlZsId+K4xJyhRrP+Fil9UNgeWUXyWH4D5cLQFnXvQJCPjZPWZ9/DCJhN
p17Hq3+/dITQN+/D6KEeJWOQnJadL3RcHXE1a+NSgS4AcznZMOTZ6+UL44n1DbVatUznGDdWtFID
mPDkOBCbw8F6JB+VWgcmzn/mpSVsS5PrCResx5OQD0LOc1NpGA1wIww4iCE57KaEaE5UUUXwaUHp
Pg0ccSdp6G0XYqlvlp02cXPCDty960ODTkeG+0cZ8t2Me8IVMMoP+OBTK6ZuTv7/LioyCzvW/rC/
Xh4LLNV44TFfJ+epHjBBmknztTAQ3wNZjclk4NbqxpVIQ/VgRI11ZIO4IXSbBhS0kHJZk6p9w9oX
E97mOcu+79nj7FG9egyf4GN46ku5uYBUNjVtFDrwY9jV0UDOkuudZsgj+Wqv/gyVSKvcBF5Y3fGc
82K46jM6Omg6lgapdKwfJ3/rMpW3JMw6bpE/fFGCCbI8CHE5tan0VWr3OIsCJ2dwyudUHAPI4TUY
G+C5j+rMf6xevrw1iPpiRq5dQUlmAwDUp/VLh+ghtBb0p07iYiYljOA64EnpOLBC0f/XrwN/+cSu
ZZnKfqYPf+L3WgSon6BinKlEQpogIbqY8he1OGAnpH/c8HRPmCWwj/IDPVQUfQHJy6qKyEnNAzMW
qnTLyKrT++Qo27BiKZMysz4EuN4TYwpWGjIYC7797tciCqIndanrDWgeSRzVSWFppoN5MYQLzuWd
+ADp1+kwTs6mX66jUdPdaiLUMwH6X1YhdtaUeSzvWVNVgaRjZwokOMaCoOJb25Mt7pf2ZH7fwDYB
a/MVLrYiluBCcQb1l1e7fnc0fh6ulzacDZfqZpcWfidP0zFiYsvPOBgEBkQ4ySxccPxWVThu77g/
bGGPG187/qEswxDtEv4G+in4B6q7rgeI2+cpzW35UOiFd/IpvooBy+k0ay+g5PQriz2t0NyfiU6w
d73OmrvvvA2Exux5qCWPaP6DzLTN63Suh7v7xgR947ytUmDeWcJ9oYFdTERsejnICQdqZgmos82Z
KoFzkt/EcdT262O7SjQifKNvyi5y0mVaDMmQj5bmOrxZ8p9IeZnHnkfh/4J3I5gtIXSFJLeTUAvo
Bgdpn6IiEckVh4/eG0DrQEx+1mYFZa3AVsJV1F8BVHfDQiwCxQe/MeroonZWaShK+gGK9e/aKmpY
1evfNT+kbLQsae969zjhBcGC82OdCZ7slu4OpRlTNUzd3Mdf9s7wSBbiTeRI6ZWzw+O4o29t0/5H
9se+RIHz0JE/nlapE8kNn8D2JSQTnxZpj/4uM0fXgosBGerKyH5FWjSQ+AdZHXssJkb3M26kAaas
zUAMyJQGHLQR+giDbposTozFC+arERUdu7HA9eJ13VW8DLByeANWhiQoONyIisENt5mPfj25NFyw
hHVFmDK9NRj0H+WfL1fSmsOiwjc7HkUds17W9bwRDnm2tXvpmOO37H6Pi+90avrYmGPLYUlkT7Cc
KLSgppEzPM4nDNEbcgHU/omUaZjUDnlBj0sYY6duD44aobf9d/QDCm4tW4dD0YHa/yQzpCC9plDE
e2WJMO+94nACdDq4kW70PPfaqkhuich9gJcb0OY1n8HDTdgqyUav9Mt6CkG9O5pkeRLiJO1suKq2
SnbYUkvHA7WwIHvW5uNBzTGEN8zN/3cS2D+w2K7u26crVlHhayzu4W1NeYZbMjUbpBRQ/z8jWgid
K3UZe/FSju3hfacY0eg9ve9CVEm5rXXw2uwVkKeUMi3fpvMGFBmsxCsI0ysd5N9jmfU3xgRY5Dci
VAuLUUPr+JiSeK+M/yjz1OhO81wlfnwUVWELVFfuH/GSzauCqMZfF/92izZqJTH/oyihsWvJiWyI
uLodVGkbsx72eiU6WtIGsHi6bgn5NevLIWFX0HpqHJq/398ldhwezfZpy3sJ9eBISBA7SQEdpLgu
meIKe4IrCOVeJ23APDk97JWgj0EEMTiJsNc/7b7VaV4XCF8u+bIwKL1rIU4g8zUsVxBj9CKfDUkq
EicE7+fzgwZt60Vrn1T+klVQUAHD8e8etz3AMsTyLXVrUxymnlC0tlY0r+LrQS/J1mOQU03qsHsN
2cxvVXlN7WmL751SI0s224XUYjxRxKecGMYI6/YMQxWfpXJkyJ5hFmyTzXj/InZrK6WN70cUJ2AN
jwys/0Fq6Pw85V+kaerUaE29MLd7lLgii84cgHNkOI3PR0vESYJEXYonDgKUSVb4VdpOutQy/Ik/
k2SSQb0iInNhilLsPAcH+mUgvFVPnqCDhZMgKwYifd/ey7grWYTSQAhm9qOtnFHjFlKc1LWae8UM
1MNXUms+zfpU8cABJMb/TAmTYy2g9svWnUYV4XA/qLa1U4DQAagyNxuV97P9MCEQZFB7Ur1gmBjf
r+8ouZuHD5lbfQEh/ZXEG0fZSm1pcuhO2mhNE2ZcphQhc3VDbE9yhkXolHp4wl8CjmPdffgUtJ81
kgbPBHDT1fBRPqECcPbn3ipO+UWCq+IzSqYVV9vGyNnb2CI+A9SVo1S3KK4NDUXYSsJ+93z7SL2C
aFrsL2gwMb2VS9q0u1HawaIB3wDGHOv3x2NJx7Gb0f1fV8qI59CC+9lhsVl8OdMC6fN1n82mbJsH
LydYD0Bxf0tVMJmtn3qjXaHZaIiL/VbafgNfQxOY5cvGte3aRgy845+DF/04xtL1oRMQpDKoaufo
AifPlUq4CgmZxbkXUwwwy0OA8brnSpswdZQH0vV2h94NJxNNRD1tco3FCjhGjC55QDWlXsq+zHcT
deW5oTBIUz/njzHrKsfBqoo4H6IVVEfmravU/3o9RUqj1jxftjX8W3mp+Nq3/f619klYk/t4DQiI
l84abuTzTwsWpTr5wU8tCwxjf94vIWAQVWhnpqXJLOzMZAQ+SMPrPWrPJN0Qj9fDVnDGvFkRLNQk
SGieKHTH8KoqoHc3mIgPWJfgnPVtqvtswhYJIYFb0mANpJhhza583HqCa+KBpSS3YY6XVNf3Lqpv
dSx/LvhpDSSeWu8LGHXfJ0aYZYA6B28PCUN3oPfEdTGaYftkREFBcwJUjPquJutx6cz0kRg25YMv
8BPWh5ZceVuGsw0zN3uRnwCksW7ZCSyrafKDQCBNNk4AfCBSwoK/EeipmAR0bylGmYxcdt8eot9d
zmeojaasIwElW9krszoe0k3YROwhf0VIR1StWO7G8hU+uW+DDfIt1zhFOhadOM1wU87CVT3hH7Y6
WwW6aImJMUUGUF2dBFZ1TphkVECFE3rbEI2ILykH2bmGbfHCJCUZUcRKSH3+8TMQ8kAuHURg6gsd
YUFINpqkQ1IaC0jtw8CZd/r3ZFnMQ96Iur7UBoan38NanrmHKHls1Y2yul3ZXfrFHLb+gR2kWOV9
/wAXcCKCEJamVHlQwGNSIDfbO4cAN65nY57E4sVY9q3cAaZxSyh2jMW93hnCJX+H/2y52u27FMll
KiSuv64jsP89bd1RazX6kL9yeJ33SRzqeR1DVxZ+c7oZ7SUswvTpj14YWUKj5xKxS7P4r5EWbgAt
ZP6XsOCYFsCj/J8VbbXwzSj7zCkryCcvjAqGdn8iym4fLpfvkctO+9qZpuLXu1pAR8F58SVwjhAz
1/iqYpgAF0KsLCHtqFsuwGuQPvsTsa5DiOqcb2vCLxQmDQ2ng+2T7Alx+oFQ1LcTh2L4TUKg67fx
bWNnhf6ZKgWn5JDWWEjydWz+nIQC6WvB0qqXwq2ogwnJwrETs0r7NREQaFWot7bcAbr7WfpDmLnc
0QU2vOQBC+hBD/omtzQJl3igvK/poA0lAv8NGkfr6R028zUeIv7WsRoCurlv4mvarXRNq3O+diVV
rIPpCCIIAJDvvJ/bebYNN2eqtQKp+QiN8jjJulSbscKiFP/XHnF+llqj7rFa3HFue1t0kYFO8dd3
YltI6Fh+l8EWSdt1rPJBQZZOpyncqTK22+HpFHzjp1CjAuMDDD28YiCQMskkyTDP1HCF9I7qDZSC
OQZEI3nOY6nDqNdMOb+MCvTS05nA508mis2ie5Hcsj+9K08nzXAX0od2W0B2luDUp4B71pv4QPm5
GEfvvTo6qLFWTLgoyUPH1sD5wHLRuaBXejuN5JTQByqcFKs1pae203Fff4T1g7215ZRKvSxOyVDV
hRtuUqRcPXQA7WOAKk1ZpxTNVBBEwuwaUj3e27t8Mb9csjbD9wgHeh+kYlxVCKbT+Wj4HMp2YR7A
y2QeijZU7E4ISa/ydMEbTCqJZ6x4FwoH5HW3L6b7opIxtXLFmrWytECdm8A8rGGYuA+uX+Jg1nSY
sDYSPxhYCSknbVbnIJVGd3YYA+r+i3VXisRaSxMsEw4ZFB59jCY6d2auJTyyDkj28rwFom0yjUZy
sR5SirAdAOCYWbIntPUVDu6f/KXeSrUUP9qoAJKtMu5H1nq+DsxS7sxY9wGkcK7T2kN8j6ByGscI
0QgzNLOisdcvteQu7tdrJ2kef59RfK7dNQD08p57AVt+Crh5KisHjPAe6msOYKBo8+Nd3smWeoXZ
uixIu6Ky+TST05PK/M8sXmcFVng5PMAUY1sazlCkf15OFTwajqumzcF92WiiQ1m+c0T7bnYzaVq+
AALLBVEXVoxngOPwJlwU7b1PA5/eOSxznSzZOO/asdoXbhf+yNe4Df/feLXMmvsq0tE/a+CuR3FL
A6g7VEHADi/VOaToE0PPkdpLzUlQ89rciJfUiaj6pdj71KOHfsvGjdfE9Pyuvhom5fHR3j4nt4l9
2xUu6PqiyWZaaFpmoYO3C4mCUQJ4O+WcofPO3oBiWwstuO6cNyEPBttjJvS/sysiCv+9fn0eCv0O
meHkpBu8B7EaG3Ul4nujySx5xZ6s0v0a41p1ZiyYZUgXDHQxKSOGs/LngPjOeyCxlYymBWFzEiHb
kz83bNpCOqmUgXrA3ZEmaQGHs6Tp2SxKj9th6N5tNGw9TBjwuq7Rg1oJ72LQHwpq6RrW8kdPKQQy
ylKpWOsS8mzTrwuUT7KtTspVChUrrLR2QW8PFKV2BLqWrT9PAwnh+DxL1ZzOZEW2fxGUhouzUat4
tSNlt5AOHT9k27MD+OKSBKrDNrd5BMCaWX09Wmr+cjNeCoijNZa2ma+iRx9FxHyNzpRDUSTIu/pr
DaTEaYmWp/4BFPqlfp2WR2c8O27kEzD2S0qHfGSz1gU41hflDahbQ9MYVNSdJAiHJB9rCcyXjO8i
GfXGdkYdwbhYujAKM/yx1C3rTtHgs2Vjcjz+5naqqXbL6GKY0mUWa2UMkUqcUyqX6U/Gg3BBBjRn
yjTrlMJMvK04fI56jz04Jxw/NrYtgULR3TNxoI9uZADxxWPLh0JG95rDGesjXEYMHXkn91KEZlr1
S0bpJhVCxCv1TGWDLbO7r/uEU+47ZXDVy7Zv0cxh/h5kypiciGxipsAL5ec6OpqvlexvRgcOADMT
1uPuPQvsEYqjlpDdt8SOOCl3MWGltzx0WpxGvqBSDUA+cxg3bgX6agClhAuFNCBewC3DbPgF2Yuq
4gRLr8/PAva5VEnUs3D3wWXetUJzvDzcf2g7B25kqdrNosyjFh57ni2nLOGeLNDoy5q0H+dJpDro
R85opy0NOHTDi4KbCCKIhmYJGlPojOl8ZEao1QkZeT1JKKh7uQwSMErfnwR+VBezyp0+RnT3Neci
3NVVLnALZJ1e2Z0M2negWVLca001e/EzRfkRxQ89yBpNWJYsLL+Fx0Jtgc1HGA0xHDZCE+ubo6QZ
w02m/1Pq2ysYlg1Dx9U9U/RBe4ZacimKYWAbubd2uv8WVRFOionSpMWL1D7xeUAq3T9CUyiS5W3o
TRwGlN3Zelj0agoPGFACm4yCaBhg1kEKDHgovafI1UnRc6Q23t1Ttgy3y6LrN0vzvH0W0s8LQ8zS
GI8KGlMecG6LR+6qxesry9m/s3lYh3dYr7QgWQqLISkAaGYcbFGiLQXUj9HH3L+rQU1yY+u/qe4k
pVaag0tu8D3/IlFKK+9UybZYx3fLGdXaa4gM2xNpn579fNTSQRoOZQNFHLN5uxXV82ypQEplsiLL
UbON72OQLcng84qfm+KpxgL8es9EdMD/qQz5/TRpqsCWNyL0rvjL4/I1CpMacfMtuSNjwKKCsUPd
w240tC61qDnaP0K+WjbLtGoVbIYupApQvkKO0DM8IUcuSuU0LQjSXwooZehTKL86NPnQQQJBbo+0
Sxkx14K5ysDp9QESgCtN027qyHUIOJrhAhTBFaoo82dya7vxqpRX1rW169cHrbTclqniG5BikAei
y3Xhk208dq9dD2QVwgDZx4ZXY7+cm+m/10WhOsek/d7C9turN70vQMVjGUoAMYV42AUX7ox4HtIR
Jg7sVof8UUkyioHTRFaMaiZZJ+pvqH9M4sV7IfciF5ZJbkLTm1+Ri677NMYxEf2P3+n6tQC5Uqbx
RT1WsL+iX81qNufM06+G2fhuy6DYMb8/ApnYrw0wepNZbHw0XSOfDboey+t/Luee8BFZ5Rr4opas
VHM9MbaDvtwuzQcxC5JWauXLoyT1VlmQ+wGI5Hrs3/k7NAWmudoG1vzPr0kezGh0nniviRqHm1aM
2knVmFwqYScp2KNmSw6o4Xv6Brwa7IQpY69lwm4j1b83h7tqaa8yMZyxQdG+PTEUvFN5y5kXNyNU
pAIEQZ1cDW9WYqStwckW1BgOQASReZykfzdLxqajrTMU28Fusy2FlOLIYeWZaNESOIyPdujfkGAw
nFiSuZqpTQOuNvwM4Wm3yM0DKXoKfQp4GEqzcBvX73Ok0hoi3sIDA2cr0Xf8xSlWwRdNlde1pU9k
QW12X6FVjOS01BDSCV0lFs4WPTbZjbPOuiS0zOip2orhmYwoFsUv+wlpBblKX0O98CvCE+IGhQKs
M2G/Tjx00aKcZujuDySc+sMQEAKodFm9THWh/ZxhPcAkekVSYShcZEQGnVWlETCTP9rzMD1/Iq9G
4AJyNUmlCWADULKaAXThY6Q4nn2zthRlp/IHiFLzfx021s6hMIecuKCTP3eSb2AcnsK8xGJ7g9Xo
okgFW+Q+0lUflTIlZJELYetIHRg/E4Q5N6e69YK7MuKxez7/HAdMiVyRA7f5BltSP3a9jvX8Rg5U
PV/lTwDIL0jepZThXW9vj06jMUTcTyWv9PxbCux4Eu9rWOsav/5uRgOWzQAvFw2I2uVQNlXCWWRC
Gq2/QSwgAyPsDhi5zjUuIcQPyaJGH59qS69o9ThrPrS3uaXhnVD5iHD3MfrTmyPafO6IFUXDSnT/
yfN3O5QTQ9dubtLoPlHN2DU9dykfIqpQylziqTS8G9RcI1btnYtq1GcDJxDdPTWnvPoUg3lfoIhM
RIo9OM/xRLyeEQVdht1a1cXt1204296hGq/kn8X7HHZ6bK4YF54SQD/eyDgPhyfX5uosYR2rYITv
iybTGmDqu4rUrw/1kfD6nnz5QKb99bk880QR/hcZ8eb9XlXP4djz6a/GrZo8IarJ8NaV1FfCri6D
O2tpbc45oRoUNESHYXmJrf8ihKtnzBJ5Hea92Zpozs4423KouiiZ5IgEsKEbmZNHIzdqDoCLu3+l
HIjxmPTd45EDnMorLYskRZFS9fH8W+9C+MVs9kLn2P2ersVu88KBKK+S6pclpZj8QXkvt0N1fXfg
AlGOaOTnrKEcjLBaPG1tbpa8eYgM3bLdfhZvBBScifsCqkddXX5Me71UsPz+FJUertE3wbHVnoob
CpHRL6zFFgrgAa+bInzBJCLwBHDEzzzRiPUveVmPoT0WBKYXOzM8sTsdmoJIaKdJ0HpBQ1gIvcPs
ps4dGPWAYe+Ui99VAe99ngTT5PK0MDMCuZ9p1gAB5H3/z3Rd9KNTdMk0ZUwWYgHek+W3NFFhKYiJ
MmdvMzdNzeJCv0mQ5/Dv9nTZTQ61J7zHMQLlCznD5eL9rr9O+qbYG8moaJ3oetnuBWFta9fJm/Nc
jy9tGhdpHsxIDU0jQk6JeltAqCe7nN2oUSHG77ZQ3dNBFnuS9IwhbV+qDUC5xsn+OzDdQgOuJog9
5tvV7UM0FoCKYfgkq1b28PZBArPD0mzQwNeA6aDnapUgDy0fKNYGQO4chVV7MO+ZELWGcL9Q4qjF
NmOq3qx8WHKDozc4nC9tQsOTQgaHA9cJnxn4keXgbGTV79WLjWnQL8PLqXxzt9KoLipnzxTx6Bgh
MB1Ki9Hn+dkl+GdfwXzSwN3FLtOMQIhKoLlSsIJva/TiK10sRpP5juZ467cNTC781CtNiWzC5u5W
MjhTsuEeKKhLVzrGkGhaEF4u//TASzKOMBmb1vAudEeidh5pSkAbGCp4/8li37wUcTc4PMQb4696
hL5rsYQLHB3XUQa0MrM6FCk1K0vzK+61pVXOEdg0aly8I6n17laNcitEvIzHsPWUHXCBa7Dvs7Ue
NdnekM1xW0Lz29KW/qIctMCo4qYdg/ymbzesXHNnwkx/LEu2NL4965gbB4JHkKONvAwNIql7ubx3
8IUJDPskGd0Vd1x1XFF3Lej+8HB6l0LZ2qmGuS6TxGV/L1LA6ErFJ/b0GWLIu/0+p9+Lngi5cDXj
LVLCD9SvcFrkhvvWE/H1TTL7DfRg6dYIop40GWa8HBNPcnIYE9y/qJULikbNuA3sUCvXX40G77cU
rqACndq/SWndJ1f9FwYWggdb/1mjabGJbempAlAPqdHUOh6cLsxGoUS8Pwgv5BCEI0ICIJjhBAmM
xNmGUoVyA9LXqXaS5/y70+WpjXVy6jO5FyO7EVnWPq0a+sB+d+Du8m73/TogWTtP1GnzVPe3vBAG
4tDd0XVFfA5aJkPWAov7WG8NxnnabfbXA5AQqn5HWEUcEHFCseCxDoqCZH1FiQLxDtpwvSGshEQT
EdMw9+4au95LFOjMZQsI7oE8n+msitiCPkL2I5Sh2lD87bBzMK6dMBBTxK4MoqOMo21m+ngRunwh
X20OdRQjmU3SdScDuHr4xkWk1FKOfW9Q+8c+MIwRRwmHILbGtllKzf8hC6LIgvm5ILkNvJEz2F51
0eKLQCzhZk7/TDnoAFI26etdg+e6DuUbkAzrroiPpn3K7Iry2/5UQfI1RGV0fJiV9AWDDfpXqKpH
T4KozlgthYy7UGJ9xDi+mNM3MBjUtgiphl71+yh5G1C1Whj823Pvawb2wSENLWlDxUTX+oDS/vev
YZTcluVms45dY+TeciPyTh+nJyKVNdO6mWdbOZabR6MehuCZqRlW1tScLWHUeX7SKxZlpIc1dQ/I
fld1zHvnlPFqabAzBRAgWbcueKlk8b3zva1oQnXUyLACpxtw2V+nxN5LWqD8jCFA5hBNFGXrDzyA
vRrQgfr5NLrQbdtlRqRUTyeRJQawxCPmpMp0FIQ4f4UkJ7EC6mjKEF55v+yqCmvNVmUD4K84c8S0
I8eRFQtgfF8K0xxpJzWyJWk3KrZDlgl/a/RSxYv8LBm1u6VWryw9cPK9CHmgmdnKo5WguqFVpNDg
JD5Vy74CRZ6dOuXz8DWiWArVaVEeP9SjoevAmFRfKJ+LsLfSjC0KKoWFgA7Y0eq/5NfiPFtZOHO5
YCCUi4tmrfCC6rpWwCL9T1PSYk0Ho1M27W2AgQu9EDVD/PRFrIUCd9SlsCVr7yteU81rBdwrKpzZ
bX6y5pIdm/j4ydQUotXgeHbRREvRPkHvymUYxdhT3mOtawLN68kuZ/GRJ+DKqsLbs++lWXO7D/Lt
ZgZtZxFBT8ZrkyaR14z+ZC/9cDA8xK1iKldrYCVU79KgAvdLsO39s8IAQN/yuRKEoLIqauJfuaC+
pXNkRhsRLjJVCOF6JWFZwnR4g7TxlPNTKwZ1Xz6OL9YJZidtxMFABtEdrIol2LWcxV/3hAbRnxHe
M6UgNx/OHQBmpvUCofm3e8FvCB0EphUWdEVIm+hsI3e2gXdamK/o/nhplgXI5hxF88gjdx6dGMFg
yaHpy2RbXs70cLw2Q0OeoU2ZzaGB2CKIc0vgSQnlxVf9X+iE3OARu1MeJS1FNkYpsiCtrzLCKc0C
Y0VnI6Tm2QeyBveBTAaxjEfnq8HKBKN0D4m40x/vjktlDrjQpqiXpYww95K/S9o20tlwd54wYIC8
6valzmpJrIJjJpURUxKkVFjRiboUCmix8fJdz7HFBA8ramtgq2a6EqOGdQYTLMqBQd7gKO2gFaGb
4I8jqb5OGmDJ6/nKNZTDgI2uLh5EGzRJ4jjE0FgVc6BZqjfxVxNzLKqmWHsyracR/Zxku8AGyeiV
tD+B3IMgzJYle7fr1dltz4Gk3QgIA/KxfACb7XmyfHYBkhZ4rSFuwkebLn8+ToLT63MWKESGrHQ8
TCA6ZLUE5H3CQXbh48y4WhCNSibmZWKV1RnkaGM8WDfjANKAAtvKTN45GTdBDRDI0WWR76I6HeZ+
U3rhIVxBinHQhHEZA/H4ThNV4m9BXK3VMVcxBEc5vdQMMS68AEKW2DXp1Lzju0iF3jNnFWSLhPKr
m5loOcHD1ae8mXCLHLT+yPvHlS/y7HtLR3wRaKS4jybUhuZ1B34Lktb1Uz1L9xKBEOKG7kDo7i0u
sgBWjVUQIItEDsKIbtCD+kV059zUoORxOKcYuCORie/AvG7Y9UZOAfv6Gq6NM38GXACWDzXONq2P
3UtBHkpDSFZauYoKgxGZ0HTnRKBy4c0LJeVR7z1w6cwZ9CLgGj32oVUc/crhLVhwYbA9lQPk9mgn
9XYUN3DqCCO0CrzhRPpYxXV5RpATrPNzJKispES1ft3FQOjcSSca+FrUPs8rrzSryOQCJT/GkwRH
FViDlALXsxK9B2LN+MVXEQjra6iQUxtd6Y9RE0kqKOew+KpsXc4qbdSCTGcSidvdGpwb8gYRV8Ms
U5BM9R9fwxcC/j1pKK+9euN9QTeBQfR8ZVsQhyjo+Zwars7X4hJPIEfKTP/zvNv5bmQ1Tgw7QmVQ
+rE9AyoZ4C5nXoKSXtcgB837CsFAFUxiKGUAKk5iFEd2D7sQIN9ITOi0UIWw83RVeRXoPyrxMSnd
i8RELHH8VOAHhp4Mr5urR0CtUhXFxg4nF/uDrbJ4S8WxqBZHjE/khPfBB6Zo7srSTOitJbrJgwct
fBucuKjUjjXEx/IF06rNrK+48zbPkd1RZRCFbttiiXalIzga7AaDA8+8V50epkDFuIVU/Gl01COP
W3Le5WD9rYlI2KbDE1Jpf5hqMWzbsYcXNBWL/PA6KDHamoX0UJAcYVbmVSrHfS1Qfi9PPGViOKs7
035tOquKPc/YJ0YaCNyb2T4PgKaY7KJJYn5DKTdtpnJH62zaSJfLUbuJsd1y1owkytt8PPbT6rfj
2Zdwq0nv6qiOrCs2BBqNGCy/9W9paMgi0dIPg68qUGVx5NZ3t4rZoK/3DGxtVv1rmh6LuPiALYX7
lDeX1ewsilHmp4vuS5UR9rFi524ZiuKnk8oRm2vb4GxWylsVAvckH6qwJR2zDD9oTh5nY+q8BAcs
mqBrgitOP/4ezCpElOJKUy9iO3WvG9vpnrywPPDiRJCaF/s6xiSaZv861r65FqxifTocz+IkR3kM
kcc2nfAmsaRGtKh7MXBrpI44mCR7rykFbBEalHkx0xFYiFxoENzbwuI/tCiTdOVzgdF9bIwZvZ1H
q3MoP0kreOR6lvHkZiF1DGxSiQE3Uyl69tnX0+cDzE7BltMHmYYIdOAdVjQZxOq8tmGc3+ktF54+
uZGgkZQOn72uyZzwii0X9cYPB9LE0LNeGOyV15YmA/zKpNi2ZQZm7IQzty1QXnrzofeJw+vtd0uQ
o1CgnUaUy1B4+NqSzxjWNYAw1NSSA+PXij/8vdh/aS7ZJooG1mkstkpT6QDCu4QFWesANhOFWLxO
8jKMkQZwoaR5S8c7M4RoXtQKTyzHRQbN8CNVP4x63J2Gr+8gksE/R7lIPDWAXqq8m+jS3UAbFEUY
yWv0eEo85Fs2OOGdb4YQNbtXL4PTIvSvRBjP3tGKWF/FZUPW9TBQMBflSGZgao8Czxb6CfT1H4lE
tSkx3k/SkdiGMe1LWJiSfGeMAh0f4Fix/B7JAzCws/zhR/iH2lWykXeAHPuKJN5D8zHkGHMj/a2p
wt0Jp8cxU+c4sqJKQg03u7SP+gf2c6owOYlxWr/Lk4wap0d5cDZC/xeXUNwMxjxCgY+l6+7rFTVC
TC6wStwR4NCwBA8QZf2T9Kr7miwzMjAgrXAVFUFobh9uU0OEInkoX8I6KG7kabI/lz9/LJsq0yOF
VS1dwzcCJhMyKNV9mx+nroOaOvZxFei4UN20VXpu+Sg+IM+xfQQiTSJ3PyvAt/ckGs9FQzeaa8uq
70cbd6APRdcnpS8Y1WwuPFPrmfDmt5LwWtcnGoB+FDdNM4T5W7l+ERr69I8DMHMr3oRhJ/TCuN/c
2BQpknN7gJ4bikYrKLo/GpkfqGBSwOr/uPoz5PEFXEDaDMZLhLZcGh8rDaYubnX5OArPUEdpml05
VpEEhSGoWTuFViogldv8MbJ022LkXRiFZeaC5kxM59kCkLBi1PqdBE6aWQgzqBbsyHeiy/SFM1pJ
846A0kCEI7oHbDicMTBVVSOyXV1xheAyfZAlUqdlY+el/GX8Gzrp+V53Qk0b5wlthC0UnUL0ac4Z
shlOxgg+AJi2qRDKZzergWPe94FMIDcnlzHoRKqPoRHApxvk2XMZ9VgIF0X+cLNisqD4AtMUqk7g
3ZxjSfQmbYcs3+PDbQmt2qw5iRXG6i2PVACbJsw/5mnMQXIsI/j5fAUmH1P/MVvTlat89WiTm/DE
twnn87Sa3tLbFcxHTZaI34hldcPfkmpR4jSyrQ0CmCu3zvXpeqwIKO2Okmx/WHa4bUIhu0ZC7B4l
sTkmAH189L0igelK6nyCpXAwQCHpjVvR19XYw5SOObK7H6wiuNZTiTUchGedESJTcGpE7PwN6HOB
+x6IlnKvjhZhBnxHrKExWiIeirVVnbMpjcGZNH8IEI/eACGK+N5R5sgAHxeoPjB3Zmz3+2dy5QVw
xQgcuoN86MekxJ0IABiKaHWVWocZHFcAq5b3QBuW6z69nDkY6FwN9W9kJlUIeTE0463CjHKbyHRs
0vdFkyBsvIllv+X0EnjEy7FTzYkCVydEfBKYoJzjTXIGtSdVQb03Dtw+Cndde25u9YN3k9YgxibQ
pEfKUnx7xvj/CyFzkd7sn+ry4GEmUtwWgGh1ZD7pFpENYEWHZha4vFjbTQkBC8woWr/tIEhznNJE
4xxCR6vWAcx2qz++9CqdA4F9aAo9dU5MLkp64s/jMFYFidnEp5xQAot5GCwlqOyPylLCFLrZCbMM
ly24IFKRdo5G9/09Q9Lt09J+ZAsGesikVGrxwcw7N3MMiBES9Rz/racl4aAPuMPccyV6WPhyod8y
+TxAc5zoYnsOhXEVJm5WBTR2p/B5XEAr/OkewEwwcxoV5UqH96EVVBvQNMxmN4ulYrYjC26x1qms
YiJIuUuKN0vvy0MKd1j/zA1MEobquf2yWAOW+bqs1GAbPcGaP8lLmJcigj7x5PJQWqbdB6reqCR3
57mF6QLyIzZokvCZrcP3YQsGu78dmPlpXiKqvVbNzkcDEgzY8UV++Z+LpurzA6K8M8VC6JCxl+V9
zD/PkMwfBTraSHuRbhtaVjVYVxVAujtFhB4PkP18HQfK0wyNyuhSsYHp9WqcuZ90hpDs2GuivLga
Ryk6p0ePbeC1kU49Wb4HUqVlv9E7pO42WHcETtS9UiQisFgUJBkzaCXUn87hGTM+0XwmKopO8jES
nYjL/OXuBL7T0ei7KnEHBTj7/+l+2lw6klaXXvR09JoXsmxDr4hhVJR0NLgYQ2Q8R4Mi9F3hsOOJ
d7CSLZobHWSVO/AqcsG0hdbju23X3W+DvR6zt/O4xGjyml48/uvWcwesHiDR82IDWbnRaqAglyGV
HkWyDeQmpW9uDPi+I3PSD6AYM0uh0KC5ArvAmn7lkpjssxb0eG2amdHxH48hBSqrK4cQYSGsn8P6
qWuCTNz0D/AcqAFowaQFwcTlwtSMbqMj2pEfb/foKLBzLsWNh8/jAzlK09mvvTKpe73TB7Sw1DOP
HoJwLycBWIKF4GnuOr8rAziuzlalLXVSVD+kgUwuK0EAmUV1Y7BWaDVJdTilkBz0x3X8YzRjJlw8
2zceUmEYgVhNIJdLv224JJPnftPGbgF7kEuG4Y/943BQYvJIhGe4AM/AA4udeEK2ENsFKhWl3CQu
7rmCRlFOjQ/TkD1SAhg07kLN5dwgki9Vqlb80VHp9u1Vb2D0808VG3uxCPZ2KTLacgDGz4YLvLfu
EFzY82FHDr+0Hwv5I2DwUX2YDkUN9zqJ6Wosf79d6Oz6rZj/54G77fl7pHRKbS4tja9EfUnxmojV
LaVYAZH0yRid/5DXysfeYvt46cNBwlO92yIQIMaqbbeAsg1e8wVo8rEXuw4+5Oy7gicqROWGIlZH
iS/+t/JMmYeEvTku+CxfbO6vcAVxpTEV1+nqK+k3tyPrCxwO1HgPfepaObUokv2BJxaZQ5LV++lr
Z5AoJUMKQdowId4tSISeix9x+yussEmFZIc4U6JC0AbcqVwpzr1yUoKXC77lGhPl6sx7tNuyDCRG
lDoms//sFxyywSBUj3qvGyiNjAGg6FgZ/eIZb3NCKy2Z25GNN858rbold7y4ya4Q2gWF2ZpWBl6d
3Afzs0atgmYdAA9i4XTkJZE46mcaB51BVgjFnmnpZILf9iv+6eU/4Cg6vSkJnSi+5wOTTJpK45F9
NP9PBPny1a3ZHU0b+b0Pv48PKTI9zVPvxeQsHAFySkGqnZWLo4z3xn2A0H6C/S4XnCzZMl47ZKfx
Kli1kDowYBB8Gd63JgmU7wkE4IVMkumGZM6bW9XOwFbYiXk0YHvjSktUlGb8i26M0WxjRbSjhZM6
p3Qo0teHYTjR04hSeoa72LnuufdzisuZD7azjEWhmy1nXXch28uUyG6gKdQnxZX6IbgXqNz8/rvY
Qvr6C3kY/9ArfWp4JuMJUllqt3nBUMbMqbi2uBN7nmORL9NvXHtbRftGiXDaAXBmsrsMyC/ZPnV7
mX7hBq2qR4DUc6Jtb8VNmuMGSUIA1ai6wSm7q5FF5QkTZ4/wdzqGf+y1R1LZO0KOpiJJTcct4wWL
v+qRUMp9JpeKC/AKp27ZMtWHP0Xuv8H9Iredg0sN9c78wVo5bW8xEBRMwSLlJR9OwHYd6+6qlA89
z5+bsjwpg+qwHqgM7QBLgFnXLUE45R24KILMxbGq1Ho2F+RzIWNvIH7mTKHrCJvCwr2r+iD7b7IU
5LLdI3Sg1vPDHm/1tCE+hyIIcJoVe8/LfSCjXO+NCxLldYygYzn9E9A9oyWSyoDYbhnfU+HN4zYw
Kzmqagn2s65gm4DDEM8cvryUbNRw5bcy6l47siGVxQgTezsU9MJQ6F+XAbwt+WxzYTodJBc/r+iw
sWtz6nnFICNh1X3LEN6TfL7tlqcBk/GqYUIXGw9FNt/dIpyXGlj+SEgG4BNJHDJsFQlCU8arUST1
Jalz4etOPwRmi4Q7auQW3YvpYPEaMDtYN22Z6nSne833QpEu52VfwTO8qQ/c3+Qcu5SjrWqWaRNy
MeGo64dPkR6r3JkInwqHHbYRnX+f/expdPSbMmX6++SiWXjztgEQlH6mTfRsJsQsjFF7nEBqeD8G
v0ORajrJV2rn05kiBpn2jxQScZkpk9FYp4iQooZYpb/iajT13dFvx3rPLWoB7AiS01ll4E7BM1Dx
aLOAE51tBAsBZA7SVXF+uI4E/bXAuwCbWb5OHmNnuiVq1Dkvdqll8z24mJ+88OmAmkx8hklBanFp
xG3NFlbjrkIZB43KGttsMpUVVk6J1UF6zP/Rve49lfXGaUVKLZGucdPHGSH/WrtYpsMaEsKboMsY
msHkbG4XzBNtyk54cdIbWQSIn32CWFPNU0Vd8URFyC6wR9QH1Y27BfGNlKcbTB34PblU8Yhhy6/0
JA0InUeqRh301G474gjbO4xyAicPKRtaSfgmDuQW9542YOrqlVh0oPIZG7PMIS46+5Y6sTi5HWtt
Y1ZvsxqM9JEd8orgToOtAHtefgFgoKDsKDd+k/HZKBS4zBJwdoO5QoA95OT0FzY1fn7MQ3FSjAix
BlkGVnnVZPSNGX+Fvf95xojYYk+JRWOS83bYsIcfXE6vsSAQetuB7NC7BZVO9SjB+jIOV48i3j3w
tbtny0fUpWwkWvPziyQYCHuG76V8Lh8KpEDcXscmwOr3hyR01L6IBxvSopL4NsUQYdoikOukX3fE
jVRBh4ex+eUmMWsIqzKvgW5x2+UtoL193JCWAr4WAJ4Z9RqzbvPW00zwMn9ev0JJhWkX3FTD3xqq
HxP1oYPtYe/1P+1H+wHdSLfM/97kBPu5WOC4iWMk6CyEnH1bRRI1ZsSCHQ0i5H3fQVnnhwoxo+Yq
yOfcnC5bXaStAyoRc0w0crPxAO0g9gc3ADANXHCOZJ7pLA7xBy1AOmFsMQDDBc1P79xWXcwaWjG5
9wO3S9jozBIUmOC44wLmeB93Gn1HU4jyh2rdBXaNiUKd8j7rSnkvrajPraUBDfQbEvhg4q+iRWjI
PHmue0IQBifgl2uCFx6Z0rTEFQ4r7T3xrPhG98vTSp5tH3EfRxIe70tr8Mp+8Afn0mW3AS+a7Sbb
g0qPZIBtp0vjavVI/TKAq9pAa6AseIzehxRfAtka+EuZ1iL4IAYJy64BHS1sANeQkplN5PKZbKLd
AiIpdEhyk6rnHe3EMSXJRNHFm2gbfJnyXSvEkaTwBv4pWohQNnDmbx9sHWBrWahsayQPcf1RrA3T
6xdfxvvQYBaCjNi34zM6Xvem5uhDDG5omisC3mVWBpfQSD66hhnoA7bKcAWYJxldoTc4cchGP+K5
u5l4uJKUs5M12hj0u6irHKaItnXggCrTnP199f+6dat4ATuVHeL9zhQ+POf+ozZv9e2NUjuTXWqT
LgswRS9sk3y5zPo2gYatBz/dqSkUIgfWLGsr1oezeWTJDkZ5jZyQc3T0aTQl+E34PmgaDvxEPT+q
4PWWpq1YRJfB2fFuGI0q2uzhPdlbaoXNE3zscRVP5BvZd/sAYjBzSmA4FWePgmEc4uXr3h+wRehi
ilQpq+Hp0ZqnfKeWGaMV2M8gHY4Aaankg9+g6cM+hBOdAnXgIq130Uh5VaQpgMfIAQRDDK1f3l5P
QBBuwIksbJGXS5aAlz4VKWH1NbEEDukyLqskk1vMwKYZvnx/iG71hvWOtLoB594fglPNcRFB3XCM
vss2SiC0CEmgn7ftJzedJS4uLyJDeWGQyfVkMcMjEl2h8cY45nXFXovORjZ6o8ZuDwo5LeTx9fss
q14gWQc902lQSI9lDhBvBWiMQVO68a3NSVGeyW4Gzv4teZudWnAnC3xLVEA8w4NwSxV//app4dG2
ZAjH5I8z2BnugUyqKe0smkZ/U8Z6y67EmucLpJhg498sAVZeA4euR9AcTGPsdDoUqA9Yg6R2o6Wz
Li4a9GZt+XPFE97vv5sArNB9T6Hs2puitEVk5zVugg1wdOhWm6tVxGbg9P+HcncMj47elLCH0QO2
KaawSmv9Td5Aj1dY0tiZo03Owxn45bON8n6V61giCSJwN9aeKcse/uVwKgF+ZveYHJXMVStz2TFZ
npOpRsQ4Nxq1ok1DKlT9Y8mmdf6cq0QrJTylR4bY5ktuMRNUyF+LrcldiMwGSkf4kzDz73dd9CNt
57+XAQDH8K0T40UzPrn7zQFlJN6Qh01rBcmyn2ZqD4Va8MWUGsWqAvkrn8WeeQ8ggVwx9aHqV+GN
8lRudsxLUeMpY/iiRU6aLQOvRNahb7nPhnu4++xkiwHxHn1krqX7Duid9HyuPr6Sq3GtZ6/bHWTV
kdqRRS0GyoJWRGcFjcgL46l1mpfJkMs4hMqEzV6ydkUPfzaEfJGuUt66eK6iui5K/O7mxHsWWHxr
Vmb63sgi98uEDdORQrXxXrAe4NQx1MaR1B100pJ6Gv7c7SP/RmRk4FE4ENMxsvK0LfI2GikES2M3
Wj3IEJjcluXZSMM/yhayZxOYZy8OrfaFFh1i7e3kZsdSoy2nbsFiVKnkbqoLn37wTTColHyZRK6c
9PYMX2qq2YBIMYOUhZnzjTpoS+EJ8HBTsmtt3Bqrz7rwMbeHZ0jgFgIQay9g258QZIZaCTUPAej/
zs/JgeEl+tRMj+7xXfJRzcAwCB7ylI/gonPRw9p0oWqqILQUO44J8mGBt7oX677tfUeN8j5IR6gT
LG7U3MOUuNUyKmLVCq4moQClSnBxy6mBUA/jUkfTHPlvnHUQwns/rReXAtQtCYCaNI3tUzcZ9oqU
taSehesGo2zHKjmdxfLbAmh29STWP73hGGIY7+IButrrW4B9v0zh9ZP5jERSddsyPGlPZSknB2Oy
uO8cpXRzzfXt3RK4nH8E1cFbGro4rjODfNjtlszHWkvfiYBuhJUX2tgst+qP576REbfUA2DJZVqk
hB14ZpY05qUsWAG2GjDopS9Nc5YSspDi7RB1aoC90XGNBaPQnfKP489vVbM/in3xFbwp3Ir1Vymq
yS1tADx6QZe2etuuCRLAfXvHWvkdAW8+AbAwaC47XseBCqwzAOdqwf00vnTdBkyCp3fjysUeM1bZ
N+eg/BaHRCmI6LtlshxoHkHflPLTEUk6C8g5yq7xCIp7wS1UEtojaabjaYO5gIxP7nJVcTIV+mTn
KW8YvnKLbmNcJh31vqhV+CCCd9Rtc5OGQHphIgZ0D4nX64f4Eh6CNmovkh6hRj+rx/Zk2pXtxX8I
KpDTCR0UgjWAd+ivNYkA1InQeLRvfboNg4w/Pkit4tjdU3lo5HjxOgDZ+fcmyuW1QFXeowAlqESI
VZ2SOsCI3ynN0ukkl8QxKeTzNTNMJ3QcDS+rDjqseEcRGUiOEkJQhfX9ouLqOmMcEIV6uyg87DnS
+ePRtnDayb7ppeUSwCdp5vaExh3XP+quVuPdYv0M3VyBkBcYV0+M4notzOUwljdg/A1z1/6/9cr/
u5eifAjAO1SV92uHCAcwYZPkZ0+VMkf1wfCwrswkvYCAi8BGtvuOVrt0Y+/bgCHYO2MIkd3/X70Z
RByAb1vLOVCAlPL26RY8Fo7wc7pq2QdtUbMYY1/PjY8VogL4PXBa7+vhTMoFOFyBhAEMpgWKrp7/
GeJs3v6NQ3cSBzogdixxm8G8cYrnDZGN5NyLPRMfbe80JJQ2YBzAFp0VMamETUSZSDF0Jc6QKvRS
dETEPPylrn031trtG1gNwBBHl6TYbkrV14WaciNTibxmUG861jgaksOwV6Gh1bGEIsS7UAN50v8X
3TPbIMxoVwKCTaQWPxJ4QishbEcO8tndKtjnr4CmULi4QwHHRITM12mggvvD2yVtYo8HycTF/r3n
K6Xb4wCNre+at7sF2i8MKz9GRU74Oy8bTDSYqpx+y1bAFNxlBGSTMCIZvvQA9drnl9MSrCOuC7/i
23VaBT6b1n+MESVU9SPRkIzgPuvdMIGcRvao6HxtNYl1S7mDCpNqEViUzo6h0tZYQu1x5l66K5yj
99iDMA7i4ZIhXjGJK4R/n7fQGd12FN04+1Ejp8XWXKCvw0EJN2QzttGx9ajzCzrmNCAPZN8Lo1rr
zE5Fexg5n213jN23HjyOwuYNoGcoOz6Rs61nYi/BRJYRXkGZNksM4r7s6Pfi50DDMFgkitB1bK/n
h4Rjb1pKjLNiP1Yus25KclffzHVXMwLBDVepqAx9w9hiDHpr/p92t+SkO86sC/p4EzjXOaelXzzb
LnNWD1igwI9PXjGARLltOGLcI5I8MmptIxuUdop75YNuNRHq4fStnUnodPpoZOpBfkMnKhLlBNqp
trdga9HqiFoBjcYe3P6KjvT/RWPZs69Ka2g6hJq8eUfMktow8vzKWBjOLpoCIaPO4kukQwtLPYW+
FC//wWp+uAyM2D5o7elAh/NeNnusSIsMpAT7wo6RX3x5MYGwIzUo+yiwP0k+Ts8sIQSO63Do2A8H
6C4jcF4r+05zMvqKABpnnjtEbkByjIrQ/7PhWI5RDTd77TXRzCI1wWfhiY4Q5ev1j+I7uvwu+//S
eD2seRysJKolH71MpTsuSfekaD7mF5AoR9TLl0PA197pacmyYqZ6C7seKZXs+AD5jFwyufGte9ZL
3iAfDv/svRGF2GK+CeKuvCD187FMozpBMDZvBJETVE3yrDv7uDWlyTSWe4ClfPu6H4H0f20S26XO
Ava1KB9CuYmNxDULZ5V5wlwE0aUb/KyPtcCce25iNKbg27wWxXHYgDE2jWVPXmT/Mid6fCTAUB34
wFF/uicGAOjP02mQ1OuEL56mVNk+w3JBWQj6eowi5/1YrwIE/wrflDqxR4vIMAUfDfk4Fadqrn14
8zyb4/PHGBnHOE+ETn4p9t+1/MhtTp4WD7HIsg9EAckJklJT/3/SA2laWSr6k7fsdLE6hbQm8SWe
vr8THjh7PJ1vu9+43/cSU7i5ib0L1ehrKuvnXB0PcXeo/jJ61/xyye1H2EXb9+XyNSOzc/w2e+FW
I9ePjfQu4HFNfGm2VlEf7EGggjuRHcYYm1ieObFqK2q7aQ+QsiQRhaXiZxjxaOtl7u0TAPgFsSqO
MXPbH+aVTqXOlDVJM+n4HJkxqg5kaOWFXY2UenewH70rhMgE9wy8oN/4NrTqnp96dhAQjXfUnV5I
ZazBu//5kS0QPXXoNXPiX1RS9Bkr6nQC3s01wqg1PB43t42lLy8iHElus09UiAQpFsULpx3SSEh3
8wP+WF/eRPp1nchkZNd2OqZPFPWSCM2lp8odCJYEKHhtTfjev65ilHPKfdBgu3+zy1NllWZYcSYo
ri1WITRD3oQiX/fHmdst72hVo32BAido2ECX20Z8BmplHhGEvHCb47yiqmMcwR5tAZrEqQVpLR9Z
CqzcOvYUO0UBxMOzxxd3JfT7WF+d6X9r+OmeSswoB1dliWKnCenaAKR0o8BmQIa6GNIQMO2V3mtV
SsvBwoB3OJ84oPMlrS6fhuY0WibgfAd2GZcsKEVmhpndYbsMgAX5CYx87XOGRQFoaZ56Y9PbmKZ2
WJu5lidNyQgEKJ2jIXEP/hM1SGwXaKfkf7OmI33I3QK3SG49RYSYRYggOKbgtG+wNSmUWF2HeGXh
ZoMICvGs1FMOQEjkfTFYcmcDSmgOJOzzf3Vk1vgSe89WAQnt+didlegZ8O5pz6j2u9zzRzhlcU9l
LdaKkdRg/n0/vln3jJ/CWYhJ2GCwIqJKgVpzxaPMnJUDQjHR89/Zu1sIt11vY5Wtcr+4ljH7H3Xt
3DP2PaXpNLfZuck9rgbFOQ+Kn6dEvt+MaPHNFkNFdQbuiHR4LxCaeKNYDEeDU/0ud6Tue3AiQXSu
9e9XmpEjRcKryQ03o9Zb0wTF6cFRAA03Ixf0WGO7JYmltKk53SQzkcBS0+sye+/tW970i7GPBFXF
SOJYkLsWdGXjwkoH1JT12Lcj7mCHqFoNRkqCwCKvqP7jOVrI3JqSb8mZEJgbAGnKCbkokbLPKgui
lPITFEAG1o6+gdK0Q9r4W2KZRDhfGgGbXIkeveTFgYL9lYUT3gUaTjJYekWdTgbY8nW05EyLM5or
Yr8NSpPQes3ETlV2L8fvsRqlhHtRvljI/Y3tiVv295SMvB0u+YSERbDFSuf5FJHgFcuO+EwoW4lt
7Y5uEeQK8QbEtkFnyNzKXOIMFluZnJEOcjAa+M4VHSc/QFueQH9f58wxiSwXsArdEczWAjSAhcWi
hcSzZLICTxfjWSaW3VMGC++tEtJJ2/+L2XVbJ1JlecktwdlQiWudcEg39cJlIdtANvtqZsbji/bO
8/ulBouNS6P6888fRDPUtgnDyFYXR0GTV9QgqjkltI0D9KG2tCZ0WG8oJHECOAnlPnZKDHjEIO+2
wUcP/UnOtR3OC87NXyA+jJx9GJyaVcnS4dDgIICj+dsOJTlXD8LVqIFx2fLBvUBFBP+pa/jpfXOA
8YnVnPceyiKp+WI0mCyod5spmoqUMnYT67YgWztg7qnP58rcURnKy6f20u6xFabIAHbKXUP9kis1
IiPByAQiYL/9BLn02PDy/aUHybHTFGj13nNLF1RNzawHXO7PoG3HQmI0UQ3YwVbMB49WkLABQMp+
22pNZBgh5fJhii17zx6lo/bGSXXkyW54rR/DoVYlZdjgbgrLfVc0cKn2/1kz6hKcDL7u1iE9qv9f
Go63yX32SdNuSvdPuRdp3FdCibKzFze+Q1fHMroFslZCLYsNb/V3dN6qBa0f4zBnVBWwPrqEhP+S
OZkpU9tuM5b/+alqJy7J80DrRKSBI3t9CX1K2IG3f3IGMiSCUIxvQp/KOLRZ6SGEwVhpgva2Q0QF
1WuIh+PJatMzZeyeHsoRnfMs1jXeEP9eVad6f7RF+FmyE3zXqgDlkHfjmUMUjKw2YurbBSrX8OlD
JSu2MO9r1n0oNC9NoFVPmTtMoFgA0I9K1m9r6pnhuZHamn+AyPJGCirtJWUaWENiskE/PV/HG1ZA
f/ZcOqUFGJnhodK3zyxtOgO3RMrsP2MM3zqOPwHQ+rcQb5gHOI0zuaIamm6rLOYSFI3ySZPvb9NB
9OcM2+D/yu5GXFlTlfA7YiEa65u71EGpfieK5uz0WLqcp4fi5UvF1miuRo3fDhGugTzzKK49WVX2
AYMZVF/6W+Cc5KqjFO8X4l5nV5LQt2kdWBO3y6l/ghQf35XpdKDFCXz/+9E2+SePmgK7x/pgAaWy
ZS/SJGFg1lO+TQWCz+IRdEqtoZ6x8tptV9ZYVrR7VQc3W3DFo+2i/8lBHpCQ/4F1W1Qojbe3ercj
nGeGyqyAfI3SPVkWBSvTHqsaHeYOwswkhc3ehp9ivOkKvrFuEo7B0c1BBhx+jei6G3ImbtwE3jDy
jqjZsuijhjjBq/Op+TmsJC74pdj9FC+XAEkH5aBwZZlMYFZh6T/aaMXi1DYA9t1Hnp269K2nWv+r
PBX6QvviMi9rvMIduFsc7oWr6XJWl3THXPvvfklfWU7RqmB9V7qadmUQ4pzKEoV7jXH5fPNMh5dl
FL9v14IXa4MABhHdDXLyWY6aKuqdz1oVvaV6Vs5LrZFJLtilvB1myJzZtY9pPKgYNL4GTSnfnPR8
87GK5TWecUR7RsUydCUdAhl9IXIadSvS/seHsYJYvP8qN5ypTcGFJnevuAxPllegNU+v1PnCdbKY
XRHStyn5SSY0SYKGioZOGuCbz9w1lHg5ySmP6Q62RFw+ZcscgLbzwtuub+ZNCJY4ecT1HAK6+NSm
l1BcfrDnS2IVQ7cJhByRPq8UMAQQ2E0JsNgvwYj8CpXlM5pYJRcLA0/LYQWjk77zlqc5vn7b9v4u
PZbvO45VeUGnY8Ik9K9DaPw7bvHScqWm6STFErEilWd+L/VM0GENdRbR3YoK2kT4hYNamyZ+ZCFf
azBkTcHw34ZZioNwga4fL0pOlp7mKFzoYcgIa/FCjksK6Ec/PPmU5m+6RvsWaFofkfaKOql864BM
O7GHUMhJ+rmwovxuhZw7L4iUZWE2sZ2F5mPAabxTv4eLDnlvEvUCGAgZF6pKZv3hS6ijmVSclRkf
bRELTnIW5KFeJPjw1+wn/XLxsYPUXCQz6J2MMlUc6n09FGP4w8FShCwk5BrE9iKiLMLmnAJoG0Bz
XeN2mdkzmzIb90RjpG3iQ7TEsSY7Nt6OMG3eTE73G39nyK5/4UUiI0IXRYZ02pCcDFMfgRXJjX3I
vDaPp1l20KjdU4JR+Kf5ccjJDG7GrzfI5pB4EyA1UeMEmIYS0in8joZRZVgUoOrKVvDmVutID19m
3yfDZ8tRzHkCH8DMDCP+uExPvOKQQLUuFuvn63t8wDKgx25PrSZTmFLmUoO9dCqDBh3rtdU8ICpZ
JpgW1K5FzTyCf+uA5PyH0nZQVIBjYvdTVG4sufC8GdEwJmo+raL+3QmGzmUYhuhQbND3VbYiAfaz
871BRR7d3shkplt+r5vZ+Ps4oxw9Q7hDohciGCfboOnQ019ZR1LfhfXLrjjgub0jouW/TCKEzs7F
vd/5LqlTmuaZ5Y2cfNVBECp8F4/yBVigAjgoTMWfdTQQVt/oNkGRv8WZV+onsJ9IStip5s1QmcjK
vjOa9nufODmyLFT/wW2C27QoNqd9czMvIZ3BbEvobYYkAKQhMTeprh23qm6oNAWax9P0Rv1klnxd
rhEbnaGnojbAyH18/RYwZ8NvXEIScBpjtzZ6bYBBa6BTTBo5qeSbamE+SvxGVeXdpmOIqKphDv/L
Gv4mS/YfiwawTHqx7PaZzOtcUjJb3TJisclo70I2FpgpTwD8oAp08DIhyZ1qmyNg+Q9BkhAXFW1G
1J4tasyWDaiuy33JmF4nvVlWZYCmifco6WD3ssfzlw+vbpivlCEoZJOUFC99bJugowmT7v6+Qrn7
VHL9rJoSIZ9v5sSRK+d9JlQlvxVt+g3bb3uWSVnAsTt7Sj6hFlzuBIGwWwOlZ/D6k8JMyHbqesJd
AEf6ztdpzq/wk00pQp/6yIE0U5yKIF/cyfUhwc2FAvtksAPHWWUmNgFn09jm+rW8wW0tkGTfZok3
kv8mKONHE3eCz7RDToGzsAd7E7qRrPylFQ2F3AmEEC7S1Gufz66pfqaJwQy+J8fxYMREMhJjYxBl
qL4VJqur91FAlgGRfuncl4vUPK0jqR9wXL09DVIvvzhhF0any22G4JqPFGEDIckEWhCuOXVdog8M
i1sk/WyNTjsBP55SD47qD33RVhTVb5cTfKEpTvyWuu9SVEm/MEKJdxZOLqipON3qdXKsQvk3XLay
IY2SakSiY0Qt7E9lsqs0Kd9A5z//xjV/2eiq8k73nllll0KlbOxN+dzsrqyXp5ptw811JcjnL30N
jf/rwnCenzZsi83kIYAKYYDU7WDmmeKim1t7A5TPpCBaDvbO5FsP0qFLXwJA/PMTKLFB3GhWmjNa
uGvYZs+uNxBa5SJF7wvvHeIJgaimjr7GV7QjK0JYCyKcfDvLHCO5mp/txA1kv7tLTGK6Nhsys6Qp
kxf7AjuIGzanHcqgkZN6MjX/Aj+PwM6oNhOcQzb5x1Irj1JVkY9zprqxjJRI2QB1uDesF9JN5ycP
/nfV2wGMlB5s0EDJz4k2jPmHcSpHpSrauJPFrEHV26aR+rIDYRU3Ba+fuvbc2RGctCTC39dlETkW
HrwqvvpuQqU3z24v7un8FmWvNyldVIainL3JlScqPn6xKA8Qz84kW2utiHMSC83eb8gCvGHEYQLm
aFdOvvCf51T8WVlI1BANg0PDVdRFHVv0sKg35Bpd1Nrg+uJjpxmDW3zXp47Fauoqnug75UT2HKN5
0hkHLhS/Y0U4MT6gxBG7EAoRYIR7BgIPePfdIWI7j5WNVHTHx7ZMUXlA+D+PY6UGRK4BlYsgNxoZ
Vb8XwDeDlDfzZzD/oilT2NTrdceF2nIcsHkKPXJRxvNft2WVNgzNPLLpbdCMOKi4NQaH5GTFdDT4
1uGSqqKWasEAZhJbpTfxoyTu7vLfDFz/sEQR39WZ1gxUl0d06+OpCAVy84V4DM5HX6k9kxhLCJc4
mDvOC1C340jwMTRVMYtYGSdv2u0GruF2NM31rIm+BMd6ZchI8xD+qIASqutu321FHr28qFtycfy4
m5gRQWD+v4w1n1ONamjedR1Ys8Uz2ubCz7nTKAoiGyRJTmjttYNhAf0eSo4xvSofGVhIZOvyAiWl
oVJSQegM8lPfVOCfXBgDgAo7y7OvtaCIM6y2iEimrv31v3pkDimdUYIl89LDYWKwoCMFXGRzYYoI
DOPN3tUHsexElZCjOi753t+pcF3SNF9F8EMMxHU36xmFY0zC+YiITI5IPHKpeFPMfTUiarShStGx
lAAVyB20ksAlnatroOCnm0KCQ13OkIaVdtc2tPVs2S1GcbFIXHH6IAuCXL0Fn07NHhATN1DPtmJs
z2+QOKznLgyYI0gKZ7hK9+r49V6pdYBSJsbRCPr1ZLe1vhS40YTg7qkwFyvlPOZWoQ8EKiH6+a5S
Xv9ImYaPblGrbNqq1gn5IqRVKEAe0G6rpD1+dxiyO6L+RVEGKj0hMzxxFbxzsmoWOoXlAkAGPWbF
L0qEdeLeUbfAFFrGDUDtImOvUaiIRqRQINkrazZ/7unha2j0nhsYQjLNe7t0hv0i6Bdjm7STuLjz
f0YEz5tMHqO8543WKC25sfhZ6O+eNq74xUApze5+Qsq497ix/FBTcA1Pch9erO8/U2LikKJJEK0O
If9oPQDaOJ3VaG3kIxEZ1jP+UdWhqYFA5wpnK/OYvZanBSQ6mRGYy8hmXkBq2BDbDb31B2s85Qjx
vUazXhIpyzJW6c68npEQ+WjvH+jS42j4JwsZK/yzwljFn5mgcttxmenKvlIYl27MYCEx2wxkXKac
VUNFWOe75YN5PO3Ee8gKiO82Ys20xiJyw/gnLDGWs6MeWaLQ5D/cvj03dRu5bAnlgdM+eG9ZUJrW
WQTVjJDji51k2jNE5DHYzK6BmFAnOTLMZlFbJ9iphWvYePU5hQAabnaDSR1F2INEUJ/itQAcAHJ5
TRx/XT/L1Ow7bD1gxUh3OO9/qx3qxEzCuRQ4TX008vhgAYMzY4jY3tNz06kdhnCWG3clvEZvjj3b
0x8ZAknHCebQsXzn2p3ZZFO+7J0siKhHyB/JyOciss+NVQ+Bobl+LjSiJpGbRKp1NzcHKH8iy7Rv
pzL47JaQJIm2b0YmNzVD58XAW/y+ulQGSrNBwfcT8yFHTeNRoMwpvU8aKjOK/xxXQxZKFIj8Xf9i
CloBD9iD7VxZkd8ctgs0ZZAvPtIPsS4uJJhFx6aydnKOi5x/znyv6UlpoW6W73dTtVrnVfeLd7wL
kHZqsK5WSnz3P+BqNbtG2HYp+QU0OjvOoyTTX3mxybySWWd/rA144IfEDMCF8f3glzhs4epnV+Gu
M2WqspNQxho7zMcVTYKSsrwfbG9Zk7LJ7dUKzz2XknjnMlSb74XwQL+aEX8w+3EInaY/jKS4DWq5
rz4MlaHt/wi7yf4U2ViTzWefIYLq8yJzjbemRAtot4fk4U2OXNRCBsktYFhAPJX8hKGFkfP/U51l
HGG4WpWoLnEEVOS/yQ+Kq/wXppdGBNrFBOMRhMrziVykp7gtrVi+ErGt4YBPfVjARWHMMoUCtNPf
NCmNPHgEX/rv155fxE+bMrTi2Cm4QWBpuYphIRXXkH0fP86LUWl8riKZSQ25ScjgV/xTX1I1Vv9+
3lHjkqblTZMFWHUcOX3mJ4OwLd7CGAQMKIKeRqDycH9GY21DiSSQU0QPb0yh6ryCCkHL692TGFAg
Jsse2KbOYM4IOXZ3QqQfid2qMe4JEsiy5R6m2FGcbFc5hqUghuYF2Md2XTcbX9AGkZy+yQTWmPAN
1WnH4pNN8xpm7ywRaTeDOnF0IPY9VXMQqnotUcn8OL0l7/qDMySNT0vZtjfTl9UuywguDbIIRVTu
0BUF7ya2zt5jr8hh4urvCkFwdeDeQKkfhIB7C+3gVGNjtYlj08KCn2nzbs6ozL9gz4CMjAfPOBXy
vKhu8tjSWTADb/Gv5FdZQq5s4yJqoMRITN+UQzEpf5hZM/QqE/v4vdB0pEBKip3xtFBjsOvdgD37
dAUhuCM512yi+PUY9VGFsJuSBXkjjaoEJy8c9nYMlU+Jrwax0TKdJS9e/ZWtYTZnGKhnpWcEx40p
4zclnzyLVXdU7hwGaweZm6bL540QEopbr+wX4PZf4uPuIsiBKSQvzLJdTg4/9ilxytG5hrSiu0q/
DTXqs5wpSxD69sH1NFjq0u16vHDYOM1VxQ4LtmSKQiFJzjgE4J3Ld5UjRWSZs46PWz1dLyC4o62n
vvtwoHgq44gor5emhfA80JvCuNmF+MuVJCLpIUwC6Q2MHdHjTLHzjNRq3ShynZvujdTi0Ph5eRBR
vqqysGECSjDUku3ZrXZ2x26pkABXsMe8yxgzxmQWdqUkFLwh1D5GMNVsn+i7o681l6qoOwBNiuDB
A1c7MOqhIGzKGQtsGV5/Z5tH+5Pj9JUj6YQxZ3Zbdrh5TxjMB10Z2PkZRLr4LwmDtT18y4nmrzIy
xdIdZGIvsr9UB0gzN//N9aO8zPlanaUxBZuy+Du8pEfV/TiIN6FF6gYo+/tdIJImLEjT/pUjntoV
e/39WeaStfxTUj4FACDZevfPavi7/NM/27e66uSIMNLOIRBAoR07OjOCwHDPy4b1ge/BikNOazJA
4pJSK+ROFQH2Rj5dLyiBIli98gaXR95K9FZ7rd+9H2TKQOthUDSUIZmFIoFrAs2iF+e5o77Szkhh
JsvatcSGUDS4HtCTjFCLy5PJCGra+6MTrenR9nkrdzfAWpSMTBl1DAxYKy3YFnJ/35IcTzDLUwJf
OKodj1fZmZGBYyONAH6dwLCzm+DR7IdT1Nmfx3MMTynY+D5QCJ0Zfw8eI4MuVVO7jEK2jo0MgQtH
+3kgXn/dTLsu+aGNBa3cRJWx4g/gJPwCVi2acrLM7Q+cpAa8JDH/II5MiNJ5u/XiDJOoojSnPqJj
XAT69LDjUgxbXmiFwMJHus1zGvSIcPE3Ix2qyg23Q6qBee52gzFtzA2hGyrtkodkooGEhdEIpCy5
dMnl37S6Vu2eqzC2am7G+OnGpxqXSd+bxPWKiZDzrZUbYHABzaJx5y8ZZkKzjoSXlC/6Ci1cs2I9
m7/OLBFRubJgafty21RNbg75eGfsDpruJGrG1dV+wJvdtIW6YOCwIK2oRjvotZoVWlK1cHVErQXR
8o9N2UHeCSk2mh5qT/8nRKtK7VqETFUNLJ4vgB7JwhHeLJ4ispKLPPGrHqYa3gDOcNVGwEna/Ro9
yU8KJwLQXZCBd0oguYYlN2jWh63Dwxy0cGAgiLnBu3fj4bi6BJzqgs/GEyy1SuzmO6tnzruVu/9n
IGfrnvJVn5ASyXCLOxfKwZszJ/WYxGyPxy3aIjtSOaVdospZ5rsI1xZnoImBYjKLmcIsmqiIej9S
CKDb9w79l4DmYYJ0ifNeU9uTmHoqpb2s+Mn3Bda4qX/Kts0m5DDXgTkLNeadypaCxJc6y4T0Fhoi
2RPSyqOJB3C6uz4VCwQYGY+YfeQ76GGfJeSXH8U2R9yfwF80e5uC0Bw0JPAg1h8b0IJK6gGolc/j
IIPrXXVhGKNyVObn+uf88tg7qtjIoebOE3xdZXZ7ANq0P86ZWY+PvJJlI7nGPRX7A73O8wZ2LcTw
XJTfzoiOYkox4VVZf878fh8/PvpFe/BEqAIZaNiYyWVPVprEVz1R5IpTBBmK6s/YgWE1O7FKTa5P
oCOZP9Q+KEfIXem7ugyyGjuj91QEnxBtaYC85b3Auimddo8lZqNaEJlBmnej90LsiowEV6Mzdn1E
szjzRd2ozCZbsxFAucoVtyZN2qd1aTiSQwRfAN7YRoduaIQCMjmkJvK88ozJSqokl/lUmLkS5ILd
NDuNXP/y3E5DGKEoTOVjHkwSM26Ldf9/SU+Ojsxtzx88EClrrnyY0h3Gmza+dR414ZNBvTiF3o/y
w6C5RvLQMs1NxzwLtfrMq8IESs4+lQ5uyBprZOKbz5AqaPR+D6KyEYwYFhrfQoFFfMZfClkH3ME1
ErJXPqoTrNGesw5NPmk6hMJKWGcb5FLFSBmapL1yrdqXzMzWazWlLrl/dO93XrZArZAazZcjRS55
kMZICAnXDRQYja00XvflQF4GA8Lh654+48OZ4TeusoUV3dIB26IrhlepVyx1LqoUAUrQuLC4Pn5a
Jd1hAU3cwEWJzzOuXVmKzVqXVurOH1lslBQMUD1OBu+pG0Xl3dglEK8rMBSWIhQrGLOztUHBvw9I
Pa275cG4ITsfiNDmCj88QA/9rHfv9cKT0OoiD3UBdRDiWurcyldoxV5he2gZbc9olf9qXdDhV508
fLnsJVXvgURVvRrTof983S2y4cYEEZEhMtmX/CWyFOB8RzmKt0iIQ2fA3Mp+GyscyBAsUjIAGWvt
HQNvKB5cOxwCdvFn5jQxEmo57n+cfnQP7bZIpFTgtMH04XwprVBPzIUnPls7AEjbSD9py8dIdZ+a
M6gNq1T5oJpfteOK7D6tn2n5AVpas+YVOCPfITbXTXpSi+Q3FxLMVgt2BKtRskJa9hJiP98eUBlv
hM/YJ0fCXtFYZTtsB7TMk35JwUiP75Bw2BrJQgSlqboazj2eL/dzmJPUB+oCgiWbOOkZqGjEtXkr
HfDJKhf4XhtzEkRk5b5HPAY7A38BlfvoIc+YKBVyMjsVQNCEHALoJ036o9OH663YuHXMPf99V6HQ
Xl7k5ZbIKGbutnZMqsvyu02JxFY+PN8hcFzxHkUpcDPos5E+N3s51WRrERQNoIXJUpUGOWJ83Ymr
ptRPVQpe1Wp3ItWdOZVDyRK6AeATq0fU4Z5nutA4TIE7uvYPLPvULKlYzagRRrYxbXsx9rmXXc96
7rfgfydgpBVQa2Dxmm5VvzWOaN2KZDvUJZeGNep81ZG+vDji3dRLVlscV044YlGswulPs2v60Sb8
vNDPhRWhjMa2REQL6G7o9JsUc7OeTWh5scDtMkkzKREl+swmFxCuWks5iiLwOtbJuTrSauyIp79d
eZmq+dI9thHTxHJ5u2IkXxdet/TnInwrqj6c4vPtYqt6j9LGORJqsEEHSDAqGhKJpu3FhSu71nsp
MPp/tzWuzvTpTiyXdBC/GPnpkJGU4PsnmclLr6qM8oTvRTX4g9Lp75lLsYCS+hRolDwca2Rn5AIJ
hKyQwaLcBwC11S6l7JS8Uwtm4cGtXbmcsho0oKEwpasHX+tq8q7tVcCZ4K0W91lvQbhIJlv+2WT0
gUG3uE0bGubhWsP5SkKO8s25sGjpzne4AsooeYljwAN7nZ25stVMl4VytqX20JsKvQikhTxAuVKo
0HFCBRj7G/4+Bl5TLlAhjMDo3jkuMvct0cciWflL0SJh0e7H7nA38sRlJyYDoeU4+vSEV1gphx8E
UjOyPiop1yAxfr+LfxEkBTF0Pvz5UDiQg2MWABcWyXIsY1oSmvmTZFIArcm4CKNLCnjDqjjkrBoZ
ExWijAUqkYhXdGheExS/q/lN/8fV+HmeR48xgLzrpxHqTddJhlcrBmDprGaGODJmKso6m1VOfQWQ
oFVa9TZFoEDMhs7XfIA5RgxEqGxpgjGz38VzORtN6njo2rsOYwEdTXXZ80dYBg8+MqE9yGL04iL7
cKlO3F2kldc3hundy0r2z47Tp3NBs6blHGdrVam1JX99KCG+hFbsewSA78HHVKKdFi6Bw7/WBYBa
FUgrO/SCnYWUX2IgBj3NmTEIp+snTDH1e80GUOfzeJc9OtvFwNyWqxtNBuC8SoxIQ/Uen1MNcte3
6D+zqPaToMuVrlAMVZCx9Mj500Mw/XehQE+cMmq/GVOeSx+BYPExoaN4v/pg9SjbUc8ahUvr2x7t
emuS1FQp1j6MLF21V47+qaysFYGB5He240+YqtGcx0ncpdVfTT1l7W4ACul0qhfu9qmdAqpzlAxe
KPZ1pi2v1ZrRCxe722sbb4iwrZ/Vz9cRLctAC7ny5wWjWP6fp1ig+GOeMFFCeUqGt/TgMqktNXsc
ZIBP8KLJVdKUD8v2uTcq2szOh/Ylaky3dQAUOskBbD/VeRM4FeBEtUCOn1V4gLCSjxTYJfSXihxi
e9I+XaEY7nSJCO2h33zM3rX0uOFSdAOd4U0VDJ82qaTPcnL4hSkaj9z/Ph2guDUe/yQh7dAFBjo+
e6L3UG4G1UYYB9BDH4uBrIC128HiWxR95IEtU+gKiBvVOoOOyVLtN47Le4dJTaxIvJE9sRo+SPHt
PCVr4mSJYHOIAuNl/KBqPX7ynNEUVknPbblIqj9T9nKizjXQd1CihG9kzB94CxCMC0FvZaB8qAdV
/5gUCHpJK8f1MwQpK8NBlGxnhC57dQW+bdxhaoUJdWqAT0mBomCGzZPDAs4hP5xssj1KeTM9GwhM
l3HVf9e82j4JoqQYBh6MYutk1/vF4FaI6tuYM3GA6GRFnsNIAc05tw0wRxMYai2hasHEnCnif3nQ
pbwdsNkxr3vCkDBWfFD6QV+5lb6ru0ky1VdBLphPjeFcld5J59pqHRuB/vIh+PiVp4J5axhGPtgy
k2hsZUkGvNIrmhmFa/CIQgZgGQEFolOdLRIdY1BMUAo2aNO0OBrlVKK0Gkuq2qoAMXovmQ9uuZN3
RoSAmRR95mKf7NI3sbdDFTx8VcMGCIKazsjVbdlJbbOyPBVHtbd2Kjo4FeBtloqnxjrZ8U05MMHv
udkILFUe5Nu9xZat9xpjy/FoFBNipBa60KAhGia+YhLq7lbbYQPmaUXL0VbaPTsVzjiUGeM9C4f4
JPANKKkB/kdt7dfJSpjkxYjqDTWi91gG+L570Is2pFy3+ZNjFqN//aBL8Ult3dtOQ3jHli6PqslP
wsafCtmZocDwpfqhkSPA7/XJABc3HaKHsRyiTePyWmMa4RMdupcnEUf0aP6brew+JcRDjMqlilZb
fd15vwcnCbofD/SyS2AYoYJzXRvrjCiqTwCXfrG1jwuBMxDXFO/gDbvdHNwZEDRCJ2932jparwh8
/gjlF5H2LwHrk8SPmn+nmRYKDjUvauyJGONTTcf5iZOZqamOOvv/rNMTQnVeU8HxH6vElO6u6hHG
bSuuuasUzCeFjIhpnRMqXdFM06Z03h4yqe6XwO32QD9WZLV4xzolKLbD1JyiISZ+eXeC18keXJPQ
1APMv7WxZwVlX9luv7KeXns1+jGwgiKAjGa3TzJD0sFwmy61y/eE0fsluhVmQzzTmaVoOWPy2i8B
loUiJzy1hw8sGMBS4O01X4bB+SWW4SbyI7C64RmbwvmTlp9oyYzaHD+a2I0lKZZn3Jq07Qa758Qn
FdjgEHTCn+MMnommgt5dwumjCRgk/wWbcXV/zIjgmrYKiQ+UU+aCxeUudAPE+ko01/eNuTIfVRUL
K/1g0EvocAPWGsQ73svYXX+vFLddq9wYGpyf/IOhKz9N5v3Dds5APYIDLpma/+pIJmcyqW2f8BpQ
QbyIWlPR2Kq1Uoak8rPsMDGhHi9dsK71jKTAPw2SGYlbxwYoYeIU+ZbMiEDGA4PLpaoKm0IZyRxB
PAAFjpucuQ5FRgmFsvGeiQ4Jm0IzSzZVtr5i7kqKR6EtQPCmSqpxG5LHMMLWYcAuhFvN4BXsVJVc
q3Y54MkCSLJQv1DHdXkVBkxOPlrUmHjblmiaTSCnFPfY2GJ06ynf2C97c5ft+cx0+2IvR/TSnLwn
00bBPwjSxd9TSQ5bU15Yc127Tpt8EuH3I+prigt9rXU5M55E5NzWvlTiYWmSkSv8GeR6ns5YR4b1
Ciegehu6s7GovNgLQnAD+fpOrPYemruAQGFmGbmy5yqDEy8ae+mcfC9eQV6+Hi6XDuDFfVJC08vu
egFa2dVJPMTs9IoYVK8hvR1CrrK2v8t+qJiqh+QhIgU1kG8TC5NT0I61JALTQwTIsEDWjtSSKL5m
X3kDE51runPhlsBjaFQyGuhFV62SUXowmaH3e0VfKmUpQrf2GgJuyxoB4LL7BjCo+znMcnmZduXh
m/FqxjEHuWJK/f2tG7PCyWZi4gy2DtuIN9N3gSXKlbljQecassc6L+gxnWlm7UBeOQXuJ2eeaBxe
GiNTaxNJd4qBM6cqKxzUfoscsS2h3cv1iMDxoVbLr++MJLM7XDKpwVl/i7wrSvvzUA/nuxnvhh1E
bKYE+9AhPh+qU+H0ITNV9ECkO1mvwNsPHuj2ajuUfTvdnGWwHxsVc+/5xV60825145T/VVQC+Nxm
/wVIxN3ZFNuFOAr4DysozAjIbEeT7l6QmUNn5AqMfkzC2ZCWzi5duAOoWfd0ENyRiJ7vcg8z1iYp
seBfEEvpdc4fCbaPvI1tNN1GRgFldzHIA+ONqDX87zsqHhfFobz3dxvGlzHPf91bBx9K1/6RUIKB
MBETpI3pe7+79JpuuMc6Xb8z6YIryOHllZMjiw9E8CayIGKW9EN3GiDHKYa7cvFBusaABbwhFZiL
xsBpcvUnRhK9RR+IB6CDO/c+CTRPaSjYS3nDffhrf34zr51dWP4T1piQzm4AT551bbjaypVNL71a
0MHgbpuWTw2jZ3qzpBat8dyy1mKJHVBz7KakaomBJC1FfdRflUnYlSs4xnd3Qm7Ci1sUYbjNveu4
GqKkKKGnvnSQCEFdaNw4gDo9/ow8E5UcT0tDcpzlCyKKno8PX+0B+tVA9npPCgzb/USHp6GAeeeD
FXpvBT06WVMGd16I06+P4yQ+/szJRil7Ae6FF3+zaVXXn5aNz95AusVgb3FCWTGyn/kVf4Tn6M86
1C3umU4P6oKwvulq1lvl7aPZRRbSA51NzkxRsD1MqTnmdW5g7BKS34KHOkI5Ju+TvXFw1AwlUIf6
FVsm6K1+J7PAOxDPgzhVeuHUQ0oLlh/1zD/tHQQy0guOJ1CwzoE2Rj66gOTdcT46uKUAIQutEO+a
3suvhfbq43CgS8AsT6RWg06pR+fZ8gneCJcSV2nQafIbC6Ii3deMN18LGVAVKvX6OKoIvYsBcMqF
yv0/cE8zSmwiZEA15UXjIII1Bw5puOdLJCex9xNFGAD7UtcfepyBF+vIZRsWGykmOq1c1IMPC0t0
1rn4qcVQddrTXQQeobro1RsgZkvFK9a1nXV64JJCRSdWQK2+En3lmMzjU1lg/GlQpUqp8eEue627
54YvudliWJpaLKCkD9AeZRgL0Vt3aSyRLNFMcU3sAiWeBBZL9MFZScZy0RemYNrnRgnwFX7vskrF
xZA34ZfEy0l8OoMLhMpzEF9Oxrvg6+db64FFd8q9poUNjmkaJZ1FIYt65VKC1amyI82FbD0YjMt3
PnPH1KsjJkNpwMIiJce7CzIVmodsTyWIEsHnKnqiwISDNU+t9W6ipSirhdxikWSnPisUpFS3lgB5
qHNGT0HmsbDPvWV632HVUWr/KeplrqV/T1B4ca8fH8g2OL/QvTjk/SMIEpydKapfCo4Lgc9sLuPy
ItLxQrZ59iLljtSAMT7oeg5ja+pVd6N9I1TUdD28RReVj5gH8JnqAdm0pwo2sM7nUysn9jg1LBg1
s8lWJ+6ToKNT5RvPe9eUl/45N+8bvuDbWMkTlESctVSOSJA+7aMtBY8I0RZHqo1f1TzXT15CsEZY
mqI8dUzQ3osjinhYFepjLwhMmhv3HkRLfRljjoXwwHuVMp9jlQzyVBgBCmhpLDCbM/Bby3pE6Feb
ZOfUuJAnYUHye69XITZNzzLMMpTSUZMZ3buTqcolIcWk6UpRemwHywfH252TVI/DrXN31J5HXCpP
cTm4odwjXRjqXETj+maIfv2bzT0QM4hKrnoDRasgyDcCtpTbzFgNOEolJikuEWNFFMrUGsImxX7G
3e+PiepRHvLPWsjGDkqvx15lbiih4r/FnTEzA9NDeLsIT+Xgt9T5XSnzLyaUOChNN4dYYTGhXfD8
9+8Hou8EL2nY+davGZ4Sx3cpatWp+r5p4TQHhX3KdXB4XNbBKbuYFmmiaJqhwJpUMw9fbgHtXDtP
lEy2hMfWN6GXKVUAv4UbSxtcQSb3mIjudRSZCnTwYT0UkgheDyTmyi2eyifhInHEgUnalIoi2myE
2Dr8X6XDqbgJyj9BYri1fEl7CmBVVYpCvgj+7mtHCgcsUdf224FxzOoUarOP5+/qsrsw/aiBMC4q
Re14Q1Nst2InN+U+c38Cnmc259EnFJP3Lf8mD6sVqvD27M71rbf/jQns2x2EWpvt+fYd1r6dRlGn
XzxtOCaZESl0MBLftlZj1zVaT9uLZJyDAh8ZWTHo0UoDXlc4rcl4is3JGwKGeNLFBz1vl/n5QVsN
Lx9if+5nMq8N1r8zo03e8VyZPnfgPZ0eKf2d+xf0R2MezvkAKp2H962c7F/S1qACxsyaT/IW+3Rw
AdqZU2wLXayypZGk4jW36pmGlySLhBWPiTyPLuGJU58RuTubiyMe0/ArxTm9XCti9xBDu/USSzXI
/FB+eB+1FXIAqdaW6egO914obqLAwpjlAJOUuY3/8Rm3gEMsFxGCRwRUQHGi/7R68CLzEHqfweZ9
Y18JCtdAcZoWxCAm5yA7EghidANGq27zCygM+GAOPPV22BOrWS0CdyQb0ObQhCxUIqXUA9GqzlM8
xRrLBujs80kl2WES/11ck95zlfcC7WM56yvv4Vf3sls60sBscSstI3dpUhane36u/6Z4Hh/40Qft
TaFupphFyGMO8c2VIN55MCmfiJT5dyqJtG+oW/AKbTFpVH9lCgI0wbiG3VgFvtupibeCxxvpoplk
mi58MESAcAqk/B+PR3tMqgE8QRf9xKjLqsqVu8cUwOLP/gBgunPvFwIg3BNEZ1q7dp8cNvCsHvsM
DFSGrb5dfNS+QLLcvO5l69gkqNKGwckCZm4DQp4hKawPo3nxtOYaKBEiI/IJ+pWpQjcSkQ3sA4te
4S+F7eIIOX6uiT7b0Pa2aMeAptXEQKL2qeBmrZYRmm3y8EGfhM8ZghAtphWU4CjQpUmSK8jt9jYh
QP7bvOGOkeQUHda+/JdX1zuKiB9O4Lfa3WchKjGg1gJzmZFVJ1BFxZe0LfNw5nKtwZT1xUT3mHKa
FVIy1bHC8HI0ia60OYyJzzQf6+JZ1d18r1yBWsdyfkyU3kMY7kTvREbpbDDze2zyLq0a6VfnD+JG
gyfwPoKCQdkOyvlyYZUhGUULo3XOlLWyFC6FJOYlrxNBvFrhd8wEC99+Wj7oPchkkO20jLhAAImc
l9grO4aAbrgW/PA1IEpncs3UyvXtDsGw31e/roc2aqF+gV28rr9Lv2Q/JezDGQJE8KsW3LFhSBBD
uJm6ta4PKzrbe8NBjtppuAGO1mbQWIXnxoWd6b8gEYukjOIV6gATIpDKpwdHppJNXrBwIAmwGOw/
debAHtnlzbcxxBryNOJoF0JrOopDozN4J+ScVZp9OKvnKGxzKqKVB9wVIYBZ8RoXvJunlxymv5b1
401h2xSRTISOlfAUi6af6efsBtqgP0kjx8I7aQJSrrerfR54ayQro8RVmjwbdfdTOhfGKKzBZT4d
M3P7uBsn7ZvrpllyhimWciaaywBAXRMf/Qn/jkD9YxKWOlJgRhlmlwT5Rxu+zCLHQyTDkgyKi2qn
knxKL39E2+D5OcubS457ZMXONlwIJTquBYwie52HV0d4zdpTppQhLnSUewYSazR/0cnpgfULDapR
BSAN/KgSov0RPZqS8LkoMZlzqEgGAZ3hHCtUmvzZ2RitLQzRhWVIQ1YNhjjAunDqmUKSaIncIuwb
PVnluVroNw1hQfiNhQphgCBQpS4f+JlOYUwttlo1iQ4orMkSCna6ae6YU3oWWb9FJm/SR6Kk3vA4
1mafxaq8qOKKcMUZR5PkNH1wlQnbp5xhj7jJLnVGuhYhgt8ROH5f5wUUt+IpfMGs6xBiTEWDJtob
4Lcy5FKh+le2Z6pK5Kybg9BFrWthhjn4S1BAJIKmnIbNFiWoc6KYljHJaxcmZv+1CvLZFyKIYFHZ
HgUvfHQDZTudOacfVLZr1/FhKLE+t/Z4Y13f0Yv/iKlHOfWx9vL/S4BL+iQbOasRRiF48jo863+x
ccYboV6QUyeR71H0jGUI/CN4/u+2Y8K7G+Ov8r2f+sMebNX78b6Vqgk4IhG12uNFTmNLUPILmptF
hdJ31KRnICdjuDHR487pIfI5GRqyXa0vPosJQ3oAScQhPOlROELMrBUro87LwZPKtfnZ5RXadBr3
vbP+nQfCaCP53iGJvifdO6pAzNbm64v1egmqo1wqcAdK3AludS0QPSOmQfxXvy1C9uBoiDv/nxUc
l2QYOAOWzh9g3MaO17Y89T0bA6NqoRvnrEKFckdnBffrknNgiGKTy/3ORMVzwFaFZtEO71wU2/b7
kA8jZmDnG6Os5IAlXMeqqXOy619ewi6wQmvzd88xSRfG4+YropodQMi+01CaVnZCbcYmWjbDQhwF
9DAWKKfqdU5/Gt9iSbV5DDJl+hZS/QNXE0PxWfMuFSR8C2QrGh/cTGhVNnDTaLiGGNwEmDtTKSKT
FQ+dES+uBZWaohfiF4qBbZOEqsNMjcYDJjz0/P9z8pQG3rMhD/bImnibmsooLsC2vXKZNx5s5pOy
8jv/hKHAz6QTOkFbSsnxZ8GIdw9vhPMxwbBf1pzjS64gt04XuH3FUB+/lOepE8KcbAAY65nrMHfK
jbGUE/ov0zJ65PnRjTQgtyJM14ESORcIGJfmBKsX2inSHePndHlIZQP1SNtZdB6yBhNvEuGUqUGm
+5QR3E/Ha25zlWNNwnqjIXEgLv+OUXZsY/bYYWINa3J1YBqDt0MgTpHCFGd1C3Z6DxiNTBnZyjAI
KTjbzhVWYWI+hLsq2AfzQHhL9xjozpDLKVjwssRuVieBqQxuKZLi6MnwnQFwHtO7wbuOJOaYHl9v
hxhL+eW1BjF6Mo7mrtAIJSEHE1I6H5dg/Rm6XMdaQG0x8ZDJgjpzpW0ItLcdMki+1eXjOgJ7VYzh
Z5+Oaco+rm1qYu58KprHXc/98OZsUiIM1Qpn7Nt55Grzv8CaVuSzA0qswh/jnsdVPBJsO0zu/kms
vjnXysxPDwkimRVv1N5R+sMtQ+AOX1BJtbhMtFtZYHr29IaZu6NY6FUaZ9QNJZmIeu3pnQVJQXfi
sKdwBig2D7E583PLcAOS5WBkajbwgl3k7kbWINPHXO6bXtywVV0ii/U4IyPOBYF/+xQUKYktFwkM
FyqDftAzMCMR7MRkgZgLbk4HFgk2CYScyp8u2PRMVystplwvKCaZZ8SpEEhxPBp32ow8wF2gyolq
FRbJK9Ohs0aublCMpaTVOUj1lDN7xjdBJoqKyO8K/pY2qKzWiiuu6Jmo0GjIzPzaHKsG1xiL13DP
2i+FGS0H9Mh/mpMBh7JQCADtL9ER5mT3YtHc6L+sJSSmdMyRl5/WG8bnTzUhuiFXW7qvbhRFCn1Y
teEF2F5a7dMcTorwF4QUtMJXFK8dga95oCf1mCd0I2UD1ZxZdKUEI76SAMHcIEP5lK45mD8p2sjp
zUCdAysPdv16zi4xA9edk10YqJOwcB9hXN4PU9fRjLSF3q7DshmO+ysJ17+iPm+zWnfRbaKU7eC9
7nqlDQ/o4L21I3yMjA4iQpTeqAIOdYBDk87FCDdfRXS6PqyzwZiwTKFOY1aYfdgBEWqaEb62St+n
E3fswBU0DSz9GKyEbfiNHXqfFA/85lyB8sG4NljbZhXUxHQEhatgUeHs7NV/fBzcR0sxCyw4CoeW
6N2snUOJl1hAaCm5IMFrGZWE1gRS4iys9uvLQbPGBU6UReFsD5tgFebUq6+3lk7D/4C24xzDiM+M
y3aQ2EQ4xz+l27LxVWkDMkzKoocqOjVp6Ui2B9xY3EEoGfXJH/n+NL7BaY/ph+4OcKX8WiSB8Kj7
AixiieleAJdTm6eechSfx5OhuV0e6yDpjYAscpfgLiURq2j/FtgdDqjD4hpN2N9Pt+9cQf5gl5jk
G8GZWS3d8kefe9Bo5b03zik8DLiFn4bAY/rIKMrD/27YoZoN1DUsSil83guriz4o9d/cLcnbGYLa
QKVla6m0nO2QkgkOHcXkabTx1HnMTknltFoiLAnWB0vLPQdVj+xncsQ63zZxrpwNNIiSvyiPCkZP
sg+ssKWQEVqyEG0N2RHuumBMGS9wANBva8QFQBtRoxuzwxGg3Y+2Ogr3stIebyOMh1qj3xyRk2bj
7PHkfyoNYtzzaKGL8GbD/WeYGwD3JhXfpSVh7UVIwHVTX6AGY3+B8OyAm16cB295PYGPiLFgztwm
u+ra8Uqey/k97FEuiXw9of0WQSUwnePpiMJbFcPFkyZxal+yvIJMVumbFGHJ4Icjc1VnSGyQR0MN
O/fbpslOeObCNqFVzWwQllxh/pAaHT8wlku38RCbcwd/DPIIxPzCxV8aDQ8IKtZ9vUx+wfoNtWJt
/1R5zvTO5p3FkgvtpNcwyyoR8+ZQRqwCiWM8esdC/RfgYhnaGrnojS3Avu9kCqtZcxtYsZi5t6JC
dxoZzYWsvYLGzi+lHYtJpyL0KnVM15O0PggCsMOZUMEP71oarZgsiuCK7qTRj9zj1Sgkph/RCeyk
3E6TI2h+fOKrUrIamhzxvl7fRduYty2QSFAEPgUDLbgFOEARIl2Z232bErsMpOpsn8K0924bJcKv
+M3NkNFlzzCmk5ow7RFSViZwpAaInDZ92rlY3RCcbjMoWr7lQ52gm2VrQfZmU3JtRGmlDn06uaFe
Nf/jdvav2Ua9EVDHEcOtEiBKxnH9jmGTeszXrp9LZ5FOfri04FDLdOEAMq2kFqtNXgTZGYy+0Ue1
fWeWESFrJbki5U9wkDaDe+QXygeo9b5OC56A4tU9FQT6EQJPXkWOX7jkyx7Rd08Zpz7qLcdVsVOM
foFLOxECJ1zdsA+EBTzdkmW1PDhaVWOWkfSQw4XsHCPDg4435wnmFIfW9bh3pbDugbVzPwwMYwKP
zq3OXmdErtkyOXSw81srNy3D7H6YMt+NOQbM7FdeNS1P6Ph660IuuGw0hbzTgxkaC+OYIB8vQ7AC
Es7mo4Ur0kT5IJpIOqYszr45HpoYRCuQhcaNvmhlPxY2ygMZZgRvtTT7l/LUtJ+KwM3L2VTPbh64
mo/Zc9EXSp2vb02iFyT5qKZWtEyUOVLMtYQKlJTzunH1vmU/lqYdiddIGonItbaDkbkM3GJAIBpC
PEyUoNWIqPZ2Que1WgL6G3xuCNYLjHqZmtTIgNze92V3nygtAfnxcgcBuN5/+HCzxkSyJTFg7Ytz
TBNwc8LwKlA9SfaHrefSOA2/WCLx3eexnl+htbs64b2VbjNA5JOh2xqpQb+HoXizXPT+FXS8Z2V+
v8veB6+is8ZEXRkq6tTEt+AS/7VRq0lV9aZjPoHLsLYkeJ2AXIbHJgSnnbheE+7SKgue7RYEMPQo
IBU2vSZuZrNLVEaGDaE3MKBAq9bZwTuwuFpJ6obdqcw12Khnz9l1tWiEoKDdNv+p/UV2N7z2Iqr8
d89P55QeeHv2w80eyiOdyiY20A1k7iEoPoGCXbbX+vZa57SgeBZMJHx2aVvvPzMg65N1uG60OxqQ
eUml+ZO1m3AnGDOTAYYr9hvykfME00UaiUWotaxuJUJpAV0LLOv6gdwCHO61uNyLJCT4lNVwZL9i
kHeuJMwi92H0scIHeTjSWpKI0B5UsTktb0SUJTcXlAx33wN69KQj1Yx/G6cQ48Q2kPjQp5iXGoaZ
NmBn1FPysM1u2vGcj+r6q+EVfCboKq9ZvkoHxRqeCemxA3lP6QSgODf2ogYLcpA7tqirjI2Qhw8D
sFFv4aVjTl+cWQ2f/7jJYV6RCqEPi5/PdVyBFfkqWtcrgf1cKBRiCRXEk28uPFLz0G0UJoCFReh2
Z7qzhSrBXqiclNNQSCUX2qwSxxIg8iUCznUJPa+R+BWVmnUiYf+17Lw0hujmZdeWHkSkRdY5VYeN
e5ctLF8GTEKbKBSvJxkkczAAK49q0o4Gl7aFosGgt5X9gxq3to66BOw8JsIGMBtaUX+kGA0ryl3g
jDj3k2AaWA90eD+ehGbvgQWHcchQ8YTGSxtNJZOPJ5z8fvUyAYzFSHSBvUIi2pFuBqed2skoluYB
fq3HWS3a5l/HppT4UiXXgSU4HutrqYoFDdU3dRZg2T45BRi5Q5xtLpkhfYPuu+9XiyXlXIQx7HMb
l11Opt4CaNcIwr5SeAxfd5iGtI4s4d03pG85GyZmTaelkNEOZGwQSE5ehMlO+vqixYNsvcO0Meg1
fjpdnUTwFK4+gWMuCx4m7imNFbs+UF23E2Zi/7Y8AOIefThCmrW3w+HY4JaeSbdOOg9KT3J0FANN
7enz2DGvW/ILt3s2uBWalapEqb5VghdPhDFuViZI/pN3vK1REyprOtA34STlOQgCSNMxAGvj18WO
NczBJ6c/4td14BCiwyjLZDLCvQ1ZiCXlRZZBUNM7udeDCaklxqaQTnDy0BEAMLkEoPs+DCEAET7E
Cy6VowBa/Eu1H/4dlvYGnQ7vo0UDoMPhNrKG+lAdSbbYMR/eWSOJpfnllNFRi/2V24AvDsfhvIbt
QDTYAUS3ciqCuq3V57+AEmrCua7IqZ+mcyCiD40TDZkwTScgsYlFN8Go3JbIQDLwCHNrFFl9JzkD
qgL1Rj1r+eU/qxVnLTqXo+FsEw0NThQyxq+ZBeEpvK86eFHGUb752DqM4zuu6d5mAL9tmisC30h5
yaZuybCkXbC39GmASFMLOVzYiKkGus7vMRrh21pkhd6m9Pbfosjh/4VvEY+8B59TyOY45Q+lItdy
OPkjCK7S5Zg7tEDj04j4Xk9bCHRU3OOqF0oPxu/W31qlcR5DqEXYP91Ic3XBOE70H9hUNd9ZVUXE
9NxiYqe1PCD3ywAZqiUWbP/CiNALl1Z4NR+/neaDepaJEtddg8dzNnpEhBgiruNDU0AAnqbsEBkp
tnMCcK5H6FqyzVdF/Kt1lMLhBwK0yJQF+ycWr5z5tifzkS0t8DjV7tuUpk/GNLg8f0m6YnTNP9Ak
tgE/sdglpmr5fdYWAEnmAmGS1YqikRAbQ4wIvjfyUJM1UrtO6MzF7Dgbet2uHYSPtysm3EbM971O
cQ8VARIvJo9NOL6WudjbplUswdhhywZmEY9DQijH/yBfAzrx/pWtbnC6fCggvrxviCiKNqUdP6m1
jcDuIwOjSq3UTm/3Fgadz+Nv9MZjwg5EtMiX9nSFtxYpzw6Sgg5BzzVegwWgV30sktg6xttzflpw
pmfJL/Geg79KBbbx1wEmpe9/ajuFkr27XOt5f7HTO4IY5/NqLk66kVmYM8bMCNfTOsY5cXa5OTWJ
eCCBu+SAnU5Ys2ABJ+dnSFhFx6xJ1LmB/urkG6brLl5kWEUezJf+DKKPPfq3BJtrUIxMLnvjriQ+
/vdYo+2ilXFlQXoqd/0YJXwEBR1NGbSc6urOByWF8N1IpOcXityAJZBwKjG8x8nlD7YI2yn6lb9l
AtmWoN1XzMtOMaEIhHGRehBFUrDNysNk45I8tUXdfKUpv0/0KL+SnF5Th6GGCDRS1Ygk/uww0sRb
BOhblpcT6p/8v8kvUQ3t+cd2zX44x3K+DcNoizFxp924hdQo91sqBaG4/De5ZyV1Sr1YcVXUnAqv
lR1dBR8isxgyTCJAbHgAOMkUTlwZdiCVi8ZhbVQ2lmqAYLsjBf4aRTI6p/+YS8dI8Cn1nL/vDpAm
5iw08kmNnUkIGuXb773enkYVPT0q2402cBaiOo+8TeE1Un+UDfFE5QNRFExzxT0NApCu8Je8OO8X
dbEN1nFq0CfFnL6W9jOOY6gz2342dSHndaSS52kRb6msDUXQGRHXEthiqwNHdnlezV4CqT5oVJKO
JAD19tiiaclSLSNOxEKlnTQt09GZc+Fctg+wT6c9JjjdFtHiMgwPyNI2MWLi93sQIdoCheoJuqKA
vN+bcsIiHtDpujddSH5ajA53RMwJY/5s/V8EgGXpI9mIulCw415zTAl0uQIDIAodvmxm9MpwytDZ
W8YrVTy2d+VHPqHVjhQW8VoZ3S4HMi253Md9l3lXtalcNlPKwhlnLTA2BfwPCx1GJbWP12WShisz
I1Gm+GJs2xo7O33vsdl4UdehuhusFJx/B9wJ9BUM03Lb301ICXYD0cEgf6vsumCn6xQF9K82t92E
X1RiumHel+3TtMzLR7mTOx8c8v1k7FxlLTJBMIpP/wSS5kmBPJdI993xjbtuj37OtuISZPmfYnhG
B6XrUp6fYLL/uWr7e2PIeL86oVOi364e7/SIkkNMS6F1WlNNBwZ6mkRjX7EuSHyNPAIhmWlyLJHG
9XRVrPD4c5huMOeyBevoOH7G5pSdi6N4Ion6rdBnRUQI+vrqFyGEuYvN6qP9mWh9xlAE4Yil9PQs
g5gECZlvVwuB48whYBSNp2OBKeiWvTtsat6DRZ656DCsCpagCXJ1XdYaJEWKi6b0PgeHPZcXBwXV
BmtleK4UkLP1NPAgVco47jbNUedt8rxpvbyCGCUtRniKg34TDs7Tab+DCYA6vEXbRoh2A4QbLFJ5
bUn1fjRkaU8j/AuMiS6475ktdJf9/GlsO8p8H/CK7Cmw7YS312gzLk+t46E+6fOb4hecoGcb/YrQ
0Zm7wRsBBeJZzhKtzPqr6yvfqTVIPRYlHCIcILgsae71BFXvhA8cNGvzFV1yzZVT48uEp3cEwrTK
oM6ImS3Q7GQrMkvseaCqQX86JA72o0Qu46rA55/qbkfOTbiNZhSGoPSa1DwSYI0HZxb/4rti2Aup
r8wVhcgdPlkV7fNwzb/mJh81IG2CoU7WZ9ccfKruzH6GippjhNRjm84RUelvtqIENPX5YHtmlA0r
LriYRz/KwjTzNv3VEgoDR9O0cLdkBlADJKw8WVo8MD+yrirvQfRigI7kGZftcyXGYV7PG/F7YGIp
arYZPyWvNQTv2ZkBT7jj8N5SihZ8k0w4ITW3mf0q6FZXdY9GizcM7bqBsTNtpvBnZXVeOBSLUjKe
8Y/8DarJTPEk0Jw2eFXhGVk4x7dBYhQNDCkEwVp1T0k8ebQsTX6Aa17woW5Vy0N76+aPhpGZp5ZS
3hwsoMZP3srWQd62SGbj/kQH4LicQWURjLTjmVoYEVZIOmzXm+s2+PvUir1UjzFtx47dWyKoiMF5
6pO+dkXzxGdlA5aaJhWNhFNHy7XNrZLiHiBAwrUatRXG4jrOgeW6GqazDRaM6fWXXG6Ehp7kRgP8
/V40wJyxA6g9ZUjsea7wpMglOI6RHzzVsyQEldGZN71yllSLaAzezfDLYZGMmei+jkLpYq0dOZF3
JXxAQ/C+/iuCoW/2Ax2H+N4CtMzzBx0gRdCZv9BtfIanS6HRzCvMpnFVqFIf1DTYCvuBM7n0w8CD
XQXUwe/xNopftLnM/wznhyETHPhP3Chcp77y1NpuQMFtANlRBe+RYwsS++9Aq4jw47GehhHshq82
CRChbBtBkli4OiV1tOMumX0X3jAOetWnZVKVi+RWyWmQhPVzcKh9ErD0QU6tGoA62NLYbyoy+coD
tvxwEc3JtByPFSsn/iXa4KvXvEDfS9XaoD+qMsl3sivx3hwVC9a0lTZPTMOJC82Ot/0HvwY7Go8k
zYD+EjXPn8gl2qjjFbz7/XjVRR+O11IO7wcxvb7c+HCNXOCpFjxp/rbwsHlm0SO5BX/+Qykf1PQs
4wUIYEPfkxwY85lDAsO7hAUOtIV0J8ygaSSVpqH+q0EsN/2F9OkY4tZlvkWuzAkq+UEkiTLjS2hz
kSXnBLz5PO1UnHHOlpV9uprG13LyED3Bq/Egiw74RBrscW5lt2T0Q44GSltdfzl9WPtMhwQcc8Qb
26uOA84W8pC/P/vcIABEpkAlW3UGc0keMKW+Hq+CrUvnFtJSdyp5YQZBCrtSjwsRiF6qDn8pQwYF
0h1eck6JTpCzTn8pFGZhATdt/KurJKVSXjFMcIt9uCspu1FFpEMfxqij5JDLvLx0VMbCWsAnthqT
3M8TMBcWjjSRuFyuaqwmZpe3jAj1/i7Zieuy4Hm1AAfjGO/uu54puH94EZDW5OozyawEIEP8F5x4
7bJrWXmSXzDygdAjYTBi0yYc0s5t6itzOTEZrZ9FHZe0EgMboRTHMelEn7fMAIJRPQ7wIlbcosMV
CEOAngTo4GSxmXUCpbbm4ob6biw6KlIQiH688selEJ3p2qTVQ/buaZYPL89IVhgp69TSd7KxDPRF
V8CGWcLSsyBl+9D+wWCLorNkNhQVP7linGLX/+aKCWyVumZrUdM3Va18SiPgW1Apswl9fBaLlRBb
TIdEhkt2b+GVmP+BQjKqHvMV/ThozZ0zWJn1X0JauJtrs9KaBb+rzY0lAWITlRwD4ay20KqyrdSE
ub0MdfBfElWVDOk0S3frCJboBeGWm/JLhq8BqsNawYy4A/tDIRvo39lXJEFf83P0qd4oVRB4//Ag
K/S9f9c8UoY4Lykq+rbFNKPnTJWp+tYbnfnpPZlwa98gSIJwzemjDbqiVgoGpZ+gVsRlYdxDPmiW
AFBOKz7xy0LwPUTy1mtYj2EeBRUvEcDNt3UWo45ZAODFVEeTBFeUXsI1v2EyJHWpVZVg2xMFgGSh
k8Q/Ts4YCfP4oLNs9HbLLnwDt1DbPr/tIgBX8LBtFQbgmYUe6jdsXQgJ7ShdMnlvvUFCiv7BYxDt
bCVI9xPSee6CVg2GwNMWAk/8xIPL9Ipkjccdt5e3Y+pRJv/ez5SsJZnD+f+b/4hA6kLV3sTci5Lf
ebr3rGk3KNpgGjSiEAo0GSFAl1cWWYhGedvmE+oU/wWxa1VdulGcSt2hVsRkv1yOPiYorzb3KS8T
zLrhBmEh7sQuIhs3eSbxC7ewz7QsBZRCqge/CqpkBGTc+saa6iGfdN0kfLeNnR52s0573EPpmEdS
DJVegXCADi/HjMVACm2gXqOqpOOff9SX/VxbRdx2Ak5Tm9849GBcsojC5mwFHNB2fzu/tGl5VwxK
bIYaeMFCIfUcQs8vnPk1lqnQaZvCnGxSRbrHop6GACLGDhi6FzkyDJ+0JBSEmLU5K7mh2Q0b1JyG
ehbiLgVVuW2vYZzxdRk5wzF0U90ID3Uymd3VOqbv9c96whgObw528zuQSB//ONqJw9ZbhutZ6sVG
vE1uqEICir3zG68To6xxXE2BLpmJSqG74QTbpK8eYhod/8XZlC4AJZnKR2usYtaDrvH8FwYrxlZj
+ZApulqvr6IMJAoEGiPUaHhlWE/tWX1v/didVkQvtdbL3k7bhnOMC8vMl2mLqGMxDxBuO+VJkIt6
YADkx0LkghyTmlViJLwLEYFYpyXq+5VTHK8rU1Uu6h5ce11Cf0kup5pELUqWQRnQKgeLC+XmR+oI
YTBUTDLxOZFlADoSnamiZD0PhTOsyRi4yPBnYQoud1y4QDqcy4WPd31QXbxc9e08RWTyhrp3vwAq
fIGZAwJjMQmHRodPeTcLZhHOjZTy9o9ern8N+W2KyjCcRTGkEEn//xdb73zIvgNnNr898HyFV/Xx
T69YnZnsbmLfmIUNiBx4nkmLsjbMxJLbgnzellr+PK/GBajbXZTn+by82Q8RM/Qor80ZyoLywR4x
waozpwtFlRd6rjQBw2QHO74iB9QvJDx7PIsHpdN1WCiC1jsQ9RNP4MfjbNLmwSFAKgn4FU6F548H
Eo5nnV25X1r2vIw1OnzNRhndlbYThUwTLl6Ak0eEpZ614JEJVRiOpyJ/ARnmUoCYytDDpJ7H9kMs
E2Q2zOH8Tg9FaT0Cm/tGi8p72NI7WXv6y+SZWmZ7Ue/aPH3N+BmXv6dvPGAwG7jrYXKc/rr1zaVe
cJg0xVljD6nsae3Bvp2HfpM4lCS5zIe5iOh+UkbkaZF6v37HMt6giui7V4pt5QFhIr83k2aq2lV2
+PNkI2m74SxJf73Jb4xwnzKLe79emutaEm9wDnB/qS4AQYETBeD3P+YQtNIHB0oWGyA7ZFWZjD/X
n/qjNQ48AfqUdJOCM1Hnog5TZD3BrqVaAftXEqQpxKa210D8y4Q3MwC9U5xz30JcpCbJLXIistD1
yDR1HKTwHapTKdTCHEdkFhaIrFbv24rZx/+Wbsmf1YZRDvzR4PGSjyWRn7trZ6uOeugc4Nu6DQS+
PTduNoAArx6vBVvsISfnx+aHZmby1O1qnChRgpm+KT12NY+HVZ/l5/f1RhZIzWy15zeMeM0tCjwr
HNgdSXn9rABlPsNZcEO1VjNzz1Ev1UGK88BBd/SdIfOWIWr/m1BxmRnI/vNG5odS6T7zLtzITLBB
lULg0AH/LvvLnj3IpSE127A6LduPNVqI2/Phwtz3A9VHbQmbrVG9iC+Ekb9gq+eAraUC+yfitRpy
c+gJYU7FY4kyeYSqa5UaSPvZpcnAk4xhQBfPgGmz/LFg+fmy+GctLPZ/mqUYUdFwhWBWv0MJMWuz
OIRHpsFkfDNBNHRdNduepxTP0AZw8FZpqwYz3JBw/lsIMWwzzHB+NGah5yDyg1SHJw24QlroNHxt
gwiXrwMl+uBnvXbL4ovtXjSWFVLWonEZJ1bxdAb5x66enjAqYFmRgDO/gB8a0s2sm1XnoLutZOy1
ktRzP64jFIQ7Eg8FzlzuQt8FvDPUIiWhntA4HfdMmOoUmALaiZiJlOA2kkFvvtWshhmUXQso+Lbz
HNuFrgaEbZHBGSM6PNIDJzjVg0WpFiLZqRZDgBGsTtE2MazbsXDxu0L9VX/DLN9oUGKtpwVB8bR0
At4ugoTynq6Y213qkJBgFGVc2/nhk9G8HBzuVLbk/QpgqepC4rOR6GOIErAiMPlKuqoX1inuI7bp
sdZS0vF3Ox+c75e5icgmEeyAN7gjYUe3VbWUvVIfdq+Se2UiWRf31MDHeBjSkVKHo8VBYcpHv9uw
tdjA3b9r/4JZVw2foUfajw02xlQQHLSUio5L8qquwv4OjnC22+uaGUtlNLdEY3I8Cy9DZ9xrWp8W
ffLhk/S/cqGN87LpUjs/sHZvkvU/9kozmCQ46d6FsMYTiFJkeilr3LWG3dmc7ifv2AGnAGIoJQtu
GWh8rE8bXnn+7Avh5FYuMHWC+yGzaBcKNyrvf7EZlVPaRXK0QYpbSD1iUpWzCtmUDeCeNgDc42z3
5LqBqWvdl/mNtBbanu2/2PLi44WcAzKq5Y0E8WfWtfZyW7piv+7GXBeA4tQRkOQiYfafLhFsr2tt
8tp7+P81okeNjEAM4wh9ehjHYsvOWz0X/+Wr+rDYTiEzI+Oujb6H4mz7EOH6if8m4v4uX4w2ZhKO
hdMzrGalaeVP9NNE1hxegmuh8cnPvMDn4P7izfhBYbhMIB0ioPkV/rscJl/J60xp9nSGDD14s5NI
u9fO9qu2whN0zEkvjwsaS3y3NRvsJ0ixpGlplTO3h0evhfXpeZPq2zPHmBBNGDUGDa6LlxmSqANg
0068AF1IxtMGeGUZHdBHunM6qIPekorwWO3b/xSBb95oWU4SZmSrDiY6DIHyd7axk5NSCq+Pp7OR
KJiu6c1sqiGFu3bY76VvfWCk8ecj8+oV0GrcBgdZ2zk6e3NlKCIe6iY9yJEnPWDBaYkiJciCQ3bh
itgpfXVviaZ/WOk1nJGA7FznVrLnrlifPu12pkgw1r1hqhnu6WQrgPWpgKg3U3DX3GEUPxg1oPd1
MCOxR9fUOTpWjD8T5ApfCKUsT81GOguGHdkofHK6RwbLuVtREm7mD+6K8V9W59fkU0x9jsV9KlRT
Zf6DUtCyZqnSjTpiB1SgtVnm2NZfCq4Rsag7a52akxQoyGgROzl55OAEi7dX7k6jNeVwI+a5sx7a
YRrffaFZOQEdr3U7CAOyQz+N5ElZtvVZ9pKsnsiRpHlQSfjKHsGHwg9k+ynkf6GlexO9jSSID+4P
+M9XEBleiTu2TGgCaauSZ8iNakHGGB/sv13+btUUy+DOjrSZvYgOPxZmgdhpbKUXOfcXeF6VqO+T
2o6cBDCSnXkCADpVoDeNJovIqmuLPJpmzFIwmwFhtbFyMiLDLl55nQuBF997YfAI5vMmVPYoY9QS
LB1lXzR2cFil2b1m/5mDaJbbZ9UQVHeKx46YuCTjiwrEnENpKHi66kuQUqQcXBIudIRt3mOfWx/L
B70R2zUH5H3tErG3etVKm3c3aUn+KqCZFt3qJzC7Us2aybiwvciY/lCahOgf2SrLH7flRpJkEijh
TbM31cwjNkZlMhqCktN3bVAquUAdJz1b/zu55xsYJ/qITbnxMBOHLyi4mulSxGzn7is1C8E2RyBx
yvQP+qv6ioVuQcOqEvbNGpYADQZ3RN6inwnj1y8/JJMa+ltpUA7sxwap+AhPW2HZDw5QekdWKA2R
35mbacZIfWQR/v+KpZ9s33aPuZQV7CfYBL02CxLfOaF+c69HcesiJTtcHX5bdxmKNxhuO5cuF6Ie
x0yxlngGemJSy4HyYbchFkNGFCwzlfTNjxFe+TlNh2seIlJw5wFlN9998pMhs+wfIGO8uPJIkJt4
icUrPcC+Jr2z9ukQi4fXs9sbQov8l/DUoOglhfKSjVr7exrLhIqHG+faHt9RAEqCVe9c+u4wOdR3
OfRapEekAGvs3iZ3qjUqNiSAqk7ZSNIHhMRHYdoTabHUZ82mRS9SEK6YnEsiB0WRy+mvzWwyQKj+
leMGlv0yF8wKls4tFEk466WjeCwz9sVgiGjYsWFA38/KxKo8r75xlf5LkH15vypCKoPex87OCcIN
Q75/LZ4En0u1heseRwT/zwq8yD3XxK30dPPkIe3/3dyRtKgYkdBtLgG1gHxoHzPYBScp549m3uCW
5gkhtVMDHuyBEOvgUP1aPeR30K+F/o7seIAOB0qebv/17ndkTSOqZD0irbxb43KsecGjr3a3vAr6
0Px+8kcvTybER5fYmtFFwoY7G5x1QTHMMb8FNDj2fLkj/xwZqqifH22zvgxmSUai9yWbx74RSbrI
B3jy15c2Ab8Tb2mLttDIlH7NqquBMHtDo5a7SnIYeYYREVExlS+JMCCcixowI/hIUVUrhzykYJq0
dWiQSM0zFZk/PhxsHLrTx+XdFm6YiwRv6EBvMz2r0CgV2rg5zs9K9OKpfdkeUUaFXFki16igLFOT
TgcUPNHKm1cPN81EzSrOD19MzzqsGMeaws8nz9PnLxVXuv1+xrP1INK2Vq1USLNOSQfbtTf0TYFl
lhQaBJhQADb97xozuc2H1j1iMWcTl4jhDIohT08bBm82ZeGBc+M0GCqMkOzjmVl2KGuTxgSu8KGv
UE1fCISCSVCP5zHD8LMumGjILEED9eI7dpgh+l5c6mflgMFUqgJLBJP0AZULBsISTSrIJz9rGTlh
MeDYE4t743i1b/ll6C8yxSSYL8tJfZWnnr6yggqSAOIjfjLGO89ZDvwEXk/GI+fZdG0hf1kqEjb4
WzHLLtsBwS9sW7apW5V7FhTwms5FarlvLfgLIPlCAfVu/RU8pXC0fRqUOTj3aA45bNjFYCkAU/lK
p9s+p7k1Rz3NYk4/sKc+qrY8DI4gQfVSV67pyGES8UvFD+eMpM6EiJsJKRKMCfayt4b9lT/3+kcG
1dPeaG/3SLEC+rxm+XFTAeLANwMu770G3HObG0hpCg08IhCNJ8/jm0yHTvyQeGxNlgAe0xDYTr2K
6UVM/Ad5tIt7K/0yi87tTLv1Id/F9ogM8+rGWEyoWEs170gIgfI40uiZHlin7/fSQbYZP4YjWaUy
YUH3FW+sZQg/oi2Y08BB5avDBSUFm/pZEN3lKaYb07DShs8pl0CIfezY6RiF3J9vT8BCHUyYb0m3
aB3dLGJW8sDqd6GffVNd2Fo3n4U+ux1BW22oDLkoWstvwR/M00HLrkzErUgCZqSsftJnJk4ve/MJ
pTU8XPbQYf4U2qbtqwutf41HH8mZF4b2KfeaxMNhEklWadJXEFbghPur3MOxIedE4n2ys4W9CUpt
fikPbdiWgqhRS0GDQUd3WAhRGuVb+UNfh8Hk1+ytHS5V8AxcFzCnIRYg2/YvZDz2tSFPEXW/9WuQ
/iYFnw5cp0XAFASU5pVD0u/QOpgmdBIgPrcBXDVjt0RkLyEfV5RaBqUGPGblZkjZjpZHHdOuVK9i
QM+MdmgKXY2UBEn3xzcWw+biFAj36UnV6SDj6vb/NGcCfQtlI//VWYCawYa8ffjT/pt/hJZprKYD
PvOiD69JkD6U7jvjr+/qWsBg1XhIquraFns0g9Yj3WtvOy0Car9DOs/hT9y7oIflhMZF6+Bcr+ZB
fitkQ8ssQ2ogPWCrlNvhcavTMhH6cVtidB33KkUSUnVj4GpEaGLhYxi4uuREFQ2mxdOaCzU8onTW
E//is7w6DOMRYoJfNxVbqBkoIEHD6ET5WLlQeRakhlk0t6+woKj2SWQvsaXORi6oKaCk+o79h764
4EpiotYYHaUkq08lLAI0m4BBpxOMNQHyCEHCaZq6I+yWsX0EMXiogc/nt5RN34VobhV1gWXENaOX
+7usGsPKTatsT9eCWqLHIdBilCtO4z4ZqpvvvsnGei99nRXgM6F3RNTM/IAztD/vnIGkk7OHKl/g
DEwNCZG6p65MAk+ykRVrWuX7bxdExVs/iFdCw1IS+7gWEc4GSAefVAX9rOnwoQdTZ41bXTKlLGg9
0Sudz5NH6+sQh3N0S1KLqwuOY6e2VuDrrw8vUrhqrMG62WXEXR+27lFeHlMPWjqC0qEOr4IjkVfC
QoMxe92lXfCrKmVbhfE4XVVNtjDmHgFe4miboalchWuyt2FIiWYCzh13rXN9OmQhUGoPCs9Ij+1H
cl3CPoPrcB6aKMflQyM3axbQxz1c5vVeLhDqxVsvM94ekAR7tvJUwF3SQIPp+aGLsfGZSksMRuQy
REe2aX5FeDd61qwulLpVQmvS9NkfGcJhFPk/IYnn37b5KxHdPy8OWrGxHcGgcxBVrjvnGky8eWVK
KudkAMTDmeD2IDucJoeMfy9iCJZczehGYyMGHH1N3yAT7I6wqSQNAqtUNDAhBAu/H8witZGZhtyi
u63K72CzlnKpWKgrOA4a1oJ8eYkOGa344oeMKnog86l+RmBIulR0zegIaiFBRTu12BcPj4MIbXKr
cRCpAJECwy1UaI9sW8zArJTyL4aNVxwb7EpxGYFM7EmccOr2DwWgXhFPF92X+tind2mQcWGsWQQi
PXT43fqmZ8JFUnlNvu5wrPXCCHrjgnPL+tPpotPViqlwHDMFpAQq/1KRu/EmMsURC7bpwmv4Ljmi
8OYuG1PYvRY4fMouBLacXaK4xfNDBIfFPjDIX5JJ8njvv1aZ0QnQo6SzFIhoDX59NbajHU0TY1iz
O53y0Dxrk7VSwhmHROALGOGM3dcWjQnUYmzZqhnUgbXX7bHeRZTNgEOzcktAEh3sFceINOvObfwS
qSSJUKiP2Kzx/oZnuNegV28tnWxyIVBNgEpApDZsMB2Khi7Xzha/RNvG1CLDfb2RH4olNUWdUjjK
3wBSZkKQCnNyDpnMwzWC4PlV36GUfyKgWw1+kWM0WUw5vFRzjLUCBE5ZsbrhY/9jeL+TOtWXsRs9
GPfxUhzFv1tjg1q2vRxL961A2xcy5pNmUXby8JyzxPhJBHVvCBg4iehs4XzbbdLKXfr5sP4wH+3T
wIJfnjh/kJnoP2pD0Kjnq7Umd5x/aQT1Y4jy3eOiG61CoKG01y+iLndKV4knVCypKPvxnxSRlUZq
MeF1cLK6vvMuuA+fs2F8Gn8WfGXPQnNr6Pfbx7sdLENcCRTL9kQs/0KF1AIxIsLvy42R9iiFcTsp
4nNl+7osVc0t/kBiM2JGR1/BbCkpbWTb5eE7xrTQWTuB+jL9SW6X0HIdjPk3Sq9n2GaBc+99xB6L
UdreosHs/U0o7+DjeSo4iZC+gQZAY8lJwH1/DpAKcYEwMdA/37GeXtXLphIsj39arRKsl2fMhxzs
94amJzSHoeH2szmZVH6k1YUKXwMZcX34RzoDcGSVPrsSP0htknC9Roz9CO05Lyf9q+GXkEWhAtWO
XKlIvVF765l/CVzfS5HxmlhN7o09Z86zmB5kPuk74sSbMnyyyB6BsbHjKp1N7NUoY/qplDW5QSci
8k4ZHtielmVRRJQoJS3rbGlZeG5qdaanLq+/F22qznTJUJP42d+hVwBeuLJJRflHu4nWBwdy34mP
lsRuwpalj6bIRYQCfdx98sAZjl5XB68i26Ne2uwZnhjY0t8Ixb9zEnnX9G+EfpwFlZXDfkiTvn1t
TqUQPpeENqH+8+X+ZeBFmMYxBJEklvSteYq32InXr7JpETo9tCbiaeok9gJ164eigDY51pcN193D
l85b39dJFBWcq12cNwkksfdYxHU7arXLpsQYhH4JN1pLNTrjrRg/UzkffREKpaysHbrFuZdbV5tG
BwEQN/jksvGlIQdEqHHssj2Tal6UMajbwz+yfHvzy4Y1Dkysn35LJeWAkOqlQMabTt9jjXN8xuQW
I+LDLRaJO3K0cVaJpoOyHOPwki0bKbjTYtqUJhOygJ6T5+XOoo7EiqisTR/Q++rsBOiVNiLmeyG5
ZQDFgPB5WJAgQ2IR0ltGhNmhAlNsyBydPyk7uz+DWHc0UVNmBm4ELgm18T+0II2vj6jdN7BUsVj9
Jrb81YjaNlXMasoqiXtHWelAo5SXC05Rhy1eHI4efoMdk/A0VMvyTEv4Q3tigUf38bL3cOpps7Q4
YkufQcO01l6lJclM//ZqBlJHpOhigP2r5BOIqrttzn+/nCATcVdLiUzy+Aa11XXaEpDmAU3YXTH6
lU18cnm3imwT2/732nI6AajOhIEDR1x6cDAbKFUfgJvajDX/c4V7lNHRfjaWAFHHPKpr4AEkhT/6
aPErb3cvWzI00ZpVmuxaNChwMDXrOwDCWPMrrT7w8juRE6r8RYSm0NlwpwcFKUfWGBIqaXsUGRSu
p0asaYqH1wyDN5BzuAVCgrig+8RLx4BIlC6CpXtw3vClorucCItTYp1HJLH1ybgMdGFfHC8oE5O9
PyQOMUtH1DzQ6IX75STMrccUg985iqXR+Of3LswahAED6Szv0OTsTlIuSgeb0UQ1iYwN45NLlgUY
uXB72zbI0CwHN1iQ5rJ8aLFgdW2P3jZgGDXwJQ3YPo2+dCxScqe8oERcUh8HVqNMbqLANQl/GnC0
nVvViuqPzvF8VyRscCPtOJ+dhlVp79yHjRuQNO/5W/sTHV48AMODpUInVCnFhEmR66gWhrtPAbyf
Nil+bgjgGVN1fTp4IJPB0dwjy5JDCHkx3dO6boAYXk+huZbzvvFaB3AvGbGv5Cknc/mefkJxOuMc
h6eeZRG6KinLxlSl9libK194C5J8TgTynD1EfY5g4AMcJgOrqPCJvwxaAKa0+5uDdxz31+fx6/Le
9400OcqbmUNPxnWx9LQC7ls+/na9TJFlt2cR6r5qRslm9CUkZEKKlhvrfxazeYxH+K4I/Kkri1vA
h6QWdBQ/vR6pfO7P9KfXEfwVA6ZF/Q8hr1ksnIzloO4LFRWkBi586JCo23R/1C46jNynT/r7mlNL
x4v8tpgUu4NjdwAYdwMBDrnCx3AVZJMw3j+dpxhTnFYXEAtBJH38a8X0FEAIQIaQQOXQvW/ad/eH
zb4VBXwdoaVL8y+5+PdTjVRt1108BpNbgkd5Kv2wzqv50P59mYJTAfVuaAXZNZ4X8yU7cWUBpXb+
zY8N7pdt1FpGoWWSwOg2XgcLxKbkxKOKgXzZTf8sgauwWGK/PFhAmkHLyyi/Cd8mRZlY4oodV1Vm
a0mlK3DEP+OiZozs2woNY1yu/9TGWp19iqqUGwv9wZ5kEoo8zDkUa+M7a54zJLkEQAXnoUfI/xzY
X5/ePeoOqShIpfRaTVubrtiSJcghxs5P+u8k9DklZr9+uYHunyG81lTYaM4WF9BXwbzEPpJVcShY
5EVsek+mO2e9WwXgY4oI4oqb6JohKzUIWFFKDIXO2u2vUMBV575s0+g9edCwL/7DiqpCsQXnrzHM
uhQ+wdd6HmopReLHuAb74G3ANUUTq+uIoIzntKIaWYXDm6C85JpPnER0NvFUAldMlQt3RCUMiKbI
jn+dU3GUXtbeL3/sMWt0dLHG3dRPIiIozoU1U3n5UMJooAfvuOb90PbxbXP9U8pI36ogbw7TBKQE
lzo6mNMnvb++zZhOczvBdQ1+o/zefKh9fEWBQgoOuNPOpxJH1gVg6Nq1D/bmqjl3Yz7ZT83Jcahk
bp+NquXpHR9WKtCYe2chWfjxbINF/z3Z5nQMsJT+f4JIAwbk+UxqbJINb3pcU0kz6zPNeqQ2wvUk
cpqgENfn5M5AZ2XW4wTSVIpvS4KSGrwRCIjaFRAIVvphaPznp6uSpYlEMwfPMK9cvbERRGjFzDDd
jMCPI3aEDnX3YbyP4QYKwCavApVXomSgX9jnUSfImlR6KLw8MmoM7qcfQJrc53+00V6GsBZMkJAb
zOtHu3zcFPFZuMsG0VpG44M17Hbb38PRiweUB27QYWQnIkBEv5jWNSxpPvxPfbF9te8piVAsJbjB
y4L2ht2PBtj7aTOI6CAE5OA0yT08Rpy/93T9QvIiX7qeE9FM+cfMGyyN0pAHm37RLvoYY4rYs1il
nCozzkCfJ53rB7N1xSd0KdFYq3apBMbTiStc/1gwOWPwqGaU5SN6OVhLMWJTrWvwfGt6jB8NyUQn
qYqofcd0zYezjSL24bzIjhh7gH0Y5e6SMDgVduTIzGKxJtZST5Fwuoisr5uikPHFgWWdlcNwdT72
3bGSv/1Ii/Ne53X3l1bOGOGCHEPh7ObMvsOO1Jq7fiylCeiA3NFw9u8NBKQeqYntc4U2IHOzZWMe
CMwGC3qQg/pxT8245k7W9T+pTV84NGOwlHeG86pEnUZcGdRoVm8RBIczjReFzrMEJxkZP9XHxE5H
bNe9tWqfcAlKo63V9ugqXHIJWhOcr7ky5V9R1doQZ5GsxrW1489JG6wXu4zErH20zEXkXt0P17ZQ
Pzwmni/3t0rVP8anVUF7nChSqLX1NL6hEgTIOpvdpnPNB2D8/hCtmfn5fjCF30o7EKcUJKWXg0FN
DZ9LK1ctZnduz6J4ZaPhHO1uWf7PGZTC/7WPdOtcOKdet21fcC+sY7pBJUyg789Eyt1Y21e77UsS
4AiD61shzA2Jrw2ZcaugtbCfywA/3VJSh90/4Kih4CfY3VSIeg1XhQGSCKpBcXZB6UdaqGnMWon1
fEFN7UX3riuvESlK65ty3EToVVua2RPjMrdByN6gvVlRntRr/a7ue4QEoFFpUa6Nwn6xkL7a/iDy
d58nZXiu44MYKku8mAWRqpBALlD1ELr2zVr71Yn2BRd4PjS7zLFU0483dnLmNSxaaBGRIuDJk4sp
HUikz+72FU1KWFh230VkgPrbtuzDNN+CHm7JYgcK9gW/Y9Frxk2hY9EngKQvcayalujxak5TaZSk
XV8zdS2dpQ2YZwElgqLgYnpEYdJ7BQzQEOkQurK7Vv4cJe8jeofJlMn03ijYvJqVgnFGfIuhrY7x
EOXzj4wNfitl0H8AedoQw9h+KwO+XU3yaBmTVttwS9PG4NRYoR5x20RJT+l1KkX8XLa8Mc8PdTTy
Jizy8tkTFN5/+kj1lrFOcfkZUEOr6X9IHVPsnLQ/nNcxe+ckcnWSC7Ig5saON96VQLrMcUBrDFY7
CMIAxwey7hf9L7O5M0cwXgooZlvYnagkLRUtdaCDGIJadMlgjfHrjT47ZmY+b8e2zY0z/lkPZv1v
FfZ///JsDJawS/mCFcHaQQzgXCe6doYzoFbtf4WX+RsDNzMkIGLVIb6bMCAyo1/hZ6NffRlJsXzn
WqcKZoKruBOTyKM8TfPxN1clBTm+sFs2jb9pKe6OSAEtW0k6ZnHiSUcgCG3YSmTCwHSUB4rzeLzg
81fqnHoBqt8YUEKQD0ZCEKFTtUFidJ8ebLqLV0POZuv6estnDN058iSuE4sgNdOSIsDpgKFhM/sJ
42xU99SHqv+2d55F6X6AX8lonaLMOwrrQhMHiu9SJxritaDFJb8wrUPKr4yQrEXvIK8rdCRP9+1U
GlFlATvFqbq+wT0igneN3xCT5GDbWUXbt+4uvHb00cnnXN2GOrC6fXzBKni4eUJdYpjfh4t5Fkp0
XXQK6kCRZywPe4ha1A3S+ptUFOykPtmJVu20WrH5ydmPHo/Om8ZSRxSashFzjZCOXED/iSJ289NU
a3KHsHqJqCYAlagG3DsNNuTaiF6+P5qgxXXjZbgF5zMrFwiC92rppufKCDb+hSKrg36W0quV2+Ol
86WAnJYTOcIJUyhfLR4NJoSqnViKzyKLXOT2+ulGBMJ6mVB9VtKDyNbLlyGW5WuWNoqpTauEE7hi
JdLa+9r/jJeinJBqy5SoI3iyQvMYMqc5RI/TCO28RcU3WjdLPL5WXjwcfXId1sMU0BF5LKj/NKqL
e7APT4potXMTIAclstLkgTDE//HfAN3gWYLGMS4vFAcFBtNnUcETXuYMaB6wOvrs/y2MqAYCwcrM
t0fXzVTZI7BzU6wjlvWLW/AB1IzaEXW7HUZV/F0w/6DfDwweWXOrT7O5EsUb83/mBK0KD6+PEuEX
fh7EtUQT1rgjhQlZ9VD9e7p15PoUdCy9ytATlDMZtQAjR4rY+4otLU2acvqjxDy7SbfBVInA2DJs
OlZo4m1m36Cy97w04cygKlSI9ViYZIL5v369HMYdKc7R0bl4PRc4h0GO81/xdgAEjZ9FmJyDWAxl
+TDuZE4K66QVl6jb6GWzfu75960jyeD7rRqPdG37VRTmbPd6QSIypmTHwWfT84Inz15nlbXDEgxB
ZN7NHI8IClhCVr6y2JScH0T9TcXstpPr/Qo2BNVx69wLh5EbVIKl567a02vvfX8YaKqlvaYxYQF7
+FZde8oaoPl4+zLq1W5JS7euWpGbraBlR6Yu0GEQL64njS+iTfjdMNcN0BloM25g2hI4LjUAoPQ/
yGBEbFNiqRfBC4qyW+M0FAqTwhIn9xAd5f7qu7+5YIhyhYTYkhoTrondrvIvgoQvDWXue+yXFsDK
T/n4cXc5VK/wISnLN+82ul5Em4snzaCitZqWqU6T0DGxLWHoSqVqAiuA4lnbZYKz16OMllkL/rf5
s6pHaB8Nd0SmWIolDbY6IB/nRQBL3keB8KcBPfzMlesS2K9mVXYKQgcEuZZt4+n7MgOvbquTRW3G
5ekwbWg0kQpSKaWWh0M65CqQTiCXhUDGqaG1uEOGpqPZAAY+8zU82cJgv70nKIfekVnDkg5EMWKG
Jp1LgvSiPbHKpNH5VkcrdwWq+fB/ebgWsFoOyeSUxwSVz3lOALaCKOBF+P4PRV43C9UgxWHFiDWE
/SL4NytgZ7Y3VxsPBF24LaOABV09RUYI1wzrVqY603zV6h9kz1lErTzXwiI2Yi97H/kBVn7iHgw4
Za+JpeaDZkuk+ge5F/XJOI+zzGXrZiH9kW6KsqWYYHUYRUI+RWAO/Ry2sgDQglLltt8wjQ2Jmlyb
4ixXbJkjutj0ghnrxc8cyjAyQcG3kl98isbkO2SPSqpspwo8eY+SQcvMjGmQIXqpDXRlZroL9tM6
ef8Q49EMLYgcgH9ZorU296jdcrv+mxsUvkgq2u+UeIA2ybb0SJ/IL8W2xyV6JqrYQJWXZ9pwwQqe
mkZnBm3EUuN4LD9ppVmXuDiuVAc1bris9UZf6/YoL1xL67B8gszIYUgeKj0qbunLjM5OSpM6AeK6
2T9WCjbF9TKIH8mYmysHgdwJ3is+v1ZniP/RrLjC/AicH+M8sU1kPnOyv7MkB4hEPzmhODYe6V4L
nACZVieiobPulvx4UFDEoL43n1pIVwuclgCfPuBYkDt9E9cBBOgRLWeBhMY3nNti8vHAvDGGFqDE
QSicdULDO4cMfU1VbvAFz9rN+y4xtkq6lN4qliwE2ptADjuNKiV8ndOXMEPsF8eImIbEV+oAKenp
ehKrpHaMdXOz5Sni99Y69VavNbff4qddnxioHmRBPVCntgl1HN1knIe2FyC7uDqjydurSFiWs2gK
ctyGf8Kc5zRpMoyMN840Ehto/vAQQQR6USmIJvPfeBiw4TqBAJMrFYP0Mgx/DcZA6cL493ObNxxu
JWkXBWadwaeFIRBC31W4J4PiWGP0bsdRJwKkx/I/pb6Cr0tI9RBWyDQcMr19XIVIWA798K95o35X
I1aDfKMLzYUCWMReMI5/W+smEiff407opkMUI4iVePZ/jCKIc1k+O+bp+BKuXqtE021rC5lWjht2
ymdEbSx9quMuYqGCRXrgOgkOi5ghq9nsqgLKtRbnwbeORMT+9uQUaO5TupPhkrzfqi3c/jD51pi4
u3m6/rtR38SVXFg9d19cl+ayea3YvHGaj4GBvdeqGIDyc8y5hLLsbCMHIxEhzigP6kvf+lb+2ncZ
3SHYN89b1AzexjmonD+dpYnZavXDWLhiBpbM1bdGVxpE0Y9I91b/2V97jVuE6J9CI2+RVt2hIT9c
gWmgj45xjw4X/ucD39EGwg+6DmVgm3DBZSHG9S6SCEHq0H9vXXh58plBZY7OVoIdd0ke1MSZU7WQ
D69SncKcHHB7IoQzS4aL82kh7ITtmpDGsJ8MhN6Bwsia3rdjEE7tfQ8gDViQ8rhSX00SYhBdeQMk
bonl98q4My3fB0u59YP6yAHBcWhLgzvSMQnXbFsQ8q68DTOMdYB4E7SM/lLjR8PR+NHP4NLRZz3c
gyClocObdzV+2d9s2UJsT3qbuKyRFg+DzExXmMXWfnTwYKHySGvbTvKwNQCJm9sTg//i+TYzldmR
RiQv8LDYaMK08+Y7bs4+/dKImFSsIgPeYiMdU+vlVgShxDWu79vXqHp9F685qn8u0UcIENo6Uh7c
Ydx7vmKKVh0LoPZEm5XOpnlA+O41pcNzeXUwRnw4Jl7lipoT0LiQAuEmHCu0wTGfQeKpQM9N80aQ
ITjmoYAtxhzYxNsNVoLLMmE0PhG/3WndKO+q6I4WE1Qy8BhyxDdylu2uMHIwKdajEnAwvFsUX9As
MaxrWcg7LUtedTpelmdDIzo3wjjaDCxnsdT8y5L20WcqD5d0Cd/YR5EoiZHqQtfX1ACM+TIvpqV6
I4g0A8nkJCAMm3ov8UbA37Y2DwHqdfwXBWrr8qqGW4i1A4H/fRLmc6/r2EuYeXqV835gsGqnk0VA
aKjFka2kQU2N57G+gb5ZaK1rZWGTsNVV7KaclE9hSelZMEzO6xpu/2D2hTvRIX9xubj6Nox9/umS
/aD7Of5xtNPurUX8z/vpZHTTz0Q1WUJWb0ed78Q0WTQIdV/QNRA9L+7yoUNDT9yiBXgdnrgjVT2k
ne675G1kPDOibHm4yDf9CUUqriwumYlnlYJQSP1A6nqF23kgwL5BuxbVTXky6ykazq9S0O1T0VuS
iN5WuiF5fuDN3sNL6hM8BONGCsU22JBCLtYbwSAShZ7omFVKY7nbB7UHGL+C0nBTz47dfs7M8647
+6Jmjy5binsTlpx5Dq5Rs8Xejoej8JX0/kgTg1iSIbSYGZ7noKHJSr0oLS1LxYXxUm9shn9I9g7R
eG90qk+gywSk7HZutggbb+PiQzc8m760EaJFKsBFDwLdXZ5uyYkw3h99ZKuptQGBVQeI27UPlqrq
ZqznPCISOQQnuIhN4KrUQAcKU0O94TDgAH1EjcnieUUjxKswYKWc0xDYaNteHtgSMAeUrZp03jJz
mS3xVfCAxeDbCK5Ya6tMoNhWevSkqc0OOE4Mz6/JSJIUqdSvifo6Y8wj44QTS8WYK/cwxWeCiB4Q
RNw4f2CUcM92HN7jnAyxe8u+9N8IpfTJo63lFGYPrqXEvyLVBaKifkKJ6KuaaM/d7ZuH6xlVABkA
vcJJbznS+kmHi2AusFmFFQiSDhbiLDHiB5uolkPdPHR0NzVFY2UyCW3ZDjrCou4AL4w90dQtPVmu
tf7U5ZBxY3zibNiVNieJO0RhqN1/pHk/MrFpsDWiWX/hwIhPp98CeAnQlqeG2v/VnNwj5Q0ON3aB
z8j4R0+Xd19q6jgnZuymajFsjpt0yN31hrFmp/I5IOwWcc/AeMViBoNzjGyfqTRG7zBcpGcf118k
Xbh9UnUGHlH8e3EhMUaMOHOwKtjrXvh0e1EbrEUCWVhyb6ANsvJWAgsDVb1i4AWZOs+/AzMZm1Ce
rQwTqWb2pKMm3BN8GqCisidqnQVJSWMFAKtRHUIcjTtI3stpa7JFxovWoTNPhgpkv634BAScVuHx
cLgkYYnW3l7tA1vOkv8yX+jSdjMf81AEZhx2gummOJrBMvxRlQmNJRUADTLGiyb+wsnaf16bPHU8
cmfTraeZlc2LhUj31X6MN5dRdB93TE3HlItQ0xzBz05uuRQijAOiH0DYf3kYS5xw9p9vsL/qnE7S
2d6hfgYHe3dKasC9oqBOwn38EC9lwB09zQJLmGvmbAmFatzDKbc7Fu5YO5vywsQIznFXlpMEZVTn
gIjAh/00IjZJ/uswuCR7RSJ8WqEuM4OI+Y9PsiZsxzwDmv7M+gxk+5EzdR5hJNrWHRkDjiylpD6n
c8BTpdYgr+wQgVcRWLUmdOpYAJouxLZuzyoRYRb2Sic/V2qZUGsWyj8k21C8zic4GqUWuHR3e9BX
Wvwd8A3+XMn6ZTXVOUUCvBrDXF329S+D9kobNsJHF0NEj88JynQw4dn3EhKk0Yti+NLAXVKac6Uv
RCabwELaE3mhFSUVivz0eCJrDxwqNnprPWsDFc68tSGZ4NKcOVKmb8DXZu0ICKVdpQFE9N8kFzZl
vxL8aaWZkKqtptBZaKsxsR7yLARai2j3uaIfDxEW7rL+xHVlX1cG39ACvBIK4TefYPhQZXmbTA11
8kGCZPQmSjPDi6nLwG9yv9/zr4iWspB/LhoEwJ8WRgd1wmBVCFa/678UOD3levv3LXJvLXi6UdX3
cxGzlvZLMAttd3Ukr0qmPVzrj5awQa3Qj7ZBu7jHqJsl9TAvVFXzyEhL5v+Z0fGQywDx51GvgjK8
6YnibVIHRSulUPUPT0UG4l74v7Fa9zHo5qi2xctKGS3TIBpR47AEMoNdbg2Y4/Xc1mtFiPQMjTcj
uy4okf5VflylZsC0jcR4QDi+rKQD309A34TXCTb9g8y79EuBnlavxInHPuefCqm10CiLW1HPoQsY
Tz5qWjZ3ZTb/5tozAUhRSbV40pTY4DT9+G0+TAfY7hGSuwgf0/H8U+lxwMtyh8nOQfmYRFeVJ27h
jz6MRFVMimhZFWW4uUgTksPqueojH4Ij7EnwND++uCKaCECEHqKrkWSF8BZ/B1mUwfVziOtjFW+r
KVAaMb4+AoAHLPMr8NdkPM8gYSDZGkaRScM/cvwKY9yj80NFSoHq1jGXGgOMZJegBrJHAzhkboEG
ZDr2iFgunaBGD1FR7k3qwDOWEjxwgby31vfP8850qTzzN0SHmE4KshtHj3BEXMt+vZ8sbyPLyhot
CXvnXPyyOOpa+71AK1T2xrlPa2cPI93PR7E4fB0tyZ6dDyS5CX+rWACKu8qKqyydMEsdxpezOGUG
3FnBUjBCue7GaYT0DKz8fjO4kyYoPzcI7Vns6I+IMt9vKSWdl6eww8TOUD8p/3yuQumdOIq/HSXy
62T/1bkIMan3lENCRBV67ndvZaA8Nv8RVFI0S4OJGWFP5/VgPi21PzXoATwNgNXZpTxQ2oXweaIb
gp74c7yBVjRZEQUvI8mHJ5xS/83l1Z0rc8bDETxFJ7NmiKXIJ7eUzYHkO6KEw3VhL4HICjpRfJzq
g1ZYqiV4HKHqPkhIcCsHmTZF6wtzQUITv75LCV87tEkJliGr7KGLGfKqco8I5/DbjthF/BnFdtNN
sK6v9orpMEc0ypWAaU1HB99huN1+N4qPVD2GiJfDxXQpwxCDMKvWuwwHAQXKpKfPz3JLRZYy8mT1
iZoO+OfMJMXKW23fgw5Snwwaswccbm5KAW2M0I8gxggXK7cichHuBYWpxXg5TGOlyfx7E9Qmboax
3XyIbePvOi31zQB65s2GkOuE5c5TRc36Zdr8Gs68ctZQoRbuqA5hj6HGDS+pwd7BxtImm9+5zmYK
PVXV8KpXPNV41M6PlSRzKF4xlHUOtIUeIKS9j1OJmXqyVShjw2qqXffKK3I9a/MMD8zvkjuqvgXG
K6LA7P3RO/Bw73od8+IEL1SROSauOi3jEQ5+7cF4S6vBPulV1fJznTv/cis533cagkDZT+yFtniT
gj0Q8hmvRd3D3DSt0SGgreym7+Z5D6ONBIYZ3+Y/Hkag/+5n6lDCzgXRm+QlU/34KgQSlbOVj1b5
AOsxyOAsv2/+RXchYfwqz1VVANNHaycU3OUXeg+WKHsxWo1rLE73F/dm7zvmmhk1Tp/my53M1FsJ
H+aFqMpUMVuJkr8O0lCmKm3qqvMYuDtYyR6iI+GBKZ8rNIKVUF734adaNAg5Yud7pVgGpc639j2P
dvEoI10bpyCz71EeuD77A8vYu1e/lN8x/cwCQSTTYooCe2f0QUoPhbnjJUC3gBfkS2yhtLD9cpk9
lTm37tTy+Rg3swsKPJ88BEZR3z5s8uZSNPsuz8khv41D7sPId50+UVR7t88plxYGXzIb4UcSYjZu
U6jNzk8IWFBXNHusU54LINGj8I79FfyNDw0gz5J+PDZrQF0jOxvJeexxvDc7hLNNM+VdD/ZMRBXq
giYjFv/xzFjx9HmegLNpuqdbmrG0xdsinTCuZ/tqRZLGk9LWSQSaylwcC5eRyBbOPPio7sl7Tr89
zBbdY0sWNndt44SSSzJ4RSySXFlxz6zn3St3n6SXAfUlu6Si2MXpz2/EFJbMY4CKb9KmxExzyLTB
Xn/+WfydVLgEwUUxuXijMgWZFaXhuEPdoXjeq8lxsE9WZH1snwXr54aK4NyVTPe8Re15tSxhyzs9
WxlWGwt4lg7wsItjwrTKCF2sY2LtVi6wwx9T+bcBO46v0V5nkqySdtkb3C6SinZlCFqt9JF8C3PP
Ex7F1rOzAwnLfw1HrseLOHgzTlatmW/FXHsDPIl1pntfz4dKG2d9Yl0Ajwvk7fkOPQ4sEW/M5MpT
PA/CiO4gIzLRiocXIQrIgG9r+PyPNmtGtF6193v7q1k1ojxkaI7lAmzCVAKk2DbeaOQuaHTEc4AB
ir8+mh1tiu32fsIEtHxcSFVfz3JXCh0+ujSE0dM83RjanbGOPvEPaWZW4p6Gn0Jq6riCzLMWxPvp
qg/YnCIHZLNJjt3ZW0iQ+dHSbCYLs5/FeOTSes6wBbp6KFOy1baLp+mNGGEyAqhnthGL0Ul5jamA
5Ru/CGRrIBBUSTF975mZAElycOsmabW+by/UPnkKPTbHcOdUPy040+2AeLzoKI+xyoNKlzJ3ZgYG
z3kDOJ5H0NLVryRS8PcUKmVLilG0k/doyG6BxhzgB+Q+uBd82L12Xw529j64yCMutRg03dpSsYQb
0TLqvwjt0h0VVFB0kFEn3JJtQTmZ6n+diSqFltH30O084gbdoNF61VJkobSWlzC8r5yfJ30eB44P
bcsu22e5+CH8Zxxtp9cMheVUVg6EC4+XRVKwlXowo2h2xywuGPuB6OlpH2zaG7jWcnqW3yHRStjp
qDo8YL199xadSnX7aSo8VprsGJzOOf7iYLN1BTOmHIVOLZUC6NqA7Gw91AycCKd7iYOClRh+jq4J
zS1HLWW19pGXiF3aWUtYHJCed0hr0Wp0j33qloi7UwDHwUIftOzKfcfu5dgotsYI7au+AGgelCUS
2QRQpUi2AUMx1yFnNzor6EdPCTlbelMMKAue0s1Uc6yX1xiK7Z3Lw+hxp3Kw4g9O0aXHoFacAuG1
jk5QN54o+j6EDOO4cULRN5G4KL1PSfMG8eLCAFMgJFwpuKagYEPZyvxx0JzPAfmxeTsrXJ7hbdfM
p+j4a0MJkLTuf2YnWjvEr1+rZqNsle7dh2daBEu54c+95GiB+MhQ8NL53w8XpqIbXAH43t5dkcke
DSLH7HYFdWY7nr9XpW3h9/8ECKWIZCJbh8bl4HuT1TVUEn07hEOEkq+WkcR1xn1iQaOMKB7gw7TN
tf9P1d3RAEe2NktEt4LQdHQl36EoAPJQnnOh5OA2zQiiTDxj0OZ0WoS+93Lr9XeAU+Mbd9/R6nq3
4O0ax0wJWf46vNPrf0LAh5Z8KFD3dNCvuDEAsyCAAptN2lPaVn5DSMT8XJTVga9MKo4KvholRqyN
wBXirLCdaXFlqVFfauZA37IEEDQ6Q/jyNIVs7+osKQqbn9FqdRlkzsF6IuUCmvYxUTKcTcbjQ/A9
FEO8SvpBzk+YsfvDG4105LX1E0gqqbIcmNwlNf90soUpKGpKBma/xbTpGy9YwU5y5m3MKT5V9y66
rr70pVjQhWBGCLfDTiGEasA4IGC8gfvCDiPo0rkY7fd+ZK1f9FE3eKZonA2pJC4+viJE64wlHczD
rFoKHuX3EfdVl380LXSsL4liOkODaAz95+85JxQMR+Agil9aYg0WuVPi1Z+mjKn4/cZwn7FwhA02
r6lsVItGHnnD52bFv+gOuTLIYs7Q/TB6kz9jcD9yXptfeWqb5V12L9u6kM97h/8uXy0mv6JRmIUx
K2fgBvGn2x8u98v/qbTXrXqoq/4pECH2Cp3XRTbGYspONs5SR1/9lWiuvRkLy/VZtRrk0LIoqBPa
T7pchFlAAXg/eqiiOptOqOua/qd2zvYqETgIitt9fNz76zideI9mKKoxsCUPDfrIQ9Zi3XEs2qR9
Zx60eQeVFTmoSm6gwryr8j7W/4KQfjNsyb2jSPB40IXJAxYiN21xPvUrovYgEfbnRYN9Ii5uLJZZ
tgEdhttY7vVUXmaEWYq2QHZ8VyqRfCRrKgPLTutYIWWzK1X0/vJl8AHFV+weLG1Fw5XLs/eEGlNH
HiV0Q2uIG7UMGYDhtpvcnVOP0dR8J74/+ZZUdzIoT5SCcIqpQQb4KmdegNqXuFuOqG33GkHSwGJU
9yO3jS0xfabTroIoSL9tWWojX760Jqicfmh5HrmZK0caRSTz6gdeOSo3bO0bn0nrFg5kLEzxqHRp
kkMQleA9qWpDBScBoH/mEoOi0b2CVHzM7ukBOwsnmnID3bTON45NUbWPBrjaJMTWN38rHqkgdEBP
IR8bkbDJDUp+ZW/wQlPSe0MBahzyKVj5/AIaNDuSwRjCUwFXTulcbIu5Zq4edAfNcFXqIllcZR5x
qZMd1aWJupCq/u4l1KVhIKNovu16Q1/5FaITZqjUVQstlnCJV41xQ13k9dieb/e/I8k5stjfXq5R
vvRDGtrp58xlQ0tBxg8l4J1zT9CilxEDPJEGTcoE6BJx/5LhDkaXRh3mJAaanRyvOPLcUPw+Eyq9
VNqw8HZFoF0kLNx48B6eObYaCO5SRmHLYf+n4c9jC8VMBdmPyePhIkUHZThTzp4E/gM6R05HhJIx
xhQm5W3c0Ym0alkPIi85iUYrpPEHbqz3BMDUdT35O5NaCf/ICdoyNkzEa0DhklshSX5GOqX9iLfW
jbKq+LSIwCGJOTaZIvovmtmtX8lh1wcY/Kmz0/0QoiOPH50TFTqE5MajHeDvYinUsuDIxSOahkSk
MffSz+w1qY1yzrWqG9j4mxRc0nb6G3pFhfj1btxKHQKBDt/67bbFnkn9EYG9PFTgnV8l5YuffhiN
Io2GQgWxsVlri7WD1RsD2OdeyClvIcTgHNt3coClkdywECOsL6W73Yltt5QgyzuRW06uC+7NEULM
u8stt3VW4BHn6Tdr5x8HhtwhPMdgc7qNQa8m0fHLN0U58FzFEK1Y/HVD5fQXIPtTwx1bJLbh8/5g
mp1ieYW5tQN/8QGTiPS5OMD2ETebOrE608CQ0FjZ2QlXMi4Ujd1Mgu3FpYdE4aWj75MZ+3FA00Zj
fDhDr/sqDsrKtI+z8+uK/o81VO5Fh0ipjw/NfhDo9rMPnMSv5er2lbmFcCVnwnjvJfaMo4rSCUfj
bMooY3WfgsJV78o4o7mA38bESIWCRzCCBEJqa7rwXNKZ/ZHV3vCV5t4tLUMo/vmKioCP4zCato2Q
ODwkwQgneiYkvDqhexMMdtHS5PcZufqesFnVHUo96EbUEzsht9EsTl8Z9Tf6ejDs0b/k4WgtWfXz
E8csTKI6C97FwhQJtb23Zf3o0FBAvGWRmSB5qj3In26xuBD09bSa7XxMsurmghfF8I6Lifm7WllP
aNlQ+cx4ZMtntyhqV6Zl5xEVFrqd2LvK7ug1eOl8YK8gvK/72ZeBxG3LswDv5ejPQ6Ej8ezyj0/s
+MEXEyC/p/8PjEVNu82crnnf3KhkBY6DT6GMMBXRcosOFYhi7rENhpo8LAsIQkOEkiuvzsu7WcQd
hU+YlZANA3s4DASZPhFql81sb1XKinfIaTzWaN2fTdDD3HhWhOkv+tdygyXOeE52OYZ+JPEOZ4JN
F4m1ibQjJunlZJ/n3vvmdBxFdl41KSMInl9fohsvBggkdE5Ef9ZH8fE6gJycjmyCMYWlTsB6SBsn
BCDmzZl7yk+JKSBsjVeQ16WsRBMmHxmtbzi6pi43GxGQBI/E/Yo/jyWtjghnYeA74DcQHkAYyiZp
9QVO4VnPxJ97p2+WixNrKZFYWXLIXOxudDX0jJeiSi3B6XOlr0CDDbUjpdgJu6sGhLrSezTwhmwo
cXjQBdRDFchdZL21nPd85c5PTHInzE/h1OWRwtriQjZImKrHWpFKtaFooic2PkLwzI+dD71W4ZEp
rVErNyHIUiqCVym8p46PddtIYxCBJrEjZg7hXEJaOm5J8uJzL05EkpweXLEJ8P4TxVqCn4AyJHey
K/iYQE7FlNz0I9cd97dcAg/SW/K1RZR4bsLNVLRDxrGmiGFt73uaXdzdXwV1AtVqwn/bi4H9eoli
UEhOyplNfVAXNoFyGrl4IJJIrmNAx8h/AMaOKc4QquWD60gouAmiHoiqbz0YV+Tk4O6H1tGKsMHP
ZMsFwJ57krbVJouHFizRPynJPobjJ4xVYXhOWzmDDc8QCyFhk0ZqMPDRqJWQCpRsST0lJpU1PaqC
prMbUXqUCibk5GPMb97kpzH4qCiEiv0MVC8gwB8R/JDdpKMpzGMuvIBHEz/YcVO9NiaMwJ9mxz/O
2Al1XtZq2F/iymnUMEDZsl/RrmoopZqH/Gf87VRbzdsvSydXO/qmA+6p7SRLoV+yzOT6qLcQ2abL
WkMFAZpgWHM7CAsXYAs1U+QEzVTkdTmTxDttoPR9l5F/KMdlq6HZHoTPUL8TOcG67I2zrlC3+4J6
uAtS+YCtgT42RVBx/9RJfZl++WnTJzLFD7YKITAZ0sIdu7HbJIO+GzyFH5zxc96b5d/tZv/lWvZg
lrdzIGk8IUJ0TmhADbVtq1PRfgiyW4AV/I7UXn938oxVZWp037Y648TGqbBjUJ82vjJSQuTFPn8F
Hrgho/InOIVDOYFjRw75y5iDCX6IfeBMI+91UC8TBMst3pAyj5qoFcOCbbcpzBF+VyQ/sVwjuohd
B7A6Z0B/Id7HygS2U+xXoZS2MqyJkOU6eEMpLZn9KHkYKKOd5zFrG/kE7na4eJBUq2bTNTgSgrSt
mcWFSYMk/dlb1gE/CNdVvsj1v3AX4YVOMse5MYSoyNAOxH9q9MJtEegX7m2xGJ7xoj8rTPCWRyH7
RaG0szlnXmsofa3pLNsrpKxVu4iCHCzgs+UmMi3o7ATJ1vM16UXE1qkD7PFaFuXsHMyztotQNGHx
3/pZLnDRIAI5UG4gCfQScSKYo0zMrjBI9BELhC4lJa8c08qnemoYLsqSeRzFiy05/rfsRyZXI5jB
BwJRANGW3au6nqXlb8FNJZWjAsVnho9eaoePDRVGcyEEYilIcFVHFjsQrbqQC8KWpj8uxLBDWkQN
9LIOgFGgzBq31sLXSubCulk1JlzNiBfnzibQD/kI9av/zXG3rxp+EhYHGb6uV6k/rQ8F7R6qD164
utd2AZDMaUWtyPze5zw0kuc+TEKJI7xXZ/WV9Aa8b2uisLR9eUEHbkE7+TmpnlAMuBo0PRFXnaGR
cBvawUqu94fvdMudwyHh2IVx0XtDQftR7pvQhDIHwsUHxTSYdRjbqtGKPo1BLtPO31sxtZmZNU9D
gxdxTI2F9vbALQeI29I2R+5iMfBCBMrUHalSktzf0BPs2vvq58T6v4gakmBk3fLwgD3oFLvf+vMe
mg3jxh0t/SXfRXBpk2bSrhIBSmAlyxxDEHx7WxDPz2isZ4aCctIaTyoOeCy9+rxqr95TX8RnQPOz
b7cA4CmvFLT9V34etfZgNIpwg+Mmt1qUbiFwM7wwoSEYyATju7HLOU20FW08QbVWWnvC7I8kiO8R
rfFmDyzoPtELlMB/aZ7gGWlLJhzSoa62gMyX4eU/i/MzCMUJhuMxMG7cJ+0jVHrs5UoSw83AHNts
zRIlEKgkn9Hl89c3dNYvVZi44+nXEP3RI8vgxx61/ZlPF91KOyQV3ceGfyXyH85R/oMNpaDLgBkG
FWGtehH3m6YpeeDj2r01zUrQuY8vXf1B9VYG5HMJKuWelCXYZwz7Ok3zYufQpoxZRV/rUQS3Wzhr
3V7Va80ry8HBz0/ks4EtdefOjQflbiAtDbhemzmNDN2mJBO8kz6ev8D7BNYJb4eGJqT5arDbBOYX
5iDfL1jOuuTlhZA5HDgQ65Kz/ApH8Nrl1IZKbJIxu0QMbKJwfPAxfvmu0BEFJgcJ61oEfMGwQhX6
pG+npw2OCAlcMRFFyu+UK5XmJf1LVVIcqXJrVv/X0uMYIh37A7F0z3uLNYmQ7ceu9bxE1tgAjpPP
rn3wEmxnsZEyEDbo/hd+4mZxp3joioFrvtlOlD9wzTeGIvUp9swIP9dxYzC8Tx1JX2TtLRXfxbID
LkCdDx0a7dTFkWMj+c/ITSMw6FwV3ZPnNP9Omk+LCycGRj32vH67Lr99rv9F3DGmAvsO1i1hVzPI
BU3gwsupxaZw/a/dbhBBzLHMlCqmT4q+WFRkyADYhUyAYl93yk92JIhDYNqMdgJa+3u06hzQgrLr
DNFUQADd9LsHPYc6gYIvXKOBxXdJAJPtd0F/PaRjSZbd7lm05jAQnzgy+qE2wk4mcHBlIKx5TS8o
vS28QIEyRYEiVvbzxyQEYSRZ1c4gZgHxDtgF/l+deplscPgQlSSfUMTLFNhdgjHW+B7KSVNV7H2W
YzAVFdjTzXJ9+vtYC0gvhdz0mN3Q0QjBWgvALchxwHoSqhXj9j5DfZg84LoWGakM0MqzYUM4nAIT
mL2hc0UbzyQvVoOC11b+9a8GIotpVOAqITKiZCLTXx+x4sS7LXY4TdKp+VX+x5dWXPOhv8uqrzyk
dK5hY+s5dA9Nr1U0OTXJgkacTyvrP59gPblaz0cn4xVRNZLBWs1+oVgwOP1xq0LNO6riWPt4BFq2
Tt/LDOOw8ntCJPA2d0qSEr3YEd5CSNAgjRd3W9jVaW7WBQmqf+gnKiKS02DFUDWtq6p8HJoDY4UD
iKFUiSwehxNDwlNbFeUNEbxseY3ApATFimfOqfsdHsNBh/fHgua7JdQpCKMYQDSeoyeA8W2O8yEh
plQY4P/MsfXPmkocQT06JToiKqRsSnjWOFdLWU51XzU6VGQBdOdxzUe8R7Bswh98o8BeMc94ygAA
t30v18VHS71dzo/itiQPAkDwVLv67NBspDO98pyh/cSMddux/qfz92TBbagn/EXdkXXNtCdbROFY
0KWbQqa/AcgcfGX6WsYUNKc+sl2R1WE+TiPH5zjhtDspgAE6QNSORO8mQGJEd+RblL0FUZhSA56N
07dM/axCQfz06JQFpSVRlQdM9PSB2o6+3Szqjj47fGHlfb0oqBPqcOIApUi90YA6tsC7tHlGMxHZ
Ld+ble/e72Cgi3Ra0zJ5+ECMi3QgfmGwPsMjXNEXIZQ3MyWYs9l2eP6MJogMYQIelRdiCD9Zndb2
V5izv8WCeTOYUlF/NS6AkfUHWzkHx3/z6EA9OL95oYkb0gkYlTpez1F6BhOke0x6BGsS7/MG+98g
QqlS1NAFn4nKd6BKoFhsGSGNdgkQk1xVtY1r9TqRXmhMD7kVFx+56Mko/UDFVbs37cQsn/MY3/5L
N7cs3pIRJAIHTrhRv3Jbco8rUzU6lo4DJiqBy2nW1kp+8JQdqdAFrTgJ32e9TT6w0SmwsW7TI1q/
r/TrmF5ersjUqhPlDOql4E33Jq716rLkGY97u3El+JnNRvjnQQ7jdluvVzrfF6ImDeFNQtrIJ1YX
wLOAcqUhsoib4pJYgN5XbWeaL1amTBpuQ0013XvJZlVFhUCPfSggL4nS6H6BqmI7DYU1dEMqJ/pA
kfuoaeOJ9NK2LShu9jLAZ2/Z356E+uNqLUM6+SQB0We1dSaofLwtgpZUcILYz6tJslBlyKiLwZv6
uIfKyVKWVS5Nnk5TxrlVj3E3x81M/BeLvKdjm8GqtIgEArLDqATtVjbaBY5kTJx0Rp27Ww8flm0R
s4VAKY8mHnBmpOkukcnTgwMZCsrFn06bv2PhcGCWAqbt/FeczRJVfgHTiPifei+Ef+q5T+SIhInZ
o9NK8faxUuhmAl2FfmcjX5qxiB+PX1iMX6zqnRP6wJWREB9tKKX3cGYIk1gH+cD1ushDi/B/42Vz
KItGbQTzPQGXpdsd/1cWMPoAOQPaYPtrIVKCG886RfBSwl05Iwx3sdAX8hnxE+xl/+AvUFW1KZPd
41wNubgnLwDp4Z5F9yzFDs6Vwrzk91BfQLfZylJQ8YWTKtSqGjs2ck/ETClNPY+ejSvWWcXS3r+d
Dsa0afQ4hw+6hPI4ptudxy3VYrkUYVX0VMnioLA6imhw4cOhXoswK7EZ+4eQL4CF8vuRAVizoQ0H
MiuqpFj5f/khT0YAhg4oP6D+zeyh56ObfpuU8lEth6433fsqwqjDf9y+Z0vVfrucPt1sHcmpF95I
+pG5dAZjWA4rMhgnhYHwnyzCjoYBUgfuOkcO1ndk45sOGf+jkNe52iZKT6xM6QciUwmNKDbKM3Lw
2aCM0zlYaY0BeclmyS5fCgwS0IxNqAoIOthuwY1yvw4xv3VthNuGoOM0YyiSAKQYWAxQ3ZDFSCVj
KJrLLWW+kXD3uPNAEzP3hcNT/rQBCHg5nPZpQ6OwTwAeliNix2G+CBsL8cgNaXxs8dG5eQk+jbJP
/Bba5PRkvl2l+CqTWb3bIvyks6fycMVxRKSdg1L55TiK2c+YJsOj+54CX5NiSWiLKmkNSYCrfwlY
oaiymG5nY5g1PPeVNGzKMcpdYY03jOp2ld9uJcQ2Z8oKLZnrPACTdcHKHS0+Zwa23D01fxAAB7MG
arBEUjsYsC33pXF7Ru6xSjtZi77BE/qQjeOyHOEgqhrIRQSkhe+MCkdTPYQhnqUDNN3+B7WvnL72
AfA/fxk+TY2FtlRQzvviVs7eq5W7dqjj0fUfqhrYvDI5IY2Wfb8e7kr5rOH9OjJ/XBe/ie2SaybX
JoCoAuR+p06Xtwh19p7b//oljkuSsoIL8AFHTUO0brkpoKiJMX6MhHd+hGmJAmZas58mkmgTmfg2
JJ6Vg0ebANvJrvhNRQiIZtVKPyC1ODc6OgyN8Ipiy+o43D5BnOfR6mwly6p22/eRnfiUT7X+mZMz
FKOASfH3kdX0aVZcWOBi7GkI1s3ygbrvTTxq3vFXwDS2IbwIJWm54k0hkSmA9pN+Od4IeJCctBip
fz011wdkFXe9uE5ZcsA3s22TLmDTk159GukDGizdg9qRYtY8TOKZ54y3KLMbxPXw9w0YVIIELvYT
0Uxq0IGKGuDFIfVCWfNKElvjOQ3KiXbFoixDuNtjvKC6PM1rn7rVaDxViR0jwFHlmCBoqePwoDHh
01I8yYMWZU93cM5srdDw0bKLLgcRmZXWWUFR/1pS1l+Ojpq7c19/mmFMmALFjt/MswDwUn/p1IOI
MQf6lsXPca3mH2PTs7LsvDVKwccK4BNjN5tkLlEqwJYMrLkf0OUUIoMNq/Bu1d2QQSHEZzC6nfJ7
4uje0n5pfNdBhu7VVe4AAWzyUDCasEgbAKMqeYYEnC7stIvrnWH6wlsXD3HdFBlTzHY42ck7XlaB
kk/vvy42EQUYnA8WTD749kOTtl8WR4bH6I1ywRjHAtIuHFqicSF1AVGxdhJuS6kdwltNPlt9TqNW
gftr7CcIjO9LG5M5bBzF80FNipektc8whWH9AzBF7xeH39CJ0AWeYCireLBncIRZ10UzZS9lQLbl
xhC9PrW85AyntdGKCuyo6nzkoQDbCjVi59SCoDfwuDeQLCZ5bq9u/i1Iiag0U3MMYbnKjiSeF0nm
5NAQhczJXFnqRFSMZwROxVqMYiFSgSwWDyhqFu925bpR0+tRtLiTi+Wl4RWlSveoler2+YmOwp/T
sApZum3mo7AzzrYBX7oVsW3ZxJ83STuwE0WfIeaI8xoc8lgu2HaVP/Kyyg5EkgHUFNbcW5yfWQH0
zwJtm9R5OqTMfeGefHJgl7NTt8cCLaZr5XcqV/aEGDEa1EQRvWEoRJ+A3wvOB7IqIoKNQOmV0Wxo
7Ll+XC6ZI5Fve48XwgwQHuIyf9Zi1hK0YGIxYJa4XT/hs8tGf91cDM+g7wuXkswg8SghlhHDkG4p
/ZNbxDNyh2lblKlij7hAcbfjn9T4nabXBYg+OA5rojIWvIMnkChm5howfOH430+MPDjO8uzj0qlo
SXIhPM0OKW/4f6RHMUlBxwA7V6yI+km/1SibGEloZzacQfRsoWlNBy8bHKL1HiFSK0p1BQfgqIpm
HKufY9uI8VhviNXKzn6E4/CZv3bzitJhrYOOAiDzFnP2py6sXeRuMSJY6ER3lFiWZ8Tsba5H0IHD
WmQlUs8CWd6vf7f9tEUAmBehRrmir0JV6MTOW8o2e/f6RXvkXbI/TYbq2NZG6lzmaB7q7iR261YA
4A2xSuio78C7zFKFPvcZaCpkZLObwBAoE5jgQdK/M/+C1Dg7H7ZL8nPM4gHHOplF+KOQYcKmPQ1R
qrFySLC/nCYrmf6ukuH55KxPIA51H9D13b1BtXto15FUTkTwoZsyNqY+snbnEpHnxHs+uu6qZHyp
29/jxGXDPzeK69JF4qAqFm7yBgzXgbK2aVCA03iLoDI7KuOMAMjrG5L2DgQ7V534q5D0wML7NQKh
/rAIY+IIlb0PODwItcyL4+oDC9KKxH+EhCEix+Y/OSeQIIZoRbQBH5dfIvr9ULX6tcK4ponF7fo0
gNEYjH5UHYSeD/fTr4oxZzt31U6q53uAOP0zykIhxEY5nmke2W13uep9VxcbYco415JQ8Sk8Jm46
VPTYCCk83RaYc4fhdFWBXPYyz290ECIr18UjdezFHdNQLy4bn42pO5NXR7iRRE8D0lyOSlTxKBAJ
FexRbqQA6KHajD/ITfj9GSBaW28aQ9QKNHjCigHZrF2atFFL+iN4NeZW7/DedkOS+9yQM/0FKKFt
KcEaQ5ogvXxtJC8be0oLoT8xXBNdNs7P7Z9glzBwgkuaLzERe3HMOv2HV6JiEALrsDR0X6ues+Jx
3zoIWmvpG7hzlDor1V6MH1EAFeJc8EyG0oLisWDRkjPUqm5G1sp8uGYZMKJzHwG1u270PDhvNtYl
yyBVzmRhCw6o9uL3n5Sy3cHfYIPf2Yaq+UKIQneLJw0N9WVqJHGbOT3Q+XqTbFGGSkOMkee9bT52
mt2e5cyYYbOxcb8jtXcqimZEX6TFA9F+RIyPnSkSVlFG4av/0wWZVU5TNXO0k+KYBlnwape0Geop
gXtys+j2FTaGrvn5xz7frG0auFBuEdIy2QC2euDil6gPDOaU6bNDDC1zmO4y2DLq5U+g+9KBIw4F
Tm3oTh9TlPSP+I4h5MIhqcWLqJ/RgR5XMguugyKNB62J2gfUTsTs7DZGoiKMchBrlWiQi6Zhrhnw
LpW280GDXPUy+wywh4CAh/rsorHhDE0QQ99rV5RKVo/I/1/GJdyu4NQM7MrjdSKi56ujS/ohsTCE
HQVOchsCl+EbrqaNfFTh5x2Ck53+4NtOfi6cc7kQXVTkDyaIK9e7qu5I16zAwr95+TPdfl36932J
nuhp6Nbdpirdoi6GbTUrNSYzcIKamwaSs3Lo88jJnnr3XZm4uXNEFhtyOkcjCgYjRQy+D5TCZe92
jRJXnmytOkZ4NXoHwX/9ejZTaJAYHly52d0/cui70KLADQlB+FSmC6XREYGZmBdEQ2Qt+DpqVpDD
EXVtnKI6v/BbJMWSpRsQUtvrEQowQltkzmtAMRZB8E/M74UL+IzKGwtCMidlUig5Q5oN795lZwXQ
8pDCOprzusostVhPZ/HqzTyAreC4Sb2kN71l8wZxMId9RYE4xphG0+KvfMjJIpsHOfCsgVcPDyBv
Up155u6NvVxXSfSCKDK8hKKov8LPhwtOYjuxe42zJkzRvCkKalgyi2BKekeHySwQ1o2WOmYxaN9J
uG+cXS5qMluz5WjjMs3AqRww23Jtah5cVcnf21YV2nR+mGssDIxIrDcYTfhX3106Pz3mgQJKmO6l
ZvXCpnwQ9GxlRZztIqJuF2zAkRyYNnxDg6zgO2jQf74QWXbHnlHonp7lxkAdv7qWi63TIxNDyogX
cih0oUS0WD/yQSEkmBD6sxf5KZvDIBWd9QfT31l4VJMr1ZRwKap3zJpPtPyb7F3CmOJgUzIajgiS
/rc8tsjOhusb0PgBPFnQxv7zcMBKUlPxd2wiMu8Rv7D77Aa2E9mft+xNZgUp9vGtMM8jB8BB2x7n
wbWXGOV955cZSSjB0NXRfCIHrJVBiLFfVsAneDw/zFxNqyAtUST5LoRXlGFcGC8/ZdYKgqUsMcQv
eoHx+AjnBq6x4oaPLKvMZHTeUhu1LdoC9L3AhOpDJNa/fSbx1bCXy7b00Ai8HXpq66SdqX7C68vD
lH7XLIRiwIIbBh7n7+YshgSLiZDYDCzBUPwsuI8hHZjg/krkZZuhy/k1pkmMHOHe1kKuWYEi2Dr4
tEhOgTLMPK2VtwjzWFR1/ypfJjX6cdAV5Ch2Pl9sq2GP69X5qYABHV6xASHxewVhjXaj0sk+nQjW
2NHGWuOlfU9c4t4C2/MY8aAmxraa4zD6lTEps+73ZEXc15MB1Q/3zqUwFLn7gBmONLbkMYj3AEEN
koG0wzir2yeB+NzruCEXzs259ccX39DuArknOj5wPdv4Nd3i8yhLwzFaQLpvYO/puo5obb3Dm9TD
J0kSicinvLuuxj+coXg4e1X23AYS3Cnrksbrs0TFfrBj71EVnV4e6Px6OSsFG4uREjAwgomuH3Q8
w/6Ned8B3BLZEpjQ8SUu4wWUA5/Au2tYcsb5B/v5LycX5JXeJi6Ng0VhOkNVj4UJqf6i+2LL5NiX
oGpCp7iVoyVtQO+5h17nmKU0RyxRnLPna1lRJPZkGwCw7WrZOW7NlBVWQxQWvPNWR2+0s1zZUbRt
v5aIJZi+sFmwDjxgSTbTaglBCvJK/BX5P8PsciuVIv45sBcsglssIg88Q9wRXcT4+HYgXXTPu3ZE
U3GS+DT0CJsxLS1LQPvjfBwJ+9gsQBsQqRREpJGtQAAkP0+d2Ef1LKqovcr7mHl/k0b87XogpsaW
IB1RRMKfQ1icjGv5apYUjc3b9pN/1KBOo5MoridsQb6Jds49gfxokrbBKFHImpPpwrM6gWg7mHjE
yjcagmzS82FBcwSuai/poq7pO1M3IhQBcxcGD8o5JYIo+iEZiKTo72z5LxHoGL/0LPdaEA/Jno2a
TY358g+XKuVvi+lOmp/cCx4l4Z1S8H5NOKm/W0GDuqxM/GSJJsjGDJfZ1CqB2Q3U0EZht69pbV+v
I/i+IfwIfBLU4vhlEoxwMajjahmkQQZ7eKS/FZylj4y3uObs592GCD+bAz/80rGGJqgXnzHj0O3Q
0QH7nTT5jVp9c3FgJ/YmjLUxvXO3MlWkgyXbwYQwzGHyGG7B4lskHBq/0bGd4tI7On+11NEQ+eJ5
mW07XWil3alRoozqpw8zzYOVLznoJiKTqxkt8MX2dWG9cdVI1j1eb3ZZFhZ8MKpqRwWMGh9dEvEt
/ZGnv+XR5qfl04j3QstnuhX/MYQ9RoaSElDM5CMavxkXP30gKM9UpkikDO99BxBkJVdg2eHsyQ8O
0LMENwOMjEtxawHxEsaZccr+UO9zIXFDIkiPZP1rGd/cS1ADZZXFYiXXToIhz7BxKoaibyz25X1i
o7x3mCIevCTn6Ye8WMuIxAMVPhTdD5oo5D47wEXrRzpv6hVQZgZXOESi2FlhLUeiDQuBc3uFbjlc
7kLjpk3eceDQ5IlSJ3HiVkSzlDZ6+r3mLYSkJPK91y0OX/+BU6qzBUid5rDymhQxSjxgdHzKQlAs
3GR1isS/YI3nVLw/Dsue3wRi4W9muNMkL5IRG70p0QwLaXYGMMEvsKGxIdq1u6i5UdVlBVEjEYvj
QpYU3Km3pXSuY3udTyzrMmPxXhDXkWX73rF6dJT8KnOaunqzfC37KV8zBs0DfuiwOPcLsqfjGxT/
koGlTvliYk4jXgZXlMBSqI1m/1jNzaJ6kKYMlGCCDzLFhUoRr128WL0rmjLLnYOpYF9tk+QhnMqU
mqG7mz6bzKQ/w4DChM/tuAntFFKwVEfnwmxgn8e+IN+KYpG46s1eIPPM6JXzi1MIVaqqn+VfiBsV
gY8R0CHtPqntzgnrfbfD2ZuPsx0NcPpBiJglqeOiNITK7+eUw4M1RlbztS7Vm4CwTf1fnY83N1m6
1rDqxUAOykZSF8vPeXn7QbfEBpxViPBOMvDiAzPoSYYSrmhSJZw5DEmLDtDu3FJTTqc24loHHbPG
nDgKx4us5Sz0X/DWVwpXrkzo+YO+u0Tmij11VY5sE4s6HCllSWceotVe2MX56WlOTJU1MeNs2sAu
+sZdASIkysHutyPrPbrreHl83M7v6+qEP7K3xHRgZlzbTu0kERtP8H4k9p4ZnGvHO9GlBTwwraDy
24ppHJ1ui0nEtPsJY/58PKJVBDabX7N6KHwKmWhdrtFU/1YDmgdwe8xtHJpiIG2jxntrSOU+2hOH
cLj+2PJtlQ1/mnzJLYsylfZQxvVp23f4wmVkC/lkvINmvsdCY9lrVSSfppRDqWejr6Qb92EC63UM
NXApmA9+DNAuIc1nlTwrB+ZFRGF9lk9ZftqHH+p1Bwl16PMw3HT/9AZ35ZpPQwF3p4MGXHHdbcdu
0SIC5TvN91EZimD6c7QYLgthSZIhDks2UZ3axKnVkzX7h/NVEF7N6mq+3ikSjFcBA7gt3Az66TI4
krDezRU1oK1y34mqhzlpVdzLYg9xEPx3vs68UTj/HP6v1fIBPFGj+MZe8sUt0TolHxu6UOPgPBZW
hgPpdBdlL8Fik8/jqMKBohu7TvOeKSuGNAiKW9KoN90zixXUxD5vhQhX4GjH2i151DLjmWWrrwxt
FM2a5P/iW77B2ujBtiU/iGiAVhANRf17h7zEk9Fi1HAcV262u6CSz59gFqZgXEDJDywwABC08M9y
hkJCBmdT5seCc2aHff4eXVUBczHFExLGTbuDpXpILnt04ddOLqpugnjP3bYyK86s4l7jfhynQhtb
yb/JK5yAZCA/7OwY0epDdIzyJOiQfMzzGfQDWhg4QdZl471Whk9mMNzXXrOiHkThyeKLgNDhwNax
qjjV9MSR/iEdAQtahgwSkZtTKUll7a6pk5PQQeJBI8drauKwuFeqP1WCI/NxSfXcj/CfDtosF7F1
D9clEBCDU90ujUEpfM4CJN///sTE2obmVi25dTWQpQjIrpEpZG9319hnSSsPu7PLmZGm4RrbloME
HRnr+pcUuqmjDm29yqVHJuJtrBMjUnh7ilYSoP7dOMychOFAC94EBvL4DfYroVq5zYRNdIHAb7C5
4wto8EfYw2YYcLVFrz6tvpGQQhhiRpTOuma6Hf50gQIlvfEJMK8NlcpukZauOT2uqj40qgMAx2rB
eZbD+UX6rHQoXpxGp2nBkIhgAaeBXV2+GIfWsOhorSanLmOaL4MqniCaebdwE6DZzO2nF7KhVjdG
+XUo8trZSf5XGpDgALJGRZEc8P6VuOjeiVc36BhnD5/OaFgUgCTRGiRt4bFSttmAkWXmi8gys88f
MEGUFy7UQ4GkunN5Oo1pHrhhvHoSgCsF8LI6KcEmCurcoYDJ7uLZv7mxXycP7ZXFUIs+1+Jeid0y
SlzGdXd7o7oBtfxmkMgvkwseBLCft/oKyweSBKkq25LhfXuqhUv1MFwyQav+8WXtuitfWPrIkn0c
Xfgn+DzNdc7ZKlyyCXcCvuNuSh9Hsoz8Fi5qKHlXLCwmvMxRBCDd5kTIEa/25SK0uoYzrfbe9ItY
5dq9zoEqRf9CaPPcRFrBpVkEisRKVM/7GIadXkxKhlbJZG3vXQwrZxB7dGqhCaArO9VpKejErPBK
wW3SBcvK5DBLNqSrmD2P7R1fepWpgI4o0LiXwQPVdulu38+6njfPrNMxVZPHKq0n2fGpsw/dRgcu
zPmKk5bMFQV9YGzCWfobwlPmTTV79e/+up1gjoxyNf0PXbz+CMcy6gK29YD8gRFea8f3H96EzcSI
86w3XdU3Xd5xbMVUqlRnVDEdJ5/h11kVvJX9zpAsOKOGVo0ja5sF/Z/zqA8N2+PL8lQfadhl21aE
EXUsW/ZCta0z8Zg1APen0+u6waV08OPh0/LPpZ8lZiW4uR2rAgvjuwDhLDLa62BRTKaxNePwK7+G
vu9UPPuE9hx+DvbNTnIrGEyYZv1hVszM4hKXEdWZg9D0aTnacRov2gP7rQ1bqfFQDKfIAQhyHl6P
urzh/kKe7DgonMDrDV3LShdlfkI9S7zvN6OYXCmFbutfWng5qW7PXb5pUYEWsObORwwuEx06lj5D
rhg7ds+a8OXxEOZKk+zEyVxdUz60fggbOu6aGmsR6BEdg1khGIE9/grLBY4qpg53lvrzO4bVMHcW
0c7N9DPCQccEzXSyiFpetU8GAvi3767gD69215CUPzc6Xb4SEWN4opgFsC0pLRKzNBoi5Miyr5WS
Y2uhpqcc1M6tpV3+CtL8mVb87J1Ty6qCCyR3a5I9hPX2VBRtKymK8cP4oqx32LX9+HcsOx46Zv/k
l/bPFM9A3uFTA/jKF1YNtZ4CHI/BL/M3PDNP+aB9GVfl5DpTpgjHFZxhfx0wrpFK8AaF2kKx9R3F
UijDHtxxhWSDHU+ytbauDqZaDPyNrriYMPeQVEmSLMLQPJBuh19DcFeP+B4jDbVClTN3u/pgmMJS
fRaxmGORPY6dWrZlQ+tRmEdH9Oi7EZrpU9BRTlTgsfRlMLJCSqcpcmj0q5BonoGD0+07pjBD9NAb
Km1Sw8ZGX6sPZsTLnMNGnPstSJGUoU3afClmfOXOiWOEu5uL1lJJkkI9Hfmm0Z+EIYAbTu8A1Z/6
Znbb+d3mOlNI4qkhzZDnJ827zVI1rcBxMsRJAsQZxY5AO0CYiUnMXNwPaXnJzjCmgxM7HcHN04IL
fTGRBHafOC2lWikaXoVDCo0s+gUCxJ3GxcV54YMFPUwowy1PXD3hrHr1otX3wAr1Q2/mgr/zf8qW
d5MIRc37FP0EkFpJFBgR9VZh/apxl/uaNgmhMCB6E79mtLvXtM0jbasmy3JIA+7ilFObIQnJrqq7
TkTlBD51EENLXTl5UC4dsFYZPkGrzmrTIzu9KuKA64oIg0bAKPbOVoaI/I52mmr4a8ZMGJw78GDW
M4VCQc4X5oXUNDCsrHtxU5SystkdjR94DL6DY1GXZGXBr0vF8JE1TbXhEakd9JYcIVMmZolJZzKd
5iAGKwdaocEGYIuvaiwn1bvhUResmqw+14Vu3gkuv1ulRXfn2o/EZDtOby46Cc5pBwcYS4iPSjMd
ZpHRjJIKfveeYryR11J20D8YC69ODNFQ3U/R2RBj9WygAQdCyNagoMnM6G2wOOTfJtWV8tCRxxE1
owki9MGnz3e4Q61Ozroqqv8bDjv0jThtSP4/y3qmyPOM8tB/mmYNCIWC4k2w4hufbRsln+AYg2nl
emvDxYDp4lmZxJleGIB0H9xU1oKVkpsHT+xIv2At3FpUzYSe4pYsFmfQ9paI6DaLPeKaFd3xJWGS
GoRzt3uGt91hV886HJCPkNP+DZHrfa8KxBT4QwQhjscR4Ew1F3c2wxu96geGz6eW6oK3hKaiESpl
HUsODaOAbxPbcJ504Z3EFLcWeFn+5+CIVkxjBmv90pC4ADJJixYL/nQHjz627zcrijKe7ul5V+ks
oXFE0+yZW0qAck94tOpEKUFP5QNFo5GAIrPTZw32AhhV9/TVB0/rX6KzIPFvT7CM+kfdl8KOIqhL
N2Cg9ygPwA6q/2xI0uIQ5/p+SeU18AuaUe9OAEPvzwQ7GP4F96saVRbN3WkyEG77Gm0y6qu92d6c
wVPA2kZphTDUT4y9Tb6WI9bPtAdT0lwefFD0tgwr1rz1SoiyzT18wxqh+X06fDqrS2kTY27yNB7W
Sex59WgoxUx7QO4Fwmjnnf02Zc9BCAGc8Ll9GA4BaLmH/5yzOA8kvnGEd+k3j73SFQTDgQpGuFtI
YTsv3/S752LqbtJHFYr3PZOpy5VbLV+hoOmO4mnPJJOXKs5rm97mGpBvi/c60PCJPm5XEd3iFd1x
wJCPMZ/cIlWSYb2OuUP9UVN57k4tRK4J9FqENWQZUV6sFv11DdnXRq7yNveZOXtWj+hIBVUH3dtv
+sK9VXvLrO1Xrs1nQDfd4WVpyjjb7RHRxUs+JGegdeDc7wGvRZKXWFxGJgRFXvhh6aJoue/tU3zv
lRMJDn65KWFv0RxBxm2FyB1NTsiUdnbp3ecOLJfCErCWwRt/CGuGYqBmliFNN8UZg7hrUpHjGcus
GspxKT00GzFBBt0xAtzwjUfQOrN2voeRyy/+Wl/Pc8qEGErJHHm+BqbZ2JXNhDxKgXo6chR2Yw2Q
UU4Q/ly4603oF80FPPSCA/Okm6QWvje2DaUCXJ7B/CZeRQjFmU/7AAs26Cy4NOYICHkntor+vcQn
NbSIAWuAwRdYcoDdAYxUxGBt0ay6GEYha0qw4d1XjmfUegU5f1ycReruHcurW7aOqBpX2sbu98rE
j3NiHBmB/jYIUB6KnQxlqW2Dvd/goK58YReSeObLDIV49LK2JpHUeHK5eaA2U5FvLHM3CtbLPgLU
Mn/qDF++G53f/tjTQfzlITqV/2VKhncwv0Scr+JEas45Tk97M/kv3rWqDuzTXIdspvL5CMsHmiYI
QV4NSlpSnNirI5Bk1XX/qllthD7mZPZ5JShWYlETx5aOHBp9szG0B3MONhjVN+nHC9jA423u9Lks
p3TLu5PAUQxDYkaHQ4sc4GcFGxSM5KvmF9bod3SZfCDfZJCuVFJu9UsTmPvloA3E5DSqTBq73m5b
4rLwqfCcbqCqSFLDYlALZvNed2ImtByN4l5cbdHM9h0MrWNn38zj2aeb2FM4qZ/RTXIa7hOcJLcK
D4x1tu3nLX2X432wA2/8jRr7a5NfC6zdZSZUG1ed3YFOWUPPPBVpaE8zpKYUYrgPiaSf+gSPv8gk
ATREOP9491gB5Qnuuy5eWj8n2KrXxwGy9k8g7v2ffywZcwjcebmpsmpe592AMJqxFajLrtws11EP
opp4r3E34bpSWbIPWsQns+sC13+gSvN/Qc3B2PDUHBO/YqHeSZBUXte1lden+1zkess49zGWsDn6
kVayJgzAOd0yDBHnJK3y7p1Qaj6yJNFghYYDXMT3CHk1UD28e+vHa25xbd4IJFRMiqxWNqbQBb9y
u+1BhvCmFQ3x6vjCW5zANb3yih9wf9agded14ZihkYtcQJWtxQs3KDAooFCTH1jZfOJ+a9bwR11z
Mw+Fv0PeNEihOrBMF9Tpn2MQMI3KsfKdKU9c71YCfihiVoDhdL9s7hczhMl6uzyGbbSivvmYJMKY
1tbu9yGzBOjtpnpUKmFqbKloHJkoreCbMFKTHIoEU1hsVHqntuOiNzU+PkHQt0tPVAvLNTvCjUON
woNnsrQGQUj3gNZQnZZesOwMp0GbxaSg1gi+ydHRP395Ie++c7vs/Uu9ztUCDVir+7xdgtrjcHps
WUDd0nmkYjBUKTtALQrhwBxw+TPbcgN94MlpnzjFydhmINarhgf6m7P3+tSdm1gAVUPMXqRuWIhb
h6FjZq89mr3TqqNNtlT8DTKr6YhobtvoKCK9eAtCIAzWmS7UclLobgbMExt4eJe9OP7XRJLArU9I
8Q5Lin3k4KICJzMkYWwfvuKKEUga2WUKpLeixlVfy7pl5GZ0Obenl+t3lcSGd4CyIDkLveNyAGva
3/TkkpXVPH1ama7V24EuEjPd5V3Dkj4DhwoXodK/xG0/quEwrcbpdc+u1/jsdk1CdprcffS1w//l
+h0Ku7kC3OWOMCTNmVFkODGiXfXZRcTERaFO9CVORQfXZCLdQbs3nCYU9TKzel6ZS5aRZ0JTyt+9
nxphSQDB9y20Rh+KYAGMr1fXDQUULxWk1Ol1heIhhky0KcD6ZIdS/6EpVMtt4NdJCMHzczsMADa2
AA9tMyCdLXevt+Tjr+D2tNFMndXfVXZm/BocZ027xfcbwNq3NGnQWcvSQxAdNtnqDEkcft2dVQcA
Pb0mzMemigydqZY7hUT3VCjFcF+ogcJBlWPhMTEF61rPA5GHXk4Yt3C5DZazn1Ef5d3ZwaRkXP8q
Kmn+5mHyBizEeGRoF3xyOOmgFy3POAE3+DhPqW0LG91rEHMYLvg+D2wbCKTMbMH730dgomn8L2fz
4Hr/g1pvbVx1OdVH9ayWoUZ0pfBeV4bEBy9P5ERCsnu49t2fKQVjNXi4+jamZvz4N5ymnciIPCCO
i7wbubseI57atAzzHIc559Ec+NB2VG70gVySpNsqzJzhKcA+8y9dMriSRGVNbNeu209b4jNS5Rh6
LAzgwctBFkdsk5Ufosqm+Vy6fKRvOVGPf13w3T72rrJlrL3ySc6WYkF1VMrTd2Qv+GSlonRIhA08
H9tgPGQJ9chsr8AiOM3QxKinPXY+LBP5ADlyG3IVP+potykXLvEHGmYA4wKn8rNtKow19wq3GUw0
mDIOXHwHzoOIQJLmzltbVg7gd0OZ3Oks8JmyCBLI3RaEUAEgHXGu2iacxSkFzVJwwioG7P/kndMd
CxopdhhHmeo3KoZrjqaHLlR7IQ2rEjD1aPwMmBJsn6zSkzK6XgY3g+g9IMG9dbmF8GInH8fiNfhL
EHtcU5uVX9+R4HpuQfVn0yW4HJqlW6ijc9xVPJOQVgNd7kLAsWxjezggIXt7r7cvfEBLJi+Yqz4X
3SvIOYpxvinU6zgtDGx/eSAq4JTkdAjGS+0TFuddfPxQQlRIrTqRKq5cZ0uV4zE03f3OenNU4+xD
NaDdIvPNU44521FJeNBu8qJ8JYkEc4rzP4aAq1WCV3h0rlBszhBR+YFvMpih/t20PlMT5aonTCxw
R0qIql4w67wdskSgYNCK4gzFdRlzCsMD1VN38i0w9AK+rejQgX+cPLIIXgLb1DuWeDEin9wtREWW
peQ5jdX0DIUDzM0yGBqrq5B+fqZqpsn654emZCa49cWshKl8aS8+8T13jwjCroVKPc33vdqW2mSX
91mrjvIpvydZEt1O6xEAhfzLHqyqGDyUMnQPH90FKthJ5BXkYXfku0dy+9sl6IfROmssEWh6dS7h
PuassIqN5BWogne7NKWAV2o8ncYT6mw+b0OSe6gHxeu/Cng0ibu1qrZ99NMn93Dm95yr1/KKJA0R
FJJ4+faRyYVhQhmx1PK8X4UtzzZYyJKsDe9FM8u2+hA3kHCFVKDmVv+B4jU8r6Md7cLveK7ttFC9
XJncm+5q9cqyFMq2qz/GLxCXevhIIH4n9TnXkNscanTqVAHGNMDp+LiFUW8dFRAnZ6amDMjmKsMa
WxKXaR8JfsPaf3KYQSHkmnvlmYE2Pbk6eqXrdybT/MClTGDQ62kga3cd8uLOOVVCdCMaTS3BXwHz
brtgecOeMR26vFQjzqw85mu4cAuI4PBgR2bkfRkeX06/FLcu40aaZHT5kzUKOsmA0t5uaMereUhd
oSvYHX5MyhmQaLKKmjlHBm908AQ+YsYXZitEVeWBSdFTSFOgHZI69rR9MJT5EfDIg/0t0ff8iOMJ
qpZCn2WvvQOh8JozICvuCBgJ13v0XnuWZrlPG/ojsW6IDMYn/SDTsW2s/2AqZIX4hA7L0P4UprUn
uvfj4KaGqyD8jp6wqisGdkNZ965qLZr++oALjcVbD7K11/90OlbdQLoUJqjGpO33gKz54YGplpBm
jSqwlxi98+VurjZfUqz3xMsyDv1cP7jLDkWULwUWAgq/Xp6zGJeSJ7j0/5P6/8vcQYc30D1nv9GJ
0n/+/h4yjLmqPeSQDjjEDtGA5EIfgOqB1lu2eJ54cXV0DFmUjNd9LEhU1MJnOH4xNDDzljg52k6i
wPMEn210rzvqo5AyMgl/ZV07QYOhpHG0mFjPRHYS75ZROfkeiayPJcdLhH0YLnAxsZaorbXptCT9
9vq2bEjdzCBPvZzV0xLnH5eRIcAmKNsVPiQ38zfk/nMbA7SMwXjo5YoN84cFOxeR8D5TkBFv6dxl
IBBFEBvLz8GKzVE96JsRvAonh57QoBO0k6TZn/mDs3dAzowaWwxnqV9uiKzxgIvMFjcgr5iWCr+v
OH1D3lLPk588b7KWTDW12Gd/MH9nugMOljgbO89zUODbE857j7ezWSRJraEKFe3oLYW0H9uYU56b
dtbfA48OSFYFUCGU3GO8RlGngGt6DTTOKki0jv3kMHotg/1b1MNVTW5H8rQD4mH3MsHGRewiy2vb
FqnL7lsosgYGp5dQPgh0IcJWqabiTBq44PwIOSoBKQ8lvI7FXhtO4qyZGpwLWL7nemL3es28ovrZ
vnvZ59jh9fnSw+e1q1iqF08MedSmWcC7ylCeIWqOxeCozMa6QeQKjx0kI+rMh1VsmGKToIuLQBQx
PPbN6FfKstdNA4y6N3qq0ahKjo7G1rjlMxD48UWA/TFdFAvPXjuzR5YEa7rNLv7Kz2aaJ0Iht68C
SXwifuess0FsxQPdJPDHqgdC4h/a+WofeWxVUl+YxFS7oZapVjX4MEbZdy7t9IXnETXZZnpFA/jg
mP9O/Z4sTTNmNuAmmi51T8+9RpgvPT+2lzta+XerjmevaB6ktNebyVaHadtkLPH0VnUjj8n+FJTR
8chWwipEp+0c4VVhgj5MtFkCGmDA0DGaSFYEbi0rgihb8SbzQwZEptVk9Oay3EttLwlVPxHWLDiI
aGYPQ/oLQB82RhcXu1woh2sbo9QfDIvteQBE4sEEEncZUumCzBMKYzbvK5A1eRmLjsOJTzQvlsmL
2KGDeH/57SbuAgYCPA2JjKL+5hjE81zr8bHZ9xjTcOcC3WY1JBuJsNWU6UxRG7pavv4QWvAuubn8
vF0uMkILgu+lVwinrb7JgdlRFvHLBw9DHJnC+V6F6k97k3mP0czYGsB/8mrzOHKygm/Vf8oR02yd
CXuSLSKCAi2I5TigR8J6az5wwzwbsKfP1m4SUc6cGFbB5UdGYiF9LDulc/H8V4lCOv0FRbm7hyNd
v1e0EGo5gwvYGbvc9Jungkhis+oZG8dFySfCdCl56Yd3ARgcEW1/C+E7hcFys69fliiol21KqtPk
eXrVJdnYhHfJEEl0PcK7rFhV+uPU3C/aXKMW8ycj3SXaCaUhqVOubOsMFMC/KEnszGYcvNWBqhmH
G9E7nGP13OGyFh6h2/DtjUlRn+K6vTO0qGanw7Kwyk2NFXvSN28ZBPWiVSfJ98Nxi1Y+6pw2EJQo
7HmHAUGKutfPScQHzr9QNewnwem6LROBFt1f0BARs8lxCPxN0RmrxzEw81lB0Yyil0NGKqLfRwGL
6/n0FAQnYgBM5GktyqoZD6Xu5ULAg77eEXR3K3Du2Uii+hfJ3aXf2KpzCwDppaWpFq62Cm7eWeYR
7+kWqzOr08xN8A1kQdZauzvYHLA1OZOuC4YgADXufGMpWm1IMGxHDc3RTPO0oh8N+Ww1BKcy9Hto
ulykDs5svu4ASNsrbrIoHzBY5Tyv/k+202zQKf93Gm4msRugs8xU+dkhQnaoK6MuqQfXodZcsdII
jCSfRaUWUKUg/71fSGrpWn3sp6vT3561DIxjhclhed9ASDGNbLkkpDTMz9tKy0DSIKsLaT3WPByP
FNOoEMzZ/sPFaNdw0lAJ7I6t+hNKoRkjRra9+blyglj1VFAWumQWOsG27kFFPD6mLroeeRvJg6Lw
IqFxwtWD/mJ7rogpvwPftlnH5fY0QR6ZHImPIheh2a0GgyP0kIzvlqtgvqyLH0I3NvQW7q1cYLry
CUZvlEWiFo66va8vdDL8QKYwTMI/bceczqrsHr3ivo2BCHVSdXTrHfduCdecssdWjIYRz6CePoPT
nXlX3OLlrdABN00ICB1u8dZISuajNat7hA5VxyELvT+nZpL4fYrYz5nRkX3tPMybt9jXD9+DkAcD
qSZYLPpP+CkTvtMyK6yQ2QsqhhzaSJgZ6vXLojCp6ry+8Me2mcFr7fEiAmzqtAz6WvOifIhzChaX
5CEqXvNT/F3LVYm29ZqXo0SuxtSTICNfxb6Z4K84s9NxsbY0crp6mineJvalnow0L30s9FpGAfp+
5hNv6kJUD6MJ3zTScM7WFeXuRoIY1INmw90y8IV+azgP2/jN5P9P28p3/qisNLggSR1P/H84Rnco
m/eE4uc/83IzynTmgh+dhuPVE2qSReUrJia9xKfu/YmRux/oUotmA9llR5746uE84crCgZwUF0iY
ImEeil8AoumUtslqom4YWTaao2xt3iA+qb7oGrdI6fOLNc3QtEc8B5xWCJ+inZ1l4+FLBYb4pUiL
wzH9sWvZHloMtVEXOLMaeb0qhBl8czfZKUgTF8JOm+L2R/DBkuyeqY0tfbAYcizc6Z2qepa1k+rE
ODES4d+vhe0dzfCv0Ga3X7ZE7rdnps65VZrU5DNTy5HHJ8lQrywIdkQYt0qh18fhzagt6bs7SUmI
hiBkIlIg9wV9VrrsgLzsflkjXmO4HD7Hh9Lt/Zqhv34NrlQrDkYxAWtQQFx4kDpGnMaE3YKpXFiT
lm7p6/xzhorY7GsSHETzITaQpgPNiaz6QHDrIX5gi/zEnQGOpgCDg5asYGI5f/Ug4mbBxMexrBgw
AswN7qLZJJD63TIisW3gj6kD9W4z4xC2Y7QFfa+UIKXa6VtwkxMOuDrwU4EO3UfL13vzyM3HR2Mc
eui2y9wVotVsKfvrRlg20AWeQP8nMrBjfYXdbWPPMlBUp6f7jnouV3rIkdA0VUzJGqxc/1fwZ/D6
FEFQ7Kr/LFb+lV9/jylDehIDtVp1vx71IX8bvq4+nKS1zneyMcXJmJNAy+d1RM9lZgqNTPHpMRkC
kd0oG5TTBlngv1YiZfDmsFL4RFKKk361ZQLzfxHcfEjNHaAL0S8I8jra0GoSzUvpfsY7nxrYW64+
hw1RSP+s3ureHt/mslAeMn9xz0eaYk/SbuIqYTXsJkJFgtUYl7miwHteyrkrZXmcTr2zptm2VuH9
1tk2ZVZxFQEsE4KABq50NQYQQCxO/FvXxVCZkCxHo2yQ3GE3p4VXePJo6Ibj4D+YSwfrvvMZ9OlY
YBrOnkAm5hMEODqKqOY2iHDqwsb5mCHxdHbO+/SrV/HrVuomes/aaw0bVMHxHQ6FxwBzPypSimbt
UpPnnJ1Nry5p9CFPb/ZljimZhwa+mOQfX/Au1pQXckxQ0qUHklnDUHGd4xOI3HFyEaeiun/6WE3L
SZFljugUqo9h6rEA40gpDrmukrBIsFDoqMp3q/rvsmJV8i8WY7zvbO+4VR9k0mNOYII0NmQpv4uQ
E8BuHaOr4UYXLgbEZcepmulFEH9Hpi7bIEZ5C1XDuKzRrN3EiW+Cxd8LO7MFxe+/AmfYE9mWEpo4
q+tFnpHeTUcSyft5EIt273BAXLZHuQUwDbRTEa+tDn4vza16OiQIkiegt3RNbcCRE97u+4MX6cL3
KasqINNG01YYDhi5oMe2Iswi+pcUZtrSHK02Yd18uzFYBS8igomvgDcxcJ7O1N/nrosRxj627ACm
NiaX03EziFo3anCYlSRDd+qmn82gNW7ThaTQcqRMCkL2ymA5JUjDs4I4VgsOTV/oNFXAwrrmY8Rw
Rv9aGFQTYyaCAKZMsZW6EiAJrK3xXFl4+6oSjlMCXwo0TnroKu1QM0hsfJSnDsvbpftMqgdVt3hd
96n3OJ9n6zUQH7pX63M1mzQlFHwbB9aVV4Us5z5L2UoJeQGAJX6TmlqtiyKw0kf6lq5DtJDGqCtC
tgAY5HLUw1qTA72mDykO8IvC650sKvqovC5oWmvinWJmDy97lbHV1g7BIdOcepSEF/wzsloyNXIC
3ecTKv9cx3kcCYm0WSi2G0m40qudVQdgVRX/OVLRy5oD0XAPatMhi9X3CNsGSTEN/72XA/bL2sHC
BLsrLJeGtP88caYDvSBZeb48vUVwAEOjCqyWWWNAlVoPBrFz9pPg4LgH8DoXaFHmWS8k8F18hhBw
dRL0wKKJP1mgv6c0LakPHtfmuyFGY06wu5ZFTtdB0KneJyX7PS8cnWXBm4mGOe/desk7nHJNzUsX
rwPdjT0RYFjcFuvwRPavp7u6KiXh/mdmYeYbuZVlTErwaB7esI8Qg3zC6/pkzwMAn5JMnpSCj/Wq
ZQ3Mr0F0A2l9hM52hq3X1h+FqMut9GHoQxV8KNMIQ6UOZagPI5o1ZXrIQ5M0sRnsfbzvuPV3fGKB
nC+jm9KNLVLRpFa8fMU1vfRX82+UCAiVpleSvMBgSo+Xyg54rQ7q+lTLM0HpG9g574oDJVBADSYb
sSmxGXt9T1Dr7dvFCR7eio85F7pmaYkzEHdAzFgilq2XKVa4kSk9WfTSIP9mp/zPDQ9I71z7LFiB
xsrB7wzBn6C9ONe4OGkIFKuw8nUJUIewa4w9hQaG3qKSmnhU9RVU+WfmvwKElCv87UIm5X9EHF4N
7OZxadYdx701dNg5eUgp48eerm/xaAlLXuuQKJ8Fb8t+3yZfotCDVXQzbN49tzSzGsfjdlYEKtCo
qU8XlofKWi0WncPEz9YeWu1rn1ws5RcfXyTt69qZNiZyyEHlJeuehKNuEEscAAtSE0gBxsL5V26u
MBBhRV7xEJkpYWuBKsXo3HKFDk2JwigkjLwQcgp29eYunCFrGR/3DiUWmRlSdPu4Vr2wYc8QsDo5
ghKDc6tDq+2W1DmT6IhYPXrFjYeEhqqGz5DcbZ6nuMh5vUa+t7osf8E09yMvNn2hrQUWz5xM0QXH
2X7MDGUfBIEJf8YZLWeQ6c5GuXl9enustDaHIVUQOUfBN2dEILiQiz9mrDuOXAvVxjV8bOX7t5/c
Q2fa6LBq/MGMW+thhkdoawv874LCeTa4drGLDTe953d56fcEpDkUtHYptAi1HP6/t/P53WgCqdCs
SWUMvrFk0+khLXJpfReNl9PKjDAyFStfbPmAy8ZFmeZZEm4MeMQr+jREALqNdHf1QyDnLSy+eZ6L
L/1LEVoLH7esKp3DRettYRTOsBuTnyjZp24H6qKXYwpmsOQyBX5mQkZLfMOGqgw2U3mHSXQggY9e
dxVzXio+n3DOKmMVL3PF8uNkjxZLg6lVbUHOdN7jccL868jDrkp4YyYn5kYKPk4Y1NkaWgnf84f5
pGT5TlZoQJkZey2heSf68H1apM0McdoXyAdYAWdn3GBnyisQCjf/OwQbCamduxhM0oGm6ZpQIp9l
m+farDPLaCWQCBZzCFYtmimKqFer/YJQEZOYGkj652dnZ7ga3W91aZN7vNriZL5bkiUUK8AtfAKx
XjOJq9b16os3CuWE8uLWPFawFlOQ6KO35QkOLPvK/UcZ8pINU1kLFA1JtlfU/IzyFVgsy7wzdCJq
Z33xsplQnKGV9BdZbF5FH9plLpNiHDivje5t6YyKLabI2OQNWGS5IiiPnsgHzMHInsNrSnO/L0y/
Le940TzvDxlhHGXN1p8fNgPQBlgdm2O47vdBML8BbZgxd2dYM6AnWhvq1aE5s9/5yyNjPinEyZ4s
Ul73caL5OD8ywMvdDmf6hmdu1SIMnzAEg8nhneCkO2CHIjrQW3Dsm0m+abUewrgiQV+RSE0U9zdb
KwJ4fegaS4fxa+UW+XCdCiBkvAFJS6b4ab6DSGeJfNZb+ORkwkMkZzz0RXhifh1tJM+2DmNv6kTp
QjG1cnj4oxlhk8TCrWTDjdDuPYzDu3QqtYGizv5WRjmMeUrxcmyQCf9TYJ/k1gzuTqq/z1yVAL+8
EUioh77z4kKuTH+OMthGutAHIipvQguxuSxuopnoaxclhobME3oEctbUHVoSoeCRtgo3UT2UOHDP
N3XyIs/E91bd/4Ebwjlwer+ICa58zWgi+bZdrqDCpq4L0i/jLmD4twrssI+nue+12tAShVPcz4+R
Om3G0rzFdJV2a+KffljtHbCfFKlm0nMRDiHNdTlDgQB7UF6KDmC2td1KAcHknG/dta8D3cC0rdrH
9SW0qLllhns7QVwzuQVDUZfCHEXBHKIc/EWWavBK4547NK/AIlFiJ4wIllXtdmbiDTAaFjH4HSyR
J3ljOXvVF24a7K4L/uTAiBAWbxlwQbVLmqKS2mM5aTWL9sxuV7pd1d1tXuUoCzzbERv0on6q6T8V
PN3FpnvWJuDbrvixeAR8hR2Pnz8xH/9A4cCbzw7DHcDRBFsL60RQUS2k4clomc2WxSEr+gY5UMSj
jXIVsCIiEhN5iWRfhgo8JC4QFijfCuE1Zv4TxttjuHn3dsjzdyTF0RVAjI5FHuqVmvuMNxYmfVo0
WiLOU8lM1nxkKL8h+9w6l7gnMlOJLqccFY+jmRh+ErjkCzuu1rLiZG+py4nDgKDoJi9v7J7DamDO
ME8xUoPYhCiCjbWHd8eZqpfBkOXh2OsrsTsDr6LQ8n78WfA+JuSNXsYFd7eX7ux+/BQ0exim/9y7
/jfXgAa6nxBi7VY94dYVhcFwWAX/3qZEwlCnBtZ3blO7zFcC0xvjuVJ2O4nwyRdDxHL6L5/lotsv
OqZJUDk/33CBf10feAOjQzdA3C7W8Pc37tFVK02N5DYNr3YhK/6pDy2gBKn9Bdxcobfb5xdFmBq0
x8qzgLopUdR+5NeE4LUIeqEfL2cnRu6i/gWapOE3IhyqlC5FN9zWtZ5M3OGxx3Wk+SJV6S0fuS3q
svxL7+P18uAMiBQQdJ1IVEEYhn5EkjuHQKnQLROFn7jzXZN7ATdYI7p3SRtgfcynaMRyCIsbvR29
t+5PX3TD22NBp2cxilO6ZEfWuO+CCmIfva8STWBSRZbWg7zB0qVEQgTbIeIO9H4ZE0tRV8COYxuc
gB+HkZjIwlcwU53UGs2jbNgmL4R8AcGehXesAZF48oy5aGQ1RofUyZeAsVA4ux+bqTzag79jXJ9w
xZQck0W5+yHRBAt8NtiOy1vBjHKvYS/d2M/AqpYscNzGn163P3hiX2BFUNBBEFxfJ4KW3OB/+Ky/
eDs6v6W/a6DZNMg99OTGIC5CfHR+wHVi++q+hrmEbATSLSEO2BL4OLOfCHpEnKUXVApFa65J0ixQ
LUcnO47qzipRrOVdXfsIYU8sBWkUE13SI04mwmodmmnMn7VKi5+dZuxa/RNl3lqXJDgUn2I3XhJ7
oRFRbuwzvqaTvncjeEJRyVjm6FV5NdFO8C9PDSYLRjWm8wRjIehdT8SQrpjt557RiSa0K8/bTd7f
yECs6OSKOGITTrjpA7PUvjQ05hFqwtHDBhF0ZwwIj8TtwcGt8F4TAsmT3M7PxgBR7DnrQbnlqTcF
KlNLshOSYUXDS2JUrwtigqCQoNosjjFkr12Iriqi72El8vD3/5mFgg8bJouf7bcdXeTeY6rrjwRo
D0HppBs+9NSx/7JE0r9WtqdF343lQsYuLG+01RCZnBbosUr9Mkx73UW4Q2957D94vX+GFT7A4yIU
yBDrtug2j2cIUL8JK8SPs/iuH1FNNg8nHOy3JqkV1S5kue8h0oqkW7IHKo+PtpdfRdFgaSqPjzXJ
Xf8gPrpvekvQ0JuFtSMBA3zPCLwDJkI4JPQn3TDLQ0HDP/CyStSB668Ro/hiJaylnBL0wScb8sdE
cp7cTozNbd+nFIP1/s06KQz0AqgdaEuyf318oRTaAk32gMdR84iUzgCy6Li80aLpOV/ZLGt31zKJ
G2WekavrULUDitstfXsWmefcv2aNqYO18N9rncMfE6w9p+VMvZOd5idbOhD4osK8lt06MHCTAkmA
JH/q5vXxnR51+gp+fiPYq7KSTu4QtAuVPVWEEuuzdov3AFBlwkF0u11oElyEF9h5BwgQ2QFJ4K8E
DiT9H/rsaMsmzyuD1HJIXXgHspOvkMkl4RB+7TrZeg09NTasS2XhrltmCyZoNEe00GGERdZe0qqc
fxxActkj9sqgsuXyYekDIwcHx/uRjeFvy6fccmY01RmQrL+nC9dPsg1PoOwadZ620iCTG+wtGtUL
ZuXKPK2bA14uWjzF3Q0ZjOZdln95mm0R3s0e+yrWCqcGl6Eb5N9LkAk4+OnN/y9ym0E4ACxTW64v
uIYoEZYv8T1hbN3DrnK6lH5PUUz1+gfQCrINtMIwQ4F9XNoxi3RsMXSPWvFpXqZ0HFlvBlfuqMgM
ozwFYAOxUhEzaZlDGlcT2t2FbO0/5tXMBRZW64N85S0g6fYnfP1iJDWjYRsYyOGuZbCKbTk7aLNg
WdUp1a2LCWRs+kQ50pX8HPa/e3Bbdrg0/eCNUv4bOJ6yJMMkUPp7fiPe5PYOR31K0GP78kw8MEQL
6BfZfzICQnT//7Vj9Ocm7fZtLRHtEzlZhYPX4gJe2HfsqoIFiFtN/8mU39uV68PSZCLwd5tE/MVY
7ZPuf+PYo35WWfmYfpx2+wnSBNgFgN6MrIgoOKSymm+8+wOapqlTkdIe6zTwe5bknoPotESR0TSF
I12blbZmZ7BsZvP4v1/ghYrm5R2wwzJlg7UboFdmRjFTEunGe9DTUzfe5d4CtHnMBynfQ1lLh4cg
/2vu2t7H1aWc4ui+aW1RK/kkfk3Fi5oB20j9VK0LH8AQtERptigHgd1J4+ajcchTkDZ3QREkfts1
0vvk6CkqhWulPfS54/6KQ6B/JsUG2fh2jbXcyKR50kw8W1DdK0NIUo8uzTVhEtx1Ral6IP5DMzOS
Nx9WgxPmEAVHWdjgKQkJjdR1RCwH4huoJ1qvQyxlAwAHToIcCVpAeQQRGzDcfM9VB3s42olqHPz+
5o3xy55ADBf4r/Q9VgQ22U1KEIfK4TmNz15v/sl3oGKC8GYVTQPGG/yYynhs4Vyuy6qpMvHdDkBZ
UJJ1XJZiB5vEWCRjDlOCz8eKXLjsLkW235mimistQnFZ6x6ufaycOfkKnKj/E58aAxIACikdFxth
KpKahwZI+/e+BVEAKl6SEapE3rMGthwEnGnLpmUw+TjaQTGFpktWsB5rnVmmx5PEmQ9Y3lR8jpQr
wBd7klUXZmr/v4a4FE6RIfR4CmkSMCcGJH2gpT0JH7mMAMdEffCIMZEh0v7B2bQ2enqC71B1SGUJ
3/SHs2zlpCVCxJQahknF/zGk0NAaIxlOJBq/rcxGg6XcHAmmUGc6rkesmVD6qmJEujPFej6/dNmA
pNve7KLH7q/orJvhxhUCC7RLHn/Ny+Z5RyKyRIFOuEGGTlCVI7HWdu/QmRidyibF+8Qfsy4lY5Fb
yuY4X0B66Z/zONFQT8uBkFI1kcWgILHYizeUi48rT/vL9MrFrAux39MGG3dUn04r0AdojXvb6N9G
jZFkeKYeA1BOzgdLUYF3Q9GvC1Wu1kJ3vSBUB1AgUV09ziQb7SsHqjj++5JQrkRlx7LeLlZzEldQ
MBYviakX6zlF/CV1pek5MLWjOqSbCEeF42da1fN9X0D6O92Sr0hJ4if0M1i0rhAsa0kpWO676rPW
PvydHGfGjiQyf5E7JbuDH/etcvBQ9uqwUrkRerY4QOSmJdOR3ldM+1LEXNPiQRbHOjpGFxTxkVLR
W4tyAbKkG6QuNx6rQ5V+0F4nfwpYtrPKaUlbJv+Yb0bXjYt6NCnDRxqGoYIJoOEWolSAR2MWlnKJ
ohCaYyq4/zOhGFLHIn4f8LJxzYXDax9zkR4pcgFtg/9bWJil8+uV0CyWrjXL+E5qn2Ee63+J2jEW
HGC803Ex9YtykgU3jmJhPut4ehdwufOrlKqxEwRJFcgkWlcWjfHYhUJzHuPVtwDD5fTGcE13Tgwe
ltTpvI/sp/FtYvQFo373da+ReO7Gm0fgYOLKwNGO/uNBDX9sNxBDOBV0IdWufxd7iUCy521KZUUs
c8WV86wAknjiTbKsnECAu2G4zef/ArhZflweZmyoMv06OLZamfEornbcl//80s0WQqnAohCZ8sxp
nybBIak2x1s6xEoKs1zRk4QcB91haQ0O5mp5EBqgQdPBhLVqHWHlmtwb2rsyGlNFHdxeZzPxlVdI
R/lRnHbSvaR35/6FwhBpTuubNacHMIY0lqoSQoW/2oloahZBJtegRaCIypTS7dEf78sEQQ+YV5/z
srZk2Xsy5vtOxJf0FO+XxWjXVTlcu4bxzyMumgSPvdTipduTF5fQ6vAoKXXd8rCgfkBB8IHhY1Uh
NJ3CqFBjsezmNNjsKtWr83JjKb894xCzXsowdgtuf+/U7xcgU8MumCj2Sso6qNBZQKwRnvSVzxSA
ZQpYihToXG6pIeeFDdbbbUs5a3PsUnyRM5/nLisYAyibwJS9JHWSNI7V2NCG4okXaTo9qmjlAdsz
MPbW11UZaF0WYz62XCOp/apK7HFF78qvR6XG03+v3EvUTzJJuXn5xG2jKlOOACBMc1BU8mQw+l+o
Tz3yoMFwfF3msGpVNiy8OJ/83CsSfNKHH+WerL9xacSmD4uePHo7klB7fhKi/PCnEOeCa/kjfG4f
LOm1SWBCHL8W9DXYTId73G3ZZpSdf4m+yS7i4ZKIi3kAh8goizbuUKeiwXd2pPc1vVo/6S5zrE1P
EVu8GJtIQb5aHSr3Lv3ps60so3yW9xW5x6X3/sMUFPmwEBcYIldLvKSHDjuYIP45kZreLUGHsq8n
OPhaTv19hdvK5VGYUC/ff2mKFN/juqf4rymfI6WNVZhkKa6H6FTWzVK9OcpVI/T96PD0Ij4N8Yr4
ZUTUXzsXo4NjB+UW/C2fxJsuhgmfej8otZ5y/5ei0CStR/8ljZ6FHtbHJ3AKFhbv0ilgbBqq+mTW
tgKToXpBOig6eCDkxOfhvP2RW19OqQZI7yDJF2Xr7JUidt1UpJARlD/ItEpRCrUBMrXryC30wfYY
72PK81r3lW5eX4ovXup8BLnNxuUrV/TgneWLSDPBqyuO5r17NVhe0PsMbfnevKyE9W3ZQ2Gjs+7H
lAwvZK9huhrOzQ4dwHJH7Y+/ruYJeOkFWt/JZdN5yfSdR1WLEZTasuJqvIf7HlyP7bS+1fPQXBd2
mC3jXQAgG43un6axXtjJCEMst7DRjQwShuZXtuob8+9704HZSrFcmWBMofw950kSsRz17mwGnF2b
3LBbgSje9c5+X19b+CC60d8M7P9hXFFyN0CI93K0PFOVVfjnMigRU2HCHlsGftZrlXVBww4y7o7e
ybrLAEd1DXKftFjE/X+i7DYAOnmJdDyahW6QEPjQGdOwWOw1aYB4lxbw8/ygUBYEllsiz9sN2hIM
US5TA+2mkoIx3rwgwSloPo8/iMUF0mU9U3413SP6rwHV2zlQv5p1xAqL4u1MfKqnem5s9gW8QPIA
tHBomQmus4RQSzxXe+yTF2HpHToLsmyykDayeZRaNWqtHtTuxxVgLEsHL/cNL35/kafOpusZ1QPn
q0Up1kGceI//FGf+gdofwobW7SvMmfTj5NrfGz4vI5u4/aMQnFV1X/e51dExLNKv8WqsEu2CoOh7
YmE9sjpMLMkwJnhE3tH5n/WLOCR55hwC7Xr6hUq5D6/yGi0409bpnn37IANvj/5ZS0JORCpcusYo
d8jyvtESlTRjFNOP74cU5sIYHBZR/3xcPQ+RVFuYKTdcKY/tJFpeADwdj2FsSNsCTgoHouyHZp6k
LVR2+yqq1mmQbOWY7WBbqEohMpyQIRUFdXi3845j2acTRJdVWH3AsCS+sDHKuypGDrdctT4gk/wQ
VPWy5Kq8Xi0/AJPJ+0mcxPUMPts13yH471k379DXpP6FV0ZKJeIggInTv4Ffd/BgcsRHXFdsLmXO
bUU89AXJ97zb/mvxKCMT+fZ12mYDREChDCx8MHMvCuaEatX385fLIW36E05/TxcNJ94XQne5DMrN
lHauy8/McRMN9g4efsdKntPlNsRlYct2oLrMMH17caaAoyskzpvckJFG+QSG6NeP3hf1UstXT1HR
oKO8yYd6cQC12ABTHZJkUxyeQb5ccslaLv9jKUvz3ljZSgSxnXyULLHTZOeBL9qhv0FK+MljbYHe
VokvDzJVoY8rud1C4YaKjb9VXMygDPKXhjgT1/jkeGFk6a7zhO1ZupNNbiYs8jDiYCTmFlRqjPdB
7uMZ3hEntmigfiDoRkN3FGDDFJi7yO5vsv8BN3NVgDhulwA23i9RzMKg3hc4LIzT60DM50Mo8dyD
UtUDSLDvox06EYZScGtM7odz0BWbge9TkKz0BtG7tztq2yz59B2KtCINB53fwo9e6+nhuA/DZx44
Z3pU5nxrtCNnC0JQILKMBf8dGl9UldP3uW0B91Qopf9XY1djrm2vF40nl+ZsIhiGMJpsud1GrAQB
o4O9iO6afRwk8fNj3mEXZwJwgf6I1lYWHcOQfj2yJK9HkVptFk8GlPUNP6sPkMeDgHfYIH8VjCaH
VUQuwOuLEnxlEv+vObkCZFGsTaeu1NX/IMPIKHDq3vIJgUgYehFklTqBwopItakdIk9PIgFPjTqH
USolsjOugBPoTDPywrJK2Jq8+a5Cz5D9j6dzLcUOd6Pt07DAy9qyxU4iYarixcdMNZbzIft2IK9D
STXuVhNUsByiS13uIpB1HZFehdYFM+T/+d8KIZFibFYGTTMZFsue7ju2HS/7tBYokAw/BslswX4k
FT6NE/doYw0FsgFZfIwO1XV05Dvn7YgsBFdogZqP42L7DRwl5aa5SCCRpz2FUP3I34KbcTxk+GWN
bA/yptOqF92LyBnVhzR+jNftLBXIQDPZ4zC3PMeFm5IeXKXXg4DAwl5Cmk4ZxvIzHfMxfaWEVt5n
OSaPaamYtZxerZdJrVwHFa0uORREQVDMgSwebHoKllYATQnnVJEP1xl6Mb+28TywxI9o5aH/qxe1
kozBmhh98vS01EQIh++CVV1XOPReTkU3FH6Qr+Gkc7ZnOlIOfpRIUmn963f25GHsgcIim5kovZP2
sD3S/15U/EIbtYPR1+sALX1SPJIX4bvbUfAhJNhubhujX5uKji74c4cupgd605SImdLGahDUbG5n
N5+FrViGVnxe2opujyZmSN8i8jlL8wS8o8WbZRcMHQpFovtMiqH4DVXECxFM5j/mUsrg1wRi16Fy
Ht+0+qRP2uAFgQkXW8ah6fEotdm3/KiYnq9FSqUy2PXk+JvU0wTMdn258bebkjKXAkVSwuLOQdz9
UxYrdfqTAe+84ZuFwkQ/HH3EWLVNIyvkxgr2iWQvkQCoGN0sG1kPhRHWdHtVoZBgRyWdx0bQjD66
Hf4VpLwhvVXgXYWkWgKMJdx7iZpBZ01YWJjJalvJZSNXgrR+1BY63ZOBFs7wBAbhk+1YmW4q4Eix
0t0ya9r6Iy6Yql20aLEPVaUYcU4i1ZrQrYvJoCLNOP26GUKVCfrjGQw4+jJYIRqHzbxsoLc6nloQ
rcOhf7karS8P4xAJQ8jzZSjOdOBo7nWVuy+BoETqodEN8C1lqkR7S1wH+3Bplaz/n6zXepiRI9pu
EB4J3V7BFHMq65erYajB9utZddx4/54qMkqR9PvBRHGoSur/gRvy6XL9LRu2VP0mJ3dLE7q1q4ri
LZDZYWlnHs9v76pfzkRbVjSn7sZi28CdMTevfBT6MUEHlXhkOzG22G6QydYtZvvBGF94QTqJFCYU
iEaz9oWQiP3s4VSSd+ecl7PV5VEuGDMFHmKJVczTUx6ViYPPqui5b2Q+rwgEO+4NiUz+J0gJ3Tay
nGkmROcChLB0YnLu86PrcyHjl6RgEDFM57Xa45ZWYyOrtQIy6KAtz1CXUf2C7PDdvkCsVoO9SW90
QPYQZQctuRNddkTQVgLqbReHcRG38OuYf7o0AsVBgDaa6MylraCZlta4V/xYK5KJEMbJnEZqmir3
2uOrMgY+1sO9LF2IyI4/XQs1QGBCwWpSjmCfnWCkvJdz+K+0YKzQ7xA4/T2ColnOsn7oH7AZQ3Hc
DzzDPYYL3Eytb54YfP8pITn2LM27uRkwl5EYz42U4lJqGaNoY33xUHrokn/xF3Z+JnWgS4/ii55i
JnCNHOPYUmYxgaC8Z81nTFYWVW/3C2ILxE7wCkh0PFqYL39ACfFDPypQqpvwb3EDe0VkKzC1e+hI
3Y2Pik25ZvAfTUqfDJkVRoRrX9iOF4p9AVu64uxW1KY/x86eMh6UWCaRSVTdYPlTBBwWu9I0aAWH
hqLh3wTOCioFtp5i/XIpRQF9W/0SyMlYV6SwPUfOL8S58DOO7RcgrGLqr79tKPg6OP5/caEcfBZ1
I/zL6Uwh/h8YX3Oeqg0uuu5gk2xQK/nAk91wxCqmHiawsofaK5KM8DlHvbsfIDbH5Yit+jSyOtAi
RaqRvixVLQOEDZJUAymQ6GgXuA9DWVjqUWMyOrshZtVxNdjshUQjcsw+yRYL7B2jKN51sBguP9xh
d8aWIVJskqdh4NtM3yF7S/mlgVohT/KdLKGl7iGCIDV1pHwSDOX4+/v1gViVe8CiAnrUtVKAqeDP
sjR+XYvz2Oj6hgIkGw47lpZeyDLTrYJePRLImMK5rfDclB2Ou6VbKixHxgNLOO3YO1Sbjp/sFx4b
p9PMa+N+EI8TvAoW6wTsy4VFgXmWM98OhNU6Dfmf1zoQUir26AxB+K2iJhqaDshXkOD/MDA4c3/4
G3jU/+kSRIGsfVCtebcic6ad5el4ciO7KF4IsceJHT2lx87pdKon5Me3Z9RbOsOkLchCEKLi+yGi
unnQ2IukzUQzVdMXyrynVRWo+AFKeh9iUzgtQgJaUlguxHRDkL+rOBFR4F3GwMVSrScYnwOE+BnK
gX4tSF+9WZHH45um9NMIGcf/VCE2BqrUay0MCBXnmoFO+z9CzDWBIDbi7H7avTVrkNhPILDEoYoi
p8pzbLSD/O2iDZRTO0jHCviwO1T5FlkPO1hDL9etpa3JwjEPDEm3xExnqY0QLLYnpoh8Yz0zm6ZU
NHVLUbJ6D8xf57VAPq70Gd4BLK6NC8bm7quKvdEw904nLTE8fLtpTsSmHXlbxI/VsbklA4/kQ9ao
dXU1VevGVLJZeE0I4MPhXaYZHAAtmDkzbPb5oV71ceMSJuSCVaPrNxsuSCUHEdaZwEVwVf6WIirD
YfQfryQ1awlNbf86BU6bN7q4uSzF+pjsy3NDK7X5hToFUcO1coiX+ddkIT/B2G6KzsDzPlQ/G55y
9MsSrTLROyXKQanjNeynFWfm1RbCiKsLigqTtKpI2a1QABtrmLl0AXS2XQgXIINNIzK/Ns8Md0Zx
NmMx2RRQb/giQWH5QMDJhWioYTG5WZPEfg+4G4h07ZfJepAw8etjggeGisdkbHUfcDFCDfQ0IGqB
hwXwHtBs7Agc4zyAw4lAOTidnLg2yMi/QOh66uni4KovPeZsZlAqyNDdFUIjuUuUTHuo2emTNFBA
eMmkznSYWiBJljnH2KrYM2hpMYRt3x5o3joncxnpc6zAjGv2SLIljubGkrMV9+FjPvMCZ9eG8y5J
b+G9qo3vlMWodEFUfh6q1SSo+a4Jg3MdIhMtjxpcshT857uFTInPcYubS2BHUWoA8eD92z1VJp5x
/b2EcOGJoqvjvqJd4ou/EBl7/qDPYahu+SwnOUVccA52yeCl+kZSPwyjHGZizzpzqgRCGAvtbTMK
7G66NbPym+ZnZARml0KH/wZkb6VEXFOCUwq2OZzdVI1Lixgc9+2k5rZE6IXkc+GoDR5pC7LmVcA4
78DJrE+ElPtSjhUiHt0aitRkyAUCulqF8JSH/E2blTeIJKXMht0DmQeA/Vtprv7XLgT26A0kh/ru
8XQE5Smb5pcqG/roCQxfL64wiHMgVBGSmCk8riISeUs89DK4QAjPEZ41dnkuVs6KjdujUIfhX/b8
GkYYQiwn4E/y/jiGTjvi+IVGw8QZUqY5G5k1E4BnhbvmxxkdbNNo52DVuK6A/YHUS2TTYXHPoVNx
dxJafxtjk+A/VGVlxeoj/4vgbpY/09nJcD+2dz5rff3JDndhQKp8k6xMqQKu3xiqyQUcm0P1BZMh
tFtOlrh7h7nLO+kxs/alHN4URAjtyuW49QoDRJgH/EWw76VghcuM/mgz9VSD1st9Wezomi2FzJ3G
xcuNMDS30uc1/hmVBMgA71RaacQtzlenYIk0ElZdNyDeGdvJ5hLoVycSfE/ApzGCdRWlFyo4dqnT
KQfjK2pKR/mqGD8WSEFVovf/LFEqniMr9gt8CC/aF5PkbzXqPiHZx4REEW5UTosV9TXGqIGxE5UK
cok5XEcUDjkiZt+GGPSlGjXL9/LeEt9ZKx6BNrACnsGvAOVnLjWF5nmhjKv8hNmxQQ/OaW4QZHT2
AD1l+drCPhHQ4BWWRjwUoiH57e3vMbtijaQe5RrHS2BCnfI9bogEIyhQlPayoDi3XKmvZCNcvdxc
CRuBF4FS9+tKk73S7Z/dd+pNOEE+xcEz7ArIykJdxJIFlgY20K7EPZZ76dzWS0TinYnaITbzz000
vM0ecSgkZV/IYisyV8Y+LrFM8ci11CRG3sKzItgUnEAFulPNoy1wo+u92up69FiQT0h6odKK4mRp
sCtFcdyIYqqSZW56txBlJScTE+oJHZ9jpzVDMA2trFDiuTEW3CN7pr7kuJz907uoBLApwYJUwX9/
RFWvgj1Bm0cdfN9E3w74Wbz4peX/7HanYrKt1zHjQwIV4ssvQI0L9pLJljLsCYjyauNw3R3MhHAu
/b83yQfPyEaBkisHl0hyW/h92SH6A4dWP2Ll4JugYgS4gpf70ofzSx6dRZRmjndxFk6YGXwxRL2F
fQBuFAPnmJXFOG9hT8FE8Lozq0Ipb/WSQdUBz85Aox1HHMAUFXWWf2Q30rbHs08VbDUmsSsnxGrt
U1PP0l1eCohTSBc3ge2xsQhKN1wgsXKbAV8B0vc7JLJBZqQl4+YLJjo9QrwfRzDdvyIyfhF5uNTY
vB6K6C61+LRkBthxp4ebs3fMOE6uwoOPwyqLYTW3/ySbCD94Ir2elMfBCJVoHfmcHptwxIPGM8Cl
Cu3qOY+G8aDZI2fEFxn/KGr12VCEw5M116T6xfyqDSqb3JjiQGIEw/8OEXVkYv8Gn5j0XtCHfQ+7
prEJRWs6iFzZk2m7qdERwCwQIa2amFso63h/r3/0fe/6wc4Pmepi8I+Lxq0TBiPww8AXmIN/GOc5
wJ80s3B6Raus+D/rSgzsGmtEva2NtUiGgojjlEP+c7ynt2P/4d+irNTh3tPTWkgg6Dkkxy3p1ned
jHaNBMr91blR8JTxgaXPasZB5gjsMPdGXA1qjM67Yr+rBlTpFh6k5aVs1N690W7M6yUaG4zUYQaP
NJ+wR6fePP901A9iBmCUcMNZNPfQvvDsgiJzQk9x2qSo2NyyPeMbnjjAngTqh1gJegzzYM9pB789
CqmIDpleK49uouIKVjJBa2UuPfY/FZiof6b4YyFvFWylClYo0RSdfQQErecpODdPX0y88IGYbsgv
1k/9WtmNgPXHK0AXCr/sA4tK5mtOsYErDX75X1ka7Vw+JSeLU4bwyqi6C136Pnx640NcQXYHghHF
DY6mJXEQ3LFCrlHO7wqDYAFDkNmqywKs6300nlA/sbHnfyMHdXzNEKuN+TobPYMVpd+V02rThiHy
K98ptokVe/38umuR07uZWTa+WX+5MPhH/24JYf/oF5xM5/Y4B5Tahedq7J6eC5c97EKw3fiOTt8Y
jOzbLSZuR4PBQ3GW5KUjtuhBqQQfMLNh1LCKMojirIPAkg7ad5saaADlWd+XsGA76eOUTSkWq2ct
d0oqcO8m8aMQk9GM0VHIWNXtrJboqzNGR8LIPZmaQzNlLCsBaC2eESOyptItR2ky+1ryBq379wPe
v6X33dd6a2SEbunmNJ2pxzOrZNAY0WpNisVFSG15f3MIlLdgihDhaUaD3v7tix1nmTmYynK4cre+
4tE5tfYiadDTxbG3pKguPmWZgiz1VxrS1K1k7mucULP9lPJ3NAnJCHXGKDVpM4OmdG9EYYx3wAVs
xX96GlcqXGcgSb1UEkfmzXkXIMht+LjZnVF03qUoCxtQsyz3eWNvg1n+lSQRdIBNufj6D9dl2TQr
+nRGmLl9kVt4alyNtfv0rL4eCPr0aVwqU8E6PoyXxGwCR6FzWeJrJc/f8Moj0/lV1w4g2To2Hy/4
sKAU/j+yMjVBhxPezB5meTYdxHSar/6a64FHS7YLbWMkuukvw2fZBaTDH2RgMGr6wNfW78WZvXi/
NPCiCX3GQKutbFpyftaOgf5dVPYCTP0KcQEe1XunRH2WMRCQ8u79RoFurd3Lz0Uo++P3FEfmbvj6
jOO62QqIdnOdP/edv4FLGthrkLGyCGov4Tfu2EnyEdMdAeQO3ezmNx9U8qi5ZqnlM5rYUEs+cjRO
qIg5PnzoJ5KYmM7DomLy4C5p5b+hhS3G5E5RXarnC6rkWtO7A9uORLIxdFFkG3T1GZO3NXjEiwIN
LC/TGirZ9wTbhn+qcRRfYzXOY/MeIMVovxj8Z4aHBovzNQ2OQv6REIAeScyKncM0eap0q0+MtcRg
NZA1S5X7N71SSnUZvnaulZTx/sofgWsBDZy8laOPc8DmmgPkGmJU4v4ENGdcniws4uGuQvTznYLf
VTptO0jrXkmrOv4PESPZ/QF+RBiU8OnuYdfUgA4ZKmKiIbzdlp6z4IiqcG4OUINA+xBXf3zb6KfU
0s+lpUck8+Ucbxe+MBULH30P45GPYC5qStytCqGRH5jcczq9wMaFItH3ZLMUK3IIMPOAE9XsmNlb
EQ5o/N/I0ayLcWRkv6Q8nzXlLA0ekfvIgDL9nXypYGvpsvwM9O/2iZZbAhhUeke+f2h/Z6Qe3sr+
huMJ3Ap7FrxFVc4pZcDEV0hPLirGlV1vpOCfN2jGU8EEO1d6YXEjgRG6nUEYXM7DQQEIzERWVqYv
NUfYb0IzsJM50MKviUm7coLsw0shSQQYVfPCgES6ErY8w8/TXnD0rr8bw3iIhed78VJQttxywm3o
1bE1buV87o/gh55OuzIWPLqTph0d/sQcO0xUxSkxTdJe48dcSNtx4II7G0InzY/H8hSvJI6Nnh4U
Ca1HaPP1n5IY8vLEMPQ7GIBHOxj+0G2QabpT57rE9JcnT69H0PNjkan1Hk6nSFYs0jxar2fy7g2V
MymER2m0pf73uAM/wI169YVmDF+4cQfQVxxxywsr10Gy0AIMxsMBegTJhSygqvZrbTxo2O2EUY0E
XyEcrDsbS91fr/IM8HcfOYupnA+XP6oqBnKfXWqMhMSongecUW4oapzn1G2rFnQHj7J5nfDzAF0Q
uuuQ1EjzAVAM52ogFxCs7b84w2xstfc8d6a+pymoeLc4XyGlELSnTUSLgRhT4nTKStuL7mBTQGdC
fa6dhcxQcebqgdWMHWBUm+fjL/ojD2eTXu0VlE18XT+t5XVks2y3LBgpxG69vNC2Lnx1jEn5Aen4
WLdtpt4PvmZ+JztH/PNNruKap1wOegfI7lTnTnI8s+/T6U05uUCe//jaE4YQmbmFw6I/gNVa9RmN
iRbyQEcfj6cIz/dTxdDw9y14JSFqFQX2Pz8EIJSXvbxpMLtamglwWreb4G83yYyHRTsp8Qt1KuwW
9lCV1jD21HbMvff7fUnkPAdoA4OtIU9AxRZsc8CKGfNU0fsQeq+MvNF6oD5DVJtb1CIKI/5J1Ian
eeg3oRTXsSF+qK84Jv3M2bnNLr55NlAYOg10FbtAN56dzFZFosOSXa8pnC65Bg8OJY5XZfkCqSmf
MuPwl9erszaamvZH3nGA+/XJh+nrvwAqOEacBiMKt/792F3mZbbatKA+TlcZ875PeBld02ycSvS9
0ybCjwftYh+IbM3cZzPEkrDUpqcmfinzxHKVQOKvNjFbLdn7OXXxOAtmaZ37mTeIajo8+3azwyvM
zs8odKE9DEL/7WWwKtvodJTEjl0WL841FcLHbA4ql1/lSE7A2YjrWwG34u7fWcHJGo3G8KfYVJM2
JFejO4+5s59OytxUu1Hb2g8LDwkt0KlSNy5vJSq9r1SKwheew/vZ+5aGVUVr4f8cR30JypLOQH2c
Q/9GivY0v1rLgHWxf6+uv+MMbulw1gBtOqJ5mLoMVqkGl/a8z9Ef6BSlS4f0vXA3dFg/UrwTmgIm
OvXAdVmhjijmoJMIHLeiblxxy8LWEsYR4z1v8Ci71K6qfKUg4+yeFuLEtrkvqbx55pHxPQmnhO+O
G1OFFQYPQR8xfnvIKyR3YzGMPtSqGXvd6A9VnA5wLdaEJNX16LRusCXo/VtSAOLRyTeYJylHGSYs
HpalC0mpr3n+CF2QyF/c+YGcGSHCPUMTzKw0cMVw/BI0J/gJnzP64fYGlPjceQw9ISpsLd8vzNLN
jyWkC2wJC68rBSxsutKKrU8YMVe5eWh6Knoic8oZo+yss7s8ET+Vwt3TWEuphIAWouNYRsttjF2O
jSe04yS2n8bkJ9LsgMgDHBN4rhN42y7XKRHQOyK3rTW9lFMucHSBLkz3BrJrcUPZiSxgiWahnCLW
OqstOJlO3VfvuLtKPMTbzlaAPJGaxyeghuMTt/by+ibL0mW7aVqs6WpeRvZ+5uueWw2N9aJEmYV/
7VzMaEEHBRh64cind+Cmi1GZSXYCsk/Lp7GZrSP7pV9vW9X1VN/QUQ4aL4QXdqJ0+aKgOgOtAfLC
eNRk+Z7p/VCvWBymLwCwAr6lxxanYnA3ASIYPpZEd5AC3hdzMS6nyXx5gLOr/07/GPqBQrjZETsY
f5xpUK8Yo6Ybx7QhGLm2vnCtER0Wu8xzLa2eYAtF2bh2BMwffXjcfOvGQN1FVQT0QAT8bmv9I1wE
gB5dWsXv21DLrohNr2hUx7pNwTc9gVkQVp+36HR+4H40iR71/zb0e+BHBLmZojlhQbWRiINWk97O
cKbAwUlbeX/TOmTEw56dhncXv1mYV6ecllZXvCad2AJeB9GMEJ60yvkdUY/Mq3KOWeqxhpCLQQHr
nNUR2uhuzWV4VR4Qh3DFeIYU2+PCWLyv3D9wuvo9hogP4+AKtDdS4FGhkG6YnBqkWbCTXh5qzZTu
y+/KdCCqeWuNiOfYIz3fAbq+UchbksIlbb4Q64ZXbZx9gNy0/qtGwIaFhOVHewUp1YW0cIy3uw+V
aKx2ciqUGcBA50pILtw0Cg5JwcEREWcW41uGkXrsLlvtDXJLuwWEab02oqwW2Ho2OZEHk0wBPh1v
KuAx7CSmOTntkhKpecnDiooYUQCqcV9hGSB1X53NzxCXShLSYAd9sYASIoqgh2er/Q6bCHNkeAKo
IoeFEJoHW7coc+NIu/sOBUdb5p+v4THfh9DmxnJ5FoYQpj2s34ee4LScDYoEGKNXlEWo31JKvcmz
781lLuK48Ia1bZALcAUzY7htrqYC18gZUuvOJxYfDwqI6pz4GYiJWGfwv4JbMO+D7Ukge+5FjXSN
nQBsTsia42QKkn7h4inSn4fFLJj/BFlsdZvWZOz+bkQXGAjbhQNfZrpSqGTbsvy+jlSIdOTONFDX
PUwMO6yMa26HC6/LROR/Ge6p4DE3KL1MF8w31W02XPyI+KhZIjHAVrEaxF53yj2NoB9uvQnuxghB
bI2SMlpBGj9zeiJaDMmRF5VboFqHgAH9lXnzlU8jO1VT2qGmDysgHemPQHv1I6w/MBtZx07n/XKs
vSz/Z62bWUjGewHaOpSjlc4bMERK7M5NvoaSWbC504gP8bdFaJpa4aXRtvNZfhKMA8inNFzxEzYr
tkC0S2ZZtUw/IX4yY81JqTh/9WQzr8D4hB60AM8HUoeaRXow5ZhLwW/PYAopbMTi1wDPOUeuYSBB
jgecG8ySXikGUjJ9hycuUGaZ0wsk3PY/8PCzEHWDDZ5r8LonNnHQzYXyL8VhSzDxmm47ZD0kL6eF
8U3pgZrlZ1LiT2AGRNDK98ElKFpjGTsBgbYiMyp8i8HihbJ+H/kbp5mV/IJmJMjDVdnUgmWXFyO9
1Bml8m11LsZaN8S48a6L8vpww/xwYU7VCAGrduzjks94BVU3F+EJCdhwUqupiTvmmM2rIPqCVyfX
S1fJ4z9WW26RS+zBqAdYPwKMXoLBsztKw9Cu8u2sA1um+K+LdFnE7v8KSfV0uK1UgYglyhMNt9hl
aBToFhgKY9tJEHJ3QaDGR2aNOAI7kLwTGHs1reTWnhlF/PwiL4TT6xfeNbZRxSDCwmmK32DtID5j
Qefj8MVn1qmle92X6o8eK1Mq84dpPHnF/xsTjVx8SEAaMvNDTXqprbHXcMCPPIwVPKueyP5VDCyc
oDg9ipkNEyL/bZYFvkbLX8t+0SeOT/dFeLXB1sMRuKPCo/Dbn9h77yn4aAtPtixVRbvP3as/w4/e
MMSocW8xv4vbRzRoKJrQJHwtrni1qGYvGVuSggDF6T/9o4pRGeHuO+QWpGMwdhlg94wKgsKtOdPs
9+V+8t35YxsXQFPxsx+eGH1q05oT30YGegRK5VCUBD/QwV5rub+KCGmrHePClwn0oFSL8SUKQpHj
h/6XPFInf2jqXfcvw+FxRo/ZFrlfTIob0shObrMiHhP3rd/mHfcn9T02Xt/AJ58xzYWO4upT3DFq
bmcEYiPx0gDkQRHsGQ/5BG2Sjr1GWAMSOr0WwIaqM9PwbpiQTHjEPOSeDN1KK4IWDLeUEkTcbVKd
7CIoQZ0etQy/vOr3Vp8e+7luGAFPJ2zQQH7ut1GEQ904Km4qclnNfeX69hhO8Gf1HngaPPYjI/P6
f3Enyt4zGW15dJV3z/IxDGo/XfOaA3whrIpi4dYoJQDecY3HUVVsch3bzJxGsluwdY4ULNcp/fec
FvpZZSzmpkh9uC+VwonmwBWtp9rh/jBUoGUTracwL8ATtHkciPfOetJFAEM3KgRSsuK5t8GcaFTo
h09S7Y8NzaL+m5v6uRl5nX7qyTumq/qIQF4MdXmJzq4kbUA9Phk0gpQ4N/oCXbPbViKokOFwhX+u
t28xpl2W8AfYpNGyOscRwX55PjyUsh13yTACQ/6TZDdcncmudsN/tNpHvJh5sM2bhqQWUSQHRoe7
yJo/6czPtQCvICuZf7WxacXyJBi9UKwJstHpMa6yfL5ghwR7g/1PAbZ5ipW52lTolOk0PjDOlf5I
3j+tIv3c+WXAAnJNRhkY/KEuGS6hXK1QR+ZP3exskEzUHxEICD/rwt2UPFlk+KRQadMgUI4xiJYA
Rc54vQoH3h6i1h5QBHjTZb6l7jADcD3xGe6jpiGonm8zYlH2Av6qj39PaQUc7GCyG0tOfIn9kvEU
692ajmKNmsJYwrh+P7gJfHa4XXHCM0rvlpwD1dM3ga26nyKXCZGm03PaC0zFy/arsWSB6yz5XvbI
GqrvVXp/KluUk7+BJH47tBJ6uDlEVMUPkOmH+rYlJCLs7iGF0uTnmPeUB4NLaHLJ0IuJRyEsNM6D
9jQe/t1iBwkL6/Jg8m29PbsVeW3rBfEqZRz/CR1Muh3Z0EGZDcagK2dPeAjtiHlH+6D63fBAJOkV
BX5AX3tRBNmq8vyRHpw2k5kwE6GCLe9oJ94WXKytmeTWhQh7u3/IRYU1249Jh60KAF/z4ZeCtGhc
tqnUhQ1tT2w6yIEnmDTVlKr0ctTYtnwnMoAJvO87yp97L9KuHn2tSjlbhP7TRlf0kEbPjjQdlbW5
7vBc1F2q/bfU1GnZN24DDuxmQedHuAiZb/bwrY/l9igws7jJLS+RSst3DXAyFmHC3yiYy14CAMNJ
sbqBMutXtLrQrnO0tedLk1GtetHOXeq84rM5w/X6vB5tiyR4kdBDUFy+Tw7ijUMJqXbJiNmAAGXI
G5YlTH/XXhq8alboa6mbBXfq2/MWvnY7nPPSd45XEuzkXwS5pu2SNSDE84lJcdcLSmYa48K3aM/Y
1t4ikFGbRd2iTfYzhqxgeF7p6JiiBqHN3e5h/JW9h3W0Lqcz5S+CliitDqIVBPHq1+bZWjURs7Ak
9V+TrNhzOF3S/ldGj7qH8clRkNTLrRYcf6RRmBE583nf397A7ST1fj5i0ILKiIsGkR2QE9sVAr0f
1v2KYlsJ6qEtidZFPWW5ibhqXcv685pCzpYly1ECozvqeNDt5fhWZ6/MpQseqDt5KoGRzvqvWgUO
lHZrzT7qGCDKkEkn/jVu9Klq614x2YWRvK0Cgr81k6s7z5KAQim9rH4k8YVBEYVXlJlpu0KLr2ny
1cQitJD+JeYz8HNA0MlT6q+JfHk0phtyrTK1XPeAO6P4AviNrK8mAk9MIc+H+RxTnrwc/hdR3IWP
n3EkSviYCtb4TxrxK8KaxOe6MF1vHlKMXoI2nVOvz0iobmDS3FexMUy8fzy+T4RxM0wvAMd50yOE
d6aJXXWL5FBZVxBQ1mwSKGyoNSicpGiHvRrYlzRlIgFMhixbnmqrncdYI7fTMqK2nawQD2+7/RbO
pJEg4mEiYGfcraOWgFzoJeySh/D1r8tTPwCc1wrYgTfqPGDYEBZ9nSnqmfgMpv6KvLFo5ntUq5EA
Kvv9XRzkAkBBUTN7NtrV8In1F/vk+jT1/DP1T7GuIMhvQ9TnwP+0nlAQu7URpskZZARSANzy+65Z
Z7QMKiMfrVkVhOZ17tx5OE3UJpF1CymudJhEkYcDW7EyoTGZBdz+H74oPkwhik6teW1LJW2U0zZL
QMmYAfIBi3cZQ5pVSrtFW2NYumSh32G7ApPYDuMoDpRfwuDpEPu+JTkGmZhGhQLdAWdgwco6Lhqv
LwYCv2sPUcaziwTBatz3H2Tg91ZOu8qD/xRnk3LkL0KndIedZm0fibsEUd0F8b8B7fXLf+k92C+L
DQOCufuM7xkSRLqa2l5ys22zwgOBfJiblsRBjAEi8cZd/IU5bY63Uk+rNCDJ4gmCvXPghsJ7Bbed
hnxbLtzTwItJS32NL+3PO/tAdx9Pz9GXKvKDP6WZFhNCIicAkWlsBd8tBMNIXgHpvxIqwsy59dmN
FsuMBAui+Awb8+XaCB25U3Bpfkam9cOiiuhMjeGlr+DSvICeUofOR4WGVXlpRybyfNBtuQr7PTzL
bRh0ukc7Cf/1YRcZck1VQ5GmhHHZHTr6wdp+IlgNTk8kr+66J2Yy+iHV20OMYTK4ypls81CJVnVR
Ngcde4Eu06dfQckgUPERv/CNCDpP93+hk8f6HE5upgKwuMtqHlO7NpRXV3NqohjGTAHpdl4FswgI
ezzexCO6O7tHfLT45NYOzjRVxC4aR69HCsQizI/pdZQoFg0EsIokfnyhUC427jh9KetuQqDnJS93
6QwECaIU9rLxvpQ1C2G/DlDQlfW0I159hsC98UV901KWgsxTJH1XQaqQpXnLnmbzguToCYP29yNP
53barxK7/JnXqT68+QV1RiXbuWjZeDOc21HvizgUGEDZW2cZRniyQVkBoM9OD8FdkrW2caEnTxVX
1JAm/612ViPsXaEuOfUgKJ2D8JS07b3R+SJWPu2SwAoY26GxejKQZ/0sQuy6IFAd8I846i66SKQu
jzSDonHqGoYpIe9Gz1HVQWHVy/brXmj/DlvJaaRlYptw+OivCmSxd7WpNgvLdIBV5euawkgbDDes
Pct4sFPJEiCkPyWQrJsK6DmALbRDxp4uUPycU05qVg+fcoditzpOfXSqlU9dKVtIIHC6ExzlxAFS
sV0sEY4e7r8uvQ5dZLJ21X4HN+QRVKBNkxOnYOZroWvXNiCaKLSz6q2TiSreLGIoeWWuzuJdQ8rp
ruLW0lrGiKePyUxEhUAtPXR1V8rJOOpNfbWOtkGcv/BTYiTELX21MxHTlkCwqKSQ89f1x1FrkBwq
dVL/2cymXhZ+jYo/yFAZX1mPCDfIz+DdpaKkeg77nD87rRmYlgk1Mt+3rxB3b67J3SeJARosB5UC
ilm12XE4Qcbb+BQ3FylU3hZZD8BktBdpeW5qLknfT1+DRru3gVx6lPl9yM1EB4iNUlsR6D+SHaoS
Na+ELd0WHXJ67CiM6Wvt7Fg/9FnCg8Tao/Uo+pW46AxQgVuUOlTGKMW8M0GolH3uFLSEtj8hji7/
41zzUtZH8myNJwjB68tH89+d7UAf4TCvVdDkWvbHH4mfvFC4kV2tST409iwrclGgHQ0uHCrZdXVk
2XtRMTr9M2NR+ZYzbTtuw0y6B3DXl/Cf5D1r7gMe69swGCtBnGQXM5CDRTq0vM1CWw29iloLMnlK
27squs2NRh4tj+p//79LkShMPCbHDc+9q+lg+swbXsbDj/I5X5yNnWZmw9bzuWI8uqCaR8TPxDFy
h+HUGl91DmcHIqEQJxYczeFgu/H6KZqldGWeo+YzVwo+sRVresh+N6KlWPfsZ5ymtiQdAS1Nclfv
uFp0jWx+hXGX/1hcxoOZ4NLAt+csLcAVIqiVYo/ydzHh4/XVwQrSICWMM3UktM3aUhg0FtmYWAI9
XNyaNgLnXEzz1o73Q6h1w73NAbOkWteHeAaTAaghu0YjZqleNgSUuFIZuGiKsLCa3mWMHrTEeIS9
uMQNdEHacWBWfkReawqgT/sCsm/9mKrW+E1tGW4JbmpobnABV3iBZR3gE5NQkfqVpCAb2UggIspA
hJ95mqmegP1x2EIRibZqo6++JlISNbSVoI8uJx6AJrna7RCaUOGirSgSXja4JagoWUA/vFMidZ4b
3xet0hv4skjRyWMfBzFsGFra2/pJn1HWAtioi4uV5T8dxjDIfWuYHrwI66OrZPCvJ7DNMXVa2164
FVINNF/91cXHWjraZvJQzmUGZBfyxRpLnt4bxr7OhHj0Esjz5yfbY8tvZZWXQklNB9zjtWFcACyH
A1rO/eJc4l8PCwkwJpLsIBWzq5YJKr/oUWHTfOkBiemjPCqTUj6SsJIzE9r/DJKASreuMpMyfxxk
mpsx5jJ9wEY1GGmlMs+sBPwY/xfVZ2uvjXeXLc2983VOtLq2ME+076VU4WUJCzhmuQsq933NXAlr
M08t0PITEl0c+DPHsZ/ZtTnnddI13NV42YFbixtFcR6IsAJ9F0x4Idw9J53HWp4IPFT1t1lwc4yr
JW7mT5ObgQ3ZIH9QGHqJr1s/jI9klRywWxU3KxA8naXnQvU1wdMio7pjTXQV+QOfiPvXLEl1btci
krw71+jG/XowObQKbCxKFxbRBLQy7ILopQQru/Dqi68OzDwYrvntvJInGLKr/ruhVfqlohUYpmf5
d1dSrcVGZKrojlNIRDlDctlNJpKmNdLrN/BgvKm2G4qULgEAIquNldmkwGuvsuJh+xXuazz3wSf8
nF1ApW8LbjlEOTTI8SpCqNgvxb9FveySu+bqqxI5R2ff0wOk6NUOVLoZSP7pgLfdz1BwIBowOXLl
QLyWIBZiCUSaj7puk7++cA7QKbpdwtneI+ssCfeOGGQg26okbf13BRRBb22Tm16WOYktD/1cIfKA
wkW3gppzlyryEgXb7fTDneZmN5esPuK0JLmwGet0MXtmV56sChX7XO0ICyYcxQ3PbNQHNZ7eMVil
uP+l6qjPU00A3tHeSAD4STRuBMxvykwI2FG6Wlu2Y4tCOiEhvpUjmsohZInAco8Inx9LEYSkfNEA
s/erCLMkh3HkE3tlwdjlyR8oZwjLkGrLln2lh4CK/DHMUktW3+mkrAGvMvKLuH9l7wsWve9cNkW8
UhlMdVQGxHh6hsJ8GJv2E8Ow1sayCOOD624m/0IPvT0A73DP6MDmZZUUfYFgnIJ6di2rNmepMZM/
inmCaF3hIQZhInKNf3ejXvc6vYlHFcgpm5lN5fO5aG18ENQY3E/RQeVqWqCocB4+qF2gCA+aMzog
4R7WQzbCdiF1N14GNFFR7J13w9s1RT/RSsGAEpam5rwkF3zNOf5Yc5cuPHOhL+CKeB3WHq2DXJf9
Ts8JEBZlyjMu9U+9zML+qPnKSIRfBirtplBl42po7HlQJ/iBqCthsXFseg0UatlhGiFsbsZ3F5a8
jhGVF1e5h7LtD0OaiORqNHrqxD86AHKF0cvgnlCfz1+yW7gP/0qUtbuptUKxNE/ncTSI3lzDf61X
823KlK32Z/lUUwyyMcOrGki/BehH2JqpBs8WvRo+Bt3tViw5ETK6cwlqO3YRXh4hY2+jtJSO55AP
cPtHF6Af+qRwL6Ob1/v+G6C0mQNsTRhkjhqrGAeAtfXBBcyyfAnqnt9O01ga139w69IuR5nu46z9
yXLt7UTx9DaA7hEf0iJPs/DhRessFqzsSTdKfJm5I9orQAAiXtiHcFJLSXD1yiJEt8UD0kGpVK2G
J+ci8ELBtv0i4eXEJHzlIfnB6D8IJjliVtuEiAqj3ffVQ0Pwv8NJQyh/bp+zAX/cL7iWaH6IwdUk
75t/uhgzY7L55ba8aYg7GNn+Jb2I7K5cLObvmqijfU15dbO8wR9QKJ1EFL2gKgIv0Z47p7ut3qCw
Zm9vmCEhRcuQIqKT7VsJFnLLPzcKqfGAR2/KHi+L9dhIrtlpXv5Uel2ndhSWT+MBX3D8MfPuQ3Ko
JU1hodyxqeHDmaTnJ+mYf+lcPvzalRG83ebpiFmEn+SnY96ooBKIoF4NJmEyZKaicTU4t/7BbBVy
SUPaOvQLziTuNBi7PaIqOQr1RV9vAIHXL6O1NNX0Skt1P7Hrbw1W9WX6/s6+hyvj8nQFF068czs7
ZooWAYsYG7f++slq48jB8HkW7SN3c+VA6UkxWjrmC1p1uYPrpZEE8kfY9CGluBe+FFKCRvQxxJL4
mpwaz/9bqJwwyMg3z6hnQv3ukxDWwudulbCWyy+hzOk9RUj+86IxjhQB3TPqxEQng8XbHkT2Jy5u
jORlV5QPcs/+OYJf4iA8v/C8kyDl0QJ04E7QSxLB54JaDBunkHg9JZ6NMUQSYcuAMjjWxrxXrViJ
7jgX08/bl0WbApieeMAvyqQLKtlz26Tc12AIWXYty7VtqXKvVPSalOTCo1hIY3oUQQ0UHnM/hzqE
zOAGaX1URZhWJ6iKoJms9NKIKuvI1iZq3W7tsvTNf3uWx2fGlHBF2kWUvOF+cXWOXKsP06HoxYu/
0bfZLkHGvW+M7P2+TZ+BoItiuXUh/Uy/dd3smwjxuGvlXFnHEOSRIy+5d8m7isv5cy4PbOEzQf7t
ckmHuHCyQ66cLxFwMoWO88pvYk2AayqEruz/evbaD1+Kh2b9SOgpAROlY7NONrf+jBjQh+lFBYGb
eCMs5LINToJXj2eYhTCpJu1OTJ5sRI8QauLXuCk+cmw2bwc3lkbqiUnryv0f8b/LY0gUTiULOuUZ
7cRLewPiG0SG5+BuLyJJzVwkphEgK2KwxvN5uOfDkBCuveL//NbFnMvtnbDH92yzhoYqz3J0QBlD
I4VAhZffe7T7Qti0FGJUmlIfYljf3Pr1dxBh/rEXz/hCZ5IKf0JCftMAsv2td9iKnZbGwhUMFWkx
7FGCxSgzBBURhNQY/O2RNegOt4os1XT1Wye81QxLnC7U5ZcOUdctpj1rqWscxxNMqn3RRCX73ftL
sVf/NYJiJz9tSDdZI5n2zLyIMvntrgAqatj2rxfRXCJ+9oT/Xb/hA4k/Mw8MUw6ucuZ7EL0+qfLb
5HKmFDKLigpx2E0+hRcXA29za+WpEbbMoggK9j7fB5WFcMs+RphWmWjjBUyoZGgVUO57KRmFc1TR
QF80gT+FY0f3DECX2731e17VvU2bqZ3uww5vh1fnjAK5CIdforMlogAetihecqCBociGVP09cx2O
3by+1XTSPdcGbxBy6CrH7AxqEBlQtlasiqRr1hcAeXUmnpwrmXqK5gnxktMN1s9YyWVfWxPVjaYv
w478BjqXcnkoAaoSwklfkTj2jQWQp4P4MbYENYoqCmmpWjtyCMPLuufoP/HpeyLonVt/N+fYGsxP
npIJzwDpqzgRS5RxmM3whsYzdb4w+0sciFY1yAJ41fjBfuZ+sRBUv4NH4VZn9HrRuJ5Mko6sjs68
va9IBO7Q+oGfWhDyuXhf+YWWOlkcl1GxGe7mF5wTtrG9wCu4OUjZsFeP0sFD6InfCBURqL7g14jv
frAXebBnTn1m9WJlLX3QGCILDbhtHte6mNnHsoDFAZ/2eqmnVc7lGklCd+pzpIXTz+jQKKLWO/DP
yDk9X4GvEY3wvsBq+mUrmpbrJd43sn+Db1UwIxR9O4TyCgBcxcFFwbjELSd1el3UbvVO5yC8JvX5
LllNqFdF1dreDSgbG3xUaJ5Mt12a9MgCBvGBf1PMBZ+VzB276rzQFwlqu8BxPglHwXiOtUuw52Dp
9TEm2g5zZjFBzXLT0lT+WVmH9g06lBUvMcYM02IlyUv7l980BhMrM0XTBkVhA/VQ4Ktst5jQWgoo
kT6al5K3kZ+yFWNc0ALG+nvH4sSICKkf64E6hgsfjZ5iwOmZB126Fj58D6ag3W3eScRz4Liljt4e
3gq38vaGs48S9Eis2105QCpYoeqDPksviTtmHS7SV5o9veskkyumSX7B1OTIW11Bdt8yXtcb9xBo
KG0O35JLb/R2EfHhk37gddDA0GJhHNhLALIiTQdsQrXOi6VNy0YyGKmdOwtKQnK5IL3XwAvF/MAF
MSPUh3S2mKWXv3JzGK8I3x+huUu2xMmZM4TPn1DkPwUZvRtE+3s1C4yrBaBF0SMU9fuOk6KDzPgp
Xb4C6M26JdOP8Cynafd7kUXyNLFzyKzKLfMkCiwUUNJn8xfUjvGJw1NNkeVcRwsHROuk27o30D9P
gD4KrVzCBhRKABZxWd6Rf2iHF64ligVqiFunDLWIQdO1NQE5ha+zyfYpTztl8w/1h+izz6OL81xW
e7Tyt026kNVH2LsCJOQex3VjAJATLJwwXALFiA8bpet25+1BganWfy5C7ovbJNFu4zscIfLhuDUr
4qDhoGui5PYBgHnmZM3b0EolbH/DmrSUBBv8Pbl44YgwCuYBUp/i8BwpXZXr1H/gzhh4relkHRlm
yzAS64Ddz5xwr3Xm2xvPKsp55dZRO0Td++DV8D1oFrP8dsQQ3VYkBUXuDZlci0rqPgk90DLmmbtO
9Bf/RH1AKLeLhEiG1Vt/6gDLQ24DAwaePNT+QC/OqdSmJjTb7Xm2mRtMr63eCHbnZwt6PUtCDq5k
ujG8dhJSRpdYkqVnDqVkqv6s1/Y6JNRYUQKHeGZaEyU2EBMB5xDb9n66CPRxHTemS/qINjXYgvqt
LKGNTil39x8uAjUSOwJL7PAHluZouHT3mC8zrwwokWfoTftFydUXMS3hJK/+w+tMCjwrO6G3uxkA
zyizjhJt9ckRUljez3GLVjb2NPRVgNCQCnj6bliCujP37hHcjA6rHHuxGk2V5netuZfNIK2R07SB
+hE8l7gy44DknBqAlBoHd38i1dXNm7/2qEQUv2ojQdtPeydZDozB90uBJTMpqHdVKSaq76HB9/mp
0MDA1UrFbeAmBHDq3VIBp3CcXE30k63bQeYrxFqyqZnyZ4Dbtg/lsN26sPTpIMfLGY7qsXSjeJnH
O9P6/SEbSRXjdPmN2sZ6sArT9BRv0hme0NQF4vQIsSUUF64tV2mroqYN2l1+BVSTOIWgILicFf2Q
P3zCEt4kM50OfyyHCGVAEtXk+RnIPjvEa1mQKVRydUKLOFH7O7M4NiiqJThZSLvH5CvYXGXGxH+g
hh/mHViQyCEL8FaKlSE4fF6p8Us5XRv0erZm+DZUqtjI/tbfyRX0NZO8TMBDA9sud9vVdkwzOyoh
6bqM2NE5m6yn/hZUC+eA4wRJOVAxR5ZFQBp+hYMklgMRh8siQUJOX8zMKKohlPKUR4h5nW6VXbgl
s2OblugI90ayHKYGeJCRggMDwdgHSbkgaeXxZQaTG8kv6iH2Q6/QzU1EluT0QaiYWWhx9shZv/bY
4GgWC6j4FPiv+kjDJ4yCbHh1fo3LXO2N3Yict427Yofm0GFM8l7RwP/6xMTrX8TsTR0tHQfQcrYB
mpOcPblUNVGGlsO5E93ln2iBdO838wJAHSVM/OvaoXHG8X168mgJQLfMxeql9GL0HzvvsmFRtxJj
TB1G3+cjNx6eA8KglSe2sWwJ3QFnosUFhxhYw5ORMbHdVRSfWmGEeg31QVHreWfyM9AFHTjj/ht2
+T4dhSsDT8VICTktFlYPn71ysKg+43PFDfICr+AaqACblZO74F1MKkk8MhP+1SepZzgJjuj8ent5
Z028li8xWSU5TYNpneb29DqzpD1l3/gMO1iULpog7tsMsQPLvrwE8SA4Ywl13KA8fCAq/ZGhUYpA
1ohUTw0FPDLw/VKYb3O3OX3R140+60y+/KgepM+HxrkPracBpN0OOoVba2zHoI/0+DWNZDGTeFxN
6vJoe4dUabMIpIGqZL2wdfXfOSq5kBH0T+K7BTyGiObFCsfg1ShZ6txU0XllQ28tBKDwCWr7Lq9z
q5B23uMAK80vD/h1qK9sKAv7a/A4rzcpIOGCekXad99kFG/B0oDdjVJSj1NeLW3nmJYtU7nk3m30
MPRsz4Oa9Zfoo5S1WoQ4yclw/qztcrGVFYtPfH4/FA+YNc4xKJocY3ZBlYjDfLt1ageLO4cZQ9Qq
sub1TGdi2vj1neSWAghGdPnCmLqCl0Y/A0SNc1Zhhiw6a3SiXGs24J6p2Dhv8b/TCXrpXk3TARlu
d9DM/D4uqHjnZm4NyaIyj8QSSnedYrieJQXBfG41Po0Z4rasDn/8AlAtKa81K6kw7x6gWa5DfFCh
nMVCdIu/UCILtc7m6f9SQF0b+m+WyyBRgoGfu0W81fVhqhz8hBBaZvPLhKRKnt7AjNc57VjNKR0L
h0SDDC3QC9y0lYujYyd46P7z3I8PxTPRpRu+NoI08wUU4msVEe6ocXzohnmWeAMFXM0yAyAwDArC
N++ZVRPlx8wEcPQYth3F9KNmnU6Mjo7lKtkaWKebYNiPSr3C8GS1eJonNBqZAK6dotTofmwnD6IA
DuGKComl++TXPfKwcV9AHkBPX+ITnGP88ubx7T6EoYKD4LiT52xd9RtoH2w/Whatr0QBmaaWuGva
RK8ZE6q3xz38IqVylH18DOOiozV9xTmMQFbKxEVQegpsZuKoPPS/tVyzXgSpBUjmYJuSM1Fm0mt3
DfaBT7gxU3peG4xlWQhgx4E66tsRDrsAFHwp7Y6zN81vkciocbN7ECjnTnskY7Feejf85uJjIB4Q
poh4/Q20xXnI2pZw68SaOYi9+1FKm+fjKffj4sv3sZ8WSGhv7GX9NAE6vZHfIUQ1oL5yKe/z7tE5
uhvQswskes5NXwtkrfalhwOn/Pqbbs8S3dl6piOnLogP5eBxVP0ixyc/gjjsGbtU7+sRyiLctAmD
W6/CnaBt2Uvlw86mdaS/h7lb0G+n79wHA2zeY3t7anLsfyx2srJy2qtzVwU/dnlUn0+NGYXbdx0c
VuUhEsrTCofOtmgM8pkvmi5sfzrkarYGMZOLcXkdce+NOTTv2rzuMjdT1OtZjjaDPOxoVElal+93
JfsQN7CG/GWoqTDOOW8AzHE/4MJD1ZCVgM9+nQk56QU+HARK8R+biiwwytsQsev4kF31DdI5h9cB
+YW40IQSmhNMGtaRAClCKutp1TstQjudVOMkPJmhMOrM/DyXoJnZNjrq82wQ/lpLTymrEcs/swOe
hpbTKzL/l2WL27tWyfDRztEvJsVy6eQsePnOoiAF4t8cAoEE1wCwbG3ruLF6qf7RjumwAbN+c5EK
OJQDmCcRHsJc3nhaq1wgxhLYTpYdap6pqQJgKCcHl8+bT49QfOI+jjBGrXtsOGJW/pSf1NmkArCi
E1WMFxOLTLUfSqrDP647a6VR7HqyHx4/RcyOWPjH+bhp6jC17TjSaALes16sUfsfXP0aX2BZNl8L
OVv0jSd6uFsjlpmmy4mrpQ04Nh4zW73KY4SlOZqIUme/7VgkM+2q+BeuW6zzS6gFGS2u/Nlppjbw
p7I9cOKApVmxPZ220+8fnLl+pefaZKPHjB7DbAb1z8s3hkHL0mxltUDKjzoQkP3TVYwbdoZo+R2H
E8eMCWgUFNCibxSA1Jsa3kQ6q/b18fh5lz9eIYqYxO8oizDm+P3wuTOR/axt1PUnm8rtXCdgMEPa
tk1V4aMeRMK0W6EuU3+fL6rRiAbDVQPovTs6jzt7a1Xw2U1KT8d8tm8DCulgGY0HDSeL+raeSRff
pRB3/y9bECSp7kAcIroXPX67SOygysVtkrE4bhSJDzJ9oAjaf7X58xWf8+IGHEdBBqsU5tDaoRWH
VgA/Bx7f7PKtE55rFMlISu6WIsPxn8xc4TF53p9T5x+YQb3QoQwsNE2WEpv7+vyqwtBoJz8lUSOr
EQag5BLH6JEnEHteabGRYbgu1aJIP5ouTo8xD4wL/MHRC968XlazlCNLbRJ1v4t2v1Z2WTkuZGkr
D1vCmmOEqhQD2duPIByyXlKQsqoE+CGj0Lf+oX34JwCkhyPEuBgY6al5gGvNhqcqe7gNAjO6QSoE
ldLpEDTces/dOPMZIUTKvavE3zfgpyVaqc+kfynudNirOGvd8gOjoCZi5kB/DzrvcshJLJ0DbcII
pUPovXyD1q7SG38ke5kco2rGWCBFHqdJhJMviAnmhPPbEDqvPEo+mXtLvg8uAJ20Ehuoo0As7GzR
Roy6G62Yc9NfIpaxjKGLY4N7Ey8/WAP2a8pKaYpUpRAXgIrcrPAG/RSsKwZCAzp4CjXCQt82Rjlz
51TxNzQZDgqaQUvDu6Vt6nglDfEyQ2hOXBI4QQ8DruMr+tJqkcJtl/cMT0SNvMCFKJZjdRJgpGS1
L7KQPl06FpaHx5vwiWJRQtUlR7ocIQWsAe7yyTZO8kn6Huv4FZN0D7eCfszJ7adeibGM+LkD/tvy
DBAxmAqrfzkMsxbUR4r279K5rfzU1pbw1RxWIUYRXDS/jL8WlR++kuJN/LekSRzkEhPuRQBPMH7v
Z/uvrP/camJrRcDfydHM1qjuyrViaRGzHlMGK1aCxPWHNXNPpJftmGCoEs65pudCENlkgwmCDAYw
mLC0bVuSwJbIJV/evbmDL0+0/npBnXeO5cz96SxJ3N78GPD2swBGrWTyYxl90VLeTAdUvWHg/n9/
vIwziw5zfwHmNN/eF5fRnrNoDcaVyQXsyz7Inyfwa+KHB1+4wFmmcQYbFATyVp+4pzds6yM8u1CP
/kLO+vs0lItN3SeRtjyXndTrK1QmoA7MT5fS9pNGxrU8aSy1rJqQOVysbXcTBFyDpfS2SCu4ct+s
T3cIpamNXVvEiSAyJXqW7OkOY8P8e4/EGBIjvTn2xXhPTNENdkaihF3osZJj5es8d8swXQuJ9v2L
4rrOiKSfmYAxK+Zk6GqKzDhWgNUF53SwRkeUt+FBRp362/4NDsBdHi8RmhaCMavtcybIPWZTQfAg
1yK/Ql6nhlATQ8902mG6PaBJ6E10XhifFsuWmyIz55HFTkCF8BtqgNV4kTrqrnnz5oTJoNJcfVwo
p8RweCmZ4noXBdhiUecW92n8OhcTBW9HtKgBmPfS+eX8Xn3nkWLS0sUUzP5ZaxD+MpGELyeCefMp
tUO06RqEEMJ32QvnJHW1nkMqfCD7GUEmWQruTf7Ab+cAxWj3Nh672UxR9L8S2qq37WQudwQG62S0
t/GT9uuzeXfSKRpa3ey67LNb0zsTHVRXjf2rWoI8Ri+MamZqiEakQVPRO7dItQ2+ZWL6qTDIouFz
YhPX1IxkT4gmma4FMM91DF2KzmaxcLpF9SsAjcTphx8hnfniNZQXTyIMPnqcXMDxC5bfJarq7lcO
xGFRTeemmzwXGYsfGmf9SMd4t3zlvLOKxoW5opsPOgJ25FgUxRCBRK0UKPpg4/SHA4FR4ReFQasQ
JafKfZ1tlTt39L9wIsJDmdqjlQI1Nt/RJw24FQ+oKIwzS1uMzQ9KtenwcxrC9vWInPa2k4k+r/hG
hATaZrcpcyrXP1SJUfdRqwdjrPKALA4AhXMSuCOxjYvDeyGz1TD4naH4XPg+lZOcHyZz7Y1nyfK8
MUaRndFvLuhexQyYMBL20gyS1ISHsR8Lh6rF1gh+LUTZog3t+JPo6KiaIxKmluPh9i6K3EFOnFjo
DKJO0W8aJNeFu+4MQI+4epyG+9hi7ovUulpwA1irUI4iYWC8SsKbDU7P23cB3li1g9lMbjz1m+Cu
CZUefr3jPlRmQT94MSrDmYBXWOiHkXN3S99hZjRGUJyf0fCAnr86A5ikbXYDgB7RqUsB4wNPdjwO
pVrwIBTBkEm76r8i6E+Tm633uHKntsnFeaoMoqCdWoNFJWGcTMNpi1JNN6Wdxi73FjZutbvjaKJX
XIJE8wKyBGqXqX2ROMASwkEzoCWSTgTfGHyPam8ssj1/VLauzqEKvo6BZXsDwqXfP37Dz0Qvpx8z
muokFAoEqJOveIFpTyzyQsgolm8rrlU2F4COwBOVoptGlFu3Fez31ibqIh3bgGn8qpcOBFvsdz1U
zMThEBVJ6rzYRLjOY7Ts8qaYHQbJ62mWDC419V0IwhkAIeRV2NbTHR3sFW/jQP4HBzpA+XU+Gvzc
W512t0mSFDlX2JHWtwLBma5wmD+Q/hQJavtqh4sA2KUiXXOnft5GUXaaY1/nNL3aHrSWGtY+uUHs
Bba24fyfOJahN5voACQrXWrhfsM+ukghN3XR3Y9tVopuCu9wPL9t9IdmTfbg0jWFzUztMqH8uxwF
OORstfQK1p+zNEJs9ZUpJTOlqak5H/zw6zo0a1LXfYyf1sZ9Y+eiXgAs+4hD7LZ6Jduh5OL2n4pb
1EiuVmHtOgW2L9je3sgXrqLCvVwVjR/YPhjAyw9YhYDdXwU3H+DDZ0ZyTSyL3bTMRDLOoY3j+l45
b5gBgMCCf24wYjqtkoKt4sDxvQa6sJAVobVEMepuek4TvHbiagc7vxJLp1dkYUJUE2FY0yA+4JWR
z4CUWQkv4fYDipab83Wvdqd2uHM1AjkBiF3Xt9ZNhzBYujz0/xC5IjRpMx6ZA0vqOuaTpLbziL4+
3JdszoayikWpSgPYDzFTwW6bnekTlmtucq2bjibPOhHXy80cLd+Xc+vV9ju8RXyY1J8i/M8epmON
K4oWE6sDFDTr38Cyv70AvSTaN3CJxv/8rShfoICr3j1dOFBgwI17yppKEQKkGs7D+hCHbS4XmvGI
52z4G7wMPTDSzTwQmGyo9xW3+QmvI93Uu0y7keCwWQxNniqGzPBoVy6i0ojJTOIp9tBlsJ8I9yJS
8SJZvBr5IClBgnmOUXlg27JnYNqoXpQ6IL1KOmkSpxM6QmVxDI27dVhPw+zyCNUdJFVxwrygiZbc
ghIiMJFvEMru7R/n4Tp6lJzM/maIXGDsQVhny3l7G/ZQ/BXzxCRwZ8A9vqkg57t1bl7zTUTI+mx4
5FQm36j40Sad0mBA5qkU9uTBmqU3hFZB+t0nIiZ4zJRmNHQdD0EDq36PZd4bTljeP7P48nM61tTJ
+ZUjyrwTuT8s5AbZZKtl/0eYOk7TkgNiGHHjUM6tVHTH+7XlECni9qqtJBnWsIrjqVKxQIWcvQlu
Yuk7ClA1epgT6LtrK7YocbscoVaIfeAIpyOZMbOzp9sWhh5bJSiV/jsOME3z3Whih+Gu8S21pRu8
za+TwBsvH1tKS6/qGPmRgvM+PKF/KYKe2hwfs6KTWm4NDaSye4/GpKWBWZwD8frCjo08uEKmB0du
NjRt2gf+kXYS8VYGPUauB/kvql65vY//XNDJiGAuyR4mQU7WDXNDZLJT14rDe58Kpt0sxwDOpRwu
zorhkLrkcsL7QeiXcpZktbxpIRIqHDudFwJOebxWBX02/oyT70XRRAweW3fezZTps6JvwAYafUR2
qzLsaHapyYI66y6zKLHmmuz8a832x/nwlDr5DPQaosYHpnute36Cmkgx0yIGbfU2Qv9jd4SsL22K
OIy79y6HyHvinmG4XtXC/xSN7jVuaHTuQ+BgZY4cfbcok0qaLAhJTUxj1A15/0Iqdkf3h85NICl6
KHiGOCElcTH0QFMdWl0zfVpriQhzvb3ARGZrpO0DIT02rPRvJjR+TCZYSP2bcu2Ploiyml2HXiiA
zoM6sD9muWgSsTzqvoF7iWK10IUb1ff0lBGAHLIaHKbKqainsob54RdNBX3+d2d/GvRXHP/hLJK2
k2Xd7VnRsJcx/ccEWNKTDg9R6Ksn/3qkPVQLG2tvT0ZLd/IF8EX65cT1tJezGVIwuzIzX2JkkZ2D
xVwi7+vvKioptJjIcWWorOC8Rw5KR+e1koxhvtuz9pP6K4qZnOUwQWxg2W2HFXFb03PbJQ7hnVjD
QA25jb2uYh+hruLNpeY6AUbBA9vSHm89f2pAhl88sWwaDCTUbqySIjv6Q5IxD12hFJemuldTOYGr
SOhuDObAV5cX/KEp4Rqt1a+w1EY3oXFvYK7/Qf3d9W/WHa4PNdYP2RzOSulGiK63Vw2v9UcCJWjz
rpWzrLuaZOOomY/Jvh8bbVklrMdCMOmu8Z0GVSWBODEqh/jtg28O2uPpJfXBhrktvim3D3DYXv8y
Fk+RxKrAj1L/5EiXr4fCeAJV1JhJ3b6HfkiOHZx5Uokcq/RtLD2cCG48U9QxlU0YP/pn3Hf+u05U
+T17BzadsHPHahHp2rh8SItQEo+RPNAzbrbCfVYpxX0SUOSEcD9lCyJyLXbUiaIFBmvQeAppyJ5a
Oe8Oj0yPCI0SGyx9IHnPflqgutM1LKYWue3QvQVCXTytuMce0RNN8trVWWR1uDyTcocbvUxc/g2j
t4kGposXadEDP/maqlqs0PEeyhvhS8cPapNw+alC6OlmKS7zKcQvNNCTSw4lmLS6tycEX5wE0D+i
roZsC6HwFxZOAdLhp5gplTY+ssGgjRQB9ZINEB5NhTyTuaos1VrhqGmd2HrTjaAqL09FgY7afLEK
CCTU+1jkjNsbeUae2V7xpYgG0Upa1gvZ4XetkJBJxiVPdJ1dBvHzEq/l0fmM7QIh4u8zNJrTcmDC
0LqQ/jiZPE0IRxXnWIi8k3cRd8OLDb5kUQVL4IQYaovV2ySdjsei0798T2pCzBXTtSvoq9idGR+h
rpdUCS8DqeHV4bd96WmyNPGwoAvZ4Xww8yKbHx9ImNbw/Aij1MKJHkwVzi08rQ8RrPE8YqT4R6cT
dOO+rjrpz7AiZ5jkAckTCqWwd/wArZptfbSlXqtkDsrtKmB53O3BombB+CPvakQ+68ZtAQwBQ0im
7aAcXP8ou/uu9/OX9dQBRFwUzQQeWBr/bKtPapGlEjNTuHUltQH9TZhbOCYyObpC+raDZNEsXhVK
/R/UheS59aJ+ZoxyGGgQoyouZLuJ/vbZ3EtXk9dM/yuUvtnnl5fn9lGD+0VVyS5t7N/0pH3MC4za
7PxIqqYvh4uuYQgJLlz7cEu0guqIvvzFoQi89fz0Pfz7kpqNkxuBcTOgHAJs5VFzprM6EEJDS034
0QATQutD1X+7NmF/VAGyQkInqnHlWA1n/BijIAnJ/K36itxYT8608Gq1H2a72MAx5excLOGGF/sW
Pm591Zl5GjHFDBX29MDGkJ3IJ4FkhzRG8VP8qE2WYJByPXzJj37n4BHV90pU+53qHmV2TLKu62vj
9ORyP2rLjR7rg31rMtiaV2yCBdQAdDWsMu2lACHZ3rCsl8DKPVYuuOXKCQ/9GVWuLBBsFE1XEulo
ORcrvAZPkMD5eklhEY0U+s/4JZIWREbsg7efqpFedjc/DmCqaWH8Kq6ME/k3t7M70s31crSxL5EU
Y+umvEN2aPPQZzTh014ahiaxaw+jDQEV79k1Yme0R46AJCzOh16pz/qGhVpQtFjHiRmg9XjMAi2B
b05TLkJEfkGEPzyD2m9fkwWjLGGWKBy2XamGEkhhA7ogiKcNRlLLt4pqqC5Vw29jaSjRQOL5xFJC
bJvwVCKgiwb3nn+xubfQzhH85ohCEyEBgbBEyo2NZkNbEw1v+3rroGvRdgcBCXCbX5sqRBbjTEQa
HJYeF9DwnH0UtZZJZ/tdThT22wfX/1lL8srNUPxn+MGK1dklFAoVHXtcm2fyx/GW5D/8wXYhcvqg
MQsdvqW0ulO5t7R9xxVjmhL63heDlJ2VfsDcznujmvg4T1YO3AgV4Hf+v9NJQAzOVPt7dsIcCqbv
0G4dp5D9ToxBjrF+8CZnCScXfIoXWGIzMC4J89idHLTG5LyP+/395lzybszW8bQC8VWwr/+srBuB
LvOBslb6rOozSLlL0qMXNo4APLpnjvLVfIOe6tWGpdIXYcU+4dvLQ1A7VOwK1WXWHKaB9VRmI6HR
YlqobxUaHciMX7sKtjV56YWiSLMwSm2kP2sc0Re7lR1jsVlhq3k+Qk735DhU3wP/xRqiqcpRb741
52K1bLa1W9jCsmPIhZUGeR6xM2dPPkJ6NvRlhSuqsS+Z2wuZ5ln3mZdAhKg8E5C/pWBOsiuQ9aL1
4rKyjg+HeoDr1XkxfkRe98Ac8RXjVygDqKOSbmQUo0fAfY5lWqnwygKYhDW0LAr1VWmIXDmrbuXg
uK0iGEtauIYirxKcu7vukVrKCZSnWB/kU8BKKI1qh/LKol5f7CEHsfRritmkPnOrctZi4Yon47TI
5/7ckwRwQydjTmDbmtOzRqBXkA8XQB6/28E3DUb+JVyfmMAxG1B98q3vXsReNamuC25JEnOufufK
pfRgV12EORjFtBCaABZzrrSa+HqG0zHiQahqK5EmmhnvpCDfE2J1GJ1aj7cUTlde6X/PmPwxL22O
bNGYyBFwbrxpDRHRVp12Kce0LPWJ2Mwejft9VYp0iYxotTo39Hqo5HQgr881P8gokpgYf/+sf27G
2QBd3HE999vRWUjPWxr1Ynv0KxLg9Yr6cNsfTA/IYRvjBU9Q/Gl508edcVYZTkzqcOLm9Kn/5zPE
WEt7drI9xNhGf4HbxvZ2NvTUm/BXbKlaSw3HK/EmPb94CE22S9EF6zMe3wWuTKsMqMMr+oKhawa9
5vTDMHxWqG96P/TqEnaUOSRnRe1ewqADndD3swDLAiDTF/Zx2sdJfExjMlA3B7Mtbqti9qubWrIz
J+hqIKGHhi0QjKbu8LLzhVvNrwXd+KZtGbJQiGt9v2kmhU1x6CbSOoBAT/7nyLtGcc4UN1gzyCdG
unNuFY+kv20UcMtW5q3qPDobTrM62TB+ijV2zba+ChhHQ67yRTPuxVIbQoB0TgLT8/Ta2a/D5zLK
1FmXqVumrmKCoT0y4a8QxymRh8xWhHJusw4usBYF7ylke6Di+0eTACKLqp4qkW1uVzkANd36vYEk
65+ky1C6u4gHzN/obNAMPYFRSFqTW64eXHzCMry1YuGFu3U99sxMeTRdbartmPMm5uU41qDzY0vL
AD3R9c7PXhpoI/jTrhwaIweYSmNs71DA7Jo/PCx0H6kozScknB81hz0ZOSuPIfIdIIBt+HPLSwUG
WpjtglYUumv6mIZ6EAvXfyLLDRKFxZP7dIGNzo+KDjdDafj5cqFobhFgT24HKnBcXVXLrtqR2Czm
GC2qqOL4UpqIlPBd4bhGdljlcRhOSn2ODc+RNpouCRTL59r7OQJhywC3lceqjgYETk3q3/l+LL7c
OPHo8/U10TZfYUv4utHnCzZwCGfuwUT6wdl6TCJBaHqJ9GYQz4p7wFNuvHCjLhGCeFfFlaPxoHIb
XgV7+gAc+Zqf4sS/DvC+NAPlCX26OBPwceYYxtOWHeKy4QIHeyGby1sfY72EujYzzy+dpu1GA8sj
vvRd3pQKaHVtY3Rqj6rsPyuDcG6LrCWJkvlN6C+ivheeaTqWbXHu99brlctBKcUwqyTn1Amn1OQ7
o5wNoZJjL066aNWK2DJ+0pRdF/2XDAdTEIcFjQAyltzeMFGyjx8g70TnILvCKytR1TbMnN6lr0RO
RxH/X0UAF/4oBNBamylJEXAmoF8j9iNy3ZQ2/IfG6QtWjZWQGyTrIPC7cPFqYZtCS4VWy3478gmy
wGJHwsLiVHRNdKmlnW6Y1Z2QQNDmRu/jAcPwU8m1NUxIDZproYzvDcmQCNp+94khfCeHvjVwQjBV
KfBQvNm0/GpF54TT+tUhDquipoRBb/1VoY1LUHP1KScYPj31s7D18Z1SaSVNIpVArwCUdWratWEq
ixN5k6uS7/53sXVN6DGkz3zKIPpdv8kduP9O3t52J7DINjUQh/TCcS5kJv2ERMC5TULO+umw66WI
6LMbEFZyu65zQITfkXbsjMuIYHYa/I8o786502uYl4mK1+WGS2oRQcFRL+iPL5VqeKSFy9qKvcj1
g+27/uXScd69cF4xvwsIbFDSqT06gFPy4lGL+ioGDyZMPXPl2ySjuTrBQ/SWDDkHJlVU18jFA9do
yYIEx0IidtdyWA+stU/hUHTM22DO/53m53njfY7DblXIe75AYps1+iDGWpcs49Ly0qgZVZfx4+G3
e2SwZUGAOm5NFo4mNzZdXkIaK8Q1FmFXA2jD90KIWGSfU5/krqIh+A/7v/s1cQF3hssMp/+wL8ZI
neQk0nKICg55Kxr5vqR0wkKdBNN7ln+cSEDp+0iIg1Hulpy5OD8ssLdaX5ORLBYJk5rCGZaP87DG
OlPLDT0KEkimaxYS/LsnFEh1NqhM1pfRRdVknZSNucrDUI3lN2Sk1lm4wzB8YBGDJVUJqVSAisSw
vOCtWdr1GGWyhAqhSI1oncTcrCnECdmkIDu4qqnZm+Qd740YdT6Y9Dsdp3Oj+8hGSzoXn//weleI
vwuD2oWhAxflrj7i5o9OmcIJ2O8TIartvynhcCuLgYKybe+p5uLqME/IY5UhDjbRSRt2AqtRSR9D
p7B3HPNm2hMlItYl+4g6DSMBFBgVP+z5TOKIo5BoTE56wBnzYYfrkcmZTZCnN5o2ULwEYTmlTZiL
1p31XYik7epkju9lu3TQjqS0/2hsrf9yd4SdSuOz7HRSx84Tg0h/TZ+ne6ulU2CDmepmbz0S84wZ
Udu0sdYkoDZOMAKsFVgfpqZeWLpI6tGnL/xrB6JEyz+Dw8LQBcEmZnytAlpdJLjmRxYJZbHRjYyV
nFmTwtfYnMpQpU4zJqNFO2Zvkall5C7RSSJJ2hMeG6LlxE5/2DOeVPZTH24WGMrDV1fdc1IiWPCz
gxkCpwTjIrhjwTyTVDrWXYKIKaSUfpfZHIXtXCzczDCxLASeQnSlnCt3SOA389nu4JITufY3sEDM
PPY/D1EBb6rIqb3vLLAXHR5qknmwo+Xl6nRt12ZcLm6h3hM4MMhtzXFuW1OnvOTCSKf9d5tlKqGu
lGloNiEtBkaisvvPaMP6WRCDcUxahpMadKWxGFieeatydLNY+hlSUCGbPzI+tFjOh51wrxXLy/I6
f1laZfsb+ZJOBbgGcABc9/EkvzeFbGG/CzU5Y/LpJnclVJsQk71e/LqcqKNiIONmm5oaFXOwRsbY
NG3JyUiIcBG5KbjZWAok8+Exrq0Vc0+3dYrERonjkjy6DstfRMtMwPUV+iL71K/ujJsBvWcuaDTQ
1ivaS7IJuas273R/Al79actkOj2eTHkbQ4OhAllO+cr6HlXIltH97jw/hm8RSXwNvBNgOJEDFhgb
7A9ym5+r3cMj4Uu5XoiBW40OB+0b7TZ/XQgn7/SYgIs2umT2BVid/NOjOces0TfKPFfWVmxZwx2F
MyPVuaFnAGHKaCmGHAm5G9Ek0B00OOn1A/kkvCgh99N7UuvLKIYhHs/z2YUyzggzkawpot4JLdKr
TXpGgcacXBhajl7lrWiz4BRkCV7zjPiG4kOnCI1bXxw0tgL2X57626MZdyHCm2IbSn8YyEaHhSEW
rGj6c3/gcn6WD5eopfuo+P3aGVBK4+uos0hqvWaBX6G2jV5v6GGQRoWxzeJ9rkGJGyQuiBoblKNb
bU28SYEbclvLrPrNpOfCFpOlcdCzo1vFSlV/0hDO3cmDFuWkzM0eJQjdY1KaOWNjeRxV4fN/N5/r
MQVzRDj/5oahehgVCMgFj9sEx6KrXHFFxaK0ugQ634AS+o0ZYdcKvQVFxGa8DxLBlOAI7e+heGNo
6xk2ZmXId4dS68qg3kcftyZNHbuyfqMIZVF+lnDSkiV39IFObcR3Bfm1ioNOgVNn9ypDOx9SITs4
1sERIlBbrxkDmOoo4OxtgSLewUkc6BF03WRtzH5rcvuEz9HIxbcaxu8jJUMYFcVxBl35wgOMLVTh
sDb0qttbXMFeHtT/fxLBkTzzw2QKaZWaYcpobXwRTWid2Qf9M4eifV/8ojqE9ZEknXgut9KXutgV
MiqhvilMx4n0PM3eyEZUw16jytlCey0DbgSSdNSGYY3m9ZapyD4s6eYJJDFmY6WFTBjYe5cLopsn
ss7E7L1p1ORlCApKkTXe8X1PZoZ83vgKNXbjmsD6TTh87+Pi3Gro/ir3SKZjmeQrf6P9R3nKMDRg
bQB2rUUZeG8LfI9Ddy/e4/aNUVZ9Cyc+iZIIORQCF7/wgR21/QKf1iqCJTfEVUPeM9X0g+m4n518
oyEaBB7yQJA85zFg+iOLQWKl1meqLOLHvnbsEC1H/D1GCXSYExHLtbl8EbbFuHotLHuMBdGP6JbH
dH15XLOkuGlCAeh1mwnCLAf4vwTVJGhBDXPURvqo7Ugr9bvq2Eef5/AL74DNSQIMecM0WM7VMu3p
HlAHz+t/VVao2gQRUKPqx8JOHanzPl4G+uBmEKOLHF2yqJtCcfjXWlA+P1SDi/4F/xNIeho1/eDH
2r0T6p5rpeIORojZYAn1lynTu4hcP8XUryt6Yb8gzB/+JLAB61iPjpCDIEyhE+JI4JHE0bRRWed3
tJPPDtniZEOwovLPSOAdxdBbdpITWu2xd2QXgNcDVGiv8B4KXxaohSKJ+oYfMSmMOzyx9Ff0O4g+
LxkYfjlCOLJxG3jV54ZFoS5YrOfEKXbAIkZXcDgSGOQWHTg3nqTyS+8yKHpM2YntG+M29nZIT3DP
UO8Py/ZaN41kdWR+w1Iwj/vC1RvdbWzhcGqwxeIK4EDLkNbrRkbqTjzc8hqwH6ePN9lDy1H43rzL
pHwcDjxUeYVBQXplrlrulBvxnZ5ernHWqzJ80ZFkpSiG0wjHl/YuIyG4VWQwUOHIbVgR0Oa9OCzz
LzI9JiukH7EecaVSdesYHbwpSb/iXJGbN0OdhuW/J3HVQQ3gUavotF9g5JHD9C6t5+Q/0IeLfAGd
z/flNG7korYuRawO28FHsCXQ6Pqi+ylNt3X8Q862CCCFMRP7FDkDqNSaOg/CvQJW+f0maL2s+Y73
BmpAN6ms4scvP2kp6MZdCMLpmceIuRWjjbz2PEjDAROEtqr7WIOHsIPldSNrPwAnCmTKc0QayH8Z
R5K42FmDYHyEntD2MsnGMW8D7WDrVv0UiX0MQSdU4JI2daCTOK2eydUa5wSVRXA+kabaJC67rq2g
+xWYXqjkxhYu6EyMrpJzaRi6KSgOpjDncA+PpdAfYiNuw6iPmtnfezbGX17JKnT8WXJe4sT0aJi0
wM0SnXqla6VmwjUhEOQM3TT79J53KYThuxnB2ctOGa7D8qi3Wu7tXxBqa+uM45etKbj+41Z7bRAD
T159N+DaF4i6JbF3A1cPlUpPQxGdKSQwBQh7c3xkaqcsGRm0nn75EW3CktDd/7f8qWZTK1KxEEch
2HgUomLqqN6c92bfpWmVNNHeKZnJOPjvrIe+PVaNyAAsZdFhFT4HhuR6Q8LcoQ5LR0ipAsYFy47b
rMeM8g5GtNXxP59HVGZA6RanHWLt4IKsFZZL+BrwFsgPKT7ehr2jcE7tEbbeDkMLj9nghlg6d+vz
MuPVSWvL+pEWsXK+/+Hx9CTEdpVP+PLgoDtsncxFfGFpSKyomLt6ij5JLu8pHy5OhPcIUnwDeyod
HVcg5UykEaOvkk/tx7LfC8rZshB1jmHkk05THPOpFZNCx9DZg0K3ylMHQjyud/TckSNsUcw6bw6p
YS4bJhe7StuzKEPgmi2L0K9qIYgJZsXP++nMIdfR1tLcwb9GEI3/tABskFyjAGuSmWobh7e3+qPG
vIeGYHzhf3KI62Sq/37q7fp4lVzCmC61Sr9Q2mwnVYuMIp6AaOkZ+KriZpf0OAQjTNLjOvy4BY2M
DX2XEW1+5E4hZei4zVEeuPRBdsT/OkqhbFhMch0H1he+fqE3oG7NxgPFWFwio+HMY2BGF5SKMFIb
95Dng2Qgtb4IFhEsdt0bfaduJdEuDleKNxW5eNP1BMC4fhEQp29aUP6f25CSZ9tZSquiHS0eEJFZ
HgrgW9X8GZx7xHsvY1bxThM+fkU8OU8m9UsyKUobgst12Wc+TprSr1K+xOBOtp89aI5LINe6znuf
l2BwhSo3qqi0AjXIuOb91L3hiphEuKScwVVlTY6KIn+A/CIlJZE5e0WzIgpOE49RXBkUljMulp8w
N/Lyf+0pHWecgitkXmiz93EEq7azP6XlLZ9B7KJFxoCRfyZebvUG/1LCd/+cnQTfA5scykb5Q7ui
4khFgEVsNySPy2NHMtsrvAcl1UVgPcb/oRRwKyfSM59vs2hMhT3rSPWkdGIly32H97jC53Kb2+oH
GJn5bjlUBr7QBtVunf9a2WgEy9w4SR2YGKM9I6xmS4zpBxcJFFX7u6nz/zOsW5vdEENusZwEnTfX
oJUYP2Y1V3vwXZuAAcu4D+ZbM3OgRugctK3690ztYS7DV+9Q35Q07QSkAFdFyjzCVZ0KgDUWz1Zb
kt+3VtC/adWUxLX4FIZKUJ7lQ7zVTGYSTYjrzkcyOJiGdUAq8YEaCjy/8wc2rnTui9DVFg5igI36
Bswg5mPwKtpsCbn+bSV3xY9xo9JlvWpHfYXBqsDR2t2HHtAwWu9h+uGv5T6LnusSSJfwahPWy6X0
c/uwHtdHJnPSpUSJyLqQbG4aG9kjq/oFXRrkvEw/Cw1Bi2sXu6bL+9lP//5xEg8PcyMWFszpQL1j
BJb5QQPdkWlOD1Bd6c4sUzmRCRugWlP7Es2T+f3sr2nhXQqXMBxa45xLeEUI1Y8NSXk1+az8Xb9G
aecm37fdefKZNgV6W/4ImnB35/KT0NNx0MnqDONkeOoz+OLaP8PcnDJ2ICgwEWTw8SpcufcWM0Yi
hiDnW4lbhAekZz/M9fUEkXp5prEYgObK4FX+DPR2T0cQH16v627pzj6sOQhjFWhggG6Af7j1ob7H
OZ8B435gc3SIU1E0FJnVLPeomUUxDLxdArbvLuqRi1PwxCo2pDCH2vvw50Z/dabCXt1verSKMXOk
BSnWbQjIb0zwAdJ7w3BMekVbxym4cmlI8rEfKlE0WtGZq5r0ZmlRpyFaYB5oN0Z2hcdKp2W3ctkJ
ED348IXaqAEKd2VaCcZoAzgKPRMQG/Cy/5PYSBMhavtULxiRJqoBNXB4bYbjSKmUlSvAqn2Frl8x
WT+ztNSW0FuiSPUw1yAvh+kW8Id15qe6I6D/xvY9JILLSwO9IUQnZfUh1lETprU0PVm5C+/2LOKe
9VWx3m6P206gd8lOKBuGMRVEjLJDis+oYYs6bNEWCfQYTyJZ6WxD2Y/apKjZ8SFUA7R4wug/hGAu
1xerP1Mff71DLfwsywBf4AgnmdjPTH5LzmpP+pmppFem5dBcLNPPbYkSlYGRjooHnXU0mYJUHoTc
05F9dMq/d7Lk4CSogEvaUobO1yBsf4H7MLfwdBnfhAtO3ozYkytvZzBn2awSOGinOldXH2nMQeQt
KxYwQgDrCvsReasW9trm46oR5CaF4cyjKjoGkULKM4YVPTCg0/S8bMUDIUFAx26b+N2BNU0/flJM
5kTNpBAw4wVVByra0jnQ/Uuo+SvSOUTH2Qs+T201gXINCNze+EHWRM6z23MnVbZYDuyNrTEcv7kC
oB24AtVGf7XmgOlaoeK2C+/NBeSfcLy3ZLVSR+8zHxvB8es9oyI+j4NXab17Q3P7TYGZwjbmUACt
uaLM07GIQZ5DnB80JV2WNtyb153SaWWNmvDqHTH9HF1Z/6tn7HuP1n+NebV/vT2iZa311LuO9wFj
hcyLJp2ksa1YVnRii2USB/F8rBwmOeWLRHl/zN7u3qefO71dFQUTdj9fLIgmUMLtOyp+q2q7RvPs
XmzgkVQQSOvj0AYQR/YhNwQGGf9a2ooRURsdo0zJhl1mPjCZJVxDqHsGZgMI9gCctYkaYs3ne7lx
ye20Icjo0wWhY2B1goG+gtiLab6Sg+yK7KKAn4y/3GAI60nU2a+iGE50zAaoWP7TwuWTluTJv4Qo
UNcDs9M7JWyoFLoz6rG/NGVqiRv1Lg2dG0pYogzzXhmZbDHkcI4yW+4V8N5apkZztDa1vXDvrAsQ
0yKTIKWoFy9jx04hxs0/SZshMxo+h6JN2qpcomArOvlrxMG/n6cwocE22PkxBXCjquJ9ppFajQ0C
Q0xx0wyC7gRywiMQhX1sp9ds2/v9ZrH1SaVC0F3SNoGV/286OUtABI0fHxJMG06WLLsFREnJKTnc
p5j0jgh/jkV+8lKBP9YJtzeKGJmSRNIbx0S7ooABBKsf/1eOhrEcHEcpJyw5LyJ3+OlxfnKu5HKf
vQDrtvIwc4G5ZG1TJVzzfhQxWNWa7ztyw5ljTXOz3l62Z+sx1qwerH/VL/QHfdhf7OWpL+vf9mUh
yJmfY4fpZWx7pMBY4S0MR0qesmx/uNlXaOZP3YdUdFLFEDgrfNeaZxRDb1+5MWx5f70AsC6NGWDL
GQN4iL1FNeGDx9Deo7xJv+Bi4GfIMH40raXMhqoEKu7CmnYY+Ini5/GBff6PF7MEEH88+oH6GEpl
pvr/gVlIqV7yOHN7IQdOyTsoqkbiMLH0A6hw414UKP/1TsnQoVAG9kBz1fWvbbJCbP3mbyjFu67i
DSKVrf/2NZe74rVkCyztHr/+Qkqd4Uj5ud87m8gqFQlGWvJy3w+vOJYRd8xCTv6MJRGd82bXVdOL
YGg56XQGKC4tC/HhOTfFfxY4bce9qJ+dXHNTwC4ahX7YvuSJCQeUr55nDAP9oYC6c1Vop3JpJ9GL
eiOIqm1nQTEmq1kxBvikALPJRUciwx+jh6Q0Qe7PzxcgvlQ6652NbVVbk6IG5E+Wr6gyMuM128Cq
e4L4qPzk5aSLqCjNtBqmU1x3/G+qKEQ4YnUradr/vi1zNO5QZvjqPk/VrM/6yE9rf8j0civD6CYW
TVQTq1k8kr8lQNPEZnQVE3GYhdupbiTy4N276C2QQu2EXpIK2B0nWyJeYr5sHbHyUtDy75u5QZUf
EQgfLDuOlWIokQQtgVCjKONl59zj+u8t1LBrd0PENf8yDEG6mzcywAVlvm/TCJZAmRWzR/M3nbRB
k6b6i2bqPLWP+HLL9O02tlzoy/ankrIRj0bAcaxJmvuPX5oMObycDEP009YiASMhdnKhhZYs//eV
ieaZ4mpBi+sX6B5Qcpuk07LojM4SracDKwx3GkdYx/iNwdpx6Gqxyv2VJAnBQHm+S8dHZxl/jfcK
DtDVkwcHd32mXkr28qiys3BP3HGFoh3iJIALWsdPgdI3FlkA984bcwEl7vEMc8N5AvX9iVc9bpfm
t3zd81z8Q0sXmLSSaV+6AYM6UINGiv1tWLOU4ZMfpg+qSfnYk+Tr55NVXrXPepHSDyvJEQlVZbcB
eBpsP9i96bUglpGfW4/tyLiArSXlqEWxHzEJAxbhNRCDopkcaHc51TOllvUBKPqyJ674yXn2Pqgz
zdYu+xko/07S6PARaRq7lYDu+61WX7wGLaSODJP2DF7/g/pOvMul9ODHNWia7RzYIK6UyjrnCmlr
ruIPeIq+dAvEUK8aJ0SL5v+CXrVf9yUOJOz5NIkS6a5+sWFj+SA4OWVo4zeZ01EUQNJQvdxy7oQy
6oYc5Dztw1yneZqH9qf9GOPunkV0dkC4PuXYWo8/R3IAwFERLKooDaVuK8oufqff9zrxPb71jWCE
y1WNNSJ+OlsnkaGNHEqh2c8uPuqDAQLBsadpkGnZa5uhYWRMZcwZcjiGlXRiZq6Q5ywIdwcb4eiC
lrUUP9MEj20qo+hbcTcVcMRH5sEga8zY0YWfTXnqwLOYVrt5ryh8zhPdp+DlumH70xqxTW/2WrDJ
sLyV/wogsD4NJA401fd3xWUjnXLwTpdvs+OvZWXGYjHH0pBbh4mVCLk7qzrfYTWlXLWR2VagdRO1
tUckWKes/YG2PlcUp21Z2SUVjyDZbWx8glCanbqTXhDIJYoTZxJjouidEVY/+18rmTIM5zA726sC
nZ5VJ34mbQhL7GRLwFg1kYx9ZVZAXnNETJM5LaJC+j+pCqLdqMkXV95vSlA2sRBRMx5tyVFPrdOJ
MXLCVb77VC127pbQWGgOUWG18mmplacp/t1uK6IbkjKlxtwK3DPO/myzBy3eMhCBujL7IW4z3o+5
yuJrZIcTLVV2OezytbQz3U3VpnQNKNMSeQkMda/B7DDvbba+e1xgXhcDr97V4vDfZnDMOp9jKIhg
8kk6Ks6Z284c6oBzULHwFRRTHtFN12ZdaFyi2f/qgEMWW4U8B6lwZ4zOIeO3vu3VgAcr5Ptt5o8k
7qvEdoOqlc9X0Ki/rFvHR+2ljMzeXITnEEHWF9XeFwN/9rGH/Q+plxG+4/5GqQMSqXFPNQJmB9PR
M9otL0KpjjcYJUd5vvpjFtFxeOUSOeJ4L2A+s4UzHQJjpEeO65vnaCLntgoxwiVAYkt6dzWTBKWa
rO1f00fXL6pKfR13GMutSwZF4pCWyBb3VkC1bXC7QD+3HEyAnFDvBVaa02ziMX6NAkbI4HuMmVdH
NSMMzZyh77jAd6O48KlKIbACIzG4dONeuwNsKg4FaXO5iJVyMkswgU3XqZ588y0TAsjyWa4bEpGG
WTqDh//aj3pSk4dEHVioPBwDqG3VyIfyOJ8BpAcg3GGVluXplNbEgUNbSyvocVZUyDQPi3tH4Wbc
aryfQJ80yHoX9LIY0xLEm9QgvG8I+s/tRatwEpyJgqhoLK36Y5Ym/55ipDIMS1O8RZ0KZ4HQ/+Gf
9qM8oa6EakqCejv7qUvNjnOQbs25MCvJampLD6S2s6JChepDlrg62HL9uleWGqUjPkFXeseDn+hO
tTUsu5224Fc7RmcpvujpFyy/NIWLnKIf9w+JMAV+FrJjLLqxoyGLNP6/I7D1b9tCtFwJytf5OeEr
zUXQOMiwQ/3sckq77Zo5dYgyTIjCRAjfKepKVkBdsxoIzbZu8uNh2VjNXhvmupDqDMd3lJMd5nfr
Q+PdXoLj9oxhk/eTo0owz8VcBmco9UsJuz1aLTLx8nHO1lKsQPnHTevJUAPUVzi5fZTT3qyPyvlr
xH1A4aMr2VbPA2O/bvwEhfZ/dV1RJk1oZxFCHBAkKCD3X6vG3jR2gmucP+u6eAIbR5XVCLAvSlE3
LeFErc/Ygsahqcc13/Ul6KSRID9Y5uCUvNt5lwi5sGljZcNM02BGptiyhimMbt+RbZH9KE3aO+Z7
4H9wOkf+m5670jKU3TXC6by8UUGkErpZAG0hP1BUOGgL7bwU2l0/Id5/Q3NMvWDWYjAdyxX4TjJ0
bWzY5Tb1nMp8iQJvdHTD1urqavTqkowZO7ZxmMh0p8RDPgDvvLDoMB2njVhJT+N/kN14gFykePNP
g/VTmPrnzx/tCqIK8RkYCghEQrjbK9zWlms9IXSHHspaPFONfo8gYfirlQmMf6GkSK/OqvlEtOQR
EcJGsQZ6W2zE5YXG5uXVbCQnkH0P330VxNWSlXBWrRNiIPa57EE+2/cK7EVOxlVrGn0qVjsUNsM8
AQq8Y7e50a0yAbDAIaK2DhhfV1LoHzOA5vNCBQ23+tQW53ACyjwKVXijT7OYxwdsFp1OlVfW2pnG
jOxOOs8HGpjMhfQ3Sn5XhRI1jWDIc6ObYL6Ua8CkDPi66Gn1hhMJ96eKZke8EqIRfw+p8W/D9qfn
2NJoXFtoyLAkKXa0cYOLI4qMuOq7zxbw9yagLw6yVRLWQUAlqHqHBgaPtujK0wf/bNrtD9mBRw/U
Z1ZD272pCdGxPYiwSGMtczPwjemHmeEF0N9Dt7alFVbdPE0crzk4wrETx0MbrC455lBSOMuUTQtZ
QQPHkf7m42kdCpJHVIW0z1DA6Wr81mbsyn/1oMepFzaWb9yUN5Yzm/TPOaY32jdofYNGO/0rQx+H
0W18lsFPsuKtpTF8c+g2CLl/aVra/OCrNnXweJSQdxJYcXnNQfU+IGGS9HBLWXOGJ0IuyujcsqrD
6A9z1XugAtjgW0NqOty6Zu87bOxQafLCS+wsEFJMTqPHNjF7j78C9SP7A/EkFec5jK2E4CHv7X6p
DbikGBp/SKzVues9JsiB3hd1PODOKyjiBt5XRqo4xCcnKUKDxy4BSBNUVYlQThPU8Noi0FWvc9Ki
YBuDii5kEolssd7FcICiqT4LDXBIaSwpI5753HSHlMm6Zfj/Jjs0/wq/1q+anb7qcf5MZ2zLjXHR
ZPkphtkF1VUPB8oVrG51oQjNV7YV30v7bizBFJiR/1OH+gy+nBkHAPnZwYcTQORvEd2cWtajvGnm
7GfoCwRh5k1b6CX7SEWKNVAoGaAKLL4F4xMicZa9xehmkID0uveioaGzSLJHt+fLHx8KW0xgTyEQ
Z6XpmoGOkGWZPyHI6b8YB/88N9yGmlKKa3f8M7+C4ZVtauhU36qduCcdm/4D+j/Q3lkjB4TrMycT
inYvmPlBkgyiAQrhFeSFJqFwnb1FqKZaI5e3emWWYTwpq2K8H/Ek+Nrrvo66cXgDaIA3K+h196wN
JxUrN3UmaM1KOQi3Pk/Qfy1EQBDb/D3GJZ66PP7Pk45aOnDHgYFKUOHUMbKfwbKLgUgrJlRteymJ
XXV23VaGdZHyue0BCzLzXD+troGosb0XJd15XKJu/Jy1n1iZ1uzN4s9ss7+m94FfSQt6AtVB2EIf
kImg11VJw/Zvo7RtzjRfTEMy8N/RTnPw24M5uCPCMRdSonVcP+yZKVZ71RZa40xu3EPfhu+3z92Q
B7BpQ4Yubi4sMBo4l3pOW32KrotIZrdR8KAPGHNQr81bI4yCYzwGsXpK2GjoFmlA8qqdrj8L1wk2
1c77eqwrQ1mQKIxsh/S+Eif4aa9/XpK8CRfe2Bt5mZ0G9IsDyv85mNicUTIOY8DDjR/SgykOXoQR
+/oNJBD1g3n64En2+Iohe/y6zo+MKF2sbuhS9NoBePf6SQcs+SOpVr6mvxCxJkZVqsTNP1T94Hbe
0kiQVxl7vFmxBZLwGsck2MWQRDNJh29nm+EUzCL2fL5qsCp0o/gwwMv22NHssdkzy62vjPYkqjVB
svO2gzUpCXwCQrctOARI6De8IA3lQ08LTJQ5G1/PJdIrPSgMJAwAvX8e+ctJCFD/SAz9MZ87jkOg
wKQy7NbwixGV1rOz8Hu6XZtFZFl5v+KCKCPHIDT1U3CUli6jBwGq3QorQdI2CASbxk68PDtb3gZX
o/fICimmYrgXgCO6LIUkhChSkgp3Jbmy6JLwVBE1zDspF1t0cCkz344qRE2AZBe4hn/HsjZnqRsE
RKMLziyWwtZEdJTwLCnc11r8vOEDWZPcsa8peC2lDvCh0HHS42L/cqSu2DuoA6MbN9wqta+1MQie
K6Vg316w6OH1qYxKtwHTmHEYEPp2eEhn7+a9O/AgKlr/DE/wWYgDVP+ia99l4hUOz/85Ry+BiAC/
CWoieNv9eU6FAP0jF/ZOAMgV9QfAD23hZYG3BsrzzCIS22d3HoG+X4rdtQvzT7lOCxzloXK4pMuo
4y4a+9Ajyk0OMru6Sxn5oA5Y2DgSmjSigIbDQjeRfE7MUJtKRGI1IunHUG4QveoHlW3o6czeQJPk
TJfWcnkv40YjRFB2lWatYUuQUPjY/XvoXPkvEUhT3OgH13i37Lfl2EhDIA+ko0amIZIzNN46ocx5
cD5sz5MppVbFGBdqEsfch/ZosIzfc9LHPpciNAfc+nEZMER4MhjAQCzLoJGgRaSD0WewnCENbd0X
rCxnou8Gtj1g5znLpfkVh9J/aweW/eXbDJe0WnSVlAgNDSBGpln0y6//Boy1IBF6H1EPouCPGlev
h33EdmXANVCIBYhZ2RGJIJqlJe3Dsgd5zi8X7Uir0p1R1JH3kodFua3I89VY5jD/RssKGdcBvUUO
YK30LpZkOg8vN+Ri3PMzS0dYAx/veuwWFTRtQghf9wr2itdcDPvKWrCUtVnTNvNw5lbgCYWSfEQ/
Dv6LzsmwliECjN+pE5O8D3W1QZjVpSO6FNdWskVNx2308vu0PJgM5iyi1wJ4n474F5yLHS52ENbF
UVqtN75Qimrw4pROpr0IPGEbkRJHJXFGbs7ZTdDhAMyjTbBSyi593zHk7NjLKH3foPJW19IPVZkz
chN0gZpWH2J89cPRFxKprLOoYBFpaEW+g3aDufza6vMKgZ1Nxl3OH21vyhpxVNJ8uIhrp3Zk/RvV
+mhF5Za+B17pDb9QFlOl6wi0H/zYojkqInu3twyjz6eDDDfYABo47nvck5NIzx11qFCP/MZOiM/5
W0TSeYNxDS9V5X5cAzYz5adwiDEIKTtNBppSJIr+jpbN7k0l+k24zRdyoFqC/sGDpjrJkFHYtZK8
XkzeqhLw3x5V0x/u1JX22j13KOl/2hU7yU6d9XRcJdKgVm/bfM7bRd2g7Bciw1xi9hIX1w4sMsss
t7sCHCJqg3zJB+04MCJUlGLD6ln0dogRu1p0R25WIdZwrzXE4ZSkzJOnfPXv6jLDPstAQIIRg7sw
1VuwPwUPxZGKCPIe4iEJbIU72xVSkbU2j87y5kYG39RD6GQ3OJkO1ZBvT7vvPTjbuXl60c72Vygr
hwz0HxE3vRpvkRAOsBWXgUMGHbRpmy8Malsj7/tMqSUomMM0WFCi979orkwD0JoliqDvW6QlvRbf
NyGJsWEMepxEu8zuZLx7gd0WaksIgXAQ15xn6uN+wZVJNikh0N4lu3qKGVAgmFR5NnWvPuKo0LiI
UBmiuTm0l/qkvhx74KV/ACdtJB4Nwr4cYAOMD8XSDPrS8QwvGsWtz2vReqfAPrYd2PsujvEJzpyM
xjsfWPalwA5VQeVHIG/poKgoGM5IGp3f+NlZBjfXoMxaMXIWwRgCTjFHV9iB8ht1ByWJurIV1oD0
H5T0f/k0TfafEcJufoEDijsjewSsBTBqxNan6zVDVayTF3ppkffmnFF7Cz31mkzWjNanvgdhC6KE
2xTJatrDAXcdcXbwDRRxdR+iKNFowhukYAXZ7ibDQzA1tUOzZsyIJZ5cY7xc75op8EXfis9IXjZ0
0EhF6UgM29wyc3nO+YTgtSZBR0fHJeKg3mmHUO3l+GjbiqOGI1dPSWOhEzBPMqoLZaV+WMWm4DzM
Dch860SHe72IPS3PFlgr7FvhYgHiGTYlJCh6pmwVYurSUVST+mix+hqe4LdhbvJBLgHpKrL/ZdXH
zMUgOwETHfoNQ+frFGvtp6vC4hCX9ebvEvVNMp1h0HaCAMIh/99RMOlaAnKJi7xhXMgb07a3fUv6
dPfY2TUjnOcDx62z0G2yFyI862dNOur/njr0Z2HK20huU0prSOyrlIgPxThyXZPe1DA2JbLaCfmm
cXrVR3E/HAUY3KkUAMTC6M4d49eX0dE+ZgcPl9jY2zjGOq9leyPPmDgCo6h02gvJHXt9dl6z82I4
Q3dVTglel/dIqvNhBP++bVUqCy47HagEhiA4CpyM4ihEwPgtyHNdvGAxMEpmVI7xGG+MumWGScb2
5p1Tc5mmgnUR2cdX4WikAFu4HWzi49LS+4oL0SHNoXMY+cZMDmBItjzJk57OQTo1QA/TQiNuMkVe
PZkSowpLLhYUYf4/lJpm8UC6oxBNQyhbW0R++D0KEKiGT7+0PZY/PrvxZEH3gvta3fulWuph2OD1
Aw20HOGGBMJ86VdAB/ydIUjjN/fhTYBDdYD3UEAUDbwobEdg8oT15HWWBnoAzXt4kbaHWA7kBT5+
RzAO3tBMUYL8FLb7yw54+X7QepXpwORv67N+KQnmSa5H+MRTPEXxpmBKzXdei+lRny01E8Lb/tJJ
X1vi2qDgcit9H6yBExgmKbtkZD/PPVtkq5DXttv4KztA/IsyBBca0ZffaosURbbExmEiB+JVKWv+
QW9hniNED6yuughudMvXe1IXf+lnzs+ATkb2iz86/moxEOCRho4idRdYLHaXUHcp0dLNobPWpxnP
ghFopTAjOS3NK4loPqW7QK6xvoZ3f5x+ReqUTdSNiQ49wX6m2T12G/rBFSnNB9r5Rkut9zVYIATF
csc48hmS9CQMCbsjpHkK7rME9DB+s5uCOkXZayNcRy0TZrYGwHyV1ADQSpAw7stGo4jrR3tLHKx6
bHLdz1jS23vy8SGEzqlwLsEcCYJpFEa2VDB3NHesfhOIC7AY3imxeY5scdrqg8ZUThHzLeDqnr4Y
/PESJCsKJKmnbwzcZxXrlvmlirSZO0uKuZ7B8g+Arp45iIu1Vum11ZRlHMiJEfl6DzmXVrToeFTi
oy/wFexUE4CBI4IRRKW32sgk/y7WED2DZSrCC6ucYON9VGv4dCsEazXTLio86QeLkxRfVTplnZrY
Q/K/9KHz4RR2H+JaDcAXI/4LsXnxn/uGbJ5Y8CiWInmzAIbk1Z/tQ/z88jfjzLWdNAiLycqD5Zot
LvA3XB07fZmSp9LOwQzwoM4PyGDGDEzYRHE9AnvUSNGeQ+H3+lmybTaN7RNDrGjlthNedHYmyuOy
mj2vcaMm9eMe3+HWzni0f6raH1XGaoyTXH7uuPc6/kfLQo8A3F9nNhi1NVVFd5f2UypzDq4u/HFp
P26ef9Tl9f/pXw6TY9lasY2tiXE6W1r9dh58MoSr0JwcQMfv5Ysms/Jk4OGXU71sT3tWBk/3DmAi
oHz7Fpm+gJoTJkIf+I0h3QPgQo5CcE/6bADnB5WntgUC9DIYm4TcJJLQn3ZMtETsteauyzCbr51u
ptO2T6bg7egMkKcgtywchjoApzIOBdXk9rTzTxXcZBZLSQgtzKazPDYAEz/yAWgxLOZiad1quz3S
uQlorLthB1hzh0wdk07D5Qff61nSZ2p2UiVNafh39PsmpCOG+IXqOvhZuvUZD4l8dyAyys2LAeJc
o3R5OKtwcHMQNgTQYs5kclZgln/+OjDuXvBpODK+XQsDChvrMtW9tbDGpgmdXGXf/Ni8U8+5BGuD
w5Vt14WfJie4NTRqRltVylQ1+Tl04bi/7sVv+QyUo6OaFjHZUuW5FCrQS4Tb89EZzx1TTpQ0R3/x
cVaKlSTJvEWOwZVKw3ohiuKcg5EeBVwJI20TBI6aLlZjyYMqixh0oW/wwkoFe9POHd3Bf5t6LKGJ
Qm0f0x7IaeqZhz6uhK/uY+jfuwowIs/pmPaJNDMjs7YkrBGZntSgXjGAz+dnOBe7sELmYo4ro/r2
Uyfi2sZiCxwct9mDyRXjqn5Orih1DTvYAeKeAN4GWtGZIkXbXypj8i4kdzWihIYDspf3UPpWzRYf
s2yg+4N+/PtW706X3I91E2CYEM1u0B+juk/rgveASTUwJ8ZGTCGwmqJazmKy3U7wlNUTG7ldxH4V
4b0S8X6RFNGGfvWRUhEn0+XYYDAzUj+imFS2D2Aw/no64J08iH+9jgNiEnSwfRj/vAU1YFTrR+tX
gVMHvMbOTqhrwtLrsJiEbbWW13CD2KzaiRHLP7qHj9FMJUArBxQF7jp5pswyo/TOa4coBqMFxKwi
RiCG7BrpguZi4eJ1l4bt7PjT/mfUJTEMBs2JNXX1s0tq+YTHcbpZvrb2b6zaqld5V+DUcNhv7cOc
131BI+6hbCtwHn5cwjz2Xxw1VYwriAyq9z/J6cj/xYdBu5o51zyAdXQH/E1eQA5ny3nhOlPr1aa2
x3dPtVSmNFqfwUscNtDWcztvLH0YBj4zMS8PlqUxqHnnSrIe0di77etZbdZEtgLzvds6hJYDCi1R
w5MDe36KNyizD/btAqqimg+ui3SKOaXfiXFKJp3uc13chf0sNokomo8QRw3TgsEvTrhG1nnRTPYx
ozcIetTQkTfnspepgNIbnnvmyfdcWJ5vkl2E1gR5uVRcaZ8dhPUzKfpkAejD12qMJKAPHy4Urv2i
d6DEF3u4OI24479XkOlVtKJ7V7APMCazMcoXqh7CE8BoWR50psmkWVoAHEm1o/FeTi81L8b5ASqX
cqBtEyC2aK2DgnN5g1gLmImfVovbjYHdEZWAKOHeHNqLhtJRkUDiF2nBeWwx1PGqQpEoHq/nfDrR
6mm4GE2Lr/D383pKncFGacaBd0C6Fpw+Tu4jHuxH3S1DqEUfxaCgyti7ehDjVdGaHKfwIKw7Tz3R
7G8tESdrFpStZiftQgMKpwMcN5KGE1YDj28oiDKuNSCU1+l0RGttTYCz02CXfbd/+71Xz6ap2si4
zzPzdSEvmIvRQtComtbG4EiGvJcSxNDea0k4Y+66RiF8Rn44b9jKB1k7xiqhTyFEeZEolpIBVtCa
9DY7Yh2AAf1O6jjkgt6wavBPMHa+B2Qat618GKq9kpYCPkwuB04I3Z6Q+yxWnhDNE2dUaylLSpWa
UaVUkV5N30TdqVxvNX7chWI3nT4nShKa2RQZM6BiYinlbD2Au6g6KxiK8Uk+msAiwTcs0uOmURCA
oC6//TJjKs7cbrG+KBOCJSyAqdvMCCv3JYSZ8qfZdmr/QKflVAZann5+E8gAR5wVLjvzKdz/yZs3
lH+up4qeKQE4UhWCJC78j/WUEBMV88iMZ88FGvhmVr7X3cuk2wyioFaesxAnQmwSEtZTTolYabh8
yFkyfTGaRGQO+3+zNS3+87Q2fNTxscvWC4UoTLOxGdy/6jVOiGqQJyVueetVcUYddhpZj7akPmIu
E6EmIpawKgnhN2nl+wFGQWjUJa7OmflDuOiG2Yvul3XDl8zZxJA1ZOowTEO3rSKxw2r06oEIR4RI
jjj2yYZvuJEca+mXRRRdnQI8Fax4NcfQ71E13iKuZm9/cWlsHbOLhoSMigpmz4+uHXlA/23V6Gc0
t2WFfGHt4CnlaMqPMKPqzFeE41e2OF6o06X8RybsL7sWdpgRamSpMyPP3XjbBjWuPAZo1Ut54C8t
iukCDW/1u1BreDs+Q1hMZ5ddyi2G26JurUf3vDW77kg+rHhBNep/5Ynf/lGKOB07HHKYxA6p7US3
gKa7Eaeyr+W+dKNyblFKQLDd52y5POa1nLrcVveB7X3egqKnT/jAplub4Ee8IhzhGYAJfRZ1PWB7
tpEHLIdNP2+ltfT9bTJqS8ZqxhFMod/Ur+7eqlWOfxntmnBOg3wYYPZzkLvsEmmtL6mCZHbZq3YJ
P66aBJPcUd9NhF2pnprWIUDKE5SSIGMH9t2kIF+ge4wsjBwobwIVtIR0Z2A5/JzM8mubq0S0T2Ir
Nq3uP39PyX3EmR7eK6cMwNFiw8uvJ/YudCuFeBrY4rKXUoTmFbe0HjXY6bkgc3E3nJcyhnm298JJ
cHYFnzI7yKbVFA4AnFHo+PZioC5Lw4hK8ain0kaDLmneKpS7cGZquFPct68zObH9njmeycGRRWE4
3O6b7P1xl2P73Azc1GcAaiekrsbFirHB/PdqG8ayfoEDBD3WqyIROaqy82yWZCTXbrx5ooBOIrdk
qkh7IFIGrYQ+RxBK8FopiZ8QS7lZIh7YwAjFex68//v1EdqZzzjasdfYaxWSRqOCUxZJW3k1OXlz
m9xQiAt3F0pDwzisFdE3/XzLqKuSfsSZGZclU1Xn+TYREkwp/FEFEKv+Iuhi2tDuq9cfgKJJnHXW
C2KTwRyMwlydQMxNtb2SyHxLkhkoJGqOOKzBFvtMXinQQ2REdsXrYSsNdrN+quVC7UDkURIKm205
UaEb+bmHp/TjPjwmy6kt0jBTsOZYxL4Avr9hrg22EiyaDRBpdfOM7fQ66HMpK7lPxZl35Cqt4aqP
MJeaw/pBcnTJrksmy3zDkL7ZOYk26p+ddEKLqLAV0820Kvt2nS60Z7owIN30UsA6ZmyRcqUExyyN
dBOS4jf6QrAf1ocVxw5FipTqPiQ5dlKyns2oznXOEkXvBK0xR+cvtWq6dhK2rVU1l1I3K/iezDr4
/+GMnjV65s1ZmIdlKSV64+dLGwTG2++EsEJFn3bRTmf7aangJA3gDHqloWKdZas/kHI5vSdfO2eD
gV+jjsyTNsLRw6ZndoFu9+XQgyx0aoKg/E5dAiaJPCCkjQsL3K4tan6nKDUoZZ30rHvvmOvzAuxD
g2hMVohUdcaRE9xLkEE1lChaX1GJfdt9vAAAUeY9VFjF4nAXk7J6iDkBWP8+bNgF6qqNSq0cwkHb
FVnH4M1plW85TYVkVIzg4kwQS3o++5rQYv6is/ePCg7zbc4esReIcWfGgW5m/PBv1gsVwCCGmg2E
FBa8DyzgQUtVero/aeBOaIl4yE03dmgviQcLDjGswieU0D6/HpfxXednhFrGDcZArtIHQ5HteW26
rcoCnnxa4XK6U2HiHrof2m/1eZKa63omJbqAz1FukL0WC2eAe4ESfUJVerZLiJ2NVay5VGBkA1SJ
jqv7U48OpPCMCdsiZsFwC5LTyAyKouPB5uTOJwMG0KsOdTfs/hcR/3BRmiqkMV6LhG5C3ZTdBeCK
2LfY279M49HwA3TVDpXFcKfvR23Q21xf9Kz6E/zKBKRg5kvjeF+KiiXkOTmzXxSDd8nnYyb3NiBJ
0QY4ivSI1xgRSx8Z+vJwQ0//WmAdeA80eQglS04Q0s5xfukb9bnegfXYDnwI22xIAtKksjn/AxVn
dILaRL9N25ilQcDFE6bty8aBfuHEhzFTKFbf9Hls6J/OXB/PTrZb9S1tpJznDD7wshv/0Igvq5r2
lvJh1MOFHdL6Efc3x7B1Ge0SaLG36+6WD8kKsreXCYiMYMOFFRbC1KBv9/p5ztoLuVpbWfxl5EVF
kkXTyRuF1oqIo5ECKahFwT7Vk+5hffB5I7gkCufxNFtHrZ537NO00ZSzy+IvoV0ZCD79fB3Hwhx7
+c+0WzfrufQ0cNC6ldagJyH0ZXQsi80+yiyNDoHsxVFovFV4ezXThldEO46XmvIRSChziGASLL4z
6384zlNotpSY41gn6gqIhO08Fj4yXxuFb77nSE+XG9lX7spiDzS8+xyRz2pj9s39zwmv7jv0p52F
vtNFZJwxFQE2j63yqqzqPzPhMgtCIw6b0ckMKsmncOsb0Wlo3+Dvoz3o905X8tQ3/KxW1mjYaB87
DTeizd8QXngyAduOazXccOTmApNSSOYWFTl1+xz8xEZzmYvQLJ4PQQg2brPKThvKTNjeaPxkq1St
JqIe+XhH4mhs33aiZpMnbhM7Hjcj1itoKKXeKt/wuwUqV7BmY/lkyFu2y5+RjrWE1ZN1e7jPUldb
hx5TlHq5OTGiWz/8Awsaeitesg/Jtwz4JdWAxYhBkVU818l7K5QuKGMctEyTn3CENPnrjsss2Yi+
u4YD3U/HkulPT05b9psIDkTncZQr5UU7slf5Cdjth5ryP7XHnG4Tgeac7MA7R14PpsGJ0FtN8yB/
eG1oZ/2NdWr87efREkn07qaFDJrz9Pp+CifsaaH+BZJo/oemXmrMx/fM+t5PqcPwGSceEWNNuxpi
KdoZSYwaldzV4RDgFWViHG64uwtsOzQTKsG2NrOy4v8EsHeuIzC7dQVQCOGv/cd5n+z7T8xPP8kL
EHo52T0AWh/Bn6C5zQnObdrdmLMJgZV4IldaWO8v7LoPx5255VIQTt+bEwKrSi/BOsgYpdRP20xf
fyasZgLvRkkeuDtkzyy6sneMbpawPZ+gqggU4PKwU8eCBr1e56TDtl16tFSHS7DmyxwUcTI86xio
m4Dszt+V9vNrVRZggMp1fzcKc68//gZblCLW+TXoBA6wzuRb1QNmmdVHhM/zuXAO4Ftr06r4fNIU
1QbVryPgp8+vzn0zJn+1uFkRsg1ZNiSjUizlFyCCPnQegSoMJq4RvC7uKJdmPFxIpreWva3JV+Pm
O4W76qk8Y5FbE4I35Tkntl+F1P78ve/K8GrQrvs+308nxbTuYZdWpbwShZpqZjFFA8zJltpuZdXE
/u1MAf46Iau0vfaQEFFXF3sw/rSqCCgxqw6VNRzNxVn9QoKLl2nFWx3mr90a94HZPOQ87YgaUEbl
CGOJsxm77mbRXLwzU7bqouUSOIMxIQTWDjnqfhstrAx02MW8XjJqiaQpFe0P1hfCMoA5kIczg4/Z
sZL/kPMbRrLNJHbV6YMFMe6mKNx8C0PCN3x6QI/AWCNnMQRXwKPNPsI5DMKfPpE7LRGcytrMAXxv
MMT6UJsd6hj7Z1Fbnd6jFwRSmqCJqUey8ga0tG3mnLj5KOl5q9adp4FJCiZbPz5ixxcsn2zKSj0b
Eu5G/Wnqf+sxVDQXoCw6khgwFIavm379c9DzRYDhlUsDIrdbNnM3r1WlMsqjyEoae3D9JzPL9vVG
XOLjvZioz7v16Ynw0I4nrgwSnLDqcowqhQzpqeH6RTqVLqjgqEvjf5lApQtuyOJeaXBhcfEhms3o
G0h14TNNPQ/2r6Zy5mwOKM2kkI0h5s3jOtG+BAdyj8pDf/0xRShZRUGX+hVrnjSvaTHAQKoXD0Ib
YROciGyCLAwo4XRW9McXuSmFTpyn7p8bhFOUabx42o7M366LVXYZjYSYQg6xlLciPEvlQ/9VSChT
8xts76IE3/5Tr+z5CHUpMFXy8tCQFXXhQ36+ydQlwaqLEs0NJZ7C3OzBfKU59+NZ5/pCMOBSdsKi
h6fZMadDtJWUgyPZoKkvFqaXgC17cKpyKjiHFnMvDttnW7pQuxmTKm+AmjPQrxgdnKYvCOaPxhFJ
+4cA7fYTvIFahwV0uEAu+PUen8nbiQ3RCFZC85lak0m3eLTtmRNzPMlnTF8CBgXZTPRW2b42w7on
swSeUBfZM99mGTUbi9r7NvabN2ZpZuYrjXJfppbX2p0MwiPb6QpVJPvqgSYhak9yuDrtEZc/WhKY
b/YsttPZd0oLVlLuUeWo8cN0xn8DAMRFrZOlaFoyLz/xQKLZpThoGj41WhK8U74TsRRRSzRK3cD4
RkF0qmE+v6kN86+V74qdxwswIM8bTTaWWfs/Au4mcWPVX/G1PymhwMxvnGFU21Cwi9C2W4lzdX2w
Z5oXht/J/Jxbl0agU34Gqjlvkzfnecuz5High1qFBR+tI2yYjJLKXBwx7dSw+DC2H+uWW8S6rCCA
TBYiAIUoPszKTINc1L3pgix3ULL41xZGpvFlUZNf1TT7WT3PRvP1+xRZ4Ezq6n/8kWpQItAVo1EK
H80jI1PLrVsphNRNYW/DdacIZnYfQgoupMocBmyd1IMbH549p/BemFYkzsyeFZM9GvvsDsgFKSph
XarINt5N+si8DtQ0Y/BxO307P55TVMXjQZ7Pv7/YaczOv8oNTEdwMjllHSuiRpHvHpSGhLpSTZR7
dmEUTT8NuOiyUmkSodHdsQfWTeZjV5rKoJ0daxBJcyVs4qm+zb2H24AaIP0jz4hlkKkrdHbK2Hcw
gD3UuSP1plEAMVPLIOexJo9ACULELtp+sHBRqO7rnM2cOIu96BSwZE3JY/VqswJ638TwnzlB/+R0
i+GL5gITy1cv3RAgCkG8Vu4n+Po/G4cIzMO6f69iGmzGZDEtKzbx/HqbqTgx3q+N4HBi9NIPKMAh
JIpXCgYaijWUb06X7LrYDOpbP1uJW+iSjmtRyc8CfMvLtVtimY+utrCU/cJXsyrk7ZPfybEx/8HH
HIS/q7Nc5XRiZ3i6B7G0ClkBvpR6w4gYh4nFd7ik90Y9anG4sxMk0OjovCf0NMOodN693L4Ib5Bm
Uw6UA10xkbvkJ2dNeScKt2Yrq6x4B5sZrzEseJxHvq50YhegksXImyC+E/gn8+lIpzdOs6/z3/qL
8AiYQH6tWDivZy4rEyFcxaETO0iImVnVIU2WA5K7IM9wAJmTwuOKZTWzBHn4fKNvmqMvNtbcnf56
qkbK0XBulscXhIjf0GZoY9OW0MND9l4Nwj8X9Yq879/sZHZS9uAXVIyqgUIoJtdzmuXtnq21LhDj
rJ5//jjbM2f17pwcSyqu8oceWwqX294nteFkUGIVHg7Xl4BQmfv83mo6HGoi7HHfU9XkHojwh4YY
vV9WNLylizUObsaEz8vr8RatjFe2PutOQFDhV4++ed4qQSRgCjapukeZNSbjmu5/41V+OekRTjnO
bnYq6Nuk+RapTcT5iu/MT5pVCuXRo+6rfmi+KWXpb5wdd+8HQQDbBpq4SjuPNzk1sba8MWM11XKE
fwpn+kDq4gxSUXo4aRCjNSuhICBA/0ozzRN7Pv9YsDZLjUuQ+r1bxJwdAzOaTgjVon3C5/5q4HCq
1NCvx4eGRN9aPtH0s6i6y3IWePEjwldnp7pQZfkgMnBIPVwiAKRGUMjLcPVqjWR+rCx3/GTxp55+
teifO+gMMBLqX/pLZUIr9soGHIysKupdTevbd+efLdZIzK07FjfrlvDTkgHGbTGOPboQp2ia6Dz3
qxY/gJRQCBn3CkgPXRXzgr/DdgqXCeMNNEu8vBYtN9oethlpg3LXwFQaDyTTDL/eWjmZ4bL+5MrM
ErOUxCY97cqbtQa38mQYHheTF3efoVV9rVKjrjJmEu4Ui4zlCK604lAcF+eY2zYnulNrsaE4A/4N
4y9DLuoMccwAI+i11+IB4J5v9lxtW84qFOFc/COne9YPTNPT5x53OEUTInbfvw+i+WrJlTCMCirP
Bt5mlDlPKkxT9VGcetpHZEmtNV2nAxvUbIBPoRvmHSTNsIlKQOPzzYofdiTeHMI5k+pejldv14R4
3g6sGVZ/54VsmhxQbz3Fg/CrX1bafTwh0Yn089zbxrXU/D0XMnmRNUQQ3kejnw5Wu7ld6YMKj4U4
+qF2eZn5ErE+e2ECLiKRwpSCygRQf4tirQy1VrQc56KGbbCoZ/n4nbPxHgFM4jhyGVfGvlOe69Pa
gZgQmmXoqLMLiK9/NRMkNRXVvwCXDrUkwlZLOSOF5gujVCHl6CTMmS93CAygPB7fiKPsiLbDXqLq
bNaQSUAGCpTNgdcpUKIMbxZhyPKD/ErjF24ITWdZ7aD9YzuQdIyHZWEsHOXb4OWGUDIodTV9lDYW
5iEmh8/FVjBdYXazjA6NiuWPbI+6AuqMT1a74zso8PaUNAHHKXZHFlU061LP4QsVqTQ8p0O8eFJF
7rwY56/lIDf/GBIQqsvM316I+8XvxEtNJGkiNyjw0nwpOABLkvHCqLbPy7kFTso8SL0LjX7B10RZ
EU94s65cVHSB5DTd0XwCE0yzUpfdy/W9QVBVCgmcwfIk2jfnwrlCXrpFXTNdbRbCuyJF3vfurTKk
YaSHQllldL4jrCEoeeH1wB2Ch+SOlvpaUKkZHfRtpk+I3LGiiPYBO6/6MEc6vhoctNl9NVpO5Czg
4t/1quWAY3Ucv17QTfmeRwIzbQ5vManyxxYGjLVN3bLqTje+bfNEOQusLKoKxGwYR/fyfKGqxIAk
8OFPDIXvhmDBk41F0BGykIGWPygm1ESN+vMBypRdhf6VRgYVlEqqbdbtXlYiEeUr8NTBCUh3top3
vv0HvOeANSeE0FnXAta4GuMbjxUhwv/gjYO+FlqjpoG/hEuvNH0ZrVweDcp4LoD755Ix08pkx9vT
vsWs2u+P9e2j4Qw0sfppjg5/JD1g9S8E7JP4rrdRkycL4Q3AKdTcEzheRLjuvicppmd5cfbepRGo
FbabdXhh+wwbhctHrFcGDVgiQdkVDqFB6R0rwmP0F6M6isQM1PZfUEfcpJ9VK6BHuq+ofAp94rov
Css2ifftkK+bTkgbkMtM4CcwIO6Lv4j91tCmedIbMpJ62rmTj/qkqBVLeWORPp0kjqVuGky2l20Q
t8F50Cb13+WUDSZqBpbgGh0BJh4LgkRETlceisOmf8uYY6FLlEA+YbQaY0vGAtDg5ulwfaRzBO1b
nvhB5T9bfefZXAdPpO2K9YXTM+AwRVq0Azo+lzgq52AqTjHf+reYn0WliFftZP/nifNqLACbeWB2
4UOR0uIsCrEYuyggyNaoWhjvWJddE7r3HD7l0L5THB/9oVvjoQDwKoqh6H7uOygP4cgztC4z+4AV
cBGBHGaYIlQa0jy+I6vJZrah9F5WCuJeZ2zpr5A2ZhIrb9UOZtRgmfHdFskWWrv+UTngo4toPP9+
Y7mFm8hgTu9JTMM3U4Wmqq15mbMUjuLaZv4uMd2bj5884UUgsqrjSXEIe3yegCLqPwjNnlvxUtKR
07eeDcPcPT8JfTCDttNUtXVWJtrBw9cGwtaWbMf51RWVQB9gGLC37YseDrGsB/94ifOqzFD8cYkh
vT9/ILrlxDgcPICM7bM7oGZEC9bi6zolQl78nzpEiPLzwBcLTbAsDmjh+q8TlT3UNs/WbUZodt7E
GAHOEb3it2R6yi9PLSC2uswqmrp3UGHVlOUUYvnsybpLk6MIhazBb7F65tXth2kHdPDEkVHQ/28A
61lmnW7fMw3jJLAxpntl4SPHiVgts4XxN0qJ2GQr5j+osJLcnptrCsUAYsd3V/43UlIrQUx11FaI
nXEX6p4H65AAQ96p2yAkDDk7RFyx82Rw80Jda6qtbgzhVQPTDnduJoXsuv0dEMdp2Jy0VxhZiNcr
T8B+K9RPF2I2E1M3nbvSv/3JEBwoZ0hkCr7usqZnjdMWBxY4ovkgdCIQZY9jo91wc6Ck7wPl8IaM
9Wi7WjA27owuNPihGJgdhkbXVm+7yRv3pAAsnX3OtrL8CyhzL3HEfH/2m9q0NPdhkf0ldpRZupOE
rnhkNE8iernrOsLvVrHUmGKtkFUyU7r3APaIDWjC4uwQyRuCZAKcuOhZtSPFMU/fh7tuUKeL//Ex
06l8K2156yT1t1wzCwgqIvByXMm5dkfav7Qtm7zyrpVThD3pfpHnN3fkPX/MVwO3PlydO/9IAHBp
fxHc4c4q2bDS9YaOFcZnU6P/xlrqf6Ddpioj/IpVFdxAjKb53YMRbQZ88z7LCyXhxQbFYulnj2Yh
Wr8gr7mMuZvMkHHD23LBLUfUgFpNPnOt1/qlkmiudcLEkdkOGJWoOwgR9yfk2KMKAyXQ2zfP6ynP
MN7PlBk/+FFstPO1o2Mh2gk4ZeqtDpsI79ZN4rGEiXbkhCvYGMBZCJzdUhQoArPh8cNCoCo20M2R
GEZbFjbDgDlz59n3YSKs/4xMSRKwVp0QcexhwspQcRcJqE30dnKqisvplwehhktr4Cww1UuRUF8G
IBSva+pHU/gCHzl/sA0cshFXh+3eUQdvjfSg/NQ4FsbvQx2yATIQ5WIpbIQhO7pqwM178pNjd2mp
q0w0l6tuNX6SicaeN/RbeM6XTgo7/NMao8YOxnDyi1zvD4q3IGEjjKtCOXRmgXAvjKyRdk3yS2zW
D1WHvtP8Kw/wQsD1qHZOSUdotlfK2nhlEYE5K2Ca5vJez5MkfAgLl5WQMWk2QrfXXRMpbeJAU3GN
/5jAYbLa+H1BPYceM3Q2Yx/rADwkKCXUZqNfqBNxyImhlMui1LqEceLBo9jydOh/h5ymGbS71oEW
IXkuW9mRPBd6VDMOQCQdbKuPESyo/ckOJtUQ4hOjOOmi1B7FQ5oq5zg3kylnvANSzJ0F2dA2YoZN
pAJCLZEIBj1v1EoN6WE21iy5uPY1hNFSbpS2saBlUEowIlxwWVo9dXNrSPKnhw0CjE/IUJPpuXfi
ylJD2RA+X35pO7fmQg2oLPiIP5yL2VbWwnHGg2ivtVnEjGf6UGbnJZj10hJExdOBAHhAUBgW1mqj
oK1OmRbEvr4InpLGusPNx5I5TiAgjLazZKCrmhDcaxc4z7yD/JRLYyfdg7yUva5CHOve6o7+TY4a
gvhSZ3bGHsSZvZQx/aaducYCsIgKuuYVmMO16Yr5GVi9RcXgriRNlDPlRbObeh1ge0JPTAuokNSh
lNMvBRrQt4x5kZWMAKIpJqKtA5ATiuzMJxG5AHtWiHc6kykWpbO4X+X1IWE4artCwzwraoBpmB58
obKabQsXTKXgLPVRfYwjaw8BOcTLjC8LKsxPtoUXqamQ03uVRZzFavfPa1skX8hnH/SNaW7KLxQq
c+oiRqRP4N/eksqyZ2LXva+A4eHVTbJw7rWdA9lAej0c1C6ITrjZhDgzmf/aBKUA9/X25hseNWLJ
y++RZeOf6O9BH86IfDfrkqEoQxKnG/SCrWWGUv5xYi5h+uHuoFz0JG+QjzTS56/jNJLNFJfL7jIA
NHrqTdYGd175G9F/9XVq8CB6JGmWD366M77E5+EtiZNJTNeVwFkj/KvoMW3QvQhkJcNMU+rwwnMV
Qcs9CTJONnrb7m7EBZ68QcNkVkHpwfjC3qs926yPRKXh03qrSb+C3IjK20lQ73Aqz5meNVVTCcfd
21l3JcoIhqTZUw6STkYnnDJvwRvkfC7NNInTskJsdTeWo9mlKMthDnLnpWrBQJeeExKmDrC8al+8
QxaEBSBqY7F6UAquwjsCgJUgPopC1apl2seXIkrnDWl7yjUYR3OfBcDv0AnWAuPN2Uk2QnWFCdo7
HX6J4x0Eb+iqIUzn0q5Y6CKxGKN3tAYMUeamfcRaVkjkZNt3q/Sr05fB1RJG5+ZvV37JEpKAggDr
KwUunM+GoapKwOksdpND4i0x/vpzG1nFUHGYis6sDKnTRy4Iq0OyRWU27Pb9M7+eWAwmCicWrVvs
ZCYntbn14d7CA/7YdLQsDtFO7ZkARJQzE1uNAGfimnxDLd30HeMkQ2Hioo5HyOtMLWKpmhtcXZjI
vwzunsgdesiv395JHA5Q8JC+lkvd4u2YdKsfZluCopyPS+xzS3I0P7UXi1u8FzMxphG5Gyupm3dK
RAIymMSFLl8n+q1xY46jIMu1Zu0uCSuY5rmZMxlnQKc6fBDfp/HxNGMpaBv406+/SRUc4DXmtV8l
oLE2QgemTH7gr1LTFYivgPjEKENo880lwsMLEnD9btYKAOlOxCVYMTRY7wm/VKnq4zLz0s0snc8R
QGGGD3YsETwEOv1sPz0TGbSQJweHh8jjffYF8gg6ZO4Bdw50Bvg52qcHAgzJqhOZKDYacHS8OSyQ
f4L7jOvG4/nSKQNiUyMabwQrZnLS6RTQjakXx4BAfr3G6cB+Ryi27KTVCm6WaQ29LLobE3DNDhgY
t6lZAlsmhwCvr9MCXu8nQgDJXYF5VwwJiembuFJxEE7ROjkZHGPrk5uwEQTG6eJW2Sy9I4WOY2Ju
bfw51PNoiNArpFalwb9GzPi7BtLKVOVZ0fLWSs0yJ0Tiqzc6lKmfpDEWm9S7iPlsSa9EYgJiJvVq
1NiJdHid2MJVZomjshNRQU3LzVq65VTxRU8A1b/iwVJ1J/Fv9/3XNX6Y3OCAW0gE0FJt72uFJROs
ZFxGPISbV9GeIY97KRjqNurtotWWEJV4PdlvnjTzQosKIXMPJDi4OTNtvGFe6rNFG1FKL2Ch8jT7
v7I03wYiw4xwij6MkfdQXW5t7xvJYsPuqZcKF/OGKxLIDtnuYr1bNXqVPjX6nPu0daPkP3QOfznE
iWgmAdcdOvAkxLcDV0CjZDZj93kkc5jzO7YrI9p6xxmbTnsRombMAQr0rJbrymo8cgAsnsLG+Ua6
tsIycTuigc0go1rDla4EaPhAbF8a1mynwyKm/Zmv8JoD93DokvyX4AhayjANZJEA0MeweHGCa3ut
QpEFhmq19ZwESk3ivBDh6L6OFBqSBGX733cvgTiO21dYvr79ekWdUeJCXRjD4D69wjYQYHqkCG3W
FAd2DyISFXKvbucR/oCDvuJU/FbFXOxaWUH5ILf+CoLX2t7STnUa4LhUoYEnqPzv1I2md9sTt5z0
oLrveWV2pO8S85w2buTgmjXy1oYP91Ug0GYN7xbxrqAxGrwNKkRT/I2tRoGsmAvPYO/uyDPAPUH8
GGETXnP4dvtrS0e6StirQUw1wzZ0xY8bQ1YggAKfJhza5scAuSqulFmSeCI9nrpaeKgkqxi/UHHU
NCnWXTt1/csGua+4bBqshRhb23Uozz7kTQ/IokIJBGgcsqA/sqIIGiBiaTpiaTYh4FyesO1I62sx
SPzBSQeLygWMNPxnhCYR4Z5YWTd4ot/Bhm6lv/4GMwrDf1QUe25oBQUg13WJoquyrLvFD1GEELak
1qPQAXxrwLcaGQHEZLx62XqmsyU1xXTMVVGCl9Ic4ApoXC8emRxDwjSAmW8prEt6ZJonlHMr11po
/xOvEBNnHJGxaQTWm5I9crqbVq4ru4tSza3s0lwzajUO1oAJ+9K/C9aLFccBAThNbfiN7+3cEXfw
5fTTW45U/0fI+2ZjV5zW51524t/BNdxL1qEgmwSvaV3/txXgWlb0UTC7B/9Obfm6gw3WefyXRtfl
smHYtsgYlPBdPMoF3y1vHGay2ejWLCZS0WOqftjt1jQNc2mG7OiDgcXvU/haGcdPI06ctuAnXmoY
s9bB9e9mCUXAd3F89HGdtVgglsEyncsiI1unaOEOJsl77UWhbDniUnrK69QvtFobvby3m0PlcXXz
QkJhAsaFEPpvdRG8Ahy69tdRjEvQdRLRy/Y6Qn+YQqhQzIZpNxK5adwEoFItyJ/0/+TLFcdD9gER
SE7PgSukEIWf7GZWcBaV2/fOW5cTH/yX8eMUr0LDoPvhoV+O0XcmoN0Ln+8ZCA8i6U+cLjCUPDp0
2zMHSDf8lYkm70BhgMADUNHrOEcpmzfm2iPT2HkAvrWmoVVIhIAimHrBpbP27egU7g95vV238E+V
xriKnoZTnMDVm/aR7bI7I6rlIK8LrNu6Wt5i3hfUKTyddPj48m1bAE4FJlxFe/fknbvaa/nHD0i8
CnIPjYsN1fD7q/33RWD8WfzQFEvuxKBWGoN+WfOpVuW1MuujfTlaE7sv0dUPSzKxAnU93JJa1obc
QIZQaxyhtC5UY+GzIqwukJybTcnchhp4bmmbc1F9CP2ZZWyhwd6DZ67TTQK9oskdnOiLa9kfvdlj
9pYGtNleXmzvM4A2C4HWg9b7RjgCVxCVWM5xPCyoco9uBv/hGao6EPbYBMHlFpMziCVb0O9ZxlFa
WBAxzh7YmpGIhTClOkiaquulfSa2Ys9//8oCdv5uvs1pwu3gvvUYjSJwe3dbC/E7+bTxQRT4Mw9p
PxU60+WPb4raWKY/hVhrh7mPdxQoIHA4d0ByXly/+MIcz6WNPxuMYgEagIKOaKDkygLHAM8pGFYE
nJQYmRvv36p8rBpKbBYqEmypGIKa7IwcT7smLlsIE8uyYEOeJ8CzGXnXKB2mSo4/SIC0Xo9z54rG
lI+UlPQvjjZxHSV5pqvuB86ALu8N4FQcChM/YV0QqbbeJsi6k/BxecT1BWuN4/gXcMyCTZWsNNfZ
cpuLyoCqqmyV5LsSENiCrem/jP8FibM8gTzIJSNYsR03xhH4kjQ1nM2Qf/j9qLraoPtEnPBa1pAW
igflenAo0Q54v/29tnimZaiza2Lr1danr13llePBvn8rLy3dnq1k4slp8xhsP7jDlVS28aer20sz
RQed66taYZfHairIV3jeAx8vcV+A1AWw6sFrgEFWLszu7OoxFNluLPKBNEty1gPgbQ3KrBWH0dQX
etk+890tWf67dd4WTJDdO/YmX4BcaeuGg0tGQfAx1B36LrDpdD9mlvONsyHajdentYXHmq+RxFVY
56iWiTMzG3/mykxZOkRpYogyo+OtgvmZ+DbO8lrcxTH92QBAwhuDgiSWO0XEadee7CFj2Y4Q+dCF
GUVVdeC8+1W0hYZBlEysHBbP0p3UWKMuBDbQRQ8a3hcg0d0e6AxVigB+BhR1cvha3+UrIfB08Y72
Zv+TDmHRFZ3Xv5qrCk0C04BiTJYEgOK5UFCAR9TYUbiYZF4MR2ffN7iLuL0HVwY7q0xSBumGGUuz
cizcRTVrQHTFkHNrQVmEQ0y5WLlWam4HlfC4O8yPdLPRs1Rjspv0u+MWMGr0Wg+nZwEv3V6vCZ6n
dVDhjlV3qCIuXdNhK3uYPP3/CAUq/xV3KcZz1Y15OzmBYcDdKB3jBjJb+XbzXkLtLT2cTbBVBcOf
qH81W8nznkoV/9++XuE08oO7tGw7HUZt7vd9Iz0O50h3sd0ncA6WR57AEPhxfn0+XhPe00P/eToB
WBsppt8GmBAJD5KdopDhtnIoXWVPcAQbWgH+jUHPczw3RiRCwla65QupxxSnwxrz8k06Rp9lZOnx
okFhizqAsyVE4PcJsv4KmUMOsiq2MIr+G2o1m4sn3JcOyyzysBdURFu44TAwXqhtopxwNsetMcRb
th56EmJFGC5Qtfi0qK6FP3uyhN64pdWo/H/NjkLhM3YIksKpqm92cvY2ZhNUlIips38JzCVlm06U
YlKvbrWiFIdJmYOnqfZYq7WqU07Hy3BGOVZHNXeKTQocsOewWla8wW49stIsessq+oQ8dfqp5kb8
6Yk4B8KeLOIrlcPPECEvy2tm9GPBlsvzOac/Th5IIRibC2N9n5PfQRM6EVwteQqyrcDvhJB/WMRS
k3Se+rXOfdDIb47k0tu4Wf7Auo+LELVYiBOR7JttV6uhcWgYoXNS3RsvghW3wsMrjgdFjpnDBz7H
oBvKG6NOdGTrPSkq85+hrrG2b3eVGpXADn3dr7whUsvSW9sMOOH0Z6v8C0U9Gjv/JB7Q2jlCLjhk
OY43E9Hvdz27s2N7hRMnS2EB632SQmMZO4PrUifuoWzYuR3/tRiBmJ+kbCX56G8Thug72z/gg99J
64dwwWC17UWw6axAiRBBfxfATVnkJcYj9BYEosSmV8VxUf8jPHAQg7fDv2FsS2E/qOkS8YPOywak
Z81CpaXf0sJk/sdiXJ2YNzDId13+Tx+9MGifXTly41TWPsbCAMiMFUWyXywb87lDk7p47h43nl7k
lVdP9ONfMzmFT3Q/ZlN0Ed7z7HHUnHCBdAareu5QiiP/qFTXfY1oxt/EeBLjmGCKvExqsmpoBV+o
c+vY/xncRHfUvD4qc2l90a9r4++yDFNfRoYlWjvGtKjUI+Vd0NcIKFCBhvT14Ltrx5wXH/xCem1h
wvjEg4i+GM6loc8kbSx+7C4mY3SVeJ/e1iX8wu/GmxyZilSAjRf83SPI4EQMzKyJq1rZ0fbPdgZv
1aE68GAG6dnIzedLY+iuGpFdkRL1rpF2tXW+M+tFeGf5IBM0o858DBBOWu7B2IPWa7h41cnLJKeH
uyLQFpyQ0p7vfrUxVq+jozLfkve3qlarh2oCz/r5ilNOmTc/PL3Mi4xoU54d9sLmfEZOmMlVvyMO
8lfUASBwTJV3qiCRHT2iCke+Fq7K8COxmdmYPTtlq7/DuYmz7TOzz+t5T/y/zrB3LgATvwf1aWcq
/tgCoyn2cOXUq7HTrMnOOnqjK09sQvq+ndL/eJ98IMcSvoT2Z+PBw31oc+TwLseMYYBP4a4XEVvM
adSiI85g9UcDB+M5akzPEtyq1o+Bgsz9NF3luKhwgs7kPXsJAA2AglaTERMGwGzKdUTMa8nxfAc7
ObWu1Sgxspu75vERmb2KWWbkM8o+ixCBO7A+G0fUF404eSl2X7VZwzmDjjMyDFJyk6n2/MnTMXiJ
zP1UZ1Y18dctVKj7slLbkCfw8aBc8+iKiclQZsQuZu8tsWYRuvcP0AratV9t7qqTOAyBm/bdrILg
wlndpiY6/8oxmMn+vR8uHqOahTVgyk1MXqs5mbzMJPPbpFmD5ZoGXDvK9ST9iKrmGt56nxaChApz
mv7u+uM1aX8P2wX46ND5iDEb3qZVgiEsDp6g8Z01k1BmHORA1spKLjJF+ZKjInYlcvR1SiWrBb5i
ie9Xa8FWyOnTGsPFY480Xo2BG+hDgzTf1EWBgFMiMZM7emX7jqABSHs1vYUOwejeOFBKr6OPkldw
m1HeRR+14aG0rLjRdi2qObRW6rv70Mm9DOxlnA9Gj+i+ki2iF3b4AiPKSEUUeO9tWWOSmTuDRC6m
uU12sJ3ovJNIBsKBYuZ03QxOBMuoxiGgg5jbryECpR6clYe7FuEQ6fSdp55n0eR6xrYZfKdG3ACo
npCHnUA72ZX0b94vY/E3Cf3mcfWu2mG8M/aRG3jt0brNm2O4sFZyajiORyzA1pTEGDc9tLjFM37A
F/j3A6Vzg41G01bjbtdFGeeyw54H49rYOgObWyvgBVQgZpDMh3WlqUQdt7VR9YR6xHZDOWPFpaFC
5Op1hLXDMTym1eJgACnWm0IGhVP7pVzyiKFKINey0lLfgZvTWvXMZu8OLxWqn55HWZZkLR+jWbeh
l8wshTr2cR/qxlpG9vU8YekEkGjo9BTb5ljrzq5x/0Xrd5cLV0FTgbDqLVheaYdKVKXCB2zYrURw
1SBjWpNBZb1VDQzEoaj9TQPVWT9x7zIYlfsHCZnhrSNOd0gfG9OZB8zzBLTk/+bOQD1LYSwMFt7e
S9XPN2BYKTc7uBZDlmG2P//KdnR/o9DVBiemJzWQCKkIFr3kGkQUm6yx3OAkaqL67VJizFbphhtZ
vIBG01uH+ClR685dsP2aMMrANcziD8A/oUm0ljBCd+teDIxIb2jhV+eZoOSHUie0l9Jodn2dzEAV
p4nZvtxbj2CdlkWJ+q2fyoyBnMkjy9tGb+to8f978ShYkE2Q6MVtoBCB9v8RHJgbd5tDBQyzucaw
01Di8nVx8NTVzWjbnZKWKkWd+qBJErukeNCUNKBucsGrHUD+KoNA/8QUhAmRF0BNzA9nSQugJDhJ
5pPUNP7UR0m6aS4Mc49zrBUWNECTAYxUklUXTNstR+KmrmexXGUQMDT6qcXuS0Fd81NZ6ShGql1G
UW9MQ3D9c1++tuGR1Bcsn7H2u977NRHm1LY7yE457BMt2UJEWuSZuPomBggESPOLP2eDNq+/s6rI
aHikYaISkf6JqXEhg45iroE4GNbNUMuRFCzYKLrXGV0VVoWHOcxAvbMg/H9yVpeqSiFiT5XXw4Pe
VVhywZGDRavBPym5wkwJn13X/GqgUexTADm01/irSz8Z75/uofipGtz3FB3JtzGSmmET/sOrTJwl
bU5Km1vZRUKC010iE4L9FNP9HFV+t0/JSIlBviv4gjxAEAbb534r1YuFs3ze5Hqk1y9GljHsAVQw
5e2UinAmQ0V2hRGHR/+5NqcC1rJtSafBYGQieUmjHKnhUBHwRKdMscsiOaK5hD5Of5euMScdkR/a
y40dF+x6AMjAwG3Lfgi4kJnVTu30UNZngdV+dbUJIxUt6Vy2THOlg+Ee+92WMa6OAfy+H6os85I2
Vg7Oz9B2SPKm6lZOGAwWpspb567Awwc4fCCRywVpYy9nfyLoKMIoJn00oxthamfb4usxUAElmLej
Jvmds5Sx1hSBJHPTtpssS7VRLIpMHM4/Sab8CtdJ2si2vxiiUN0H2eIxtO4eAi+29YqZfIpmT6JV
SXe5SaD4/uFayHOeGN0ItpKFKsCSgNWh+/PjfO3svQ0E/W0qO+CZkF8jRkijAU1uyk9GQfphE53b
3ay8FsFdd77ybzgGmlNHYZjNRIvNUZBVUsDA+0LbYOfZ6JG3dVFtgRP8gMzwJs65NacOmBWhOh9f
5Uvonj8zJKaDOR55r3Dd3vHPa6qVU5YfpPZxQEsQ1BLzMIq14aJUsO8AX85uVSmern2yqd5TPb92
w6eUANoFwbNJOA8mYc+KiCGZlTf511qP6BrrmUW5QcnZmtif0Exm+7OzIGmmsD1QU22ZdCkfLY5j
3hFrHA2Vsv8WFwmOqWYn3EegZzEZL7N4Gs2MvnLJTxyH8eHUBBCL+Il1T3nUEm8S+LlxJW5Q4g2Y
+kZE+1aUfTVOlqGg20Vt6qYwFZMAYuI/x0oOiWuWuzejdPMeEYArdhAOxfDI1Z2gTQ0o4cWqDoBA
bMssec8rWFWFvqgsY6xDbIagRv3USPtjZvvGTTNkRf86+TANoefeBI9EHJe1qJ570ODUiW+y8gZw
3XrS0esKaCcb433p7S+CpG8bhWWuIwxYUdUbJf+xyX/jzOpz/XBaEntNeedTZmJynm1FTtPedOor
Wv9zi5zz53v6fYcscOnhX88WjGuLzy0YNvRBINOJqWWjBonNTqrgNn1LNbbDQ6+K38yELNEjQ5HI
qkJQHqYwSmAAsGyhxun3OuVt+khacDBZG4wY+HGZQM4rKYEKXTLobpLqQ4IcgQJ2y0jVEhxRkU1b
lOT/oIg+aI2e4BHNYsPGIvNANNQJ9iY30TLjDNBL9XxknxqpBZ6ckb0OnRDeTh4j9UiNLXW8hcHZ
/4LBRlP+lDOQcMPYMCzoAznx+ZlCc7tliRsFQEZeRNqgc4jyugJXZNsRmpPDbK4Cik2Rh3jwluAX
bd6CTzEaFPaqDMrsrSHA+0+M4FK7O3sQHNMdBd3zvNgQb4t+OfeDokGBSshi0LSVBK3QF9CcPHag
oe1wTpU7/qj7h7inFpoj956Uh6hyf80uQG1xW5kaaS81aAClk5/qMUEL32f4R4u48hIIQdaWHHu3
ga5qSMcgYEm7kkND95HhZKi1+/mMczZmswWsEGPvVU4SFmTkH0hqNHUfpvR2Lt/eCIo5YbRl4mv9
40nEXPoHd52jldeYEFeLV1TNBhMTEWsvrsHuYdHZtqSqIQIA3RvqKKVzEI+A/9A5NeTYEjgPnC56
kd+Z9RsU8n1WR/+OsRSsB+4TeB0X5g+kNnwvI43nxex+ksA3kkFpMNFi3rjJ+CWqxUTxUkLciMae
W7C8wM3W+vNtSf2my+4EBssx957m3CMG03Qyuz3Huck4QlqMpF125oxYu7ZAVc/TRjuL2jze8N0d
R3Qo4371Warr+b2t4mz49Sv+AdI1FwyFTQF+hbBL3iLOg0AMChznW4f8Mk+5AvynDrAz0tjgQ6qE
ztMi+u1hE53jY9SYxRegnv232MZ5sWCvlsVUubR64kxoEicc6U0txi8Q4rY/nnv6ZaFnMqANJ2j0
Z61S6+CXi97DeJF/Ly5l9HVU1S22OEc9yt2Lje7tNZ5ocTGO06Fki7lXqIAUvhSt780MH0U6/bIP
IMsizjb8K5BkCpR3t4f4bhcgQGWsxVhi/h6L+aCXdTEPUDmQwG1AQYV3FP+k/prudtaSSzr7cp0/
BBRNmYXrC3UyyJHcyRh97sypkbyPyOgNGXl5tyVc6DKMTPlCGudxk832zUA2jSUliF3w3wiPEJAE
kQW6fs9A9r5YAbDeKKn44vdPKCch3wufTntjroJNlreF2rRfDn+9mNu2uIHAo4ACGJDhYwR9cxRo
rTY4elM0oSI3JYyqbDmWqCMiOrDT1tq/brmzVNLsxc5H2asnz0AJlg3pdyRcTNmo3GHGgxkJuPQL
gG5iE0YCaSaw7xvzcMKbz+b2lYTrOA9hVgRCocP327TO1YhF41e7i6VhgQEjxSUKua8uCaA3ZxyB
VZG+2f3vF5Voazr15jmWT+R+UwcpaNx1tOJTt9F0tY0vY8P/LUXSW12YaDDj/I9++w4xfCIRj5O1
280iQI8UTqEzc7BoaK61v2aQI30oC2RTA4bRKgQ7lgHAU24hRZCRysjamKn9Qhp2PgD67296mYnr
W6m9hhzO1gAFIc1e9WwlcnfBAURFJfX/kbeQ3+3F4YwqoJQ50kPx2AKJMf6SauDElnFVHqsAsGTJ
7khh9Jxh74poq1b71VLKG+DKqIGr5Smq9yU03OAHQ63ZqvF4nN52xvsCftyMwVsKEsV5UAmanBcj
9W+IxQxz8YVOcdjXh2A6P5QcImDg23kC0nqX4+iHM5zOHZymUsiyiwy7qY2bIkog07TIQC9TU5lX
vocvU97dmje3A0kJxUSdFQB9sJxLJoKgt7/vokDKttVHgGZ9nPO+pQOFZnzJ5vcwca4hLNie2hwH
9tdsxOcz9p2/t5LbFEOYKJ92mRMoe2ahhHn2gtEbPm99C4gOXBL5sD2QOtYDGXTNXGPQCKBowaam
dV8jaTCDDyUiw1cQHfj6SLqeOvBjAYyClqwhuSnZV6rjeHH7uTXpiNBlfjSBswFgjN3ox0oVcTFP
YGrdkvWJv5AihvVlL6PMgqXZwSvguTGkp2IEuR8sCct5yRFb2VHRbkRuqV6fwGSu2wmDqPQKwo8O
9sYlVxqZXPuKhQzeK4/8/E2Rsozu+u9UqMillPm6pwH7rwenOFLNty0HMJFTEFHR3QoyA9FrhIbN
sqg9a2aifJxsK0IbvvmKWlo0TEuqWBtSqt4vm1s+iWdxfnktrpd1vC5k+dcuIkUtDqiJoEl2JI0V
5z/VjkXa4hGNLPzjNfnhLfZb4B8YXu+v6kOFSz8T/6sPEOV1zs/4qFkAYUx2l2yuoIHQnBmmPe4k
zlL4lOAj7N2VOm5Eyo3Kr3v2zWWr5fUR94qYBa1NyvZrXCarl11glmKYrKIqdrKhG1QfChdS/HWX
0LZBM4gNLZhO4knsvDRku5ReaCv9/5q5SfXP+D4te/f2M9ZjGTK15pPoWKd2RHzlDjNnuDIiMX8y
yCqiCXWIgn02QNhR3xeWnPi6scAFA8gxhDz1CeIU31IOW0mSV2BSwN9AMFzrK/wsUh0j+Q6yoSAg
6kTEGQ5Du9+aptqceMzKoG+BU5hnLl52z70VIgw6phZY0vL+6RRcMXFEF9/QQcyjLbU+6lhWGQkn
tgUbvHActY5dmkxHltQwi09ZUDKzEHBK5QNEaz2SbtiknSjAgT1fM16asdqAI2nVnxf5uYsaSTOp
zLGyUTg5uxpyg23jOIY/hrcL/YGM1BF34vQeLSTpcQIhag+IPcipKzZnvfHYlbdUZGRoEd19i6sp
UgV7PIQXmwzPrQVqmQD5nMsDQeafg+V7Z1YAP5JlgfYaJzwRDs4QfmDgIdhtPf3eIYJ1oxqQSfgU
4wNfCxQZ9bch+wYmmimMPeG3wMww7gbbkTz4y18g9xAWeiMwS9WIaT4cWT0tfr7PlKipld7Fm797
TcDYcF4QdF1HLag66Jp7i8Mi2BGdhYBqx6xa6IM/m4LMyiJdeczqwJwxNRioDoAvfA9lxmC91/zh
PUMj0oLilDtkyWXWHEbOMixWI3omTl2wh2rpEE9ML+tfcrEZABY+vt9WXEdU4/T7zd7iCpIK4Jym
bJqwGW2HlJq+e+Zcl52R8vEK3s7AeHm90xWdib2cAD1OpPYGntDZnhZr6w/X5fVWghlu0Yfj6Zom
fQ/MaSU8ghbNz28SH0yMSOGBfFdgIvKGFQP309rD68rJ9d4ZUlmp0tsG/XFl1tfa0Rimt/OTjICL
AeesHMQjIcEe3MobMMYL3sLI2UCiuYCyepd8aWVGgKn34+LOIgcr8HrsIwMABEUfTAeQ9UoECW+l
kmq587du/QjF9d13IvYT4FtJ5O0yNlpVqeqPSOEcV3MwiWzjpNYDDQ2iTjMlp8AHpsC9DWBQs2u4
7fZFwqpjxWF9iEZYjho7Ud4m3IYrTxlg4kk1Q/4YfGCWBXA7UFvaXG4YYLSLXojaRe0YufEJK2Jx
4fAsXEwwZiSaK/heQHpwm/EP9jzT3ll+p+QFIVKjN/bqvfqfk/nk2KcSP3WQVMUyNuZRaATCqbLX
MXEXbwpzq5+l+Im6E/OkBIKH6tSNl3LysxspXA6ryT0IT+c56i+lte1J1MznNf/YODSw7EQ4XXUB
ZNKPDE7qw/fX6q8n0VTHhHwk/7UoiGPYQ3fcxgJnYter3HTV9Oxbe0Owdoz11eZ6QzLAZE7UYtIV
vc9ZlDQt05VLjpjnUPdMd474Hh9AyTtSevO4vvrLsz+hl/yvlAlcPYyac55544s/J+Vc1vpo7kto
La2CnxCqZeNM4YNL+eaB5xCCtphJANm02FoTITpFIVF+Woi18w5aJW27wkIAA1wjQqXPrj4Du04t
xGDakqw3ZOjRcVyw0OATsI1IEtI7YwW0kE+Rp+DgFEvwE2BjMW8gkDcXKYJhjMaIy1f9QyPBPFDc
8itoNGB+k77VNGcmuvKvx3nWH7kEBoV+qJIImps3fZM0B0QalZGz6UNdrE0lNVt4jjPGm08HXyh5
v/CTDrLbLg/bqLq+YY+ka70mDiv1tVrZMMa7qctCyL0WjiXdC2uWaGUrbLYQWq0CJ/PnjMxnJR5H
cpxZAUPOZIh5s28hwdp9XHuQ9lsKR6GZ1KDdlwT59nJINhI9yxS30wvInAwBdB7xEDWTn2+fbJUQ
BxboKtxWVi4fw1ry9TjxGYP0NezWo6K8UdCQmEFdZgHv47sl250yUzRLiGU9PsiBoEGTBii2lOEF
3F3nsa/GPZ6s5gr2dlMI7rrcqC5yczsfeYYO8AA86P6mzvySYbtUJ0J60xI+db4yWC1Ve9gv5eLP
hPGs6BXaREF2uX7Avdv3Iv38mjt5b+/XhApahkcKvsqeagmaTnisf+yzcnphq7NtzL493gvO5gQ7
fNnrhJ4DC60fg1eqqPYIHKZLvGoSN87HczAQemc0ZDyZRn/3ylSVMr+6KuhXLizXmEPhu4HruEav
xnAMcul7/MGBuLhHO30PMTrNKCKdOwbsu6Pu7ARrWsJxJKII1oeHT33J2odfgHhFD04WhPDoB/m6
ROyt4q4sZhwMW6NxKlauKht1g0JkVLJ48SU1ETKUX2hfimNeVJ5PoECL5daGB3QEZM1kRjbvACn0
NHVh/HJDhP8/rxgFFOIkKWRAKFdXJe1Qac+vGJyoGVY3HxXJrrj6/XQGjSpcT9U7lmSecADffr1H
yONmD0zcT/x2IIyq0+oEjixSB9gd3Wzq5td1libpJ8wXEUfCYPo/yZmQWHanShBAzpKalEXH1Mrl
nVvDInBwyEHqKJGFn9BLbA9vEqtbmVV2NaZtZaEoXRK2EQTT9fffxDrmaw0454299wSuvOuFh10l
pU8d5ix2mxxN5yT8V7AP+H+dqzBKV8R+kdFiDELmWCJ7vKv81pM5OwoKLCFe/AcMgO0aa6QZTKnC
NxP/MlGl9Ge/SwCTN++91kH7AZo+F6SGVw9ZopOLZ7E8J/E33mFvVf3JLMwrJwdUFWpKbsDMRgEQ
1jXwmzwNk1e+4REvF3Wm2TJpFxAovZLcCdAws7XjdEVqqD6hV/F4tKB0hHpIJ8v3bUYoFD2zIxh2
ofrrAXmAul6CctXVOwLOlqxcBoG+/HSDzu8zZrX00q4O46vxhKDmP2xH6Aye1TEusH5oahIavss8
6969Y73N+XFZZkWTbpUtsyoObI6W1VaaclXg896RpgyAzSJXa8f4t7ozRVVL7Ef4i1hsAEJjEeLC
rjeaZiPbRVQkThGe6LdFPTsksCNTQFa6OEqsUw/fhQVRkPVTwg8egJ4g89OY1yHlm6xTHmnxdFNa
BfqqphRtD6BOcxh4ekHUuvJ7K/L70LpAIZwyhY9U/h7Db7Ize8sb1gZ1m8Umfr/P4HnhLGBEnJ8C
dLkCN+asKt/410Q4DFJlT60PCntO9ztHM06W6J3vVoQTNKHXXiYIDjscL03HHYZDbituWAnP3xDi
kEcaMtEgHmHw6q4NzBKfUMFC2Rc6HMp16RGO9zPmJOMp2jXUaToZjGuivpXeUR8CGyB+9gHVukIk
jbzkYYqbkRbjaZY4laF2Rccufkp3HhiRg2/WapjnNpL1U+3HWnX6dZqHjR2wAgA/WrcYVDtRpgXw
Mj/glj/OEmFIvY6lRqXAgGFvlRiM3LW1i4SupzNk2SpQieb2P8tvog4ev7ZDw+UTZhY2RYb1zolo
6Uiy5wqdR4MQDLtZ99Sm6GCZV8hcjeGpbTr4VSanrxAc4ooHoNkzxzhSa9cJcLdjA2g1ciPPijOb
QjY5cZILGx9FmT9mrDh11kl67twUld8ghmZ93TZk3P2D+90XoeAhIILKqDR2VAEm8c+0MUPKBUlx
pV5dWChlVqX51suszndalEQx/BJSygtyCGdlhOTmhwR+H+Ve+gqszlEW8abr8bgHT+JLpdSNdpmr
v0tStZY5oE1kHkgb8X1TZUFMu+Y0XgzhbFxEY/cXA8GkkUd2SwZ6asca6yXumFOEpPQpZcNoeoDF
Y5FbnJEu5sG9whZ5nApshXKVsTtQP3Yhylf2KccQKWBR9E/daa8cBIiXDGIsYJwKB4h96qJ12RdJ
CP/FkL5/GNSKm1JutwF6cWZTsb1VMm0d2iY84kS2dQIliJhLmfvHive+Q57XSYFIBqGePuBCaK9+
EEcZ3welrHHx2C1o7tCqf/lDko10gk+5f+mu4tJS1g/7DhYAB6aRSMMg2tHBgYcasddb9QIEdMAQ
xSYjugDFFpOuyjZFibOlkL2jzuR04XWCvCyt1v0UluFH5WXNLkt/lkFuzP/9vX1L8/WUEsUM2fl+
GE4oGt+GVqVq+6VYGhJ7HEE798PfttUG+fckvxzT19xInX0HeWKGn5ffLz1ndhQOvGv9cqjVXEah
4BvDgaj1pwS91UBgjze+gY9yTZrqGlADj/M4kQrm9dKS/uoc2QIy04jrC8C5PGb/GDInmHXVS9QZ
OYe8NznmX19jrUiQiRAaDX84E7wOfzzVLYC38nUO3cIkSCjlAoQ6JFHHLLxX2Yspb6G7NXWBU66K
q35Aa8nBsrV9swzrIEr7FuDr2mPcMCXubCiyeh0eyL0I19PhTLWyTbR/Xq59CapySy+rH2/aI6q5
WwbEWOgOJ+Ra5qiqY1H411TqkZS7tVdaqL/nfvdD/RD9i1XbgK7HlcDs8KRxKQYy+ggE4Vd9hYsE
HGemDeksS+nhDArJLrR013yBNCJZvsnZHiWqTEKCs7YSvOy7AjoRbDUfk/JhmqVbFsT+6HuU4Sa1
25VjZC0ZTqc2MjWILiGfg1Gc9MIN3JdiA5JyTOavvv+AqYHs7wgxAbzBDL+wXdZg2oKKUOe1IoOX
gpTtC9b6HmVrr3KOAVpj71f+NW6MjMZX4CEa6XSsKHcikl8GwSQxcMjNoQJxBhc7yMf4mmEvz8lm
G64TqMLwM9PZXdf/b3nn6lLxSIS8wEIiAUfNAr+rbv0LGHWsI2j+bjDMKEk2v1pBFWpl8L1WCM6Z
xHsDN4BqEzNgkN+RHo1D3SbKahdVLyF4EqSPoKxMXcHSofsA8L0OHLhFrOJizfRs1RyDISNjzYus
biwhYwa1iHKt/U4I0in5aKCTO7ojWJExwmDbSefMyLDfvyZ0gqx/sLg7+1kX12DoMr5Ft52VgpVE
Dj5ZkMgVgFAhbiBck0VVF08fLwangvgkSEuBrfTKkJ0S1aOftpSYyaQZpMp4AgNU+H4wWwslytct
V20M04oli3rVuWbRfMpAJQ+3wQQI6dT8OZyD0oh7tIGzVdCPse70Yj7qt6mnaW14EHzeN7VRNltf
dwrrOFY8XEworVwK4IGs7mL7p59dnqhvUoP430QKSjON9Qz2d9OGcg8/FJ+joWLsVo4AZVvzbxF4
riGTsb3tMVhEtaNCxiKcELZInB7mttemohKTNFIh90p0ME3wWSjAoFauk+mSLuMq9+CcgKo4ZuBB
irhuw1Lm00MKa9Lu/PiUzu+P5ZA8YEZHaM2Ph2QhpErQzvVFctDsLIyWBj2X53yyMPMJI0gn8QmT
5pzTjTyXW5gVgk25r/8Pr1hhpaBV4DkmTNOHUbJSMv58DPtUGXTl/XndnQ1GIz/OVfaAJW4bv6Pv
qnYtxiFwQB8S8R7wODn3cx1pyHcEMgXX7BJ7YgQtzv0tmBn4ORTMS2qxvRSOTZbWBP1qyzAGacGf
r33tVKfbL6SVxngPVVBeDdvMCBPLCcQsZClDuKJkRO764O5z+dC5O+Boy9/qG+XYjLXRVc2r6aNo
7Z6+6E1y/GDUk29XM6ej2YbmAkKZ9cHsiuInR+MDlE4SlyLZryZqTW6I8V163ZufDErgDgUDI+0P
nLuVN5uDthzUdXmIy46xRjbNbLqBeudZPdE2/S+DxzrBfDPibBv261XRZAxzjH+I1mBL0v6HkgdA
3GfZ+VHeWyDUy9dwooytRTXSKvgRE6y9ihUfAby4VYNIlMhU2jVyQlaWcR+EYjUSkdZhkdNwuQo4
rsm3Qd8hLsuexsd/wt2fY2APe2RxL1W/nZZkL/ebJLGvFxb+jglFdhHGJtkUB9ynUazVus2k3N88
CMGE/oolf31K9miOhdKduwrg4d57QQNwV7y3OSZPuWaOrrcY00yfhTaGFDckdAMA8kynYq6wMzPS
ATQrA9nvYQV7LFN3E2W5FpRQ6maRBkmyA5tDGrMJ6rp54/Dg4xDPmPliN+1h8sWyt9Bksc9SfSvj
+W7QF+1CiFbJXpq2cYALVo/7KpzI4du119TiM7A4lyavQsxpffvuXUjrrg5Em7hBN1UVLKDmWUDn
rzdQdsXvBdJTP0orN+NmbqeuQ+EVgKy8dbTBfhdzcMQ96Tx+IsgZIiVMs7w33G5uLj+OE2MKu4sP
kmHP7Ag4wGMggllMXJYQFAT5m0Ty/4Ata/+KE+oXuQ/pyHmzAmy5c1Oo90PFNLnVljfQy+Sc1c5m
zDNUKNPWNowidUvK/8NPIEBr15yTtJ0A/QI6veiQkXayWZMruaWti5M+gP5L06etudb1iz7be3Te
xbJLHn1hXgYLc3mlmVNWgCkew6Ia5e3lhY6fa6eL/eb0cuavBSykGZgHJkECR3GABtsEXoJ0ttE1
3egKTuLGCNLIGPPOo/AUlnDynA9UjBfmvSpbN0Uww5Nh8y+yikzn7cx9fwl6Y9k+DT9OYqcyqiMF
HBfghbNHyPn1HhjB4okCW2sETY2IZRj9QeoPvaMO6U41QGdk2sm4Ij15GmWOTSBMkL7zo6MNwboW
EGdEePo+VOaUu0WySlzuxFGhyyTk2fay6m9yIwsybFeOtXHh083vc8ONxVQlkrSOuWIzMQzPF4jg
QWQV8RxslMw4cSjwADLiaIpJn2F0rmIVAtZUhiE/73rYOdg8NCI+V9RKQ4YR7o8amW8+ppC0omsA
O9qZVKFdjwLQ7nbFsWNGIvqGrVRrKzeee3XuuPjV/sIG7Z1GpRW/NmSDnJ7ssf5FGxQ1QWHWR43a
6FS3dlprU71nYrfOBd5eISvfWOqF5qNkMjtijHvVMX3/B9OelNdgiH6dyjITFfJc/oPsnjVxwoP7
MdU0jNm+iAS1AQo30EFw4dXO1EnHasmzfJNUaizRkiBhWXhNcXQvUI2rby6Le4ikPsqB5r4+8Qr7
ua6zP/UVET8jVH1yR83QZBehP2EIvgbDUGVnAh2eazMEKiDs3hmyru3BJuVx/uiUQ6xK5cahnQLB
OMjDaoC8rpamXGY0wkM0UTgVDTgma6f6+gCa77SbFlmdcr5Dq9iFcBNn7lImOkgCMaPd4xN0sX+1
pGaVlM2ocQp+PS+5+5FaqRFBKzi0lLSFW14Z0FOn3y7ySzu3vcWrXgE3ZtpwCyWwmb/1trMqADUO
SaifmaYN923dyrKxu4ZAAcFplPiqQcPLc0z3xxtqk9SM2MpBoCneTfBg8zXz1FrMwcyD+sp9liMz
9KX89WsQvnlaQfzmahd4BJ5y1e9TrVlf5Kl7S1aBrxW01NLdtvUYbLmNtifyvXa9Zvvb1B7BFs1d
geZcpbNnLKeJ+zqU9liwsnVZJiGmhYVVg6DhngLSoN8MXOZZHB7SI/Y0GAE4G2K0Cs7dD8ni5fUl
19Meoa/A0f2dBUKJXqTcpvmuufk2NyILMhbcFbWaqQw9xGOTI3syJrerLDoSjFMHgB3P1Iwf1Auo
LvjxtFB7v4sgsWOlW8ucg+XfLiq5+ZJN/E4Z2esWpABSihDgsIQBOPmk5pcvYzC8ido0u+94xagY
oI/1Ckc2lWNS055ENnmoIR7mPR4svGZFsv1dnE5a3hTlWWVhiFGvLBS08tFZr/rwcNcGoYprIvOn
ISIOzf83fv35iASFrmf71iazgLldqQiCoxJ5pWoI3Fm1c/ngrEghYT3iz+B/6IPJLolW5arcuQhE
tzY/Cz5HcPDwMaoVNAih/jbtNFOxZHm+yc1eG1Km6VgWO0O4Ny8PC7PwnV0Xp0qYbnnK1F/9q1Xq
9pqOB7wz9lGYc/dnt0KT0WwUXsAHqos4FVvGdU/e6AVbj3whzNbCBH6zVB/UfkWQ7VA93fo4vDaC
TDzIEp9aOCZ4HLYRhFswvo2ydLOciA8xr/XgKxm3JIiDpUsZpXeK6q3deFvlS8JsfFvismo2rkzT
Q44H4B/fqhXVV8RdcVr9PzMC+Ki7/49BaHSUNx2LKmYdTLAcE85wKUDtcJvftpXC+YQZDSpAVPuy
g2+1BNwFPeyYUFQUn1md1xVySu1JHqr9Rm9bYhDCPhr0hR99UPXresvkprzV/hh7Vqzq1/M2vWFS
1tWKnHUIQDe5CL7G4CJLB7ce1ckHwBTk9fjdLBS2Asbur099BJicZKOg6QkpjG4ivT3Gn6k2ROG+
QLRZRxI/On14J+Pd8QImJ3qZ0I6XMqPU7nyrWlXsc4xZuAeM1BBjz3KX0ph8vZ2YwaVeYWF78b8u
o4oolzm8VPUMbElqLG/qRwGGJDjZZv5RUfGWs21GOJ01OtjJBtgKoEszp8OQEgJ8PKI767CqgWLH
4V+PUTHKONgo6vhXlrYbErg/KJRngh3dv4uHfZhOCdDp3Meu9jORICGJ3dK0fIa+8HN8VR6LoOps
P8EdfBGnUfjiAjWGyp+IJdAX95IIU5BPsplROAtQECB6EXfoaQYMYFlOTalTew8P4HKUiuIR9+3G
Lfi6YSoBugTQqj1YE/eXQgtOWeuZARZiVJx+7f0stzylOH+hV9MvhvB5FE95eOq9wpKmsgFCW/Vy
zHRywMHbtf4v1TXM2hRUueqL7S21jkxkQBnBn7zarpFGP8/eiDbMZqmnbQvmheVN4k2lHmWZiIHQ
Nl0lNOuCkrYgApQtRXsGOjsXp4ZlY5O9SxrFXnC2UNqigqQGgyjeqCWBXTPr/Po5HQULgFzdMtV4
2tFtfAPUQYPJi9Tai0XcY7qwO+kRh+Hi+ve2V6tZu2+M7nUoaK4pQJRNoGP/Fs/UyLWML3Hbh7R6
pEh66KtuOAPLB+X/zk6/92ybhw0DONeQHpCdJUJ0UsHkAysutovpg2OacMwXthAtcF3MQTjwnGoN
zYp9kibqLmTqlAwsBDWaOtLngJgUFOU2kETvVL0dH/liRThyE0yJnc+Q8O5v279qmfKrD9vss++Y
0J7rypWF+/w0gEiqb3pLu7cwjohpcWl0ZygmHd/ask65vQDuvhyyl837P6e6T98QocTDdnL/Ki0k
ruH5dxMAE6aoNcctyVRljXgs4fLc+8VWih8EuPz+muzFVXBakq07lqMXsn+7kc3jTtfmKcmyM9fq
/0UeGk+wqSGIrYAF5FsXdJNxWW2YP+A+Gv+qXwWiOfVe1Q0vvobhDcWozgXhWnmTzWoXw7lX2C2V
ruqPY11fgM7+hHtkdpGxsHZpzkaKLmmrhA8GmdrDLDmdXbSX6K0K4OU0Cwus9SVWmM3Wbey9QJM1
8cDLcUGNe6psKTAs01SNuAoYKunf6OUmY7zwx7426n2BuzSWQ8tlXiACqagJIfMyZvoh/2Kla0pk
bhCMbyjbcIqfjygnwbXIHnBXZsrODv5HX1pmtma62l2yKVNDRJg64xK2MrfAgMY2Hg7bWiU6zlEK
RIHp+zybPYPKHlxvx3kDz9TSzDTI13SyCc2J2oiMKV/LLV90hFpkwKVscpl7F/m8X02AATnks8tc
qNELAwTrkQvYtZAiEWKVswRvQ3Lp+NEfy0P9vUULqWwjgrD15Y27u8ajTX+FcpFbTOAOxkyQJdF7
sUxXo90rtiJBwUrK2zPsFZ4fEH+3N5F6e9uAMwg/crZQGL3KxnhCobJ76Vj3gfQRnZ/ryXvTyMMw
2Up5G0nFZyF3W6xRc3o2B2+dtD3+JE/Cwd0kvJIL1Drh4qioNNhXfv0CDY8ITs1uTZ5NFthsiuI2
Ptu5oOhm3gp1PNIOO9Sx14hd0fAoUWch1ow8ZsA2U6LFTM03RrRaf0VATyh9zvBYyMJbu53M1/qz
Di7toDxa6KUlAwqwJVV3TWPHK4qLZZJdzPKgG1mt3RdFMEkYzjg9n7SI4uXaN2Qa6kPo/WM6X9k7
yGs0Ga2+PgPuzODtOxCCvk9Y9Z3jTgRfcfQGYZFjJpXsLsed7WtB7UwyNYP0UIW4arevzwk0zN9z
u+ND1cSYJPPRFQ0gPUHr3p4o4iuXJbuKyo/3uoA3qZQAlefnoYIS84AL2/evPhWAaLui6PrfRBWa
WStI9ZrQHn5sftq4L969PcfFnNTxBRMFxqmc3h6jKgPGqwVECd26eZDuI2Gv+6L631qViYHlOW2h
WiGCcG6QKGKYOKxFnVQbsllLbuQ+Rh4h2atgHo3ZIM9FBdPMUyzHm+rk2UIL/EfEfItV41fJuDbn
f0mEv5sYz2NgigERzrQr7muEpMkDBFMOzG8Kvhao7j6+JgpsrYWOI2xEo5wqcpa/i4onrQDUxuFB
9DDft+vFe54yg0vwOe4eFUaGVRey7jX4iWVsYXidHjb/CFsggqwaMSIUoe/WOskJRNYMsL6la8nT
GxyvNgcNdLLeZw2LnRqMlvO24BM3ne79uZIrCnGbmoHZaGNbprnjQSfDNNKiAWuHN7aGAWBIjHTo
Y1m+w2keJ5KoeXZhnQB/dAV8D32o1ZeePuFMn12uaYagrtutFXd4lF+lEB7K3Gbo1TflS+l817r+
J97V9B7BuyzwvLDoCOkfbwTJHyiV64GV12aTDh8sfic9LwIxlF/YgMS4OjoSUrKSJ+t44Hd0mHpP
fJJx0X+35bPzcwA7ML7V9wznlZIkJzG0pKS/WL7Jt+uzN3IfQQJ59WpG4LREtplzGn5LVG1o84oH
DmfZXLS239isOCRSZ52e6tBMs5N71UMzkD+WJSKgdAxiiDAST9w2RF7FUVzkfjNz5J7ZhC50AQYu
otp5Jehi6F0T2Q9RHMpvW5asImIl9ChbXMLUWQKEnHOwF3yjL+IlG7uie54tlKIoiIVNdq6HU+ct
XAyLXk9uGpD0HsRHh0QuvJWLP3H7ZPQqwECGZuaVF/Cvu7s92ZCuB7cgRskNNJFCGPDTVmOErodM
BAQw0Mdf8Q7lS0BGIv2yU2hnjDJDrro/PTrTRHvr4A3Q5gECjt4q757uTEUyP2CtaYxHoUlmJPwR
CKDm6cxSs6ncOTb2E1WfhxnjKtwK5hgjrpe8nnjZZ+n6phvDGZkGO0wI4AomU0Ap8bdf7Oz/LgpZ
ehMnu80AxKeNuBNiLoxJa9Zkda4ysrqmTrzE6qbmQfgCXVMdAG2G94VIlDpZhOWKprLVJN6IcVCE
WCxsiOl+hwFl6nhA2kZUWyCqa3daoPNT8ZN2IQ4FoFYO3OQjJvbZo2JvZKNRQffCrht0ynZrrCEX
YTbqWeDG7sTs8qzkCXCh2Gu//5TcatzVw644s0Iss45B8zq3H/HSgn+Hte4RMBRLRbDHyruu0Qsz
SAJM9Dl++6FZEGJ4MGNY8DQ7KC6j5ce9NP8mkMgy0ZE09EJ34P74JETc+KaPtHvTuTQCWqbEa3KX
Ar3ef+M1AKBf01MVr/gVgiv0qYoAdgj0Et+iwvNnRoua6fyWdXFUeBzawkZLxOVxU9y1XiiW8FLf
6bfMNp+WlZV33d5G/jigfVrnMAinivDHdz0kTxyMHM5NG52+oLYmLJixolbb5z/N2RQaCLlPYyOH
otO/8rDV1+QvV8PrVve0Am7bqETMCnislysFYOpSEK/mzP4ossbO6ccESX2JLsJaXvwVvwDBOfE8
ZcsR1RNx9SiF5i1PxFT5nBq0qk5TtbRS4hmFz41rGbPuNbiPDVA3v/d3X53EMsHe7V4EgZfJITfq
xF//1Cps08mwkl2caum31W6tf8ZG8eXduUvgDr/vfVEUXV2vQnPX56yVsP+ED0VSfpk0gX4Zl6Ze
otLQQdlvBJKVN5sCb59fO3S9UQD7P+JVoyz9u4l4GOxKz6p7jKW6JfMHcizSDTwyx8zMQjlH9NUQ
L8ACNY8OVwDMwGVkPyxW08l3FztH76tP+zxqlckJOIwyEZli+YsJL6KoxZeXhBmtMj+WeFHPpkqv
9WkVpBpIFxdMQ/ShMkuAzESmyD/6ZdWikf48rbGuWZlrRAhiIhDE/HtzbVLlzf8KyIrlbVNTOeES
/kZ0LZ3WBVGG9v1qJqAbIia6RTTAuW9/WqHVFUccCxNU4G9XRwsfgEKbwHllqsFdmDbvlHMIVXyg
csdAZxZeh23P8jOjyEqkKhcUDavLMWA9T8Hn+3rlCv4K3gmMYJPGC5gCAh2yzWY0pU3jT34xyuIf
VCavG45PegfGckBluTm74c/QeiTuZM7RI0zZf6C0cPLOKOE6q2Leyq8rhxGAut7/DIuQ++TWKhgh
yuDBgE4drECoej4z8Hu6Uhpw8w8V3KcboL/X63qeYLxDqtyu5+ohTp8M+b0hMVezqOOYdPAOcCYE
u8GYAuykEwMhwOptQejIpJ8Mp01h1g1w80TBaHKEyr9wk+mQBbZuvYwyinpGV4L9858nW1D4/tGb
9eUUU9GqcdgcmYjbJ+kYI0Wr5NJnqd1uRJWu3zwCJdzBic2hTl3am7rn7YAdBAqDdlQoiiGAttdH
aG/ya6I1zaOrFwwlKRWMqVStTnNftQXHxhLeE6mr32XKatudfL5Y8/vfQHRs5AUQWwfe8Yct9KQe
amr7sqSLgDd5om3XTt7dEv/mgyafaJYSqd8xtKgO5SEVgbXbWwfFEwCST1LtS8hDi2mihj1boWUQ
3toZ7t8K7zPSqMcG3wKqm25zokeeYF2+7bMUhfO7Ks7Dit8goW+Ok44FbjIehGZowzC8zMhqQHft
JBffAgRyMWCr5TaafelrkNWGa9YBQfOiFpqIOXbnQNOUMEhWl75GkC8OEZcR2llUaMQT0gTvNn7i
MlOjW4DRkSBPTs0yvh9iqKx9kJbz6em3KzAILt2nxFsI8gF2fDwU34HT2KAXH7hk34s+1xt/rBFm
Of1OYjvsQaPiVOWfGF4R93TjEe83YUXHLDW4mOg/pNmXl0nZ5gV+nqrcbSgGmKxsWs/H2znjBSHT
aIs1Yl229YKA0Ea1l9Bv63CYKViZCf4jHA0LDG+1USmxzG7oB61sPL4Z6ic1ZL/kRTo0IVeoPBwv
8zvLfTFdIUc3gm0di7zTaEXKJWNQqpuTs16kalaTyzm0Re+VG3yA1esdCz3D8TZZ5SAKb7tT4akS
yiBlF2fbYxIqcLISRKCU3f77a4uMqfyY+jLbzadlHq0G+cPE0SN89NADj0GxhIp21AF8J44gnHcm
Y8JUiDF0B805E8PUQs7oO+pH6Pm3st2XX+hR+wLKNqL3lueSooZDb8960y2WRKmxqRWeQJYJYndd
os/MuYNWSvtY5/bLcz99dE5Cq+FFcuhiMe+NJjogLhVKnU3vVfDYkmkaDVGamdRer2bfvzYzrNhh
r9jYkCR/lff6Y9HERhY4jVTbcYUF7TjMfEkacLxIqY2trxvZAhVCrb5SxS+A8PJpmLurKc3/2+XZ
FPcKHVMdCU8NtgPBdgRUbf6AkMucBIAG3so6aejse71IsKWf73QRVHcXQ8zB3KOX0CqlNo0SZG/R
/d2gQRkTzgpwt5jZN+wvJyUWpklaBULUGT1RP7X04G8m48svyArYzDO4FUe5jv+GStP1y6VMVhLO
SJIws9/qzqZ+aazzE4a3blOdf2nEmg7MRHqH5PUgAZfY4aDXQzYHaXflq6quctWujyN5wBmoCRdf
sFD1XnQDonJ2cIxMAXDFvsWmfD+vymni/5E7w1WXLcuhRLUoEN8LKuWFf6zfWC8XxDHbaA4BJ9Mx
nGq7xrPg7jeGKB7QNlGl+dJr1YGzn6CkVL3dspv/PtX7CHAaTPnvDJX6VELz42ZScCgbUrKOCA5A
IEj+e34j7U7xhA6CCWXtFdZ/viZgLuanmfv2ga4pmS2tCzGPEWkaQFYFKVUV6LYVJSpp3h4GI/03
llOvW6fha/d10Pre8VbOscLrc4lLeAcqWf3R8X05zxlVM3+nOC5T3PMq5lbvKKNXUMrwozpB6HeJ
DqJMymt7bG1hnHGjbqH4bqlx1pWOc3TGnzHcv0CVVwXGrHVs+zL02zVdq6TEiZsdTng2VHs13ZBe
xlPhIaEvw/vZxo7cXOYwiQvDwfdoKWok24kxFVSsiiHBZw3MQdtouC2Dz72c+o/YqOAgRN+TQ7yT
YTx2oBQsM7fzLY/t49Vh6pp1M0/ectPPyAhny8Ntkx/sOEiRMwvsD7meTdITY/9SotsXXSOwQS90
ecNEyeKnYADyhXytMCG4N98qUxcHNBp5WGZfu6auIoIG76lDhNXviEwFJbczPOPpSshzcWU26dyK
gvGjmqeNy0aYsNQT494hNlOADWZsXqe5VgtxJUpiqOIoqYAoJc9GnxN2xT4lgGElivJB6LNJlWRK
UeGkA55nVzaHRksR+Z1EFARXDBPJy9FUe97OGv7kUi6yv4Lhd8R/gc7sfIhWqUYFtbkDM3KTNRA0
XjIg4t6VEAn/iT+BxebyNwSDqyheCb60CdBc8T7Tt58fyTndZ/xSjlt4j8g3t1dyZXJF7MnpRhq2
zd4r1UL3PF6DURNGMmkK1akyNnIARK4TZeHhbFwEbf9e+ZDtgdOMwOJdgOAMsw+afX3UKlJxZs2f
wMYV9HpLEum8Z8dcYv5HKnnUzKP2ztF5l05B+hfr9aQZ56ViCZayKHcqP4B3IM5bYDvJ2ae8/8dx
LtEz5faCkCoiNlm9cVlhv7CydYv+Jxpd8Xi+RlHUzdpKqe632mc4rXmCVdtVKuwqRhTe8kFqf318
romFKmgMH1aOxVbzg5Qs3+q+3MJ9/LLixZJb4FnuBCr2LrtT8pRA0n14hMg6lC/J26x4hPyVJJLE
mG+5Nl7npsk7lkIFs/OQqHFCCt+uguiJrYBcWY0m2mU0tEEIGrsneSNGrP1J9PNSLxL8+oAx0zOR
Alv2TSIHrmxzVf9s85SC4uh6TGZUHp004AxQ0mt0yW4oQ4z3jFvtVo2wvAWLyM8RtMeTGyTS8Vwx
KCohbL3woAOB3KVJGiMCWVwS3hO5xUKOrbnYKtxI0IlVWkC82Y6TQZLMdEWkDgqfXqp3Oe6AsP+t
o6HREUgOhuz/iMWYUFbG1yjygScb9XE5hHWozAcnHxUxF2Lx2QKg26Q55cpsAj6nnrfpZh8cPaEu
stU+MyF/9GnlEwtrpgRhV1HZ9KBL4a9p0yAca6t9fAlQa30Y1m2Ngyvw9+ljivM3HbS3r+pOYUf5
gFAQMOV8OFvPaWkGcE27jfffOrUliqZ+QG2Opa0GR2mVVcVwDp+CkywD7HheEYIyXKQL4ikScOMZ
Zhigcu1wWdYxMd35WoMGkICh3xsRD9/ouS8+Ge71ro3H65Eyw6QMQIVhlZ8GDBOQs5pId34kPfyi
Z18yY/aaSq6NF0bETFcpdpuOfNoYiCojN9o8C9g1mTc14tVd3NvYYROJO3X11LBztNOKPOxexriA
CYkat1SFg3eboC6sozlHNv7itMNMlJcHiRRifTA59vZUx5nC42y9YiWe2O9Y3fh0WNrytnf4Kg7p
SUJd3nanjY7AMWnUXl7kSkm9n1kQPmTKzuVtGlKyey2KpFyvkhUAxpBMbH+lgcGpSZpGuy02xh2W
9RpXfYZb65Oqg8BnBdv0V5w5Xhn7/Q0QSPiJIZRF8l+0CPoVSvUmBkLeiHhcAVthD/6ncrAtU3PZ
Cm2necnQDEumYj3qBG9OI4Zy2lCk6jeyPCY9eQlJR3lFCgEbE/n7onhLR18cSGveLggV02UtMVWb
xfHVfmeDyKm5nxJxHJymQT69zPiCRZai3BqDlAg7sqwNe7dozp3U5qlQdRJD4LQzGdHLisjZ+vMW
mzbhnWs/Ax4yuLklAdOxEFstHmxpa/gdrq8x3EN/373iwFBKbyx7fQOe3GMJYpgSNWTDL5FoQLu2
f1cIstUOUvBHcBsZbTGHLDWBc23O5nTp3rsyeiC/h1i/7yNOsAFR7zvVr48dmPXriqwZ32tT2J8T
VL6BfSNBhIK2brXcPmFlXZSBNany0MEl6II2M7TjTtNv8rPPdsLTu7tsR/h1LFshR10sb914RtAv
paOhgH5rHEHkyf+CWq7fJfUD8fnWlJJ5f3zWSB2ikGBEnFI3QTYIa/R90Hi2btVaGBG316CoSBCe
gqnvlN7Ok6biFSSlCh0y6nDuoajwFn3gjjEJ/bLhjzhcLW2n6+PzaMnTDH88nLzdAF0k/HTOUEWE
LCLbheddsQaAFsmSLr/OpD9Iy0csHKEn0MFI6pdjvoq2nwqTa26VnIG3XrTNpDZ24zvEF0j7eXNM
2t/b9F4XJiWrg+q7x+x4SruPABG1/aJoPIQI7zazeWCWbCxXayIyhScLfht2Jhb3Z1jEdJzc/yr6
toPEkASGyUdnteJNNPSKrJuWVtH+4Ps4H1YN1BSRvvrIN69JrhLT7d1p2ajTfNm2FKttmu8fArDo
SBRpt0kifuHYoSjTQKKf644Gi4F/1aCqEsBmUa9GKJORyDbmMZE6HgUNtKZy/h0eSZfhKSkhixIv
uzsCnoQVkCMZaQv1giHrVmydktLrp01Bkx2AvuoKWhsRMf685BrFuTxUaxGZK8Dfp6Lbfy6j6nyP
TwzF85a0hH+z8U+Fdi+bq+7C5CMXZuDk4EbIlS6cSVPwKTsO2epAiCsM+++tqa3TZ8OfSCBO3J+O
yItwIeZaM9BkdZvb0L0o07H3yC4xcPv98zWeMYHwyd05C7z72dWRMAu797e2U0aKBEwPasUVhJ8u
EIEIk5XjjeOkqBUgx/dSJ18or0sYhphmThMAEbCNnHJqvB3zdIRb5x0nftoBQLo5VMUk2JFNImMw
ZgC+54+gsHVicvrIAN9+bTh6UQhYtYEXEPCCUCxjOhBOAVu5j1tTck6cr+x6pv3+PiVywCtjamZ6
dqLqeXw9qu0D3gmPmPwV3NHPOzN8FnIqwTVjWfxMMjjzgokGN6/4W5EUvhqUWP/CjAPfGFX9/afQ
bTUIGU9ESIpxeMMJrEmyASqfixMI0a6SsfnW9JSQMdxh/7/UJiKfSAVCKRt8AFBLMZ1/y9rCLgCN
1zLrndA4FgYHv5L3Z/wbnXB1/EUdb0kGQcDmyLW0N4vh5XB5pcXpAuydi9tfZkhARPBaTWP7FjGU
RvDpkiZqT+8psvZDq7rzN/YJ0XFcTZclV6GiK/W6RWft+3euQNSU1jc3zlj6aYCBbTdvlFkGwQg+
An/BxJcuunwXXDKj9qhfQSw4rVv2soOvsGugXJF/Y/pcom31gKpp9jQrPyr8Tp32EsqL7JFHYDWw
Ap/CsTffFJbPzCPB8og6nx1E87LHGocoqYTo0Ki6YHeJAPQHs7nbh3snoXOX852t0DtvgbcWaM90
hWMqdvXQQOFArHmQsmoC/N/LXOYttvgmzhYrus17avPnjLPp/mqzZzh4Sx3m3Bc9lDRab6MrznPh
qKOiBLO+ZF3fTWLmzTKmhgKo9FLkV+1uwlCCnnDUxBQ9dWezt6Y7B1eMwSEjU27g4+Kk1swJ5IA6
jsb1uEQ3yuM+3yPjdPh9SaJTxlZxUbYKC7mHz4D9WEsTntrAa2z7gc+md/P7mlvYNSCy/QEgDqyo
F0/2eStSAaO8z+vvEF/ZCmOk4i38h4n3qg7Lnnvi8jqEE8WuQ89vLUOh/8RO8V6cUSTFQ1f/81/3
vh0KFy0PnN7uTR13zBxwq7W90Q72QWThGZyZC6QrUXoak/PEJ+vR0S14CGXpvytGRsT59850FfJP
8QEKaGfUxZur1p8/oArUJfYBACziRQR6FkPZ9yWsODYDP1pob5Q9/KtQf8DlJDGfrQjY2o7rdIj+
T/uLyMpm1985zdyny8qolc6z5v2fLFVwAkpsMthCddkXzWJg/5ujvDFFHvLAPxHLu0HUnGpjEz6p
u/MjWTbqb6VA2IYZY8Rjh+sMEwSzxA+9xPlBh/CxqAwUKCy41vOc5ppp1hqvus5fdPgHTMN1/4yL
V6pewM6Fom7RARse3NV+oWzVE/gqcYuHZJlWCRVvSIwRjnu3xmD7FOvfOfqA+6P+x1ylsr+OIUw6
54wkwZ3+d8vgiS2GANBZ6wd054t4Dml/7RjZoE3rDc/t07MI4J4HNa12OTNw0E0YenAC/UjdlqPm
6ia0+ozXnV89Dmo5SeeqpK9BkqUiMbVjbFVTpeV0vbWdOqPBKctcLGRoKCKRFpE3gdEzNeoxWPWr
ljhkHSYfNl6tvlqLaePaGK6UtYrEaY2KuslmcfB82bW8QFjiO9W03OpkSx5FBLgLN1CtifCBy4XB
pfA/xYUWR67Shek3vd95gBFlNRlpwTiCik3StAjGT+FFjj3AP05g5rIw3aubXWvLrQRCZUlJv6o1
LRXiHuN77+vJbkLp0gWJaLOzYDlVN5kouPne3UA7o4cXWEB9X2ZZNscTaC6rkx66ApK+dTAzKc4v
6p5m5aVwt6cpTZU7mtFJUvfu+H1t8aQsMwtkZlRsZLvUk5SF7y97J5kCubdbCDrQauI/nXmpdRXo
YUVe+cfJn6RR7iYIdPYSqdtptPz5GMrPO/yYvG7tXOzBPl5Bl+bxatQBTnPhfz/AZ5taeL8YeL3d
jjkOG5cxKFe6Oxou1dDFySh9ExgbIawMinStmisraNr14eoX3U5cR+FzIMKr/RuQaYfHWJWOvrm3
cPrBlkiDk/KL/j1XuCYFz0YwCW3ch3sbf01LuotwypNKGFukwwbSCHWtB/BjR/LEsKIhxh50YdGp
mdWslBKqpe4qAFHGUcOjfjm6FKsZLeUJDay42Y/GQm9qU30Wg1D0NiivqUGXmrlI4HcEwYzNsAwE
65SG6qSmlNdc11mE1WsL/45tWQHtHtW6WGkK21c5xbXYVsdbwqfzkPuwQkcesLuCRpBJksk6fOtP
S0U/38+QYVpARXFashO+iY8kg/pxAy6kRZNlIq4wwr5u4wB+rTbPjS7SDxN+eubmmNNxRrt/QzQe
x+NTDMx8JMD67DZgU1WGsg8F7gWcuaymTqwlExuh+9XlLcgrYUqymX/wRDXMxd7SoxPdgJdZNvAJ
WW2NoZZ3dJ3DV8FQ9OpVsDV7tE5cnoRyeERQ3RidR/1dToXOGmkkDcud8WwPqQPUqGFqjk8+fmIq
NpZcCUc1LGFo8CQaBTJZhfTQwlTpp7ReHLRp/giGxrW7KIhwpxSLAizrV4ezZXccuUeUkO4bMqlx
t5Noth7QP3cClngIxjf3QaSfQuIvh0L8ZwIIfLLqThtGNtTTDXMrbH7I5uxZpIB7CKhbLPFG5ETp
Fj+XnLK0nZjXW5Sd9oAEZ+lMpAaCJ+Kj5OoMwRbXI8V2Fb9v+KwaPTCiFSBGIZVtXPd6H0OVNKUn
D89zdtS0ialpeiv3uW8MvGVfXs3ZXQSC3DwNUTw1Uqtwqn2svlLpr5+B6M8J9aWWGNGH266j1+b3
dk2xk9GR2CPtlSHD+U20J22BL6IA7lkNlWhzmQHi/EuRAcYREW8/49mWkn18Ye4aCOTErvA4Dcfe
xLowjaRGlFTUWup5hg/AZncFdRorok52t+OFl9MbIEztiBK8EmXrEcFAAM9jhyi4hOK7Bvga7P1v
aUKxPgYLuNZb3aTS0o/mDbxSuk6OSeLcGYkIm7lW8Wj0ZvUNSzKbx3dyOVXA3BLTh1whzRoGbeZ+
BrwElHAyJ/GueQolbs8rtpHhzxPmlkObENPLTdkyOxof7s1x6oosywixlrz9OT3XMzqaUwuHnoTE
X6HK1PClyd2tvI9Q9QZ9cAmS1fm0XkYNa/aLZdkgk9EVxHEG6ZylDKBSmLZuUvZRnak4oqisjigd
l3A6KaH+i6S7SXt1PeFl3GPeEb5AWgHT/E/a7RptjrdJX8AQbTc3JTUZHkGVm8of3ZlTpa8z2yZX
GPqVHd/l/7RA0VpsKpAzr0FlTJHx0jImlpLSqGns8KLhkf1r2nBw9rWOp6sGnEhmYok6dnXIg3Ud
kcgdGBAlIpfX4PXmZIQKLMDkRApl0InLu0U/FQkHxRGJPRCkIikSKSaN/EMkJTGd3neitIH/Qjbs
5BlfIyoJNh6MP/CTotVjqevAZ2YI+U5Eqt8sWce4c0xVlcFNhgUGzJvBPjwwJc/N+M0N6AwXXpKd
86LxiRnhhPDa1J9BJbw7F5T6HkmFErzLGD9w0d4o5sHypmglaHS/910EdB/7VE7uZWF9f8iOKn5c
9gFQqUhs3mSVYN+xnU6M7MddFrdZXo2FgLMCQtJM+a2hKWquLHQ2dv1Ob89i+hmfUrwXY7LzVriW
yr4HyZ/xA/CPYDtKIGurikBUP9C+DgdIdcSaEZnVmn4V6iVs1P/MoxEfmnN1FM6FoPGZvcR2T5JK
ILidn1kjnST/bpwRNLQNtVTd4D+PzPyQB1Yb7gganqJytV98OPBE8VSv2EeiIVN4cuNvlJW1SDOf
cpA173fzBSWdq9WeWubYgRcN+bGqJpmD1z1NliwnrsgKBz6/2bajrqIq6aggjH+5bhCcTQk1epQx
9udz5hUhf5Kf+/QcJg7XWKmw2RXrlmKe8Eo4TJYG1NQNYFWiuUNo4+sJgq/acKcrYbJU+1tZkakv
/wfs3x9NBQff6UDIzA4/1/DwbDbOwNF3mpASV84tHrKjaB22mFKyxcnun3TMgkts7WiAnKbLWLjW
nlBNHuIHyY+n6ByCAPq7R9OhFgpyNbffBoNv8YbO8DH2rNzZbJuif1a5zVYFs7cSbAwJN4PAuNlB
kTxsKPFoOK2d7WaOqWyZPUr2KqQATxD+t0r/NZ8lwNU5REIY6l9bdJOibOyrReHGVO4B+7xJdA/T
m/rnDQ91nGMvQcMG2MptsPITwUr3TtJ47/EKa6qDHb7ur/n5o1wOXjvTkgHxs+TIpQdMze9nfUJ0
Zn0VC1sfoaEkUJRPHfd4cqwaiASWzZbt1yptxNhLGAHIWXMIaEk1T6RA9jKGaOabQaVrdHBUydoi
4IqlxY1jsaQnSEZBtNsiybP++0PWmzcyp8a6Zpo1HOxmU+CnTMFGTHuYJr76RurPWAi1PV2UyoOJ
HFTmR2DV54/SJ9bIntog56Kxgk1B87/4FjJ5IpfW9a1bCeMaw5rrOpuMA8ZgMlZQHjUNn7zDj9Td
leEvMhg7/GiDKhVF9Qm44apkF4COlRwVxe8PEE20z7YNdSXvpQNVchWxhJo+FXp6bwUMQagp7mZc
DIRyxi78QiLQ7ooKb76e7Aw06rkIetLjXgSy+9WJrnvMfMswrIHpkPryA1ISjXfeozWLzwBxM4wZ
mnNSXQTBlXPwI1W3zcq85ZqIAeVqkrwDYYnMtZ7+VqhYWRdbaVUFwyP/PnhuJZW9ZBCV6gsgqe8t
5F/7vecz24CGRT9CkISIVu4d3YSqOqZF/yf7CNVcaTJEwEAe+aJaI/9VEHDyf6KGg9VZ0FH84WXZ
hFeJrMj+Lcc85jl75+J8q/HbMg+C6KLqhDzLUrI+qy4o9lrwzKwdv3drZ/Yu964QIFEZQKsfzSKS
maXOL4CWU2JjyU5B7TQCpBhj+LuJTiXRTBwp2joVtJA0zPVLOJjGc2suQvmqki0CyuuHCk5IE9Pq
fcdQQ0ZYlRmb/or7ScMwl/IVnHIAM2zSslZvc4b/yIybLUNMr17QeS5qMsFcbHYpSVz1h/IiRdV5
bVwbYNxsNmjo62K8u0uQW0A1l4XUYpCuANCjZkbG/YJao/z7vCb4NWRgjHDY4eVG+BgvYUc+GWtx
a0sZMzlaR3wJRuioU6MZVXZWq7REwEK5PDdfIiF3mps+zs22iAeM2kkeDmtAQEhFE9FpTsuyCJqr
YPA2t8MggyxgyFpznBD/ttwSPAmuayKUO4Nj5VzbXlUggfiYi5OVZavYDx4v2inud0WOAkv9YwGs
hv9407V9lRuQjLJEzAvzH4LofAwQxWcBZ5bJfAp0My789Ypyx9VODLh8S8RBjKNu5ByUtoFQJah9
3cMzhyJW/qFcnCOwB0e4iZVXCfcguxmw+DKMaN2bvmNKArpQILyKSlXoqPd94bZHpS1cToWMPqxw
eqwb5DEecBVLPwYJ/EKGCUdWCoAJzQnx0mSOWJ/M9HWkmKrzUiDPPJ5Xj7OBx2kvfCFy847Hya3J
Jukv9UJRQfvdouoM986WGU50z8BGZ25GbCdidQp2rAIzp6Rru0gDLSVvTHOGmXj64akVgquIuI5T
d+AMuv3cSeKzzwR559oNswXD6BYXMyuuTvwDwvkFfej+qfd/Cki+ZJQdHTQmpkZH3zfH4s6Bq7vf
jCQshNQs2H9SSEPdhrIl+2/N03X/CNT75tMJJwE6SQXkzsjijG7iy0Uu4KUQvP1WaJ8IXHbvXBMD
+duKrBbfKX+Bqo6uVhM6twFICizpn/1XPQwVwovYmO+R9w8q1iep6HSepJe0Rqlm3XZEuFZQflhl
fcyDsoiISWRF+u6WAwMerHaJqqA2y8Kb0ag3vUfWrKtGnDxGcb7nUgY6f8U5oBFnE5iR2Q5G98jF
4dv9ZM5/Wo+mOJ1YiFmdEm3yrHbO4Z4tX4s0nJoSSZlM7jkBBM715bAVAs4qvC4OnQl1grH1sdkK
kEWMcQs4bzK87VF6sPZo2ZRvL8OljupiUlobeMo+shlAbkOmoKQJiNGwezjQ9KU4hVq7t6OJPu1G
A/kvdsn4xryLmpzOu94BcRjLp1sNHDqxDgfOHho+bd26qC70vneu/7iUYHVKU4P0BgnLpcwBfPe8
O4du/bp/Bh8GcZd9vzQXom5KwIqIwF45mxZqHCezbduxifUG4sdbL6PymtIgsgsnKrMWRZtAmDTt
z92uIwWth6D2BlZw1hp7wOERBtCr1xgxSiqX8mjs+rnjM9+hh/rW9/09Km4DQ9z/OytzyGkBFGoo
nYRaHWegAUTZOP6kmqBxb0///0v4aYpBCYVTdcmJWmTFvwesJLA+89uTagNwC9to8CUQMkjoDc9A
a2s5BAdOuF9QRqv9PpvKN0Ot4kdXmWyKOheA3sT2j2Riaxpi9NidHpBJWKiv2bChmrqLY47Jyx61
2kMYJBt+q8PrSziWQ5AImsOan3ymYUiGtDkfU0Tk334cWw8TwyiP6Dd9n1lZ5a+0u/88yXSzga0Y
9WFCJ8+8gDxOk8K1Dw31lerZYEGPYa00ixXABkoPkDbh/FlokX2jceuEjXBFLBy+kCZDxMDxJ7gy
9Rjc9e2Bq3SRAoz+ijr/BArF37RUhjvxDMOIVQMoAlOcX+A6tZ2L4P2lqjptftGqD2YYtjw3ibhE
ZFuVjSVfVoaqLnw44eAQgzxfjV/Lksj/8Tv1CV9oykEpqfeN9o8U8Wp0ogh5RnwztkeMjvTnjgsO
xUuPNUGdba5tSTFzxBO3wPNG5dHrtAgtV0rmypT/VqFfselndk6HGbdiy5kt+qVVit5LmYx7GprU
bK/JcHghGLpLYKx5dmHbiC6fl+uaPPj5yfhnJx20E6GadYzL+qv1cmugyvfBJDZE0V8H+L9O52Cd
0bUU9+9rfleVuTu/JT9irenlGGVknSTWrB48PcgmFrmBaQGHBmxjlEmhUO77WRv2XeQ9zeEV0nIL
EjNZWKQQ/Tf3DIaT8VsxgtA442JyaCHicwYKZyDwfS3Zd/K6LD2m57MmmmiojVGmcGC9JXyhM4sr
TCcMWlW42kGRDlvtcZQpiJ99bKr9o46iG7c3+o6QtYhIFrWZXk1kzxP+pusvgV2WecTlcdY/lQkB
UaJMlkEvQb9N1cpJ99bGNKJVGmURUTNJuKUzHcHezDe8cQH4StoJYj8lv0379AKTfa6BZ9XptaUx
9ITksjNGDr5HwvY67SyfmLJY0NBo0gtAE/eRWZJuunZQSNB6MkKBvl5sd7iBmWphjt8tkpIVUPS/
9o71Q+phNzoYFxDuG1XzYfCBZESt5USs6bS4qq+W7/sJ/ASYXWxgXE0XE2YUTilR93JQOb11MT2Y
qzRXE/9pXc5EzvtEtOAUY6m+puQGd9ARC1SfeJh2NiEEH6uTe42dPDmxCWgK89OjcVeRZrk+yZQB
z0zS9Wdj+2j9/f8ly5TkyBtBRNBZzyQsnu4hbTz/jik4mqirp/zDWD/rKOyye+aKJ0mHDDvihd9k
SrgfhLF0u5pCMZ+d9jdtd15AwkCNY0EHhIQwx+MpSVkLpq2aqOgV/sS7FX/S2NiPD2hVUmCzlcv4
pr8melrXvvcIfUUVLqnvSUohIoLKyFL63N08IHTLN8UylOPT8z5pSxhDpIeq/Y0CvUIbjw4IymtZ
/pBh9wq8t/WMXQQ2vMX9K2Fw3HSQX45CSCOSgbVGmviHkaMzidKnsUhj9gU7SZh9aXNlPaCl6i1B
RYJ3IUMWFkn0dmY0wPEfnznciIhQMU6SS7OCILhPDzenzfRpac/rRysMbwYltgvIQkwdAu4Kw01U
MiOk1AT4kW4MkNh58SqxnOSLpWCoSouPODZtowSIzAjqfhfbNM+5/5RcVYvfnDV7RjPnh94twQHL
MrWCu0rNJ7wLXSNxO63iHkNykw2P2LldojakIibh63U3fzdxlnRASekrZvlSqKQkFGVsLNyaIoqr
FQymdIIeFd+YsaQt2YxttNVs77Y8FfiQYPKUQJh044fVk1ISHlygwJwQTwZQW2hLUq3tfPdH3eJB
7LqauJ5m33J9Dzrz4neLz5pvNwAxd1SgbkTTwP2gQ8gfjM7z/UTmnzXV8fBwRrEu7EUw9vBh3zBJ
iL7h1L0vWkQy39wk9NgZaFtOQtxzq8pe6Oridu2rvwAnhLNk8odPqZQ/PUZrGUIdXTt7HxUyOdzs
vPsgtskp8nEnk4M0q1s6/FkOSxxGIVSW4Vfpy7j8avFz5P0W2qrtJ9abyt28GdGH/NLC2xJCdZmL
OVf6gJfeAbQycLmioXCv3gsBp2jnCokAIwjQzsZmh+DQSr7N2BUsIT/rNvAUcKDzOLQ7bNthUAhx
Qm6q87E/fBTmOF0jvX/ZbxaBNBg3rWlGR7R5mAN7il8x2WMW3Fq0nA/yuhGWbqfpFxUq+W5HwnN1
/+G4Jc/ZwJLcB4FyUoz8Ox5mJ+KIGPkA+1y1YFFYBOoRQZt1CF0VC++7ROWgs50U+0er8oiPo8bd
fS3lXVTFJUndHOr4Ohmho8d0EDBxTMZhXOpAJh01BozvEC4mEQBf/44Jdd9MeFaD6zznOEu3oefj
BzbKQpianFsEsGzfCBprEuD2SitxviN35MqYKNjK0glO1/pyeUAzXXLluCwvMfWBMsxkp5e5dkRt
U+Aid48dHV5AYh5KHOMFi56SBjLSUPn9797uTpmt8iiXXtkF0tbHqtVs4a5jQ1fFAD155Js38/mT
bjR9BsMHQYtLf9e2glwdcCU5pTfQPOI3lbQS64wTOIfwhHmud6PPspwxL2mgT40H2KDNia7YbOcE
chQqxxkXguEJ6fXKTboWMP+1yR8lFndZH17AiAGzCnB7HJmFWLjqa50s1ngSdeU7BEyOSNiMfp23
j4PZsCKnDIwCXldJtalUD+FAO1CnvUYyXy6B2NqlsCqXgdH691uGwGBHPpcKVYM8GAs8IeTWysjN
/CDuVlRyciPRVjHMYXIoB1U9ETngrbz4sRkZpqWRCShrDVb+QZ7zk6oIPxMWIo1Vbko3k9YPyi3Y
T1f9RAB718iEXfbhlT79se9lb+qwbOdPTo76N4GAIuZMtkvkIaSYK6Tmdf5SUgN5vcZ1jG5mbijk
Kp9dtJh4pozuiJ1F7t0xZKWhaUSdC+TPlhfx5p40r2yWnDSQ/BeN/d7c3MoVQ7SGq4DK6xYtPVFt
FszalNAJ/v3x/dADemSXQyRyVH0l1IKT5iisI98FVL99fuCOme+eFYi+DTw2OIYuQDBJxKfCzfHM
Z49QIyWu9FpiXN/22IJ95VN8IV3e3GYNCP2SqRCeUFjaIuhJF0fZ04QBFazAFFv3stDYwD60MSAx
Fd0ceXXmqe9kbZy3eyCNDRn6Z4eEmFLf1pchim0ggdNl1U15D6mopCFQ1UHguD7yzlKPQ/cjSi40
kLOiLuG1UZadb7pA4VGTGZtV4p6rZSjtKnkQ8t3uByeRvR1VkQ0qRj+Dj6sqUs73T1n70ymqA4ih
Y2UzUirnT1kxHBBA+rjPc26tcDhLta7dR5+hesAdWk0r+yZbugMiv2OTJ5C6KdRhK7vWPyohpJlP
MydsqgWnlNCNW6rFD9fiX+Av3RqI4OFG54dZyBgnfowVC7roegJk5bbAoCtWNCk6aaqVD9jjKgT4
DR4X7tJb4H3x7J7jDeyY2UApfdFEkVw4ZZkarFc6uWKuGKHy+VrJimK8IZphVAZAkWV6ifUhy699
18EPDjqBnoYDIqD8mbHXL0BwFfa+pqiIXrvZ/pQZa3hmMa78Ma4D4D/c5A9+Aqebw7h+622UqFIw
TeOwBZu0p6SVJFk55Gt7Tf4gYuSj1ojCnkLvsLKCiU99oDDLynpywBSdlyz96654q3wkh/hyJ8Tj
/AeASSHJ6CyKxkrEWqTXHjP0blhRSJOu0KJAw/rRICvoebbKCIMzp9gOxfhkifGQ146uAaSSjo5w
wRM06xAXD0rgu3hmaf8l54DlY3oIbRs0e3/+EN9cWSyIFOtZapQ39JvhMdHFl9a0U9wH16R3w22q
KxqUCUNGOGoua6MrIPkS3vwPpV8mocsYnnEZ4zq57oeTTKYc4++pNvSHua+o6LEawozLTXM7zZaq
I7T3XLW45eDmWkQQmWv5Gb+SZFQeBMT+1W++2e00qCXm2ZI7XbQoBiDBhM0E02eSJEDuZEz+uS3z
+j1IMNjPIxPr9x+IsO5EafLcdYjObO+kbFDTeM9/Ly8/gEHm8UtUZWN6PZxWIrafVLc1bPtibyJx
zGFirm+70Aib7OKVBVO03ob5BftiId5So2D3bUL/2aEfdhFj1iVWw3oj0/4Vv3E8173/OoG3Fbj1
ZTupXk8Z/fZULRNEJ/yNj3bL70RGXUMSXUZwK7k7VGnzVwLWo8cyzQdtveDik4s8AVTsMcSsfRu5
Rz4d3ajwYNcXrlx+8BeBv/N+ofvLghUVIGKpSSzv28rwMLbQWIrv6CmiN1HmGbAKEjvFpv4cqwo7
XYSz8nvud6cQCddbunxIlKnY/4iS0EzY6JywPiqsVnj8L2YfwAH1zM4NpaTAvmmchnyV1CeC+oce
oUN2/1uRogSbINjS8uknL6xeJg8OKiZ4Gei+6FBahzAqcxPBrzEMjtNzZ0ofhldX6d0AjfBmPZ+C
v31S5XEdLMdZFiQZ/cGqM6gyQf9ai8xS8lWJCiknAyUY2oj4CJqZN1qgj2PsYQGFginM2jxT7Jnc
VvCOxur0UJKTlcdZTYaSaQmAn3VBBJYP6h1t5BtH5LTcUbPO1uvM+Oq8lzl31f+VSLy8dnwwbhE3
8K9jtow/4wLJOwt7b09q+IBI3Z3M7uSEk6dbeeA5r48W1nsFpgqS8iGm4419xyUcltGl1Slxw8P0
RqSODjcJtmMk10q5flZ+BDfHzIP6wzf6eRD6Ss7gtBWuBURYnIS3VNuCeqWUUukQZdhxDC3n6Ks9
esdU6gcbrgfpJvChdU7Fa1VZ/5SH89nkqAcRuYTUE8gQipgNhX6++r1Eze3Dzemh1kjQ3DySDs09
4Jpt2NXNXfwv+uk5kfp/Hji9iadKn0Vbvt6j43KbPfeYSqNHPC4TQ3vucbPvurrTjq2eaQxgezAW
c7ue1BKYO2HyjZenJ7USBG2jhsrqWrdjDoUPSkEDc+TPJS6Knh7Axly/DYQ3YL1VRW9LeMGzSUMz
aPeqdWeKDJQK2z7NW+hX75AVvEnLsjPE8MVtEcAw3Vzm+yysTG6jZ75sRn1X/gGcObLbLf2iugxu
6tH1nL06gdiNEg0Q5BACH2WPh5VKX/r8E71GGC+dSwI3teg26FW7gxj57l5ZyOrContt7yDE4FoP
dXJs3mspUzWX2z1HYe9pJSOActWz1LdWzt90baPiQ9zG0u64QCxKeMraLDy01eG9CPY4f9U5zuai
9UFZr0KHCpjuKc5uKgsH+FgzuBI0Vltt7bGQ+UKJp+fJOevud7+CUgcJEY255dF82AzpUWlUe+I4
ZH548xkwCCGipsc99doDO7GWfSD4BDUsk4utTJj/hhfb7DDovwOBy9hmeN3YRhJIOHwbNBrUh+Y6
HftNCTInjj0DjJ75ELsibTOWpRRn7DgHVFOHzBTpO61B5aL9vPMpmxY+xEuM0CK5BFRBNlEtrB56
xphNint1AHWA6EysQWqtDUNEqoNbG1ZY0z2qEvQ3CcWTrj6+bjLoiA0J9Z+uZHvqH2vP1qpm1QTx
tPNCc+zsc7pDtS4rH8INxMbKn+tRpvqx9uqcucZ3CkvRNrK/6g5ivSpkJa75r4NewGYCD9g0hlmr
a1tmwQbhIyLwkcUoP+5An6w9CV/w8altb+Pkr9GM5L3BZuS/opldlanIRzccrl+5L+i+/EjeAp8b
AWqiLhb5PCR3YgC5ye0BthqKBAskIyIxb7SVAqbo3f8bsfFmx71foDFmp5PQtm0NAHn+bl+A3VZJ
xX/yMulRKrIOzn99aGJB8nvJ9fKknOhcU+eSaJADqzp02Qec+EiMeo2N5+3/sAZzLN6kSLPEemMq
O38Z8kdG72c7GVLl99O5vfL+cyfLel4jOtUFBkPpvzvcQrbmNRWkz6EEHs5np2r0p6EfW7Jpb21r
T+46libutqx6DbitO1m9wrv9Pmkd3M11REvooyQxZ3lVf8JCCKFztt4k7WwMtB/TP8yqUiwRJn/Z
i22iPHbiaxN6EVqxdPHiGM8kPvVspeoz5l0efCbS1allVpnmvVjOvzKgeLiMzIJwgvVBzOPfsMIB
6jZ+VJqYlaEDbSyGwXRyggoPPakeyh0AiECtxXdeKxkLzkXM7E3dbGA9xa0NuBZwRDROY3sFGRQ0
DN3eebTRslgUnS6gM2/qLbrI+TYwvBbR4gKB5OJ9HzQWxGdOs+qvwgtpuaov1xS8SRe/1HoY+XWa
YGLUd7Jk1iRC8JYj2HmRABZlUGSjqS6a6IvtWkgN8R8ekPSzfFwGzC/kvOdnixohBmIwDK9s5B5W
+JRslPTZIK4vf7++kxnFzmdhs/Fdazqrg9v87OzP4zeHQ6EXco85xmNU5aQp2/pNLsnO5t9OCm2v
mj8+GrJXlVqabzPSNS7Psc5sWs8bQydVwgqacOk0WUMK1nDvlZZX7Mt8wrwRFDAopYVbzmRkrEA/
UH0VnQgQc+ZkIGFXuMx8ah61tGH1iXomSPdAxxdLnDCmVLo092BcDEsd4jIegsE23ibQ9cXmV9km
PGcgOzqt1Z3was8CWbUns/0XnXok1ZXINzr+AW98YfKNFtoiCbbpIWE67KGxQW3+Upok6VZJXwjp
GrUHOHpA4zOF7ewYvE+g0fQBHsRbdyB2bjE7t1UMJU27BWz8si4Z9WuNcw4zC7MwaAXHFDQ4Lgrx
cppKUpfQdNvDupB8f2XbuPnZDpqmbwqGPBdQB80CeKZLAiRUNwYdmilTDZdZ3kJrsjDj9yOxbeod
HOBA7ideiZN6/dwwYrXrf33rkz/EVBRqLHnbemjP1jDzAUTUTId3DUoUxaPrIQCBNZaMSSn34f4s
Yw14UQpH5jZo/Mr0o0OD5y16M/AfK+GfONr0DoN6YOcRwG0UGDUOKeZL3D7cJ2ePZrWuFXqP8qNX
do6xMP6QT00gWb6e1UpM1jAadDLp3oFbb1rgrvw+pBUh1CzFiCMos9XrbM0b9BUOBNzD71j1BUha
LK/fOf7HVBH4BOek1iYkY2lKzvzid28c8EGzGJ/vDcgiIzUnhG2D4ASybbiq7e/aevogbQJRCGtV
XyPxjOVQjuag3s7iZ1stXe+O+/lszxrfa3v8sMA+DDp8FCe8SLubJNwcS4jSLFOx0LBAjGda+ElV
TYBFHe4KS4kwjk5QgrMJqJfiE7mqoXxUMpxhHsFFX7U6AmFc9GkEhD2ENb85UTLFfeoSfMzy3VMB
Fbnh2TOpSMPkfsUm1yIMYLxtoBjnXZnQcbdsTch9HKzOCDRF+IxY47Fy4aWUX+MxHDJa3Hdw8HGu
Pg3vdZRKpKaRz5O3WDWCyvb/Up7Tmvn/OWUysKxVkuSK9aP+ULLTAeAiHO9tnPsERIcGtG3HThva
M7TwBmbh+xki5ywBrgGtA2MNg+FWJfhWVLlBIPQoIazPxJsbrAFwRSrudlJGlwJnzUW3K43Gbug3
5XtY1s/YUS5v+HN+qX9Xnx3Xw5YTqJcAgrlManVPHHMV75PMJCDf+fzF1Xtsf9V3YnxnkYQqun8/
PU1nxzyQfBBzpyOwhiNaR/tkLiu0MfU4zpBWM/K1pmh1jFn234lcQDPYtl+dGCDpiMo0DKMG7sZF
PTTLzi7IVyHHw68AaRbxsuC7gEmYqhVzmVpKFWkRc3r8m8afNE2r29KGtq6GncxsCRWn2BLaSSS7
8hd0GuNWWjyL621ESJBhjOdajwu8kqEgoQn0ibmYNQQshkagSxGVr7tGVkvPqBmp9OlbDKXcQ7zU
cooFfCqLuRIFGZnF7VfzJU80Ue2HaGj2ljQow5066WvG7iySkCg/+tSAGnPjRzBkbnsSJWnGw2xK
lwHOgncpXJDwuQaxHflFC4k1gA6c4uILDNe5LTcUK7AlnAYfCUwcW91bXpmL7ukq6xuvUQDaEzpe
VcyQt1T2hdWPSxbFvS931fu24y8h9K1CLSfINmTFXYNkJZ5wglTeDcW5sJYo35KC1yt4p5AFufrg
3hpEf2pfL6zpwIHBIK/7/XgSKSZifImil3ChJziIPwGBC0JG9ZlY5cz+09fKxA+0F8lZFt31tIdv
lfHQZFlqGp5BDlS+rftHyOBgEDMKH5zobMX1ZraIA3bvkqdsmZItjWkrwBIK09JBmNKY/MFRYhjX
LYlNv/aIzOLQ269s9w/Mvr+tUc0YYkkQXE+q0WotMNVD2y450C4hrMGWGQMPj5MUDN2YVvFJHQBG
KGJCEa6KkfPeN5u3jDaWu3/UXfXEws5TTMTYcnZFSR/Kau4rVC0hNP9N/6SG/tkPyChSeZGQyfat
7Pq+w492oTniqsy2leqG6mLg/I0aYDNwSrlg+fNcQW68IWrmKl3WSBQ35rkB0HLgFj3Z/fm+tB1e
xgmlCKsUjzXxCezVo36scvv28EpQLh9Y2TYY8CjViYphhwCwWx8XezIifwxbIJns690MZNgcbEzH
ZHi+/T+381FGFzuZbxvmOzf34cRirQwufnM38ivobRtPZ79NTD0maYdVhafhzKPE/Mlc27RJ0HZ/
tgwCfXI73ud0pU1knfGK9f1oaZ/ROuMt3AxHfOA+VodKOC/7g85A4BvDo/mBqkiOGq5i7u9h+8Nl
i/7xtHgtkss0WP0bVsT1BcxafHsrydFx7LL61DUg9rTA3tQl7rXr4/TYBA4X+89Z0LFnnpmAf5lL
Y+f0JbF58DNVkiZdi2nPEH+BdxTT4P053IA5wxII31pvD/nKxdTGpsP1Qu9jc6XNNYDGFQXAHZEH
OFb+h7MWVUVqDRsqGCIN3hMOKbq4Cy3oVN3JV9bLbQsH5fcZeCAY0nFBsSaY+DxkRytkFLvnCmyU
7ehAdjrsIpCRkRw341nuQ1iTDsM7AcOHjpWwLhCOa3hHyZIineWpG/JeHXFdhCxDEuCkAUJ+l2fz
3gYgfSAdT08iQgL8YYshLnRenEOz2QAIR2nBG8JYJiOyrSolvc3SHlYHCQapnlOHVXgzNxBDhNmY
cOJhwomOgV7Tn8mm6RmOViV21E60QN534+Gf7zeUYaePNyt/jtG4KKWX8R2NiUD+5gt+uWKdsmYO
LJlREACEDO2KkP9AOIkk0bEVqLuI19VO+gzwzVWz/dAIWDY7TcgmyEdcW4jWSLJOWitbBG5g0hGF
paDptJpg7OuA07kxVOc5uVhP2D4xc3sn102lClqx5m5IcE5B8EO3eATFwxbgNtSwdCm8kkozA5UP
mDX+gVe2EMeGJgbubmdKPnPEbgtN2T6j7CPzySN/ut0o8oJQmvm0F+5f6N7w0ymSuxlAmxOgemHM
k/T+lMSPSraGqqe1Hx1TvoiFQdJtKRNXrlxatVynTl8s7S+35cGRcLxvhXqNtGB5TWpQkyXBuMdm
odYksBhYTy8ATVNnwQG0Je2cBX6Sd4tl9vV8gcjWcvpIn2hjRN+/TNwAF+GtCJEMoSR0SK0UaH+q
W2QU45EUclqOPUGs2Nu+1KEV9ihZH03nHbOFDADgSjgUhKLZ2wB93d1A7WAnYKO09zO34w9+E5fF
VdkBHlOniDAL1NCEtc6JN/rXXWmMrHFZ/7+obsM98C/IiOqrusM0tF5Y+hDl85ifFH+Wa+OoIb0Y
PS3pcuKew8RUlqMbaqbEvd39PTL2ispprYVbdWtTbuVCGsGnuTgeD4SQykEuxg+DmW+JlzzxMfTT
rs5hDwD1OaXPTg3WjFZnlWct6BzIndgIiDSQgWxTYguAtXzr4suTm38BKhPpE7jGHOPpKt5QRXr7
AHX6qfJ/BMtKRKy+D4diGXAFZCy/QKyOYC2gkS9Z0Ub5BpqexsKnwd7U1y883O+g7xRy8X1YkyIJ
aNPO3daqwh5kQuvLqRgR8gaizokfb0isoOuBJp85l7rLBVGx9yov/fLHt2AIa0hPl2nY3UiEZITR
UCT8UHHWJUygE7JlaqSD6akmTM2lgm4cJUAq4Uhem6rbeOs6xmFR/OzUs+/uNzxCfZdGc8LsodeI
G7QtgHKK+t+P8b4zoNfxnnXcPNFZKim8uy79th8B0JHTxm/+myZd4Sp47dpOWnQKLLTgJNbT6dp2
UBa6okym1RJUeM0Iod4oM6fOqCsXDB04ulE4cevvq1u/e1ZrVzkDr4dIq+aXyQ/SW0WRuFRDf7Eh
JqChcGThOMvr4ffLfsLT5dYQSZz2Eh3UzfyhanyknQQR/l1HyEWp6D0PMmUTk7URdTXTut9uwF2i
dcvbLMNmITHOYZwihTdJz0va7LIDmE0sPreYy8tA9cMSJo1jSNHm2GZ0N+TRxLFgp3esNVH4LFpX
eg/G9T92preWC3loMNLUgqp8PoEk0pzBrnoK6hJnDJZd7LFOl94Kv1IOGkm9A88kEXfGsxUXT46C
56A/HP+/Jv0n2laPJUpDWayZA3jPkNfMaERGT2x7FJZOZvBT9mnHWcNMLOxxN/r6QuyIWayNaDo2
k2Kj/Ssop333pABAWHubSfrELbfIZwC6LhShSRnNtM3iWaws+/GGcN0Rqew2F77kNuYRKiR36VZE
ElTu7A6sD0xnvn3zv3sIXSEvSRLdnDOHbo+JTPnIqfKxEBHUoszUktvuCZOqJ5ZQRvDUIojRgN7b
6V7QoYLMpuaM3fNi/ULYvm6K6f2sga5EH3+K/wJ8E7gMX9LWoJPzgO8Fc2FyV+Gt5kUAW/0yUmmb
G9XE6nN4wQKUT4z3tp5IT4VfZIEzA+YdMkMBDkRpn5Ka3LTnhLcGHge1xMhWuMyOZF6CjB0Dsjfl
E+GJBYstFyxE/w9c6U8GEUA62LVp0Hb6MKaG15HFio53K2uPCF7SpsMnZpMWwLql8Mecn7McL2Ou
coTiTrrXspbtZ+arwtptRmkzu03AoHkHolqaetExP9MoeDXRJSkPnDGw6E0lTacH/v4U516hQhjI
LXt2M1fzaLfk9gIZ0GaFR4V8UJjI5oQ56VwPkMaiccv7bL1E8Y92XwvjegBkhjSis1q6XB0668RQ
ikve6EOO3S2RgiSLPZJxfcyg5DPwV7wSumOj7j7hVrhDZirBkupJ8F/x5704ppfhI9hPs9O3s6f1
3D+v1ykfxoGnEfLefdHz1IDySx2eXtLPnc8fxhirf0p0s4SGci+pU3CuOgfP9b/sTNSjuzCqbVi4
Kk/d0EbWhMnhQV2glLYBSTcJaky1cS+RMXdvU2t5MqA5yVKaDYqmzGIdZDXBFl6l7ps6B0lvVx1b
E2SCHY5qUqW7QqsYM3vZMJSFD1Gktzpf8i8MqUJhvW82SIG9Nn+wBRTsx1OA3+2ZxYOHmT79McRE
nyFO6mO9aiO5fHujzSlo30GFSpJzCF8SVd1IVszMBJayyrQfTUBI/um/KFzlaUv0QgNW4ILeceGu
AfORXBJPsJmiZ1WMqr2LHj4feI86eVb8lPgEBN7m/4tYYEiBMojZetybFcWTTrxK7Z4zwJxE0ipX
9QBuSbSU32qGPi6SmTyz+sF3P8gHhmhyjZqp1QwcCLR19vx3iJMoXWFMteHEm+4xVbMkK3xAb1iS
eGodxIkpqGFR/9n2WwIhJDJkmSGkPO7f2E+f23UF50nTpWpb5L0PQObNJpS9bEV/KsociS+opDIt
Tq1ibKLPJqY41s8pnCYbeh1SuVDPqbRjACtgzFH06RTGA/1GrvVvJ43ASyNo18+m1LcbFHyOw8Iu
dahlIRdX+GFeZkxsz1SS8RSY9wS6IO6D1uEjNJLEmDPASZoC6Q6Und23Rpx3YQCglLDuRvz8sWnY
mfp2qfCsputS1OZNpAqf8Z16XFd9HUP7ZZDWghRrjeFd3eNdYYIGFg5QSeqBZcD9aNBrsRAuoM9l
d/BGvIi1dy7+2BNiQqHPKUaxLX7q0psS7zYnw0Wo4noqz6EQT4wQ447MTXEFT5eKJFlVxYtY9ljl
E9FUb9gbR+EH3rq/ulPh/5lG6FliP9Fl9/XEyNz6cunAo+J42YO78Heu2AB9mbfLrUqtpxS0zZwH
wBB/YHZTeetTilMTjTnNuL8+wf8QMAnQRPQrHhJRsmLnY4Z8lE6atfhm2QX8SoxnzxxaKIni6BUE
VCh/G1ehzJechhOACxBv2WKBQRJgKvQlowj4K8+Y4dyhj4sucXhV1/R6EHbWmzOvOHNDNINM1SBn
FBgmH/Czn/BVMXRHycTdqXYuMWZVp9N/QnXea45j2GINsV2vf6uTXadwMZZNYj2NnyJ123Neft21
8eXjlObR/7mMPNDv0e0r2XVzaiQCWf5Q5ooQsjc4JdQVAVaQJhIIAqM5swxyhCVgbNsRjaS8KL7R
Ww4wwG0TSoYmEE+k+BlQwBjVkj1cg+M7HkbAssKgPKXNgAx40HQmE8CY4FKEyC5EigPcHpK4ayG5
QrLkfulaxwEu8IkzJ4rdkOJzBakKn2D+alw/OdN2yuy0AkUKIdqCkdihz5ciBTM8cl9frBokYwy8
uYER9mowIYdqnm+NLQnZw5ylN0hhtREc2YnQZUrso7X0LDnroldujJRcvYPg+nhnj3o6wq21lgwt
pYPA0FDrDFg6HbS6/GBn78cv0GcnjOYPlyxQDEKk2UaB557vWd9ct1Vszly5syzfQwWq3x6FD0Wm
JLpTAiVC6+RzXFLSEXmDs+wP988cnWJ4kl40w+DQpVQWtycna+oZgaCixmhAUUO2jMMBqLOUkOUi
SrFpVT1ws8dI3MigUIFcG2GIalIS6uJfBIGysCE/uGzbai8H2wrDkXxarxhWMMKvCBxXddAp4OuJ
U2GzL9O5bk0hjmL85OdeljGi03NCH+5ULT2Y8jyarmZ9bd5iA7rsp2QfAHlEai3fEdIfKGM12qb5
iq2p5CIWZeMkzH1n0sxu1dqiwAVCSu7wnmysVciyZs8VFTPSfz0ZX6Guf1ddxlODmw2oCFBvdHqw
J3TyY8mgdB+Bkx2Wm1e5C8EL5VnkrOk5VOUU46LuaS3SGWBG1zxrkBAw5Z6mdW783gIqD/rCf2eC
v0b+i7pfv78nUueYrt3PPYEfcRr9TpdnqOhyBQMVlALw6JIbbzWHKNym+CtqIq7qKRuCREkq+RXk
Ez7MpffLGYg5ZxGG5Z4LVmbxd/3m5Xqeexer2+fuCpcEiVn5teGp4JUW6AFUjw/W4d1Y7CK33uGl
bi7Jhh7BVYr6ZpB77eecYP0ysEvUqAvva+THp4SkTFM+e9YhJvYAj8k//uKBalh4yARgiVabgrgZ
6YboBUSnuBFemf7xv/WWztlLsBuXFVrP8/IB2Mlq/H3hY8G07hdUMWtQ16AUPEqrQj7uxhb2GTVx
cXlN8Jg7j60bJKj+KV23vv9dLtB7xdM04lqXYW1i+y1bGO7XEWFLzjQiY2zlZ5cnA6gAhABS4b3Y
WpyJuUDLdsXXxJAlEW4txhW5IIQ3C9L2tj7Mxpp7+8Xh/2s/cWN4bF53eObk+msgJU1uWVAiHNp0
oDabgAkAel/7WjsOG7EBE/CD+ywwGdZYg1J29O2mOBAyT0YPj69rSO3/1fFVrgKV1c1u/L5uuqHD
NWeAPu1ETVuu8MrhLaLNF/rdhYK9X9VLD64IF8DjZvjiYZyq9Z8Kgc5lx1yJAu4zk8FHm5uJyqED
7CWnT5npP7b4RLqsdBznkyKLcDie/ttIqx9Mc+8fNeYBusI4CQbL5crG3coVVOevFNFD6gDoRdKT
ExJ6kdn92xW3F4OKhLWPfDu06+9dADpUVlbcSiwVXRR32i5mr0UzWx9Em4a/7RWO6kaALZLjfFIv
XzGlsTHjoGXTJRFerYHQsFq1AmyY733d3+mNXCP0HZ5D7HjSY0o00BPIiQ4NDpHbD8XN5837mNno
71hydMn8cmrJHKDd4+sXGBBjgrpKByIjKfGgiydfXi11UW1Fp8PUMYBKQOLJEfsw6yD/imWH6l/9
8+Tnh/gMBobf62bBl2yHVVBch2rdOaoSg0oDK7i+sNixH8G9AssVPaaAT5vA5LZjbivgbW0ZgxA9
EW5pLwmqf7t0K60buqDXCqfBbgU/W0QpLKSmehUwDQbNzP96tcLWLYC1iCbt+15OiMR0ROCIN1Et
UizgVszOgbRvSS3iEqNwHdiUXxN5bRtKWk1i2i96leo45/OY3FiUP6eZZ/oOIYQ0bK/OCNL7K2WZ
QHa0nXCYMpsqm+9RZYt1RNCk1RX0rIwIQs+8iSyWvXQ+JrQT8V6CNnD7BWGQCEGtr2mdxZDEkgCF
zwSgiD9aPhLwdYmjWy72L/EJoADNfNjyZYTAMmppKwbk4D6dZmwCBkqcjTYe07muobexBf2eTr5G
wrNCzIjTvaFMMb1hjOKvUpGECsPvHEo/y2mYZKGQKc0BZoWBj4qpL9NKcU4mC6alFUHqzKAr6Lgs
K9C/3e+OgttI/7O4Vu/fI1JUYfXfgG4mkKPBaQu2A7cai7gy+m+RYnvvn5+hCNc9W5KOnxh6qgxc
Nqv7snHuDwbjBc5CoVQvsrCNZva3tITXEybT1GFj3HXVZsREs0KPnO3fsLjeWq9Ung14TFT1kftN
4h+eYmFTtqAsFAG53yiQFbdkVt97i4uYXNn7SMenACBRgqTBesRHIyY0Zn8IvNs4iyWNfnN6jERz
oZnhiHq8Ob0SoehHM32C9KPKOyYz+TmbCa2hd8s6fdMbhl8JoWsnkme6X3uq4o24MjpOdRQuehAe
fTJzzsan3Ajtjx4ioQ0dy9a8WIRJSrLZMQk3nNUYU49ACJk5eM15pv3hHoeJRJ+Wmm/2RebmULfE
DsrviZkdZ4zfsMlnAr9XRAXk+dnE8pZidlj2JpguJsCT5GWflFG8VZss02hXfD0HEzpQ9NlzrVf/
CYaM2JTDlVCF8jjjXzq72viSnj/1UhbmK4/32ShsqsoxoKglGNtwN8RfEoG51Tto4awMnHmSP2MZ
JEiJmA5CUPsOY019hHV1DOVtXa2A9idK+Sq0eIkWEgwxKBWk3fzCe3sz5prs+6vqj8tdsCDI7jsQ
5wjUPGwsj0f5/Cb2QNCPso59thNn8ZsraWMgHCsmMQZnRClWVd96RBrxDEel1b2yoz3v8oWjSrcC
z4QvpnX+0vrGKYpH+83WrFuTVdRDvx9yvwJzV5yZ5ZmHkJC5lbxvdheiMt7JViuQ/FmqIf2KUMHE
vgKP5lfx6YGpiU9X53nlflFGeYPFJHL/kjYzfJhSbL8qB/QbgStoeFDQ3JEOpwbs58S4SBkCqRUu
yF05G95iiPtO4WRB2SzBkBaiRYzxiqzV/5YYcTdvdO7H8pjfAf5c0OSLDbqVp9LaOpG6dsfzSm45
0gX3nVrWY9+zuGSzU48aWFSSEmtSJtT8Dzonj6VSBSeyvx7DLst41fs9njUSz5HM+S0OJQBY28QC
x0y/pT2yYozJ/xY3G4Dmo22pfeXm27HGW0xBiofMgnCn+M8h9PaZ4rkx3XoRrKIT9XScL7o/4sip
1LNElMNFYXsBQ3Zm1eMVCEtYRopC3q8u0wrJ2hnIaBwbxajKh9QteZDHyIijuoijFMmYwHcLkKzQ
jP1GIQLddf8pO/NV/K/9ps0BnCtmw5pGFWSTzsmLNPG/Ee8/xtTUv4EK8E4e1FlGHbvBW06NQ+Iy
EyszT7KZbHp9sxXXLcvfW+czQ/TvpSfk/ELWOfBnNxedExS60mMiu6b3s06BKTwKLYlrYnhdJ5L9
NUGiui2mBZ3kp0v4LbjlazbPPj8mid817DiYCwj7F+UXSxgK9kHcfhXJqvEIPcqkcrFFxSi9Ks+k
dQMrR1WsXTs0R+ERsyfZY8evxg163j9HJXcrEMPA1pyYO17Ib5D+hB95o+3IJNWRZCwBu5hrlR84
89st3/ffomSuCqdPBEyxvewFOcugQDC7fGxjIBCkT2PFJPZllUq1sMh2Sq291ZxPnLxEsSzJf6tq
qo0OeLI2CV4CXMErMspX/uvVKJplVxnkS+50Xwzij4s4vHfH+A6KD5uIf0G2DYp7H3rWRMeM39qz
RoLcHOw/lZRGJy8IkbpDdJRkh72BUdQFeVXp5Y2MPPV4fwHvLCxg08UCum4cgmqn5t94jqXlv49/
YxdeOQZCBJdgaWQFAbRyxcUce4piNFWOMUknrTcnPOIim3Yj1kD1bzX8CI3sbhI2LwM3owFq3Y5R
7rca/74io/RD4rXnPVFr3T5KUuxkhUM5ZyYJWJxSTg4Yi79mz6JgHcimFLB1+Ofo3bmA/oCZ2duF
/+LB0na4eUf/LD36Tj6L5g2ldZtTkC8RPgvO6da8YxnOYxN61M/YUJV0fbTevlj8HBVulGcpmcMz
crJT++u6iubJ4fMowNpaN+LCPh+SSFaQPuONbPseY3nBFetxTINEZ/7rgoyisNZtCsebi0KDsYkx
6wzfG3TZM2mXkZ2y5ss5vOrwfVl6BdJJoGWmPRlNvwtzwfRlZ1mPNHj60VZ1PlBH+IEf1cgZ4bqw
KkAoLSqmQFVn9ivFl9jFwukqkHHGl+yBvM/BnwUSz8FHqrtB1yTMhaQ296RcmZJG6xx5KKQXOwgu
/xAGbeJCf+Ae8l3f4cPVfA0QP36l+RLUnn8suCURNyskNR9oWE/0lPiKkqNS2ZuJumiRJUskeZN8
00SDEV7M1HMQaSXy7DFi7b1qb4kgOikH47im3e6ogqAsXqHcKCyHTEC0Ku8IwATR4vIH540KVr+H
omTQ/TA82IfIE8GwulcRAeU9CsXcUF1rBGn+5EFmG4YOlZ0eYe0PfBjUKIzOjRinjBt7n9g2z5y/
nFfqj5Oh1XgHndoRF5YKx25QlZ4EnsZBhtJwvSn3LXTSTuruwnQl9fqhTEPFtSmywfmIp1RXqE0C
rqQqpfKgs4IpunY4YM3PPQcc1Ap3ojE47JLyUwGW75V1tLXeTspfqU5lE1l/mAt9mkQAtJkIpHo4
qc2UeTZpREAmOlwustVOo5DFBFfNM+RM6ZV9WRdygC1vBltecMz8IiPq1bQjHAlmNu18ZzdsqGEE
GE/JJMxbtm7dYZS42bFungYbGUUd+V+DJw+ou5g+fMffonS+9kqreSWJQoInBuioXALEjKPnJKTa
QWKP+D4EknWiIjnQIf4p8ouVSMn5l2nUPFzQZgGKD9uTbPVRWgotF3XJ8TjYlg/EDgFCywsmHfhr
phiLcNePNu1Sibju9O9YoxN3ej0NvJJ2yc/Fsqy1qBgSQuGkgRXu/VVyoBjdzi28VBmPqDpJxyK/
SfX2IUGhvWK4qLSPdzIQdcwWKXEdgqV35nfXRhKIRgr8dROa9rUTPkB7PEOqaf1ZGNwuH2pFbfba
mrPm4ZSctO657n5PvyC6XDxXBb91yAKUMBWD0tIX0ZztsA/5oJQFs4bEcFDhPGqNZLoO0UHybn/S
VvadEWEWYrsZYANjAMd8+GgzKDZD41RJAG+v1AnRF5kUA0THLJaAhz8f4hl0wXbuYg9VXAFSPN7b
PzeqC9oU5E2H8lMAw0AIG7kZ2Q7EfQW/yJmf81ipIPnMniAY9Sm6r0T4IhXF6j6EFsAmiY73MeKa
LqARjrvtoPSPAvhUKKCY1aXodPbheMZ0Km7tf76Bp20PNIbCv2k6gcThA8DaLcXa0wbNcSnUsIGD
SMwY5GEDdwRZyhleZT8lUbNj9qeMwYz7KmuzY+HP0Yf1lrr47ytxKwaMEcox4fgico+noZTAeE1x
h1T7uvXLJzO3obqsvbw87oEFv/zaH0LCmIBDqo1CPhpwDe15CD6gtCyoCZSP5Iden/El/yn4PLs9
EqpBUUFww5fGZVhdGPOkc8fJM3MG6WUprO8cwGG0qZt8nH19/gjq1EhvTeMTnRqI2GLZ7QcskbSh
Yn4hkMUKlggpezvFeGzlh+XCjZ5DFfVBXilywgq2YJeB1jLLq0za5EyAkeDhjAbVzYiYUGmqPKe0
P+JPnSm89H+c6GDAU+fA+DOPJhZ1pBBS0iPMWQMHKamlbMWQkpQgb6KJ/Nl9f9RtV3Q1SJLISjX6
3RcDMnTfYP5x75veGh+96dfZlIBNLmFS6OsaXZ+r2HbEXG2cdZEmL2w2Z3vcOz9YPBT9By03kZC8
KPBuxZcRCObpwRilhvf/ywqeIUfOg35BkptmNiY9JOMP1xJKQyMtDL5MzRsHoGJ3PZ5/semZOwXg
tBu7jXxygPM6gSe6Dxi0mMiSDY1b3/Cu5Qi8ElO63CA92grFknIARHWEvcrIktfq3GumRVYsk4RW
0ZA7+GQDe49TyaR8n/UUqsK2rmyMMuqMDpFuubLDlgCWSDt1wrQwCS6o/3OxbyoqrNrzs5k5VfFG
QT2HWw+IBseX9JmTgsbgdQnv7+FJyqAEu275RjuAfoicXXmJwQQ1/T4yfDgHmKxQRYwyP8mimZHc
IHOLxel5ZDcORUrbX4FcsVvbJ5y8dZkUcOs1eaKM3CwPHR3oOXMDkrg8YMDGCOwNd0bBZAzFi+gG
UCgg1M1AC1kASxSC52Mb5t7N3lLF+0HQenMxQ4xKj7N6VNmBhyKRhyTO2O9jXPAfxkQftyWiuFpu
xSgWqjPa9caWALwBkx8zBR5Gl2Oygg7+Nr6UaYgVA8llDc1YWGVAMlfFR/9b0/jPwrrecyogPDK8
b7OkIYPSNGhQdKJ7CLH4m8p+Ji5l/m3sWumoFyDOK2KusID5OHJ9DCOFEMvGmx3dwve//U6yUxam
m/obrmeU6heNjosRkwsURdeISGNNsG61GCZfDiydrsnEeylyohV8vZdFHcl0ShEm89ulbrw2fjrU
StQsg8rc0YlMuRIQg88lQINFgu+CuDAtq1rkCTW1Cp5s2EIEb5nw+cbXIx/8YHkP+IABey0tMQyO
7NOhZkvsx1bySa3rjja3BeIilbyWruMkim/Xw+qR95yNKZsJd7tctH+drcBaZIoBcyL7TMY+PKTE
giuqCF73raIhgIbeJqm3GzjqcbjClfTJsU+quQraGWK58ohK4NAWtNT4Ghju1SIpl2YQExKktA9I
BwRXdxdFiyRaGs8obJXJ/7aqajgFVp6wVL4Q/TRFSzJUP15EHe/59Aif6nlfNkPb7LdQ8A5hnYs6
ydmY0GgHDww2OCA3BniqqkiEez8ys/mMFNEkxV/YVogwVBsAus34S2PJckbD7xRk+LMQ7SlPiubL
uzb3XiqS9k/mfwZca487J8GIaEE9bQS915yKlGBDTfaoWC+dTSZRROsHyvZAWTxGRAU2gniKqQvn
L7Mxn96WjicvRwX31ko4s/lutgPjOmf1/P+34GbdeMJrWiD+KVahyDL9sQKEZUeZaNeLhqC3+7Lr
nr3yg8psdZUXIZMEfTMQaHRTM+3Y0vgc6xd0Enxh/3wTU+Kkp+Eh0F1rL3KY05fmtLfExow0Yxo5
aRna7MASL0Ux9gh7LwSsyTXN0ND0eeQD0iAK/83MQSACiVs+I3Mq1lAFslGXjrI8sJLWFI1So2Ux
RHY3kLWJoUws2y6VwBuqznpq2ojYOhJfg4Tm6BBfShgdKTBuAJnZBhpmGNB6WL8ZGouIZ+ovx01Q
mbldnmKD1q2/NbAWdxsK9lehhhM5EdE9YIfQwMzkhgr0r+CjiQaPxF1Bg9Ph2p7vlCG26RLQbdMU
GslhSEDxqWXyPKug9sVBkC5/CHtgTAon79rgqPmPHdabszg/cXb/bNNWkalYfz7OXB4eTTT1IJAm
6vFne4PojIyK+nyCCTs4N8yZQ0YB2crogSvGA+Z3KHIDJyLSop4dF23Zj88ikcYXo+oGPhN3qmCT
redbCpNga3Ty5A2Wqo5nTa51k4LjbhNaI1OH+eQvGALpUEmnkBUqCOkdfGN+NK7jURTj9A+4SJ0L
fReM/m111g6SkBqgGzp7amCIvGKvsKL7KQLC5VNrND9nNj4ztQolygJ523HW0dGAiWC8rTH2TLHn
TkogO/YAIlFS5lNFHVsK4Oj6hphVHJIJ8q0m5E7LnKPh8n5gXeIj2gg6+37nsQMoXW7p61buRCcM
vQaa8ZEbMZMUAlGtxCTZBAq1IpAMFo1twIVJ8zo66PtCcldvXuD2s0kr4pHMyPGaoCY46CpAVaET
pSWDV4GE0rat++KcTPrENS8qfGyEk+AbcdwxEBwEoAR3RmjavwkNJYYC9wfTQ/b6kaFqxy24dyf3
Vbp5O3BhvzxMARYH7ajCKk6G5bKV/JC1bl48Zw6/dyZXz25JKui9tbwZeEEweRvsse9Jz4aVHM+L
anpjG5MtDyeW5XFLzkD4ZdX4fjdolMfO+m6Yr9qbJql9lz730YguXlpeHiijKpSnjM3jJJEz+N4C
nCFiGu0IYFucMSCmX3ssJlvU6KXMY5LgFaAIJsfupEJ9NS84q6hdDyjoNFwr+8xqN9PoRtm8+cbv
k7ZABiRlFg6gRjGqs9XwYXVPNf0lD90RD8tLqQxSozniqJCSPNo8qdFhlbOVBu6QB1SOQhQVKJOr
Epr0hu5J4hw1JABo86XW12WI4lH6AskwU7gU0jMF1Jax1yVVpvwmncx5meoQPHVWkWl97X/LH75H
Y9xgz7biELPGdlkmwkIyWl88UxFlbTssRAPCmCQAjrk5e8+KwuNxAPq7wAp86zfaQZJp+sG1ILEk
7KYfNKY0snDrpA2Q0X5E6+WvwRE3vjr1i+EFtoTB8nM1f4jwraMvDz3hTaSHuNRZC5zGHtWj+ndn
KdpoNKVY1DIAqlyxCK+sPvPvbl9FGMc0OEII2yBvYqfifx3nRuHDHvzhPEqNdwZbwhlD69EJ8+Ml
GLu+yb4VoEJpJNa+BmCvnrhSvh1R02C0QUsZb7PbPPLup1FI04MfJcV8zDgAUwGo/GM7QcTtyp1h
1hFl7hbcKWaE40ta/dS3WnC1RMDJsvmIDceoRNEf8fIl9dr0YojCxzpc/lQ2fObB5nG/bnlD7bPW
IBK41fA+TIdGvlVXQqZmhS/I4QSRwb1iX1DKiuNCkMHEusyKfovzJwlM9xLWLcfvrwjyNskoqcAv
s9jfa9IRxLYT5V8mj1+/z3pZ78WdAKxXvZkWZenGymLW8UEShGXrcgdRac+kE57IqSrittsD4xZR
vZ8RHO2WgD2lcQz2zn+/Yv6CPcvMzkUOKZK5xVZbCohP9vT6cKXaf16UC1XDh+sYYhlfJ6HJ9OKt
qCPKC3HBc6kjoUKob1H56pxlRvRvoZ1FdPvI792cdrgkaPEXMxK8IPsbX6mXssy8n0F9Gj+kVneh
sdA6T60g6PCfbMQaagLOquTTeLHFkhXueqg7lkKJvrQ50DRwiP/HbEK+Q8CbQc++rhrbgUtI6IAc
DXIDXxt0FdqBeO5gACm7y5E21RCiaKa571W6ekwaJpa/iB5SRpAJQEbV9rHYjU6aNg4OWlYgvbmI
UlpmPeyQT82Hdw3H7ZSbHcgHaEdR1LlEU908WnYrgYW6aXrIxAvgcHMggs919HRc3NfRD2KJirfp
QxSsdpjK0EEKlGDeCsll69QYobqc6XKhukTpcHwHw/HiApr/zC9XpJmV9gBz+38Op6NpVKhBkrZc
0QQiOERwIED0IvT9AnY88oCxH9YaR60H6eK/1NPYGxq2uTMjKlxq9u/1PhRH2QGZwWDPA2MuCnHt
hhJx9F1yvbKATsj39zLyPEVVMlh9QipNMCb20OQhCrgwrqKdpAloEzlxSPb3mkzKvO3iERRy6LOR
/MwK3ujRtGBUjlXbK/E37Kp5c7X1AD9zW3G1g/lh7dWK9tm0S6XxmeszXdIiqLMKnVp+lHmGZ4Pw
2HGQvzs6YyBXS9qrYqS2WERhl/uT0YkRFR4vg81Mi92Ok6tb6KVsfrnLx4Cg/P+8TkZo/lYFgejq
C3Wt5XG8yZcaSEnYmfR7TU3aEvVoORmYCMxjecJ4D/B9rc+J7BzDwanf8SIQNL81gOjWEnBjXPUP
gKJNaLbtnKj2BchEWDnhALVTaOWWeXoike2LjsMtaPxCA93AYb5s+oGyQLXz6mR9aJo+eKMWikK6
f5aoZ0GFkOyc3BlwWWt2kRv3Kk1atEpfS0HWdYvtc9ToOo+a4WTGdCQSIYXVovvQbBUh/dJLXU+x
UvdN5wr46IAzQPayRyvoOSU7Q+7hYQdN6AsjweGoFuOyrCS1po8PQlvTS4aBOLJA3SZgYuClUjAr
v5gZoo0iy+AdLfmgrzQhNeAs6nREuCwpuvbQLL1pm+y7nu1oQbr6uosWdj+LMNCo0c668YmRPuTc
JTVl0eJKNAHrMHjaC6ciyQjHfNIPnABXUPV+C0CnjLQIe24bJLvaKHgxyF9JNduoxBtceLyoN0/Q
U0z/LzDB/1ilQcNMcyon19iswmNAUbiRvgnchWqnU9nzQ4sBL/l15GibOE1QC4f8bE+/EhnJhxTD
91PtLMuHmglViMDcZybCdwnMqtHXH/d75FNpXvB/XysROhPqQfn61mfe496kiVT8p/Ck+bWDgV5v
JHTfJTFTcyyxHlXZp6CDtE4aHH53wAddo7v/BYWe9T5anrYHVJdbBfNLNTQYeqjikxpILw1kHsmV
fCBLNTPlPmk/hKDagbAZKEGQz9F8xtc8+CgtFzFHQlsI1a6f0qf1780+bLpsariY95TkLImdgK6N
z4Rr1iQaS8R5GHYiL1bIxR+G5dCthFl7joOF+GllZqiFH2zngfBEv3rC9XBGL0IeEHtS8nCBujMy
hymfhwV+uNj2Brxofja0oYxiasZjYitK63NzNU+jl0yc40JkdbcfH5laVO1TVz+O8kiFdBbBHyUJ
oXU/QAO7OhyXRjEyvMpZUrHWTRcagItQXQF9IRc5nVL84tNcPeJPoI+cD9ZkEH5a9NwBZ6kD9ec8
U8rKlRdiCxiLND1DD/fH7xnQoEqCo54F1Ah2BZ9vcPjOde8iVBKWEVArWnPoEnVQA/ODMi1TvjcM
erkN5x3SAhZJK11DfVW6CM5Z4+t340TJzefuwWbigaqNJJTQpxxOdlnkVj7KlNWwUVZUVF7992Sm
MB4CuEEYDV1eziIghXk+NVk8JnzFwoUAVtQR0rPwuYhQuoPjOoDN9lkqI4bn6DNiQjOCjeYK/1xS
zvGeZjJM1f6qxPW5IkZmuE7undifl+YVb4YMD8Oe7KMUvJMVBOQaVH8tCE98LWLcG6UkD9O9i+zC
pUuwDjPXQzeHlmPdOrRDdnArq7+zFCk4slzT2JTDCwPCNQbWPTk/fwolsPEyLIEUDY2VXl+Er27j
SazlC0MSML8oHzmr1Cn3+PiX0WakGKiUQbu+kyh1+bAU73CJi4vILyx09F4g5AfviUkSvEy15XSo
P3cWBv+cNdZgYNFo0P1NJTzCV/Waq+5O1m/pAJDmSr0HLNLRlEbvBWSbvGpk9WqxDpCOi2eRWj7x
gJzFg23RgN5j7uHz/5gqmhwxBFm5huSWtqJKmDNaB0yeMjeJqXxKiHRkUBuzvUXmOxdesL5MtznB
Dlu1TCGQJ2z9zb1OBpsPRHkY4099nlYKEXZ2uNmzbxYF6snnp9OEHX88APVFlPitk8BtFuPXLamM
NUxNXxuvcrY/NIWop3tMTxYYXVt5cPYIU02J+CTSp/q2k72iy1fSAnZHlXthCsGc8K6VjjDCSwvJ
ozmKaRKXYY6mJ4xl8iXSKhnihCGZ5ZILz9ERIwSKT//rbikhDmibTHfUUaPYRgT58pbxTmZMOSYU
nY7SKji+Z4Z5mI/SvoI+/jMkNLidxA+hS29QwjFemipyq8kKiXCkYJ8ELKsgKekA0oIWnY1/jKxO
t7D2hHofqqiMTxW8IO3aE9trGa/9zWsujaIe0UQ0bwInbp98iaraLdzjf3TzwEsi8j5F+7g/nQVd
+pf+RTMTPHeux28bFhg3/IkFxGh4xz2pZEG7D7d7dLeklMmDGC9u2me0/q+3ECE6U/qXdNL3y9tI
cNtdqb+U8F5nyMSd2iaCWTeEl32PjI1PXjIhPhnnTBZL9Wvjps8q4NcFNYJ6MW6t38EMMugp4rKi
MY1BC6WklclVjg6WfXkKJFGKscUOZsAc7Ji0pRqNLhyR7ki8KAWz0d8foBdlObIDsCoN92C1dOju
9D7l6QN+D6DtQ7NklbSHt5OxqW7/AFBiMFgeXgoFXCxADNCDaCqe3DtOa0L6t2hmW475dRBlTY9l
rvQoNI/cDXPWA1N6Y4wseLbWqGp0uRcP38g4lO7+ikY7iBaRh7toRkcp80yLfItCtJK4vGmsuEqA
QyHIBY5fRfsnqrYvbol5TOufxEVZOl6lRQznczpngFbUrxxiV6Awzx3UJPN+M3zEvO23JI4oHdkZ
o74z1T1aP7e0BEHiATYefJtmOnk5mAcUsfQ5fde5q2uDvS5tdA9pvpu9cZij20RePm4uo7BlEBk3
UBAWHMO8qEvff/6qyFfNx/EpPFUrHpDSlpClp8UnUZuoQ/MrZ0puV0nPvEvz4qJqp8hiCudB++ei
LLHhHyjFdB6aXVLWQScnnrD9+sf7cUsq96wuhUo6IT6GSuAbN5ShFPOQvFm8vz/G7bAypukbqpk1
mbvkStGOWgFgF+0iXT+J8CeVER9AZhzmPx6rFXraGD6mo/t3cA8ZdpgzLyIZ/oa7GjFv7KFi/Aol
bn8yTDXSVavJiNmjGJNzx8s791YBAtEQYjOqE6mtnVV1pTpGoUF1vC4ftVvz+jezi+FKqzigFiYZ
V5h/NfNquVLAGKBH+K2cD63jdVZ8iOGs+/Txye2Lu0QcnONVNolTboFvS4TVQPeenMl96JE4e0J7
NQpjzsQMNVk4wDkkMTuGJyEPLU7X3hpm3U/OL4ePQfQZML0On1mR3uWlMilDYqOu3wu59aQzyisd
uf8P84e4J96tZCmaQ9SjO9LiGxf375A5FoEFzYcj8WDKaUpELivq334/lYBWqo1YRtqWJEIZE1H0
pzxBrCZix3TtN1c4TsjLFnifE+Dc0CT45NfnMgXtTurbOiqtcNVR96HD42f2PujD0G2pMMiZa+X8
XNWm9hdtWTiUn9v181gE6V2Edx0UbtXzDEOt0RFlgguvtKfvhAzh9xqlWUWQaEJ9lL7oukDuV0s4
+JpMVuIHvnj5ANdlUV0XytrOdE5cM2+tgAjHMor+MRiVIZJNHiJNTqAUWY2mSrEv42XQLYS8DYTa
KrcM1cVL46zp1erN+3aQsDNBhy5811Xbin3eX5SdPk34YsBXMvqLI8mc2Kkf9DmrViXiafE8ov4M
aQ7uQzLEIsC6qwBq2JvZ0I8eNdUHZYkBJ3yayjrPkgdmNAJjmPEMt8OEJj4IFlP1jHN8j7svwDks
5J0tyfu93UQn/89oM76WjQOW2K6tXfbFoCUPl66kYU2eB5C46TCE4WGmoyAeJcAVTynA82MCERLU
fMRYDzFSjj+U2GTxNugMEplHR7ezhBlFwbh3mlP/Y2fEQ7n6pSCHFSu6acNcaR87AXCLXU2xzcOd
UFyeNVEz0eMxZPWQRclBoznZD2pGa+RDOtMN4lGwj3R5d+dLoMOC3kZwqcLNkBmh3NJqQ3/MtKRB
pbzFad0GgCBkxufwBrLpGas4P551lpSx5rOjC0QDQQPsG5FrWi/1MeRrVGwerwIVhIAFZdidZ3Qz
i6/59NQ2dQqIZ3RsBMzB7AV8ilU8RGZ6HAmuuWc7Vc669Je3mwpuenYpySTTN9E13VEk2RpNFDFd
SgnaDRVZH4FzfFvSAist3pzR1wDxtP3Bum4/pJfHiM/K883Mg++v6AOOhXWQpV4kO+RtqlsVtXqh
tXZeLLCvUMC4nBdkr5kjYCjgvuxfb7PkjZloxEfATkJ8fb+8O45ORR5hwY7aPaV1qs7xrobwH8A8
ShmkcH+TcgXjhqq7Ce4L6/Ipu1bPJyhG92D1jbDjOU2pdSors742kDH8zYEQaQnq/NLJhzbckI8Q
kgisdaUXsDoMJq2LWjjiuCoifRuxBg6vg60iUa9lpmbFfR49t37luIQhuXrUS0wtI6Fkrriz5wBN
0rcIUGdGn/Rwnr7MTp1d4b5+fYcuuljSRvxSXtqzn2IH523xdVt7gOzKI6td70hFScidmMfppgmF
ODi9bBvqB6FVLMrmJIUrPTKOube2el1PnxkzuGQum0/2z7QuKbSZAxNEePryL7cssvzRp0Fc6bNS
trvTVKmikpQiJBPj4nAQK8AurBeOafOayQyeIPdiZ8fcKYtfc4PdL43KagpV9hPJZM49Rvg4dBRL
Ezr2kuU8ddHJAkSriJZxqQTC4J89jH45I0CJSDx/vftrVUtXO35um43cEi1rWHbnB0wLqtUN4qVd
3zJEM3YGCXM9fZF54Vws7BY++ZbsFouwFAkMMv1oS4IzfiasRZlQwkCbm8/LbV31bqRGUQ5CFbC/
WMNMn0frIBo5mwNONNtqF2W3gT9Q/4SPk5iAysnr1/2yZIC+S8tJsQMonFF3/JYEO0sydE2u/MIK
bOKpB2qcGwr62gIQxDMT8MVrdZqhgM4Ih1wE8YDjfO7+HKYm5FqwjlqqhccXXM3ssp9UTh+WSX6/
UJNt71tGl/kUt1r6kQxJRp0Zs3PqSfBgO2rZknutONm1e0ZiQwPb+Da2C+HazJRxPsoLKXZX/nJY
VIpLY8NFwyje/MBsfNvX9e9UpyagARMNyDna0PmNI0cct5N15s4xmex5thxrSbjB6gTgfUrdKY2r
zAXbC1fHMboMTz8MKfIYlZXYZnl+I142cunJqKAIjlTBZ3qQRbtZA8Px4Wunl45G480pgWgM4Lvx
lkXe/n7P+WQPWP90Fmq5rWnk8CwlYBqDQjuKso6ykQPrbaXaEbazn/nTm18SIqbDI1e6+AAiEdjF
n0CPTWUmGWW+npMo/3T44pCtHe/qxeBm7yd+Y0KjLmqaNGsWtXoFEE229WQVJftHsSO0yVzdhCQA
+ZjkdhI6PNbxwkw05Bagn7Y5/q9igxm69QeHC6HtuM5yPw1MGUco1Da+egkWsK+xxpKBMYVh4vqz
nDuPSNFyAi3edUBP1JC1Qgv3/QMPg+32r6UyPzj3H/FVlflOiQniwmgjYGrAW1/LeSTUp/s/xFZm
NWett+F3WYdF1VcZXSHWRJ4qmCvVYMvc5+atxpfn9N4GptjasuWtqAqxTgwtvAs03OzOFz/1xfMv
drC+Sm9i1hmRhFDnCg6CD0AkD0gG43/JRrkMQM8LZIACLBTx8GzSizm2cq3mKWy6TdsFbdO/AebG
m5QDVQCKY4u4UrLLHvbOP0zOBy5lI749trtJ9AkMIac8k0pzn1QxKlYpZLAHU0xFah4B76OX1aAc
dTcElFbPfRQZ3cuJRTX/IcPe0VAqTZlT33gf+0UCFQaDlIWhk8lulQPYiCjhRLfBUE1yk5Vdo8Wj
GfU8J0B5m+tuNaoSVm9eZcib5oSDnLupUwhXJQUKfzGVOlO43hB3saVWWg7LN8TohmCKT7N2V+RS
UTkKCtXjn8U+rSMwDoEgQJk4KU3B4H6+7qgQxM0+18BejW6solbhjGSks1UW+wMRgdKhaVlo/WQ/
TQJnh37/XK5yDTiacdxsLOOZ41ftVzcdRQxkGiJ/sPAmosg22SO+P9K08UfbXBgp9zxarGweNiP0
nJYj8iw8DhO0P36fXfitYA+MpqXpR6pmkyXezJ+TO95sTGUp3xbfVhWTbnHZwWpN/HVLmEWRZ3il
R0eyzTvZJN+TKEUC+u8CBThxwAK9SKTqmQ+p9J6vWW3LaKyQw7Lic3CFMitd/gN0hR2n2Wr2ikYq
ny9btbDAp/Gpn6j7ZnOxWVFgWPOtG/QvjsAi/j2RwURCqs0g0Kmm10x7R8gLs6iUdJ5jaT0mM80T
v6AopeWCoe+sagkrFSARDBrJKpwnPOm5idHXy1H/jzwAj4ddI5jBBEpvqTTfAZYHe9sc2hBonpwH
jXni7y7xuzTjTbtGhAbxCyGbUZHJkmCKWLa/80kUIpbvBugKOt0yqHn0bAksR9vjQ7GTs8BZheiR
U/jSss9/8Wu1k1KQGzU56Cc756yVwtxjAzx/WTTdkBblY1p6LQUkK88J2Sh3rwIEz8mtJBQFL+5r
d7wndTdMConzeIGmI7V3hyL9OJ8xI0TUdFhoWQN9d+VsVrQ+QerDHjw1NKGOCoqkaa7NtIRNuQnE
X/JWVFiV12JbwiuTSv/bt3als+C4ryBnNmNFsSVzC+E5bR8l8exD14MUwCf0QAtU4TdJmOsxd1dT
EjXnpOLxzvN5qcktc9L8/Zo9uTXTlkR63vf/nTFunBzA4/nFW2YDBz7iNh1eVXuMLjwNIrGBv0qZ
Nf42UBT2qMfIkyogW6aqGrncAJRhcRIFPrSF0X2vt81Q0QVkMVa8VucJntL95t4KnvYJMoOZFO/m
K5EooJ1drRQcnRfxim0dFeU3hcNtItaVGCVAVKVm1nS0F7oyIJYeOUKiE4Eo0oP7VWlVs8BWkC3H
oEhkhf1zATkOP+idJj6grhKSc8eNFw1NvOUETTyrYm1Q/O0oq4TmY+nP8/IcbrA6QdD6Zz5dh7ag
esvL8cVQYHRjyN342TC7hh9R2/h1D5bffcxmKqTgXWRyDv6h/79tdLOHR59ecA+howdDJjAXt/gI
oUAcRZZ5ZDsS7i9A5l6JfJSBZVC+Tt11dKGoOOHpSv0Kme1cslA6A/5Wvyp9QSiG4LzLvu2HyLfC
4ESj+i44NTJwCaUR6rvLfrqKR0CY2iV1GpSIKPojJISdD/FTOYXlcftQzRPl5eNiRAXYGbeH8hmJ
pMef/GGVPqB1MbUmkklzhKXy8tAeJ5t/0PNp0woNPqCOWNuWZwegvYtGQ1BcKiNxurkG6YBTXQz/
FWzqwOY6qbqg4kYARPkvzIKfuXIzvZFde07c+ERv/Acekp+xQxhnV9RB5RtkSW51wA37kTrYukxz
TJPuTryXbxks512ldKipmpEDkysItNQo/+yAC9B8ayeJPYKiFLN+ywUvEGdstnGVjXuIl/NOELTm
0oz2IPX6O1hdpgOBAxyIcop0FyvAeKzccyySyFhaGfeeYNcbUKoj/Y4VJ7+s19Bi8yNIdCBYRBtH
8RnG9vv2Wio6CB5IdP7jgMGn3hiRXgn8ecwitprwqutDUTuCPCPeXFlL0Fik8BY91MsmCTcocL6T
R5048D3EPBD01khm5sYKz7pziwFlmNSjfBABR1gHyHvTDgoT00YO+GHj2vqJeId5yBKuIpYMxvC3
8XL0Q0cCv24QE2g3ajs1x5wcUZQBB7uYXXCY5j8pFv8X+RrLVRbYHrxYSX3If9gEdFLpZT/Peo8t
e1l4bb2qaaE6mdmt4efjV3/lZFeGLxiXkBMbYyc8WAOwEiUhsRhC4IQD6DjmZLlpqW5rPypEQxap
cqWbAxBh+qYIyQ2AtoVs6icUcVZU+u8sNpZ/g3X/2FvjjLBEnLxWGX0Y7+AFfTir/OY8Oirh069/
ACBuiI3K9wSwVOum7YgUDhi0VeKq9oVIoGPWCbeq0vcANiQiiw7jPWQtVG5csXIw3qLHYjpkgrTm
MT7Go314Mzn1H7qorwf6Q08uQ4rsan9VvtmaB+CE39o0TY8k6jZRJoyiwdh+kW2ujJV32r22nyEI
mJh26r+sQ0YIkdvWvZXJFAa6WxpkMUURJnplTf5E3MPS/z48DsG1MbmjJ+EUrYf9JOxmPgmJWiLf
RV3BDBh1Dlf4a2eO+XTZJeZ1OiyVaJ6VkwVzj9jJcJmrT1VctV4XZBTkPinJentX2jei7JuYb8aM
GFyzdKW8Fnn7hK1ntE6L2gSGgjOAUe6c1k8WN56YjlGKzOvRz3oTuh9m27DAxr9RUcP2RywRd5mg
McoW7VMYpdWQD0/lrwlNgzeWg/STKslx/Iu9PCSVgLnBvtKf8rqpFMZbi5hXZ+/itHhcrtqhdOi8
0iWhjzQKJjWRSY4zClDcR6UMtJ4xhPli0/IWIvnJicGA7P9O1OnESabim/UewTjiOQ0E0M3iDEcw
ozgNfPNutn/RwaAObAjQg6KpKpvfAzrzAeoP41CFp7PiEZm0YrNDIHHHBGwKefSoPVwPyr9cIE/9
c+ic/lPYbxiCl0V0Q5eZfh3gu+psYsvEKG1+d0xaA9WZlpBouroquBRm5YsWPI8qScNd0w1NQizk
EPQ6fp7P2fv4bFmK8TXNoJEdUNTqwV1YHDkFM6c3IfHQwSkFIcEA8Fokzf89oAO1STNq1XYUErDL
2KVQmh0c8SdAjQbnYzkCpN/zMDPt/+UA2L1E16iqw1CI2T6cw9k6pCzKEjXUiUNjmLQVc7Rl1C64
vyiFO4eYckHX6DF8S2wtQ5onKDxjI2au6ATvIEmJ8qLZlmnL/oOaVtRrAn+c90GS798zF0sfoZvr
g6AXn72jhUVuda8Gs4KiZoSSka5Lkt91h9gypbYYnqObKbFF29MOLiAeJQW0NAvd5NGATKFpfmKE
d5zghUGrYx5yozjUVuwc9DTSrJ3hxA8mZAdUkSORvrAkSq6iCY+msr39Udkz3ri/uBxDHRYO+ApQ
nNuBObsKe53x9kx4wgg8pbRNN7ixL9ysvuADIAuGM4gJpRaDmuwK1R6u1QCC2SWj/BGfBgxR0oLb
gebAl1BIXfw7JtejfnZdqj2R3tPYq721YHguiVR6BFk8sBgtcaR1D5kgjZqYP/s42pa2ZixvxFKv
pl76xS0LkmG5wjnHc94XiisSnIPl7Jc7hpgqzArURExr3EY57BGaj5qBJbPWIaLLPUBXaxwR07dQ
O/UfMhM74vgMsVnWI53iMAhwtqbMaY/YYSj4QJOda7the1uOjbJdQVK46lBtO1pRaWpoFkQftS9e
vHLSH/7mnFQUpyF0ISZl7sbagmQI7Galt0ktkbBx2CfdZPq/4JDa7puL29FLKeGuAbwE2NEInMoi
L0U7zmNR1nZMh/ZrenQe3XFJy+YCNTDD110Epe5a+oxFTTHvwvJtLI1PAy3UUVpGwYkQITUyhv6u
NT8DWfPRMP0TPx/V38CkZU3lmbR1ZCc7ZfvU5YP1qu+cLfzJQjDqqnsdBvKlU0dlm7yyVpVBlwT7
RLIr7Tm+K7jEufHKqqxI0A6ba78jFfAhap6vHC14lWG671nP/UJGht97Y7mIHOqijA04BpXyP6jb
6D2CLX2B8/V44i4NyUKFaHbnpw+t0Ql3+cUe0KrEZtmgUzHEhGFujK5CK5hh21JDbvPe48XNJ5AI
si9oMCxV0Wb6N6eYmmto/QnmLtiPg/JC9SkaWpZ0tSAOClTun55wnCd+FTnicgLaLUhYOcOaGWiR
L23YO6x1mCRQMz+ZJbVRqRWqVPuGWQmBQwjzEpvGRU8K8SvJaI1aqg02dTMaTDrorO5odkOuivh3
FnvTpGDroEO4Tbja9jGb/a99lISC6Cd2TT+DchaE2Mx8M44mxUi4DEslbHi3bpaDC8QvPf/VYfYH
+kAkCWnHSnnmN427P5p5xnZ75vffU2JUWOhTH+GZUPd6FxRsGmT299JiThRCmmCBoz67bShdUYKz
EI6A2rpknaNMktlvlUVvKypifv80qK62YGWfXJKIthYWDrJEF2QW5U7KEmK9zdW2A2LoHvzVrGBw
5h8cX1vubA4sjcobiZn8xY2t9xhq+sSmGNOjCwmbIVSNtR6MLNM35qwSfxIK6eM3SvVu0mnlBu+S
5vdbphasV2Qt1q0vCmtTWr/Znr0h5XwyvEgp5Ev9GZ1G9+ew9kGIr78VY+ZHiwVvaFB3CiQLM3U7
nMGhfW4+S5Tdtfp5HgrTommbGiXfr6Nq0efLFp3YlExfwHH8KdcxX6ytEXU7IP+bwSQcykHq2fyq
kBMZTNA5ekFLoF5Nj4pbfmxqJBB+d+ANq++4/RXv9qF7/UUMqu+nD6KZiOWvgWFj20NT/2m68s5y
aJtRHwyFAi6JavCiUBdNqENazYrN/+S4JjfCcIPkg6bcydoBgumtXxeg/gG1FgNHsqMrBzSjXMxe
xryy5vbZzkcxr2UDKhHrMOCRkVVkKVhiSXxVsrlvnEhgY8I86zBEr85bKDqnfdw9TFZozDL0CyEQ
Wvd1A9Li8AyekpRAwH7qArYokNNDSinq3DrN3fATRAaFPaHgbiigKeptEveR9rEGscgiWsJ4W7i8
YrOGrHnj+zaI55ORd6RjLg+23IVFfEZzud/2ViL0aWsH4Zf0VK4/AeLDR6x/+76KIWmC0RkJ6uIt
aMlCUNj0vNH6RRC4+MqEk1KFAV3fuOL3kZujTQ2dIddWN9kuKXhTZOyxES9ZSDCVQ/m+pznWqEIk
YmcRTCMWaM2u1lMDv73il4sVqmROHbF7ObFW8/h9406hn4l/QHLTc+7DHocoML4kxLjlvuxg+tAw
gZ38zJkwtFbn58wsGOz9edIZ4ATMmSeg4QdO/GT0Lms48TLu9TqzHmv76GrXw/5/FuO+1S63Qul2
MzsN7ft8PaIcLLO7fKv0np26v1ll27kESkAtUr7Pkj3z5GsMqVOGdV06ao2Ple5fysUxHCVYRBua
U9ysAfifWg6MqH67Tdg2R+sC8hb8HojmgYeyqsVImOBYYTPJV2gli9gKdwJk8TjGOiO7VNFlWQvw
H1caKVqui2BnTWep2oCPNUqmi5kAiRzljLqjw2XZmWo0m5c5bKPKjhR8uAJj+sQYSLNDjH/bQ+Bu
IMeSU2qw/Jh8nMmG42BcAvK69Nxx6eGdyl+b44uD12rUfNUcxIhZeYkVAkoHNH8QWbTXE/jVyQ94
xcQMTr0JizwTjdT5zilvIC34pYECXIQyPx3G8NOSF8h4YhwOmkudXIZwqVfXzTm0mSh70NmcVL25
zkoldviuG8TiuzZA5pE62hdqPGi4GdD1NXTkguBkB8ROk2GsYJhEi2vR+Y7D5m+M5QjYcttfVLts
xsKGu33Sq/vzn+rzCGtyakk/qUJHh9cWjNSoA1Ed6AB0vCl3XBCrqAdhMPa6oT5atkKkQ/IflbHC
cpzw8ojFcHhYbsfXM/yM0jC6Axv8C3j6UGqW3Di0Meam4ypkyF5XMq9KBGCfNXeEEA8i68JP46RQ
dZL95P2LVnirSrxXAS1vYiXRaLVK238QiLkdP+vpTUhf3gYB+Iftqjl2BeISgzfyuwBEhf3kczSO
2Hdm7PDePIAG7H+8JkF/NZldGZ1ylDMtr22NCG8LmkQtOUlN+VuE43fHS/MkQD5kTpS01iXT87Bw
6CN2MGAw5f1APe37hdGCSVtzzsCtkTQLfUZpOopax2kDAEr/e9ijrKKu1uMf2TqfKPqQ9byZ323f
0mi76N7AlE8sl7xIipg6M/WXxhlvkLrg/QHhkv64KGuT+Z0CUSi0q7oO1C7xg6NvU1w9ijPj2Iel
rsZTn9xhg/4B+TgKFpKUQPICloD7YPKA0pURs4MSFxj6F/hFpaNa7cAtODKjDqSpKFSTU8ZO/4qa
8+9wnvimDhh0ok3dTbYqCmLgdG9HhuX9nThlTPWt7Nh/ud38FBPu7Ici1XlCys69UtqdL1OrBIP5
OghQm/6ady+PmnWMZVUTtSADWNZnkxMrM8I2tjvHQ3Ee2tzl7UlWlzojGUPZivP+86oKglaqnPEy
+q8pgB5tfwFOpMDeaBal/+6XbxzWmhh7+LnRSvp4/D/q1LBPn3auDMgdWwbhN0Dp916JDnDcmdHj
C+/XxxQO5T0nIv3H0R+LWoNxagueqy3xdHbmq20Hhw2iRzgG+FwnL/Z5+HbuuyvuWEp9F8vrCo+t
5czWhrUiuwJfyYMdB6ma1WBnLkhiSm32gpzZJQyWrC7HAFlexwKRdYs2RhS0ydP6/CGy/siOqZR0
3XpPPFetQI0yykvy9JxMy6IgJgztVBQruHCDbWwdR1XzrJdA/AS1gi8wJhtEZCcfyQZq+SYiJ6DL
leWuLpVfP1Y4fOpF6eUpZxbLToCQgoQU9+HZWx8CMr5+ZNO3jA4anrIxV8FHsxtCYfvTrqYjHzhK
RYrhUhTqA++OLyqYYEabnynfk2hERY3/yomjh63+Mz5wumfMzS1dokm0WotrnlfCDV9yrQJDBAdA
+GqvvJSYNrG2HYGSNySGGbwxEwgFwabNbvwSXeqc/Ef89LSXTGIfIDuRqxPxrf5eFKlqGmtjlm4V
IKT5sLADHvdH4t2p3EhuRgtAuW781dmJwWBLdw8XPHeEQiCdKMhTOdt7H9YVPBB4Oo/DNRnW3E/t
/a8VxhihQMJwiNORT3vXYW1uIQG9rupPcXAJwPYPN74LwIQ6M1EhXoVTMhEJULFXl1mOG6Q9yl4o
v2tschFn0rd4vZp0lO4FHVXlbpABwbMfM5XRFiFcg6djJkQfSEWj07Kq6SRlrZS9wCPSruqQaTFZ
JlUkH9/fQ5dJSSMQe5cFZIrK4UGSZS6kOausnbfDxS9O7Ws1f/E7xa6qYxuKwkghG2MbsszNaJzO
2MR6qhfQrAE5FhBtmFeOiP888u3UnF4i8m1P93fuj5d4dYJ85CsnWg0b6s2LJ30O17qhHPfEsGLZ
ABSqM1exTC7VlOeKKe6fdV/8vdNFxYrhTLSdnhoIP+Z+2U/aK2w6a+aQLnqdMI2RF08NuL7ZLwUh
YqTBCBgjU3xyyBU5lohrd2Sw9GNzDbBVSbD5lUWbqLvD3FNvBuoF/AFJ+H7mvmkpPJ8e2Bt3JrpS
whOuMlp1x0C9QonTvWY1Lr3PjPUWIxSaMJmLo1raG8appROxca20suh59ZuZakRYqk4zAIBhUScQ
5/cpQ5EUZ6j6IH/9JQWizbnHxsApruy35wY0q/oSRdDKJ8bByu/HThJbg775kuY0O0x+jhNYuStk
EZNrsi70gbg7iqo2sC9bwIENlVZqszCLfcBgXbHt1T0Bjw+q1731iHtPq2s5c6FD6FBhd+i8+eE+
RquAlNApS6vms2QkVYGUa22A4MstrTjM8x4GudbVUQvTIaLIEoTZiisgETJO9SsvZ6/VyghhIlT9
4/mzO6dJ+nUBao7SuVn+T2gBwTvRG34QqJ0WhnlhPU0AhL/X9JN8OuIFJn1DqjENCfYhw/Xe5bOB
sywNU08m8rRIU6+xrgbSNzhOrt0uFT68LzkcnalnCGRBvZSRL7aTeVba5rLkRjBuOGvHYRzCFjie
ilTZFZVSBlwg2NiIyhPR5Qfn7VAJhzqPsteUGVAnU6fmLTy4FBatBbYsKNhxyGKaXPyyurraAw4C
RrvQIIQnrNIlnV3RLRcWon8hfU9ARJO++DAsyBMCQRFQaFV92+UlvQVsrur818SCRRui2QkGMBRI
WQigeDmkcKeWSOYfBsUCAOKWC/3c7Au3RRUODscm/BvRQVaNLzNCQZ/CZhNTb2dYG5hHG8BgtDEs
fDfJyTwe6D6GMh1NrhK+uEkQ8ZJ4CAKXz2lDpDozYuUj6u4MdV30IEqITiJGYhrCv3gXTI0azgiP
zRjhFIurzwb/GHAolK0q6ibQvFALPkrqlNzmaMZsvNNeBpmnujhF3xIvzT/vGQptH4ALA21mEzvi
/1xGbZHLXOZRlq8j10lum89chHJii/SD5Uc6i6j/7g0tM9m0Rez851T3+Glm64MWUvM+xOWmTv5Y
mPdkADTdNu7hjWASRh0EDE7sy5S5H/WEpAPnGFf5hIZ9V7lrSmbdjYlqmLpTABNOLFZ0gksqXasb
f6hS6NPNhniBGciKBe1rmODlEyit/Js7P6c2pMXgUTh6pI8Epf+4HrZQYxP2YTFmq7zosSIcQXn6
LTntze8yBhdB72jE4tBulFDh8xW9rmaLOfddsag71uB5iUOnsXNVz7wtpR+zDpFH+FfJ5gsXrp3t
xXnbrtipMTN/wy94y+1zYRGXKfYEiw8MPT/ZKNLn7Bf05qXjroU1W+vxmlmkcXzAJsso2N0LptHB
c16vIuA34HgQOWn/zTRLybGmBGVL8VuVO03t7aexgyVcnU0rHdaxnXFPO838uFdrRsXy5UrY8kEC
y1E+J/jss2E9Jojzmaymbq0903QPUZPZ2W3wJKt6ezkc7uKKMkIx04GrR9TXw4iWTVvZrH2p6Z37
6opcr1EfXBLv10BHseNjawASQfcGyRFJpZkJdsaCwDEPqfpAcNLsreV2USRoxFk2acxIagjtkZs3
XUTX3hjTpj6FCO813PJPL12uDCahRYSwKEYjvdW6eB9chBTRHDq+J3lSWsyEjopJlLkD4zLFH2BP
VCD3KRtu/EQGoyEtrT/4hSoZ0VkT+0zJgW2zbsCw5AaXAZtFcfbPcBaO1Kzv5qFiSdPoVLZvVUwC
FREuZ0d06eMGhD6hGpH+uPMZ/14k9hTjq8u2pf8zWMQUND1WiNZzzzn5ueUVl37US3YjzOZSDjjv
oq17ja9PRqHLaVYGEArVQ47vSk7X2aBVncZHISgKyRnwv2/Mp7XKIlnk1c0afaKpRGprMoS/mNb5
Mi87T5gOewKEtKFTDE1IgBn1+3kMslcfbfMUyJzsWyWt5pGqsSzOeDLvN113MIykruht752Rz1A6
byoHhJYaRdPTi+SJQk/o5fyGRc7SZ0dNubXlWjZbtSPfuoPkBZ3yW7YJx5hPdEsZ3VgTur9HD4w6
Ql3uKev+OS/sF9aJzRk63t0dafAKfT3+gHKdkdICGp/8Iu7Q0m5KEmxlEJpPEOtsjAFmnZPegT7o
mYagQFqL5Sl7u1qKAc3OT7dkdqj1I+8Wn/OHa8jN0SKedX0hO26gcnAC33xcMP9ScHRY/7+gKUlF
peUMr0FWB6IUmeiZTn+u4VbIxeYSeBVUjLyNKRLslp8IV7R+rhlG8vovLkwh37n8LLHiNGcdBaw0
KgooN9C8e54IA7ydMQtlsqr7QLdv4FZ/NcVrakspsIS6ZGLotnEiQ39NvmQ42w6t7GAG1ONpSY8M
h8nkCjVq4uElO5FKbmMxvLtayR9AthY2HUTgiG2nLjJVmIVPAmTYxlzfkT8mAZCG7KyddthNvBtD
8+/dq+rz8W/vtNUyeD1BfqfWNWcYGVJhcUdNMOj0NpCbnopWyfe85vfTqSevTfjsdW4+RXw4WOlt
FUES/x8b3ShWr6q+odTlXq9S58jJqN/MaTLZxD/931oQ+oQaT8LIcqlzNxrBka1HS+JFjcxWYwwf
luNw0mfyWBypo7sdJAEU+Arr//98/L4yfl7QKuYyANlCJxneDMQK5EBUtwSl2GI5U/jQOx7y6IyH
0TH+lhDtAp9Rtp1BXo51yUnynWQr6DzTElzjs2kkNaII92sWxYlIjSVD0fTPWppixJMBzcCglfSF
+8uRbCKMNoB+DypHYALJeclgCrsBKfvuhqaFLJgG9BQ5EHpune/U85GZ6B5o1m/CvPhb1mXrbNEY
c5IQg0AkYIZnGd0FN5ZHMRc8PxldSzzaoIG5llYaHRtn5IiQtVoSyOGJwTUi3Sc/PENGWpCqC6PG
mqtRi5bNvhmVF6zdP6ENq1kXZ6c3sTnM7rRxhBoQVaDBxEUKQ0PKz3iwmED2MiFStzUBWFJyfGcC
T7wYn68soT1bwQG84S5mmOaoAkbKAbKesQmDrNTZzRg0ECCdBlHQxIYJkq8Yaste0rhNTA/ci+5Q
8u/qo6fjyhN4dWZ5fsJF/GWjtX1VqWFgfHget9kzMbKux0czc4/wgTbOokFpH2S7LH2GR5VHvuFu
hhP9WzoKiAVjDXmMqHlciolPBiUsYxIiEteMKgcO4u2KTiGka0LB/vmJWF5MbxytIi2aMUYFwDFk
7mt5ilNAFlz4RqAvJh6u5lYSngAKzBB60wJgcDjulhUIor7kAqRNUU9gS7qg6pZZ7PuchTz+vKsN
DI7iUQ+HxEUZfJ3i8rF1YzyKHpkfAebszDKMElQqz/uAQWOt8iK+gWhQT6SJARnOekyzpmoMcGxT
tzQZdFVW3yj7txQI3vP+MGVU0WEuZVrzD0AbYoU2eC1693F6h0yQK9f63prQRw/unEDMorZXFicR
1o5VryiaayV86B5E3LLPW+4bOwwcApuhEapveQUhyEGlLTcYp5lRzIXbrFVXJJw4Jc60HYP4ArJP
y5lXhdJ71O6rZWZp0BZRxDhfEHcBv4oJ16BU838YilEG36aI+kB7SHjvokSFpRyaxBNpOGzTOdIc
V80lpReoY/BS8SJFcSK1LS0eRdaaMQx7/PBArpBGsLRqNGvYZfbmiBYGqLYStD4TsEmJZGyzVzc9
QFPNwbIQd7fBsv+SBpcdUxuEtVflemq85epcn1cijQ/zJQZBOKM1f4eVnAYNv+xdXSOaKWoC93yO
r5eJFtsHQjBR82XIYiySb6BwA+Ey649PoiUX6bgEYZvfEp7IYLyvrAs//yal5R//XgvljFFuPvFS
MVm2vzZMz7CtSJwfkYW/o04K+C1fD52+tulfC8B5HVYwjCByIyABAe5PoJH3TnYo2DhMOQ6I51D/
YQl5MSbCgg1tr4fwRVRjcNuytPF3qGe2NG8veHuUpbHmGFA5C+j7ymbhIKt6Az8kD690Vx++03vv
58GmpCweAsDOicgK+C9WXWXpFCUhkU93sPvwTSndYO8k2/En3yhNMfaHSIufMSo5ENy/EIgLbnZN
tzEggmG/7xvp9sSkg8hWSujNinXs9XLvBLQXNXh8bxWPrqCIUgcwhDCgsUeZmoJ6fJT6HepDtvJa
0AswL+T8euh7BtRQlgDIfco7QCs/HIMMzgoMYBPnU4qqvHxC+gos1aqE7sJanaC6APd9noKSlJFk
a2B7HCWxSqb5UrZS5AM5G5GwwiuJd6GBzRZlaxvYpjzmw+5pF94+Uj16gLlYOerEYv38CUZP6iw2
owU7Y30AGtLOOrMXd8bQ4eegKwrVkIDda9Twalkxce1OtbtWMcHtcwvmm16wbRUoZ1j1KNbWhCN4
sBCxbp0G3cU+0zfXHcLxW7B41gzE3wXp/FVlMa6xIcuUzgBfIceZqZHH1AXkCjpGPvcUHDBsSd4K
Tsu13uHBoWIG7S0nO2UiCg+DBhVKZqT00IrvWpNx6YDNVddAyRqLrNzf/lMsanQasaMF07Ij0K5l
8N506D1dVUtCviVeZgFgsB68s0pNhnN7OJJuVSlBSMaz1wVMOWOdk2kLyH8gJxU87Jv04+8Ug7K3
IMXaZThjeK6LhuTVNymCrYwyUtaK+CxKxPg8rM/lYBsBzhSqmSi2GXWv4KYKbuOFJwUrr0EhswXd
AxFAKjHC84tP+miORL+ejP735Xw4lg4dhPaXlYYpYc0XGulYI8xmkSjewmhdvRYiGiFDPvGFjA8G
5YV1nWc9GYFfOR3i6eP5nqGjyXjFMcsMv687u8TTyE1K2CzZdYq7f7emdcVnySkmPqs+uRnYvmCN
rY3N9COb0zu1sFCSAaymeD0OC0EL4VAWymerX9FQnn4wxAtgSgz1UBsTowYO6QdtF1asApfLfj4/
3rRfiynRUesukuu+AvesstRMyDZ4GNpOFMS9cVtMA/Lrn8rmk1if4/IY9Ay3usGBhtZihPvwT+/U
jJfj49fVh50VYLU8Ci7es+o4B/1e4zjy09adiDWUmtLTiz7Iscu2Qa3mUha2nMSSlgNrszeZre8P
LAnyT/7zdlxvTkqZ4XT3jB47HMLEE9Z0rlg0Ko+BvqLZWFyPBEsvboseMXJJlbg/7GtQGGwwNi4b
iOkKFNXNwyOUxcOzLJirlhhnNiBs+TOn+eFYpeNJpPonjVrxIkXU3/Lc0UkW3MEuRhmqGbbD6mEt
Ixb4PIqKIm1W+esDMN+x107YBZ5FefyCskCTZWYvzdS1rT9jM+60G35L+LB/9kFaaQrZoo6awmkX
mWL7NYdCIv8EhE/zHUk5iG1HdK5hl0m67kjwgULLvW4JFBoiG7222YubTZPfsfgAERKc//lxELlb
sbNkwQQZ0abmu8EzE8J97oeOXwh7KTpl/itKWTpm4jrET7mzkJroOjSGpN3zXji1GIVtFY//5gbN
HUGrzIz2HdLA7dNgJrDc9cO4gY0wHMuLjvc7Ylmzrf6/xQq23B9rIso4Gtdf6ritQO0EaApmBp4v
7s6I0hmJW8sw0Jj8BMXwZM/W8iMbA/U/zmkHBHo06Uj5bIJ6/YL/QjAwIaQyJdwODlSQHOEhWcAj
+wx19RkfVZ4Q2MN0zHhUx7NqWzOX4RJTHHzUqiUs6Ft8MjhJ9+VcOv2P865v7+pDXXieiMLH+h2S
EOuGDkGGxl0wGyr0nRoIobM3SC1u03FFkiq9E5LxXST9JzqidL6q7XgNlL+kLQTQUEdTzRUhHTfJ
onLKQ/EEuNMHp9XtYIBCaZ3Qk7Tev/Tk7/lifpiDRQt+cYoFiCdFJbFVzlStEJ/6u8HByrIEjuA9
9AbnZzrE0A8grzUauRP/0RGRLdB+BWDoDZx5NUK93/UScgIRuL/3ZONFdt33vOLjQ5HqzZlRY58t
RKWAsEliLR0ODDFjYgPiw6s8aK/u3aouNU0l8BsPznIL0E0w1Z4IJm5CbEWp33HCEsJk+pfEd0VT
kbdhsMh1UGY4sdN9ly9n6AaDqhujeIuDXssJEBCpfiZxSr7jfXkN31svIrb/HEP4aatJzkUcGlx2
q2mSWTN1fZ4wd4Lye0K7nTtqy07MCOqXjOXRFjpLVcHC/I5ZPZpRY+kkYYx1Ke4XtxHgsP04QmBw
Azn8X4H6qhwasMi0UrlBul0mBrEoC4OnK6s3tk3FG5s84SJe9LX5k7EEqfnnyaEcdNq9ir35A52C
0R1hv3av4wEa9N2dN8JgW7/nA/83f1btxzlftLkBPRRTWWc0yNymGG/YKTWJp2rWLUy5r+8fThwN
9mIMQyUuTMIOG4NoLJdJ0UEW4K85Ph1MbYChdw+J3QpjMT5AS3p7VsusT+moNYYDaFtnzs7elFMO
x/UVZ/u2tjg0ws7AFDIGJrYwpCrNZx5W/oOPQQ3EFqRKTcTH3SnwbuudTL+ONvHXKwjKGa0cntEt
1XB6XG8/9bfWPNBIOFxQOXiuCZWascuw7j0lt4LAsDfQnabr/NqCh/32OomuDwmbYz0uv2jtkMhp
WhvO67QaxEEmAWLlbzjjQ5SIi+bCJSUC7T14tA683WHPl76wQkM2HmJnpvxoCWsa5jb1tnPH8BAf
jeWsmXmHqJ4OOVTWNTThWDjUL8smFve2cvIFCHtsH1ih+F4VHQ0ASNhCMcuh58y8q3JBolnziDkT
IiBZxJtd0hPHJIud7MF24z5ipf/1bnM2MaKtL60npWuxcuo08z/pizIMNdae4TeoCHhBpGtArwjJ
jeM+OBjSfL8AUPN95LDqjlFr+qF8R7R62nxdli099s4800rWTU9we9LX0nDN4q4TF3/C1n0ef6CY
qERw4oeVgVmn6MNjIoGWpjfR2JTXRWlL1KYGyOIhGISTjlisnNIFbWDKnrtb9f8346d1S7/ezInN
c/ZcleDrYJyrCG7+R4iA/LVzHlwWQyrmFnfrcuzq+vzfBKlRlZY0Ez3CIx+W5Iov8gaOLeecvc9Z
TzoLpgfydbmkR8JRzAcYwyXyKsfFsZn2eOANWKJ4faqq9BtWjt/L/t+hLQrm3FOuoip3DKvmV8fT
rohHd2xEmE5Ja2ndVWBacKR23CcFBoJT93tlfhlFKILYxGkoPXfwM+GFheLBQwPnxJLa02C+1wFX
HQLVBBtwvERGbRM8H0DmAHIBJResESgUleQhjnc0Sgm3W5j3kKthwtPe9L9I8RSX9zP8nbBpD2pT
GzODkSVKoGwWElKIV60FvIxNQjLLo2kFWIakNppcMSlRi7+V/O+KxLkjfnRak8kiCKdD3wAf4WqI
1ecF2X1XeV584b4F95Dq9wD7XCGoY8s7hAtJOuOk6EzHmKAf3xzpQF/BhXSO0Sy/887IYQmGjujs
uiHI7qABUL0pZznHFCf5ILpqGoRRwtFEur7stkgPtCpGVi4qjbDDhFzEgOUJ0f1CmJB3Sa1O5C1J
AipyfmZrL/9OHwRo/+qfWD9tnGsV1wEWd5ZhyjzbRllLkoKPKz3cCQBnl088qgqGIR2kuzEoqz6H
WCMMmbf5tJHivQ91s4OrSUjUZZlV4bMHFe0SmWdsXO4kz2Lc80164scp4ARP7NY554TsCxtT2TlT
fXbOgQj2PyFm9DlsrXa5QVVWuaje+eVRVIOIRGR9OCKkqSH78LngR28lNypjIdP9+ktFJDwhlZpN
wXsexXC4Q6LoRsulV+1gkUg6mHTfdSzyLrK4kkzA6y7pQsmxVQtnVam246ZjHWAO8t57nHMskSbl
KE8pZRUPnWMIKdTv2iaf3/KfU5HQHejjSSij2mSvN7Z5b+KhPvaxQRUn/C/VFlkNap4gduxIP6bD
3IhnUr6puNyGu5cDdp5Vkqv7Sy8svPJ64MbFbDEOwgey+ITYn/5oIHq0ZNmORpwV3yf/kmDuh4MY
Jhnu7zzCuM9LeZUt+5nvcN7E1amIOr7BAwAIVnO6sBEM9qd/rnaQeCfpDaKZoRTRcgtEQRQMbtIN
/M3Ey9T914JRjJjML+s5u1O774BFGGYh8UYiULwszhTZqR1FEdPt7k/lREw++B+7XHJnXW4bj9i/
TFJhW2zbuIqe0kMT0R0irEKLhMb2yldXDrV7G20Q0r5pteXQcLk55Wq2Qr7e80CBvxghcrjG/Ye2
15L6qTXmEUKrD4z37SJbPG2wqCl5T1n9kipPYGm2Mcks0/oLVO6S+l0+vZnVNOGqsbE8HJvBkVAi
flZTep0BhR0i94+VsuajJZZ7h82v4grCktHL0WtwmzXQX3MPpiBq7coYudO4gdHL26GCJlGSYNXH
zLuS6nrjGsZDFPdrrC8WhPjz5b7TeyugJCgy7Gra1tOec6beY2nmvMaRbECxVaHbfK8F/68xWDMU
jzy0ibtTPJvRIsw1wWtKaD6YNbP3qWm+Q3zDv6xw39IOstkCDdSiAM6Zj9WiWPjtZ62L+ve+HMGm
IMqfx23v82fo9coslkZF9wKi2c3bU6PbiHaZH53Zos1BWf6MbPGIzW/iD2teLcHOzYA9evcHjtUy
fvrQmJtzJZngwxDLRcBdKzZWahInFiLBKisonjBgoHHm0aXK0H69cbu98QybPFJq9vpS/7WMrG1Y
SW+4dtJaddtAZAdI6vYmUvHFEYQBz0+TExSENsRnZykY7PKYho8RjMoPyRm5lCEdWjCP8EsAz+0N
/6Tp7OnlOm1dglM6oEji2TwJCLKApluTPhZl4t0jTAeqODaaKsveUTfnCCzBxLomIUHOBVZVNRlX
VMBxoTVMC1Y4oU5t9fndAN6Umxlgfq7fCWz/u+yztt+lwvlAYkmg/leeoVUHtVfIN+eTAyhyJh8E
tguerQ0oB6pbnw/Y0onc+8KlCOQ6cCKEWYMmC+VfX7M7e3M/0TO4SjjGVkXwVUFg4pS3r0vv+aza
1kfp+hrEsdhokgl4P0KMU8K2id1yLWQ/Izm3KLFBJltH0eS3CH2QV/Fdlozwnojlpyo8646IR0ty
xNIspkhOMHbeIO1d+znRgY9tmOABcjOji2qJG/IO3RS2AnKO0OSxTlbqJcZlGZk26Dl+nAAjHTBN
fCQHp0TPs6zZOR6tbXnQdKI32eGymBhVrIrHIgV9FvJhsA86qY5/Dw8+2E9qdQrnUPm2E9d/YzM9
OX0DV2gOie3Jwt/AZmEg1P5+VXunOymgLvPRJldhkhJyKIULyNpJ5Bqf34//8BHQDb7cUTk0k7f5
BcgNxRlHo9umv2yEkcFgEZMrjjj6v54WTy7k5CT8WGqZNsyo8JhjGi9JBy1WuaNJFkrDWeQVVM9b
fIarpXT2CZrMjmUXUyeboSTE3toJlv3g48gLWO8IfFer2zTfuVd87ux/fbgbLE6XEzznNh5jla6C
l9rEtMjbqx/l3BJZOIQt8s/O4DVeMkzJ5uow2VeZq3VbYpSoF80gdRL25NjXuwtx5ko8C3iaOmY3
J5FwQIBTAFP0qRicPNd7IObYW2uuZVKdnuuw/O2yKe8uhlZhD+IdFZYRYKjb0nZOY8G0j5nUfxfa
GzQbTDdXNlKKWX11vM8Oyle4r7JFTngRN2JT+ei5D0xxhmDCAYf/0E3jCu/nlznmj0219YFXpXsa
7q/mqc/GE9066VZseLI2mWRQJ5XDHGHcP1VxNAS1LH9Xph2Yp6IEoJV9+BMe4BR57DrJnv8vshXW
ZxA2UhG7zw04VmMWkU1oNMtmwDnjEPhO2PXZsBuGvfEQAt3VmUAr48zJntdAjD7g28pRvHTz4O0/
G6t6itIDPv7pqfEqmXz65KSAijq1KTCBoM4roPgPWN0LW4DYiq2ACtYvXpQWIxvRepLy3rCEEn//
zbWLEmysk8wRHkyBX2FtWYae3QfRDlJ79bO2WpQF4ugVJ98UNKlexf/WO15GcrkzGeC0f7Vn4MWl
9DbQ0y80J3VKjE3brgn2Qtm0mjMbVi1SCD2IV5yQEsuXsr1ACXCbUJ/oSFzFpcKkfYDMvknwrDLC
Atdxx6+h5OxtLYX0HWZPDZUdrAgnHQbRSpIfDJbeUAaEtzvvUsDJiFG66M3S0nBt0txFvcjmUJB0
qlnbkL3olEzlh7tgQukcHVt5WNoqGvb3EcB+mjzHlq0wh7G/LjZRW/rXEVe1NMce/o7tw3K8cLHd
AHw6EWvKVRcGWnFJxkvbsavwq+r8t5GQhKaIMRhpHlXGqYGmJWi1w9HojOXZRPtEeB+3zKHeszhw
RmOCBpSF/kBLBVvZemPdp+nwSQTik45n71QgGyb/IdydYAvSv6HdwdlxZeoVbxSY+8XrF7fpMhFp
7A3M7znJeBrTMUo/p8OiRw8j92dbt58v1nPnjFw53noaakPRptn9C18foGQ+F2sXRNgd9VWM/unt
cCyLGyV21Z3tU4AufM8K92+J+Dn35ct0A3ORfhwEJhxbvx0okAd3hNO+1vDH8vEcHeUmbBX5Ba/D
ruqXaunNHOhsgy+XQugQD/BFmYQ1ObArWGncEhQd+X4M8gi1KFdUq6VrQm7z1TL4C1f/M6Rcv3Ov
q/BmAU9wYSIGIv4OpMZHLyE/VwRsiFb3OOPU81GJ3AlRbmn7v6MqjrZI1/mXXJ8VHCYxe9z/Dh7T
hyDeLJaSwANM45b9E5rt+0/YuSh/L/j9iPW1Q9UnmcxLxoNCvTGiXy7t7Dq3JLb2FTRgm7EkFIpb
/vvPDFO8QeZhKw40VZXOV7SY8x7QB4Xlj7t6iGb7ki1Dnhft+WSbvlfiJ/9+NHKUBOWiEK2DwjEc
mvQeRdBB2UUpzktW83JojtHs5pQ1UFbCPeos3NueJUU8evEJT8FoHW51gNoPzOC51nUuTFzzJsQA
dLQLEBZtwRVDWD4JFrA1gHYmiWLlJg014NzHfu4DOH4C6wmVW/8qws42hNvJPl8X8U4I3orv1ssd
oYh7AA6o2KSIDG27VUdQ0KVbtIoskxeLHKruHBUe9Kl6zZi8cpoQkPVMww18a0uWM7eLJlgV6Oye
GuIcBjnozZAPX+FOB9Ol8IB7qeCRDaF4pa0bC/3V+mVXG/h5XGhZbUfTZv06REDe/fo96RK6IawT
k0ybARc08MnxTiragPeaaYxUxeuzxP4sAw3uZKhg/BhQAEy2sEvZklG4RVHoG5p7yBODphDFRQQs
qzdqAYIeyVtOFB72eqS9XanjEI7dWfaUV20Wj2I9SX2Rb44ODFBi4/0gWtOOW4uaf23KKeKFWIq+
B315u+NB6+c/172Z4us6Zwc30S/mabeIH6I3C3aqmi0xP6Oe6lfAsuF4lm2EojTaabVimConTtnk
X6NMPm8ti96hqhErvP7O1D/3s8fAHlrLFGbXG0hhEp2SIfPG3Xctq+41YvnrWN7BlOYRvmlHfAnz
GYlJZIleEl2Qi+/Xpe074NmLLR3h2tDeQkCkWub2Ua2/ITy0I2Jrw3MJUpIflPaB8xePJujQhGxn
xmYnybNouZpRe4EVa49s/tQQWZF4rBbXMArWiSiJhmnNuy84n2a9RdVZETtjWc347vIa/uRld9ty
geoGiurReDGTE7broAryp9DW7HWJClGqrcsiqdwSXvF3XMWB56NvYUKImpl03ZVl7G+qRr0eFHhr
4wBR3NePndsxaSAtluPe7u3ENndqY1/ZF5FT9/D3rtgMp0xAcOjggmy3kD5qR2sbpurt8fsZ8SiP
+jn2LhZrqc1bFUl/0UnN008u0xjZLi+CAhODWFQzysESU2OIAfL+hPu7tLfnCtwoPrxDok9Ezt0p
7pWrN2IT2VnyIIRLw09eQdYAQan5qQ3a0R1mSy2qy2XpXCBoQqT5E2AuedM0I2/t0FS+ATu+q+SY
/H4nxTE8klipguB6oXdagn400tkT5U8xbSHp3yvvcVuKhNicg6eqsaNE6NnYalVKTUPWHA2NLbB3
T/pgpA0UxueA7EgYIUa8K6dsqN77HOzY5xdBBiny1YHPSaGX0Nf9kK3TOw2egaLfjVdw28LIvdfY
uEA8nvjeiC3KV+4qJpAU6Z0iTKZj4dCrkDcTLOgI4UbfhCVOZxUg1YePNWdD9TPlhLiASPHSQlq2
50YQSMOJod5FgJ5ixwM8j5FMcmiSIUYGNUtUTIPkPiWYL6M8H/HhLh2bJOk3Pv2OYKjiwerteVgi
KYLlUXI5j+N72Ax9rMEusgyq/ot4JWRI6K3kOrfHoNYryLgrruJR56LlQ1VvOoayVK4AmClWjyaO
5XYkbrPkaopwBssrrGF/XTDpNxiEr7oEA/0QvA4EXR5IhoZFxvj/7l0ji8ABB8Z98vcOHMdHF3qa
/SA4NeGO0q5cSLHIc6Sj78CtrIyyf4ssOzrnxUnnKX05xj20ND5O71DhOQTmVzFTI7OgvPqJ7mYT
3Zd1E0NDQMRBL5t3Ljs0lrsDGiKpPwemob2jvipv1oaymwmOiFnzML+MouIdUgdPnPVNhaWwzGKB
IzhZwBElq225xf5cDEyhqRUhAPZrHq7a7jhVT+B469hCaOgvbG8FNyf2veHcGXs4OnHOw9dNqGln
8vGvMZ4K5+IMzxj8/qy/f4cvcD4u/gmOQ5yWSQoDg79zDY3yN5FlOB4G9tyyZGXAlEQbhtwQs0qq
5mocze1lnfjbz9jCmlgRp+AZmwkPLkbTpUEIfNhtDPv5B/dEarD88GK17JmgeSN5BjrSXTLSAmMd
W25CqCOnnSwdQbrJozcIU39tkfySRDbHWDvZNdP3fIegLZkpWEm7CnNKwLXxINEnzCjSDYbKXv6l
Iq7gNxC+1LOh2TCC9MF7n0IAC7e8hMJDnYOunsrTozXD+CaaSdH+EQK3TQtgVln5Ar3A2Rdpbath
8OkqXTwdwEXnAVOEaK+/EY8qk0RuwS0MqJA6C7ebVhK+qru/1k+mQ+BhkwXCLvRbscTOJOCDj+Ch
wmQYlJ8yorTg0sCk43oQFyAQop9AYqHlPVRD9ln8rZQ9JoIlND4S3nQK4+pvktDkMk+PlrWPDPnO
Sie6Pu9FZBOmiS/U1zUWtBc7j793LEgbVIq/hYWqK2bqm+UOMw4xUBkSleohyQREqvKX1FllWoCL
N5H8Vye5pX/WWiLIbVS9FoF5UlSqzeJIPxdXXNfFDyedk+YAPi9rvnCZkBoosdKjxCcu8loyv+tM
QwGP8dgz2B6fFqiwlpNqbYpdrvIvY62HF7Gog89vf+4QAUv7gtiE25UHCfjueNoOW14xgzll+cyr
lJaavPD7iVmtdkyRoY0uqi06Gohf7YObxfYHPEzdsaF2FqGqanlA22uT1nRMN9S3CmKse8wV2K7w
pnzTzcrXtaw/hUzTNH0TNEhk62wQfuJEAS+zg/AdcB7ddZsf+8bk3timsMSrfCwRGqWHG1hxgyf/
RubC0sNNfpCmtGBw4NqvSnNVBVWvkWxmzSbYN99pLQF81XxdOGxZKa9gcrD63PZ4yJtKStNI7Wex
p+mvVbffUiAuhB8a7H8EOuA9zicpvQVakAG03u+6XRJpurmwMoKDG89OQRjGJsGhXXHtRQs/Hf3/
UCHVOAOiBgS0iEsM8OwsVdR8Y9LfAj542C2JucmqqxGYGv+c2yoD0Xbo3aVvgy67AnJQBkQBcA8U
o7J85o3IqDQfjqIsO9+CeyXoJTZ2Ft8pkawrzR3qdRW9Rf6J4PBtLk4OuSJQB8+b9arrN4tBUazB
aBooROtFcL/8aoYYLKyo6L6fJq/qcEIGCBVVsHwkNksdDj23NMS8hpO8BVIPo9vEaLIWrCmipnNv
JdlXJ7QZf+zXdxXZ/f28rbN5f8PlZ4Z1ALQg+gTci90SiQKClnjWUqA2hvATao3DK9Ma8xXovV0G
MpxnHSGuHcRuGgvD/zK8KUFeXaqTQjqmFJSdO+hfYkPz0MWpC1uNyN0eidARwzEFM/QqyLzLNKFt
Y3L2Uu2uRqkP82ApQuwr5OZXzgn7noGoWwztZxgjfORVEEX1wdbhr9ptGcg440OfaP60suxyaLpi
lQINwP1W/XpK7XZbEUDaqIO0EdhAn+433MxL50fe+6/bSImc+qhRfXnL+4Nv1tjUc/6jCSr/Dm28
9t0U6xye85Z7imjHITUmwNkKuT2l/oJr+lo9CAh6BKnSPYaAj4YBpb0Fz3J62UCNIogcGJ9Ly9FG
rCEQel9bQj9GBBudVe8Z0dOTWzxU0R4PuVhokQgddx6fqD9LabglcwDnfH7YaP9ktwBE9RwknmrJ
EVdl2iRYnNtbO2V3JPpYStxEIg6kqoUBAoH85qwg+yyE/MRVDhLjqKE2IJlDivjWOmpxnSMknEVq
BfPvbnh3UpKJ19XZAJdjdn95BjZOA+JNI6hORRdVxU9d3SDDOMRVTjcaU801N0zUoKmPWdyCYXQQ
8BRzKWWWCGgZ8675iAPP6Bz5BjJ3wkGamTsGuHdQMyo2VQkKCB4SgdV+Yf8uHKQWIKT9fUmlTmR3
Zs28ZUnffZsji7RFRM20sFL3unatRGU1PgFyiJUiFWWLeT5jFE0nvZuPUw1bD+u+NgtWIGbE8xhq
bsGepucd+HCfiyPBZqpBH49VaPecvLDuMYCNOl2bbBf2qL5wcJrNIZGUbVG9+xRP4C63QpWfETCk
dD5mDQqfrBalpMsCjlpDOZZc21DaGJyyuKgfAvLVCUqEEb+RpWHjlaUuqo3U1VjV2Da+m2kN1peS
ST1sa+X63Xpz5/2w7J5dVmdk8YX+ARh+/+F2FRjp1/3X9HFupjfbZDAkvaf5EHXbS9iJxrz/sotn
Zc1nLPApjQjxBA5JyXQZ1U3+w4sJj7ZJJkL2Ad5dwE+obGvPC87V3WIuk52LNd+lfSd+Zds3+Jpj
L36XuJyMmEm/+svpQBb37OxuakKMsALAfsU9oNPHHesDj6Urc7Hk2gT+SGNDnCXSp+NpxfZt8s0t
Ee6JmTe4WhlplwP9mDbQYrOXu51nhJVs8CnAuI8qeo0wtL+lTZit81HQuH5GUZtZkcR65kj2jn5b
CE93w2Fx5+xk+XnrYrHtODt+ZXfUFqmpFMrkx/+IJ1XG2mvg5DU4MTT8ck0XRgaUeIbAVyfHRmHf
+2yqHSeGlj6C/I+jFfDCJQSRLiMeR185sGa9fM+4IiWufw3SRybU5th8VYIey4Uj+amLc4icXGgG
WxXFEj65k+9V7qsMwN3ZvCq9VTogrlXmQ2QyRnwm/b2ctLNDmz7o+2f6Dn6Hb5V+e7grrZqM5qZy
KS+Jz7Mn+pWo3HxwnaZUDmXh9MTIxaREGREBxnpfG84hBXOIQLmz4q3VbdklvXs8/Eom755TbMWw
wxC4ArSZMz45sfu5VGQbl5dWoWYcbuOLBjzwSKL7QMQyGDTVG/ChMvzOakW5mVMWh+L5SjzpcwQa
O3KiLP2AgayNIr+PEHRTL9JFO+AxedAiyfjA8TTKzGHTDVE8Ufs2ijWjtK7vc7mahjsiCYJ1z4/y
yZ3hz3EsjAR38GLVrrM/3SL9FrpEJ0cmovZFVUrzJeuJQ2YO/rTQRlftdAz8lP9WFeEViKFiYQ5k
V+yWuDW3QIxXejTitRHptr+eWCnO/QNmYE0uNagRgpqcPBppxPqgTCTPSQ03xUR5U43eoK40bQHh
FjrV+AByFkFDxRdt6egXi8hHACCEAkJ3D3KJ92Cb3Sy8VZSqFgNxLbz5iIjrAAcVtUpMS9dqN+zq
H9l3JvN414Ex+Vwy5zEIF0L6xbPUTlqpzOc8gaF4ELde17/vyrIBJYVXOkQ6jk/lsR+ozalmPPDE
0ztNm35+dJNhzl2esLU40hibPaIxUNtZDDjLQDmwLK5UcRff7cWP+kxljruSBsvPDPFylAkZEUe3
wV69pD+yTFoUMmK3tK3YBz+xlBM+kwf9K0Mu1YtVjwxn+X1Y89p4GyUWUVR1exhwyz+5PogcgEZ0
7gfjmaiBEK6yd7YHOy8KxuDszCFU8hDeKkSh/z9ww2BqUHIy3xK4DXyw9ptbMZg6e7Hl38w7uXXq
DmVt/p3EfGNQsGsvR+uE3Ga5KeARpf6fsdKw0tQD15caAN3S1ccyz4CwRsZV1qgjrorZUeKswQOf
KmlIYvUi4uzZqNcPZxQhM1FgT/uQBJuLTzHzOKPw+rxQoQVce1lEJGv8VqefzojOlfpAe4QtxwP9
YahV0e4WqDz/go8smNBmRAQ+5/mfPi3LgwZg0XK2ZoX4nMlSwY46Rm6COutO1iAPC4zSs8j42xsu
xr3OA9VeiLRrcs9ZZAgI7TlF4lBkUiwiVMN/1Yf/03QHXZgqHvV0Q+hWlVj7yoDjIKlJnYR4KHIo
diQiyzvRxPKlfPoKoM5Vbm3fGtWdyLUI75hgEPq1bcnY1N1ERPnhARgwbk7kaTh03W/uoLlDRTzG
W5c8q1gtSdPASMTudW5jS9tl6ChWlNBqV5nV+srpLugCoxQPR1ylo3XX1yneN2lk/bj/Yf1dXBw0
iLVtFxe0rl0sYUMrn4Er2gJJcVmWSeGYpCV2WWy7vha9/r4Mtpjvo1vbLvVIa6zdY/+vauQJpQjz
G/xCdoqQpyEguZZzps6+qLQlNPRMYJ4LaFJL0PduAZHszTu7ryruRg65qpZnN1phRQvdb8jWND8L
oifihx8lcO96Xq6JfXX9AjOlde2X8yFfbJDf2fcWhNjLKHmyV3xiLo80XV+UoFk9iYFeUCtYUG08
mOsMsD5ysg0ceAHm0a0zlUF4RnaVPYa8zLQ57LKhU4Bqktk5rAFHJ9gTVQLeiyjNySG5J1cpaGKr
hcmdxIbQ8029FbiLITCtnHqcTbcK/1AuP+mj1+eAM1CDo+wdleDWxXWfoubob9RId34ZERykJ85O
OlEW7WUYtcd2jqic5uuPXCqPzFDTPogfqCqODLld0NK6R46FWXvv35ZwV/jUSH5cAChXdaZsMJ6e
gkl6O9D7Z+jEyCurbDBrMWtYjJ+wYncZN1LJqhFx3WvwEbIEYym3AvAUwCzQghdNlTJx4UZO+7z6
dN6oNBSdNvdi1sTD222V4sZuBSOLipOJWW98LZownDrpew9FJLhKc1VeXd1c+qhPTdRoKve0omYq
b8yyFvliT18lfq/LYZVW1edOStRBDQvRHQM1sEm5c8PQQ9a5hqufPq4KYuWsBrMHMndHAKp5isIG
nThtviworSeALrDiN3df+hdVBRxrtJi7ycBJWQINHqbQxj0VuSyU6EKRXUWhtkeFzcB5dX+4QcIi
gQZ+BkXek+liicBh8tsk4gYx9aHfKqaDgiXDdsCh0ybrW+O7oJAKrWT+L9cYdUYh8aDOMOr47MnI
7ypthdJkFgAx+gJFsHB87f/QsVQmMp8/dGfDoxmsUe9LffYB4h3SFl8Nb6NUuF4OlG/9xTvVIpza
Zz2L8L7tXEs53chL8Vo2tIHZIxKTgJSG1z/K/yJmKWtBVkokVhtLBYH7SBF4YFXJMlIfSCjWxj/y
marnhRWibdnZ8gun0iU1uJ1SgdV07eP/uc74PLXMlG4Q0utSPPUUjgWwrFRZYV4YwY0qmlvo86Of
sl5ejkyWRZMYMicBRa+LaVhgHqstAoZFNT2x5xmojQKOSYjLihvZ+6eE+VfgG+hLLxPAIHE1V4KH
mguUzHUBQnHTl6dRnjzOQji/Ahwdz1+N2iKf2dFupfqv2pN9CYiRzNVXKFC5IBuqfHmLxCfTurCD
ssEuwCC6aHVVRbX3IMvupv8p/0Yc3EP+QCKky7SQ3jjhUHGChwV+/VxrW1IVJBMcm+8lmSRiXFs/
P28cEFqrhU0pcnKtRrCG6k1+yYF+wcq2vGV1AeLcxCzUWYVBAfklfP7uJnBkWsMU6UK9f1m+oO0J
zeUKZp6QlFlw549BzXjiLuRJ9xhSlM8TeTsAr9JwwJjHlEbAWTToxvlbbdDOtFOlitxP4m0oEn+F
N/izP8aNxIJznwgTc5+1qGucfhsJ2pP1Rm9xkz8aD8cdpeQRc2aaoQ1eQ2aK9CkH2NJuSwOV7dGA
LGR4OOpXabYB6uujPBVHePd7NuSRg+4OgEDymQhoX1HOFyD2uc/PAG+HyRHc9Q2XPE7+UO2wq/Wb
5l4K4VkO6wayd6SJqPW3O2vU0kqI9Mr3/9tzEP28UtLwSO5sictESmbA35YVmsoayc83u1uJcquf
tGE3sWaNh2bgtxOjduJ8fe8Pbxeuti1GO7B/dVMPDgGIeBv8zTV4hXCjfZs3pGwXq6Hk6S+8ndGV
1lwkTX3Wd0Ypsjnd9CAUJzfpOEl4kGA1eeB2kf2rfxjWDk8bzL3jklGPUBf7O0qcINgtN7D1Hz8U
nsjWpfi7+TrK9fingR5GZjc0yLVhs4xUR3CvJRw7GauIpAhMdhlz0Mv1LYWV0BH39TBY4pFsacyV
U40fjcTDib4SuVq3T8+RtoEm7iLcDyIf3YYlh+gbDeYws/D/SaVaULh/Lczy6nj5moGdwsPZeqkN
NJl6DAOXYAFDDAatLsAvwMhT/5bPfffAal0zr1xYw1rBHJlDoHGGLEaVqQvw4cKGOmNVYC5LYFDT
9XUHCwCQ1HwaUqS/ShdonSkFjfL2ZPIOl3YpumXjTrW4R0rAn/KwUB8HRHva0VUCacTnkj/LXVvG
XgA4omUu5BxOXMZ7XqQLhyJazk+cSli3lMIe87ek23d6rvQC31Mx0+pJBZMl4IFq8jO7mm3oEIu5
ffXRgPkzQ1JER7BpaiUYQ9QPpq1s3jeTd4W+ujdQvW/7HjCZ5Cv3NJoNRTMPq6oFJmTjeQJerSfc
mjS8lRvMCu/wyA/8TjXXmH77nmISMccabS1TZejNQBUDNswhU1YJvC5M63bXN10Rg5UFSYiHDRBJ
m72lgrPxWKD4QkJXnG0wlNVkmZY6lRMkeKqTMsNN7pMSqu5i190PGl8R7QOIbJz4fUHIPSj7n3Ou
nJvIzC0A9LXVsNY5VM1rGfurF/yGthKsHEhcCTh8iULNtbuMBj/DF2OJGS/GJANImRU8J/U99YkU
N9YzS3UhApQ9jnEplu7PQUZ3wPBPdv6V1TQRZnBVArIkbIE4qWfnCoUpwcIZIncOoRmwCzPciPOa
e58GLNgqLP+bmdm3L4lQHSd+gshNzH1fYxbjttoSzimdeC3Gz206ef0mIazDj1MRpanKLXBO2D2F
HiWJxttbVSl5naJS94wK4wOIT8rIWykuBaAFjeO/hy9B5DfTRhwzHN9kK+lGYGgGQje+78lF0Cy3
hNhQWxODSv5PfVczgwajJwZgww9r+4OQIC7rK3DKYyKe4aws3qv1N9za4N4pXQZOlcWkxtYEYyny
xHTRieHAt3K70NTdxrPwgkML42Od2c3/lL0l0a+Fg3qfDyglxV/tiYhaacAU17cENTzAvRhePs+P
XvDDqfnunEUYKabv47QJ+24/upz2Fjig+g4z6tB47IUk5Q0cuQQHzX/+Mv3LzzXBkSKKiYipFRA/
SEGC2ffzRoG/7s+NjK6YtZjb8C8TBcskH318KxIkmkD5rrMxwd1nibQanm8DA4QfR8Z6jSdd1KwZ
cKYWvoXLL8DpT4ynvvKTdiRaEqVQ5zfLX476iNNsSm74kKVTopWeT8YtThwGcHdszKQmZPOxNh1B
obsYHugK2EWynRh8BZtJs+kAsYQXaqWNAA0o0NsjUF5TZ3ITiy7OOG4z3Gb/3kh4r5AZwrsg7vnB
VNCPFYRdblo4vwsPjpCac5nKD5tOSO/KkT5zTgWiogjX9mTOcxXYqVzr9Fp1T5fvLPL0OkdHZpe7
vKQbUw1mllBryqzsV8e8Pg4yt9rQKkp1SDOHi+IpmJxJYUlkdVAzOy/Rl2cWhEwNuAsNqKAkrEwp
i2IJ90aOQ+ryIr9ABNuHkSrPS2SlH96a6NnXLBC/ddKLas9VhunSd7tRBHxwRFE4Xz4xm8HnP4c5
xV5RxU9zzMFFjkJ/cXnsVZ3yYUzvIVRdMc5dTh5XytQCDpIpy1ftho1nyj3AKYbK6O4JFhbAdgsP
XwK6xK/GnEaGGG7PUJcX6PAidRvb158nCd1g9wtQ8mfGClUIlIt1UKK6uqk4esCCjdVZ1VC94tv2
rXJRS4EaDDsjyHRwvgDrzyM/Gyap/UjyklsvWdInSEiBb5zI/0cNIJf6nZGbSpSmK3Oi+8cV2YYg
ip4CG+KGm29/LDZqJIYKHQfbqn0nhy9pXddJUr6AukfSjRB3OVwRm/L//SvbeaLOjSQS1BxqC26H
e8o22WO7emYqOmRCwWbR52YGHaZ782tqvJzBkL3PpCp1kNfvsrx1Pjb59R5C+Wkv/VgVz21iFS44
5E/Saqxud1V5NZRk4rHIGjZzhpUJsK2dnJigDsTobKf9sF44UHqII8ktCDlx1qNMoCqL+EmdIHpR
cB+MGPHXVE4MJyNKPXfygpq0akFRtC+Kj7+bWpQooBKb0jcEedPDAXPliHYevIKwQa8vDdAF1/8R
WvwsmKrqo53zhU19LhsW7Ph10fWKY6TUaKFo9RCZB3Yf9O7pyvdg1940omdAoLcdx6G6b+53xzSC
HxHwpVEPu3SA4us9Pp5hmPUazXG9qnM6EApDM18lPZG9i0Ju0Umbb70YAVOd6ElCWGsKftS6SD2p
DjTyYOAaQD3upvHSOduBMp456C/KKW83ZncGzj6aXOpwlG/JqlRc3B75NTNeEnOYeLitWMBwLA6Q
pSMbvNhdWh8vayl+t5H2auUMLg6cIF48xQN7WGrKhWzrf9pA08MK/EGPi/QITNXainu2s51Xhj+j
E65xM06YmAiYsOkiiOou6p1nDkmjsWcoqczKgdstxFjaTgKgcIiQMYnwj9XzfI1suMpkP9cZtZ0X
SuXvGL47+MhNt0repUS8uxs7EKlaBf2uZjvmLSv45cA4z6yoMLLzRV5qOEkDvjkgem/IUFVhtZfb
WYYnDN2pc4sWlPIFlQnnFyJ+OFJRDbQFZSB6r8byWk375dKSgLIMgKgzPpcGAVkwCpDfYwZENs/N
6ZGB2pk/fjuexZ6dTRDJyyWD9fbkSB/bErEOWZx9pCRQlVwTnjtHPWP45KK/Sr4xX+i+Tm8mOufZ
dsiaVkPBTvqVbgIMefuMhaS7ZJGgdCbN8GjFGbvw+sahwWXfCKGY/xCh69zo5BGTWolyZfBBwizh
7rXwsS+V6dYT7vTRr0iojR+Wjkoy3fnKGTzJfAjK4VJpPpS0qdbsILelhyMZZBZ7gepXsmS+1Ds5
a9nihZ2swPHYjHSFHB476W4DQuZABy6olCy6/TcJADkvEyneWp+AiCVdrfDVc4vaGG7s694L7FVr
cd3Bd5bbzDxlHbdMRqqv+y0zAGq1w5S08rFcE4Vn3mzWuTj+BNITZnjT6BYurSvUkPOH4OaTIBnm
HE5rBW5jk4wNJs+4biEmN/W9Yi/s4zRu88fDa8vzykXrQhM4JIVCzOdHZbtf8QTj/rsHciwDfLFh
gg+rHAcN/hk4dsPQRR5rWFLofb9RSwuM39SvSXtVZdU62Svn3pOiBbQSgk+8h1XTrv0Ly9qWQw2z
jzdoeQ02uZauOdjDB3Q/QkodrznVqEHbYGQMe/xo9946816jLV+gLRUxO3jUOlyd57Z4nfVJERO1
X7eBamlhbBPryx1CgiYq1KnD7ILGPV0+/P8F4fXs9xrRKTL1whAIjECAezMsXWz9rP9MRpjqTldF
hGun/du51QbwE7hoIy6ADo0bu4sIz21H0OqVgX8eDmQwh0iGtjlUQbwuO1L0WxGv8PFA9paJAMsB
mp0Va7QxtsrtT/nrDlAxl7ECIjM3FLALbAEWdm9scxtXZ2BgJbp12ATY6Wlje2GFsxSQntevlQC+
LFXLJyCPDkB7367UdfsjsUE41qTWkBhQtpqbd7ntw3Yzg7K1b4N+lk/rH6rN63D7HrmKlenB/aFj
GUGHvk8I5i1hD5VhdWllOMc1RCrYYC4fshK/MIVNTWp88xKplrkB67cLj+HJh8hto/awxy2GUd/6
COVqr3WpF4WqBcjuJ75BVZNDdoIXtHRLb4rea8W6GJNiYBOoI+F7osDzNoGaZos2/0UkExjszpdU
OVPyNnZ7g3uNDNBohsTkv9zBXSGWsUkcJBZSdrNl1Zswr2pahR31BGPbETrcEa3iibp0w2MJNETM
r6G0x5R37jN1euvYZTJEnPhiR/8mMF56xCQQP1+LWLNd1EyVxufRFsdnurq8ZIqbZreyOrxAGXw/
Fqw1ez+WFOQWY+j71da0FMn+KXfoMRuX9vGw8XvSlVVPGF5jU6P6mXurIWYL6jhtQ5RUTYhTpvxZ
iKX72jME97vPuWP4WbYWHE1N0OYGum+QBYiWf2Vga4oetKGPni2zB20PTtMIKFRuyUqna4HqmhYy
6P3YksbyC0AYQYSgdmhlhAYD9ByfaZertQ7M3P+iVgZWlMDvGRCDHDZI3ws3DGs6goaBVvEJphLi
MLBCie8POEKuY+R1Krn3XVtIRSJehRLniHcfUbVqA2NVPziiS379OlODio4ywO+P4MES8So+DqF5
fWVNDOxauLzLwbq+ckkwLswjvLbpAZO52t/Kt/0wGwoz6Eq6WzAiUrR1l7/auxJjzaRe90pVkQ//
/Cd4PG/Wfm5bqkK2naKh8A69TP4wiR2Q7s0yjrFikKhVVerHUitLzGAnPjcGmJueyDQp1PoZvDsj
okrB9mz0eoc/O7fecwTg5cgiQcqGnf04pS27LEOp/ovK4a6hgGytSA7dkqbORbI+q5tLOmjFB5xS
9nn/NXoZunrW9AfrXGULPsbgqMmm1mGXZ1I0L2DPXF6vt4EGlKeHYbcTQ/4baPHwRUC3r4Y8171t
Zu12q6cVnlJBpl/D83cxX5Xr67LwR3ebCT68rEIlY55rlc2ryiL15lxDEA2Mk5Ac/CCdVxWz13MH
lz2tevUvzT3lr9HJ8tABdwXKFN9EEgKau0OqGY1YlSsg5dKtK7XaIOjHBqunmZu4gHbEq2FdUTTu
roSckrYH752ctxlyS9qyG+FaZQTA5/9WWIUyF5v3pg3OOwbPxxTtn6lv2j0hjxFX3kuxiafY+IBi
pciyw3eGLWPnuwPmG2tmaZOnIASPI1MBPjrwL0dJTGG+Q00jUuhnL8IcjeraA2qX+9cL6k3DJ81Z
i06McIUXF/4kIPhUNTZa9OEEoFVEJuxftN7B600XNsGrZ+TnvNi26dSZAAVp2h6+/o1mww0DgBTJ
u+TJ8PZXH+Klm7E5ZKhzQNPCVX0nhnq0GFfhHpsnLoE2dlk6b39aopQHkswO1lbYuRtN4o3E2cqf
RrAgF3t5tMJdbYWMHXzlvsjPL4zV45tIHOBuwrn2CAWDlx5yNaLWyglNUkxt5tfIpp5WsvVF5bRo
dkkHrBCXxv7btxva45mIx7ZGutRxn6qeFQjFEh6QzzLpkVwIQVeSgm1jLQsMRh+tiy7HgmEGyxOu
O5spy86vfekYHHYbpccoFSaSzjL4ek9LKL2MKN1lH+4qZgQ7PMwzXa5hwZTpT9cjiMk9aO66oYqf
tEEGEFrEEoVnecM+Tin2YuWRBml5B5dH687Ypx619moQVvd/YZ2vrBR8qw+dV14LA8FKptbJX6cX
od9447AVc2iFAGoZ/Wh1e51x2UsELPLaexs09JHHFBVWaOVly9OBcHWF9KAarXAkaJD0C/Fluxfx
Tt1F4xavj5DJwnJuS3w4y0Kl42R9TTnGFTSZPQRS6FNmL8vpZoPX1tELmsaLiEtYgVPoPD/4Cwnb
M//usQW3M/LHRs7ZV737gr+oGRvQT8nEYTSq20eodDPchtvESWP1Odv8h2DxAG3QKWO2SgpuuCN4
i371/tLWApXA+r7OGoYrfFBHoLOxpRUhzBdwqsdHmxVe6TbteIu2RvYW6Hd4gSJaktGYMn8jQeeq
ajuprRMqbU4w1y+4gk+/twDOejvfmQXNBgp/uv0+v/ewE/L0gdU1AWTlqyZdFmTbmv7f8u59JQjC
1ZYTrwbU9+dvo+y5yMGlKoHhy48KqSNfsCSoKHHlwvQ41Q+o25lCt/YkL43qMgtXpxDURW4JHaMg
BbtykIGijpmMG2P9CWurFxNiJ73xd5SLY9nenJxLJ6kk6qV/FrQvVldpC7au6OfdepkpB3/hXf9H
DT1CuPmNpGDvJvYjWHSo+L1d1q+/TWZikZPxa4gmrKKUOqChFSuYqnXemTwTvLoJFytK9zGDeHCS
cVDAhuUjV7t2fPjir6CKDx4RmfK8spSBpDv4x/x5CeRVDa0ydvPPBuAOhTH/fs9MBd006MA697lx
rVLWc3E6I1gO5mYDAQPU9Bif/Ha9buvvVKUszWorxZ51S1J1+olGAN0PpouDSbtnEH2dhwLz2PuY
wIs9S0rlkEoV9cfjiqwhl+lUvmorhurTsic0KiMBTRjtVsfUCvu/jCEnF00whIT19Dgz1kkVZUJL
QVxRhL8E7zEwqwh/aFelvZR3caQGX7l5QgUi2QQeQTIkb58CSJw+qWszSu3sbEdwxLFaw0EbT+FL
MCMEPuUnsc8cdWoLC5Rj7J35F3gnF3GwongUrRMToJeQ9P2PRBMeOckCODQgy0yx5dtRXWhZOLZu
WEi8w9Rvmv85R3ZMlSRQYjrAfWqt1CbpM/op1QYTcSevvN5c5MHPqFDXRSS2QDvjqV0eTPmDgYCF
9+zWwBJNrUOgkxvw2gNpgIjujOiSB/QqV3TIVp4VUJYSaVw0+KWrERV2kPRuh2dnmU+HVyyTMt59
VS/PXcB4POnFJa9p4s4VPzwrzxBsSK5DE2NgJ2YzflRzc1SuIbGv1gdjAgHLk0Km3yk6GObrlKp9
OAJ9aBA1tOTgtZ1q0GrlmpGrOo7bLQfl9ApioDHgVTqchpQ/UboxnnZIv2KbMxnmJqHZxlsfRJq8
xj9fMI8I1ZEPVS031DpS+pdvyLejsi+im802PNaWMVRA5AxMXRXZf6nD54Nn35vZ362CJMVnHnlw
RPUEoAbW424kOg4Lrj2RBiRTc4jKi2qd+ggWNLVLFQ+OzDolDdLrpuDsJr/1AhexZDD1WHzMTLYb
+K6sMGguI7pxF3scFaoURSyQkfFH1dwxQ1K7GqM7JMTFOZwAqhnZeX9X60QXrOMBl7Knls5kFD+3
Zfm3KCsttOV8a6+bE70ezoOVcyu5aL20XWuWRI6lIksTUOkk2q7+M0UN9iBRWOoNlhGHfetAVzhH
H1bH8RdfgxI4UltMoblQrKyYa4CY/uQxvGrqdxjACqnPFXrdZ1paeEMROM9YYdbDlyhA/HZOCnzU
YZCf9sS4QWGBjbD98OPtH0OAwGg1npTquv11uDxj1NKEzvkX82yf0u+P4uueyAZDDv1gKG6bdPH9
vTZI21LhHslc2h0PTtNH5ksvnFi4z9bpNEO4vZm7+iR0XdHQj0taV06mZwyELneAP26pTfvp1SM6
YSxzxJCbz4YW1RdzT0MKGtTR3mBNQws8kUZX3P7TYTuZLxla2j0EHY+6O48iirre0cmTYgXwkT6u
DCp7AgHMw1L88WI1OWcwmljDv0JLz6fHxn+J0Ugry6+1yOBx4Lebv8AkJFomDfjWeSymKAJ4ycqU
/C56rkYGvz6nvx2rpXKH/ExWpQNIA7MO69Bx9zcKT8I3X+STxmnDdYD9jYOjCz/OdkxcYaZyh7Y6
IHEPutnx0GdT0iqMXC+o4guBRAQyZCby9pX5HNWlfxw8wdJtlUTVKt88tqM0z3SunlC7J3iHVSnS
15iJq3LckBnHDusTsy7F7NQQ6lneIcQYCK5n8fJxQV2G3PTaDEfaGfScEy6L/HxqvagyjBVIPktv
LW+JcajWNFdcHEi5RDag0UaIebGOPi1GAhf0BzIHOQhMEaSj7wARjnOoZlUMNFsnZrUNbln0qwzC
w7oDj2V5qBRRA0oournKLYH0duvf8yG05eJHO3J3cwQ2ZqpbRp+egw1Lc2VpVrWqTSrgn/pRoEci
ANyLOyrUFOdb4uj17PClF25UEyGd28U++fruq8OTpoW+5QTgKYmO5VPxTsNabjyg+3xn5eK1OwWY
soFh19Uu5tLXkrZacklS24eU5AZYUkTIx22w0kn+nUbT8yQykpotvbXgUuy3It3Aj5m17Fne3aKQ
bWLQWNivhnyw5st1MaNOx/zOupmf7BNa4H1PUj4fqha2xq4H1veEDMXTa5nIa56Jfhh/I1qT/s3m
jlL+BEdvISZ0U0hBgv8Kbl1J5YoAQ1noCOirwa3o2FRQlolErrzh0/xYoeEx3RZcWb06pgpcH5Bj
8erGXBS40DyCMRl9QTHvL+XqTusFEYVZDsKJmB5+Pqad09sXieLUIMY5wpqgQFcywG22Ej85ZZxM
4RlYa0RGAaJwOttFLVL8NhxIXh0OhZyjTwnOPmldz/Wu5pAlVLvMGIRDJSnuzqY8UYwYtoXu78YW
O+xdUORE4z7BNe94MMfbFFBq/7eQMX2kwBtEul5bgQUqimwGV0o8aswsLtwmCBVl64NWNqd1v7j3
HWkzvR9IKoidTHLtU1Bd9KcyoNh11U2GqD1VY6E0Pi04bxm4WyIPnvQHEVTEdrW85XC/QxpBYnfu
xyOQVDRPCHXw57B6z8umn2ATZxZdhn3KdxIwJATIB/BXyofWd1qNiXLgRHaYRZP/ytI9VmePusYw
zggFCq1jSX3ARtE9attIIXtTdv3yoAVgqXf6/lce7ySPf0vVXglPLKOPhj3IWBXf1ANY1TOX5P/u
vYFbrhpLVtVGYrmqH+dOShdgEhD9WO0ctT1Kw2IfwURX/EalF50vG4GvuahNDRiXf5L4hZznHCMr
vA8AP8Lxoy6vbLzYoYoD7auF4GpxGGR91z63XALKYdwZB4xGuR2V9UFLdLNDY/qw6qnToAMhJILO
WkzcxcxLjot7dOr1LND+PtwJ/MX3IEAYCI6ORH2A0J2eWWWUnNYNxTKkTHZH6Xzo3fI0HkqEMKwU
CxzCWIaOqQZF5lGujblRiSTCWZiPBY/z0aYLci0tEbZueRPM35W4u57xUSb4DcHHyuaLy4/v3EIf
q5UXLm6aBI5WK7gzRDwk1jiEO2dwZf3cfpK4WNJ9xaI81PnFHd4VcyUcKtUEwxmHtw8chJEkvb+C
+srf3X/4UbfPPW+ur7wGjlqtORKNkSK8dlvAkvyTMw8mDwDRwobVW9k6oe2PyNZMYOv6BtBCFIkg
TDv7ze0SK8d4JTWOkipgykH2qYhaz9H2jmeQVca9POAHjZeMZs+tE4SX9SzOc8uYcdftWN8CzBgN
wtgE1UXXZalikE98a+sW9Q9hv/hJOpbyro75IzliPSlSF2smqhIXLZjBPMrNu/kKzgSBVASDdmEV
AjdL3tc7lCY+xMRQWQMg32a6+Iw4VdM5Brgc8C/aYlxAuEnQ7D80PtyNP/6ob9cCuuoGK3p8T0ew
+HWREPz8DDpezAaxj5nIdeAWZN8eJC4OZdsxp852hFJPePU2Kf2v/sDgF9vAnbtvV6jymnpDf/0h
Wal8B+5soWcLOxzq4ti3v4GblUfMBMBDc256FON3YwHCD59YiIQ2DHfSN/kVPLTCHYU9oftfIYmD
RvwKx4PVl97SL553mu0TiSz+0Ar3GMPVIWv/NUIvBbgZ3Ul+XQvqvCOARYLGohQNPhBbwOgAjjcz
E2rh4vnDWfI0p5ROAI1XuQarPiwo+0j+DydhLjXY3ABBysikdZelV3wSyCInYbAKTe3dhXXCHvw2
NBMXBSL3SOEFZ1I9oUef2O/DhTd9/KkFafHw/N3DKeVRB7dCqGPU+kRCAcU4zKqsToHQ7IerDGAc
voGgsKw4MmsXUduN1MZ9xmE/Qqo39xD9GEcHS8ybaxg2d6BtaCRu/Wra6efRVyKKUlzK5gTXeaD5
+zgMc0IQy2MIXrg8iCrZ6l6SP1L7q6ri+pq/B2BGcwztzG6i8hLT/i/mw0w5kzB9ScCLZyWATsgG
8+16tr+pqwmqwmUvMFO042RRRot5RbwdgZqpsQJfnrX3QbNtWfqyt6pXR2M+tjoF7CNpxyPs4Uob
gQ2Gql335oXkDBIHvIkrCoJ8s7st0IZVnhcK8rBxcJfftibe9gc16pslZ0jeJFAyhjA1sNenRl9Y
tnLpmseB+yKXZatPWRunnfDX2HF52jUVfhboV5oeNj/oZFnuQ03hpuOiMLKMqQDJkc4KrwN6quti
O2FWhqSWf057i6bkpnxq4zN1lX781oJwgqVU5d+9nQvn0jNLx4QfE2r4Dn970UvKsKsPC49nN5Er
vvNZ5YG/3bizsDeqtxoRpZsNyU9AvmT0XPmuIbeA3JI31LUHe971/glULj3IaYEuDAtg/CSH+MDN
8mNb5xFLErG1J9ifS+W6nOw+Bs0EaEwaKYmDQjrWDTCpA91zUOymKSW33NYGXkAL3XCBBB82IilE
XhWUy5GxVtnQ8naCW1x92IdYRO3r55Xa1pc4IHsu+NoeJwi3BRWooIab/wQ7CZCQhHyIL+pLUhba
E1CKLif6fZpQn96W2oK73lcw2jPLPRKF2pOooGwoKgAHoPYyeFXIA6Xth3XY5FDQ1WiRBCvdv1LR
wG6CLt6dfmu2OCIEAL/K6iN65ahadqvllN50ByZ+mWR25MvSfQABIOeorMLKEZpTHFBVNU4lSzQV
aKCxIvngn02snEFWAmr2qhLEPZHR+SMLe2Mv1yAgKmPOXQhnpVGVA0Wm5qhnLk175V1KjFW0RtLi
VU3muDYPJg3oVCjQl9wsQkTSKBqRA+tX9iRDoVZbaqHOwCQ2ZCIwaadSE9afuXwk/YL+43OVSJRO
F2MyyezYbUz8Qe0pz65yD2O+iBBP7Mk+/MUdr9ENalhBx7tjYbj5sJcsUffdzLy/CvOXpxEE7FQf
Xxo2Tdk4LLj34x4dpYG11I1gyaL+uqieRfyKjUjaKfJXzb8WT0VDTi5HMtJb37ji5UYcyDw9Na4G
EhDaNXjYGdEs96R5Q1k4+49NSIvpe/oM+LlOPFcYSCkTdtVu6+lqxaLPtEC/M8jncjN0oRobfbsb
T2B9nO/fpaARP3TMhjB2GgnO0WRNBWkD4mxkJfcAVXwYF0znrN4sbizaR49BNUHthMf4neXcb8xJ
9Jl2z5RPc+QXCPeYvuqeniNRm+ZOeEuhb0FY0FtTIFV5yuXGrrUQGfOpon6HT/uBsDz6DG4Yj2R+
mIa/wd7TMlSPLrxar+mxVK7yhZzaX1NPv+77RvIU+wDHxwjlyb5yTANQKgO2DA+vKauBPPZl6l4+
hXZuvuWguzQB6hz091O4mKzKbJpU/Rsbsh3PNa1GAFzgMCaaUlilxZfuIypMuzTnA245tGY3HrJr
VcckLb1lSfaezMg8jbk1/AVRGEkrsvLAL1mZoDv0vP9DxdtcqXa9tjONohKM5GAjvPgVL2SMm0C+
qbz58DIX1qcwoEdeApE/VpWlquNYyYChwuQF86CdHLBNbyvp62SnuBRGNPZntVvCLyif33MTaAYU
ncVToDiUm0eAN9K8ZtcdgjXk+OgodJhLiWEtlznVQRpoPp2FJY+4QqmdKIsnipAH9oYY44AwwAVx
ORCAlR3JqPQBxl07dxnKPmcRE+u6MK2a4iyMajN78TitcOLlzJaZjdkRuIP352nSuRI6pc2Clsa8
0ZhQ1vGF1Yg3j4B/q//5IzXJYJFfcUQoF2pUTkcPTp6ZWzmoIjyWZK/lWIuqr66z91uHcRNCgc3C
j0AbhAfVCY4yDSZ8/8WSR+wwyWt28pAR+H3q6Q3RC9tSGL84wQcp5zGIjljHisVf0kDH4dnj2IsY
rVODDbODdfyjmtGdxrf0p7gO/L8aNhpJ2SwDV3zWJx99LoKGpZhPBGyZu2N0230eqblSUjjVQebX
F/0MEASHEzC6NjlN5mNYpoIdzgcozCEl4D9ld7/fAU668p8T/9G1i+65OmqpHiJHMT0ktcj4yC4I
fsRqqUS/UCiuL4BBHC2FWoe2LK/9GSSxZZDdCSCCTFtr3t3xXdUhottZgMx1YStkTk9zc6qcve+Z
g9b2xWe2VqMiUK+ChYTpawwLydrsdJCrroYvYTURIBvLNFeqmfnqGey6g4pug6rr6FY/mvCrFuWR
fWksBmC7HsreVbT7iZVv2bKWxC8fpHDJSJeuGOM4Ts4m0E6OIj65fNSfeAFCD20ich7q7a9Dzlp2
mT7zPEhiwmTGSzaHQhnpSMYyHSfuITtqTwjve2Y2PwdRE55njlNuiQqq89LHv0to+5tbRL/MSD/j
g69CoRZhKwYiEhg1T95V0KQRsyHRELNlhVnl/MENjUTSjauS1FhMW8OJUYKg77hUeHTTKG4hSQQJ
1rKQ06MhV9HxECicCiELMnR93Xy++xLXsA2ZqdQPPfsUHGVBUjyRm0PorJJHK70azPqUCLfBn34q
RdkHP8RR/5+IEYbK83PpSuvSyCWyMqjIdHFAO64oTeDxm5hAhI8LRZpqidxDt2kIHbVrOmzwwD12
Fwgt0WMM68r5Sa/7x+Rxk7esNw+JBZTIjM9b0d/sSfzj10qHMqGYDS6iydocQGXJTvlv2YSX3BBb
tt2qfOHKt2G7QZAScFrH5o575o56Gx3qf6lOMRah9PlbjdZY+skEMHHrPgHDGkZ5P/t9x+kDlIFj
13tNvZ5UqARVusi8P4usuZtu2qZM6fLur919p7lpkC195ni80P7kqx/E/GXxtsLR3tENcHsk3zKi
KKL8ixDKk+PmTmuinPjyDPUuNpULZzqfht8YR3XBAWbKLCg4OUoeCL9UzfjDdzItNk3HavifhAbY
Sl/9hqUcea+WY7Ldp1J061XQoS5hX+hAKEVZ4gyVSNvcjLY1Vt59UWqg+Z+1gwbVC2XmqxCDC/ye
XeB5cr95BhcVARLeLiSl8kuhXzTEHDinkCpazGgBz4nfebZJKGN2EYziBW/lecledojAMkcb9tvk
e2ynbIr/BEb0uzovgAwcNyBiJC5ZmqeWdVogOpDikI2zg3siA83jVu5+53eWXnK6o8ZVJrlGqtcd
UgmGTDMLHAVrPsLFbzbCO9V6QR7w+HHlsVwjgEdA2PM8Et2vNgNKxLGPYHPg/huYVqCUOkvob7QI
3cD69fQZ2F2ut6y14EcunSMqjC0XvaY4OGdCLvYWQz4GHp/+gDUZBY8hscnrPvxHrFV6Ae+0oGy2
3gBpInbo5c7nVao1FjUekX/wZQsVbMhO/BjCIT+hU6pnGIx4xJoE+I/kVSa4EGUMpAM6xTMtv34r
mijIH3nIKnV0Te4VnAR1S2BlcR+Wv0s+Kqw0BexiJxQCWAyqdO5rv7Nlq3hfeX9yAjZeWIdH9s7y
6pm0XD7ghWa9x+afQJaP2AWhb+4SYSLmBG9ihqQ3zg7lFGWG+F0YsGkSEUswnCrdLc25QuGm3faf
tLDLlxwom1Dtc1Z2nPe1dGVhfnQ+5JU4Q6V7mpdxD01EFElAHvvFBt8jPHGyZPlT1jIlTB8VepbP
tyGu2m9BjvBi1p0L09z21M7hh4dDsf8am+04tm26Yyysqy4AZzlNl/Wr1s2TxiD2j3QqLEkwbrHp
fl78z1thQrIGxjAUFs7MqwhQ8yjMr7NBH2Dy7WZztsDGuStlAhPUqPcimLjLa0Asz5zuy4xBWcNb
tXP0MO5dOTNbqHaTFSkxJH8j2JvQuDyShN3XEHa78vbixGvPv5Yz+M49PS45UUBLsPLn0oBVLVXK
RL0N6dEg+Vk3k+9WNs+Ap/VuXMv10LHxD4bJUjS2bXGpFHwnRvYeM600M5Xc+hiAUm0xqgmxa/AR
saoF6Ptp+4bgX9Al1rr0yicI+psQC+V+O3wJ2HnklNJsoZxdFAVhkoNYcI7m03KVxq77f8PPwRAa
xtgXdwNfcqc0Y3vqUW6KGuLLBa30OG8uW1Z86suFXB174U0Yhh7kzmZrPgnf+qtY1I72VVmOySEK
OngDWaAumSX0KGY5yq1gnAZAypdLYZv1bfv4PYfzVp9ShSNz+6TPrbBN4/KBMzyFtUgmCJ3zmEiL
L+TPVpECoBxMs6L2EAH28evlz8EtQ5doE/2lQm4gmsVVLhhNAbm/26REzvaIpWiuSwCGyTlEmldU
Z9Qv0f+CfdJx6Qlf4Pq54ZMlnerTM9d83dp8F8J2DXeX21vdcYWNaXihwRBT/0aGMGd/zGCwop0E
+w+MtEcw0N3jPh7ij10gPuqCXOMNxKirgfXZ6G4Q5TKOgL6PRj2VFHrjyksqCNUj4zSoZ+EjtDvN
8+DY2ckys2FeJvg/otgPYx3O2uv5F1kF2Jm++J9iaSUuYJ1TUH2xaqsi/dAozaV5EcvgsIs49tQg
WN+sPddvrVvIhsrVzATNlHBWhS8MXB9Bb8wItMf0oxngAf3pxbWFL8OMNhqXh9TX1OHjlFYv+8bi
8B+PdgDiJXQ5E5KQj6Dqe5pcvhYQV+Y4U58zGxWX4JRg6NesvMNlZDgA4EokaGY9vd8JmPHZDrMq
FUqAKFz8OFMmLQUNZ60IuC4T+kwhpLW7oMytxeHz6T0OzzN49ni6GFe9O08Z3UaBuCGjMRduCMb3
HcDf6UZXUHTPfMn8S1gCJy/NHPo0YQuj6lvNbDtMx116way4eXA3po9BjFYdKL7F/IrN/sgX0eRE
7aABKwG8SJ2GJFjNcOxmwe3V6ke3ml1NioFbGrBK5aRaAv/U0W/J3eRT+dM23QEvyhg+qNhsZwYb
yI4ElLKlz3GB1ImDDqH4Ne1u4KeNaaM7RVmCxIKDLi0q0e0htpUy7VR7MYMlBPdbZy80IVjO8b0p
PbUKyEYa31DHRLfyvXASCtv5TbOOriUm0AKJ9Sc6BAfUAU1nkqpldEdfwySk+Q90tQ1fFX5cY93h
KX9xPxVUe/z9RVZ6M9qzIiODUxZYKdlsn9MSM9QbejPyR2sA4cH7M8DeoCQDTXZCKANhhqp1Rnzq
RxnUO/qCT7dzsrDZANXZuQ2uQHqXQF9kre02i4owhLvSCGYYO8pi8H+F9VTutBqCnlPoDamCNJD0
lkMx5qghTbktCFpkCq27gnkZ6RytTEqJR8fh8uaw2MDryIt1f8rRAZzLV3pJjAMnKegjvhkYzQjq
HojdO4n2l0anVccp8W4MnRLvms5cR0DX+kKe6VN4L7Mv13rlX50bJ+mfe/cZBHtMoX715qTXeRfB
oc1/dl9opYJGeFqWXPhCSMfrs7qhI4uz2YEvh7PIDzw3WYqFprlBrww3e2royqpAtliOsO+90Eez
O410FX8QLzho2pTJdHS8ONsrL9nz3qzYy/SUAfvtRlBZ/cF9lvDUVJMCDqPh5O9i3hWWnCSh/lEO
dbd2eV/k63zx9iLCNdsQyURi/1o5jzLPEARYTKH+RJ0Qz0QcbZRwL/v6BmZew4QZHz+Hge2wZwHc
P2sRtpKHkjls/R29e3ouLmn9qA2ucOMF5EXi+IUFxq42rlh14kxslZCWD6PLsJMDA3HTESBwpWO8
tjspWrBnX9rhsZj5b58Hnhhy/1Ogs4TPmHDEl/tlyazIQmM4jlV4GzSpFmyfHNY9PX4G07PMdsbg
fwkEsX349H5bKSmNLVWcdGDTb3VaTCiq2LgkKtVcMtq6W+fEI6F+JVrZm/WHnIFjVI6twxqJ2a35
3SawhFB1TcPRt+xEwyHLt9PijKurTMSmq/8Is8LupWeG7VOAU6bbSj27XuVgcVKzIFtYpauRNh91
DV9C13/Yp988nV/VcNCMwym6YOH9YY95MqfuoMLKSGgZx7BOGfhFe6NBpGsVXoFy7YJ6hVzDyzxZ
7Q1s05GKripfTxZyDezjSYA7vhAoXejTkLPoisiTegMzRZsBV3fR1N1aohJeoFFPwIsBhWt29XIe
bGZjUGOJZhMF4xxak1gJNVvO01U9i8005USGn0XLZHWqo16jyWs7a8KSetFEo/G2LT7djovtp1VT
CSes199I8WCngmgcb0tIJ3AeVFtBF/gJoIoCr25zLsI0vAn5L4gkR/7Lcn8EncwCZY6jWoph/r2+
ZNKxKIK2/T1a+3s/6gKxgZF8aKY1RGVbzWjoeJrQ9MV13dbXvRr3nGeCfRb3fIfzAxPtBoG7eW2K
/w2yjq125wFiypBi4094qbebox+jjdhYWEJvY7iy7rgLwIbRp98TQJqfZZmsoI3OG1ivQ1APfOmw
H7rAANmFRQLBUbeRHZXoSRb9DiteamLdbjLCgCMhqKr/bgrnoDvN6dtGieUG5bobNrvy39WMHHFo
CTE+s/q1lRJCIMOLWJuCMpEIFnSFbS5y9WBSGHoIjdA0YIcqFn2Cr2M0F0wIyp4dA7oXCcYcKkLM
m5g3+V4A/fPhD8aEY5MoAhdvZLO/kDNdHd9MdXOaPC1HUeG2SrYrYZzr5mkeiDJZGBCHp4NddAU9
otvnFm4bYyPpuUwdxFzi+Tj6inTlo/3MccpAfv92RZAKWFx6lce36WLfB9+4LgnGJ74lVlcCKmCx
5sqnzYkl8DmeLllANzC9sFDU3hOuErW+FeD8waN/5u8Um1KY3Lg8lynijRkSv6sFZKk2o1DTdO87
xLp2gJxARPuF8/wSjS7rfnW3bvI+5vzoo90eDZBMYzLGK8St+VH5s6yHcSSLpbgbesP7bORIFSEx
/qVV8lQVPYSamgpRzqKJcEcqS03rfQSIvJqXyxaCdy4K84UIh+MUIwGm/w4sgJpJ7wtqwuoA4syw
rzpUDnKDyGZywnutThGbsE+2BDGSNos4lkMoi0+6emIbNUjtwU4fjKtt+3NcwF7cRupOSTta0M9s
/eY7LLY+oTeYNRqWB1QUhONrkRQMP6uDpkQ73A7AkEXEK3TUBwRsZcdmUJKUG4ClFqXs08SwnLjy
mC26rRm+B1CX7uBPUpBiMJPP6UYwddlL+n77UiyztIasgDZbKkW3KJQL2KjcffVzTFatNB8oZv3e
0GHz3HtTE01FSqu/XNQlXVRpcRtDkBwyJ5QE8LhWBHHzuDyGg3fFX2XEP3eGtprh8nUz26A+FFxk
WYf/JUoRURjfOTWjVU4MqSbTxEruDMWQ0PAzJzqUI1LdMP/OKHbUPk0X7TABnhzubE5XfNI2Jrr+
1IMrdKV8HeD7iEpfuHlE7MTuRAPapofytohQHd9whpUZ46soZCO8loR3qohlZxL9KaV2uB6CQbP0
SxQtRs/NOZySNjEFAVCFoCWKQR8KnVn2ZGvmJxrMekq/GHmWLmwdYTko2x4W74xPgPX1+SXGA345
VlKwThE65gFo4Lre8lDpEp0c07aWjzn9cFaoDsf8l8xVP4fd9UEoqyQitAg7sTp7ZaWfhSlduwqn
S4hljqLLdpcm4ER1UkftDAKDJsu2a0haswjS3cFGWDfHsAFoaHV9yf5f7OpOxYcuG1YozYaQ7vdH
sP3XqNYJ4CxFaNqtB65Rw44Jko9kBhtkiOmefFLuRzj0KMm+RV1w5xqYyuInmb3zuvjMpHHzTMuX
g5e7qNObqUC4oTlK+UjMP7Jhwfxp9iuD6pmE7MK0G2V0FTOhlopmkLvt9/x/4gICiYat5Dk4S1hb
AGc3gWe8ztV/QLFAsRf/UN9KfuwVVrzalCk9AtbHWqwgUapHAZ2IUzJ1rpv0FXOGESlZA661+Uey
fdX3VFBDegTMAIy22vfNklovfgkTcaFwEkggphGeBWdEeW3QHEfUxntXCSxDkhINa180rHSq1mwG
Q2HTzHVxWEHtVrDO4/CAs6BYnXr9Q0SgckcZLTFxCiFfLWNlpU3PA+pfbn7cG+mjQDPs0nYNrD93
3G0lCOD1QcnwoG5NXYKm3l+mtTT3EagOx9SndeiknyK+s26mSUYHuQyxMuCPQvq533qgO2MrtqVM
GuDoIBfKaRXvZEgLPBID7BSL9PFqxe9itn0blXYB8FFiVGXsoXgHBVIS07rEnpYa+CiF1DkVBQdW
ABnHMpE0DkE+d/7JJxZbasjkKJedb3XLS2m0/k7Jk6TTflXpLMCuoxGXbWoP34BK6lrcU5OF+y+d
LX2ZMnKFH6m0KqlYzDSD2x9sRDlDC7zwxZWL0eNFiJPsSfRrZwi/hGZzmLuaqQEvJOnq0vOtFG3P
/PNVeirrUrzAy85zeuoAy7VQXoowGBBu6ucRrMHnOODLlCPK9ACa/oSs+RuVlhVHtE2v6usxGl2w
3V6F9LNmRE9FS1qt74dp7+avD1tVP5pPbs1LD/RcsbSWcbE0N4KjP1nAmaiDeYA2xg151o/jcWwz
FLtqEQ9AMwKFXhLKa+/r5aYS7heBS4MBLBobKhwKbStfa09ThMah0qj+0sgjqpUg6DttxF/nR7/9
LFkNH7MRJChy+60HitCnVv2jcbnlpQJPSPPACcJsfS9NYsZdqzoRPVV/UcuxXr1hjtoAbkO/jT4F
kubMhSHqhVYiImJooVKjGxQYDfXJ6mINWTcfcR0c3Nb+VGHB+NNbsOtD8cqj9z1c7Ds3WtiezjIW
A109YKVQISfqpHhTTuBgc7Zby8IJBacekRfOMZ9OZrAHloIlcx9Sclw32D0JsqGY0c7rmW9DqZi6
/TTClsE8Bx51B5WhWjmGGXDFLrxIuGvaKN2sPHzphaWmcJ4O6tYet3RK2VxoWfCTy3BQDFS1bEU9
SRN1ybj+rNE07PptL25qZV/N2B4N4O1VkZho1FLvBsAHv76UHs0vtWPfODG12SGuhvczvsBizYUx
KOaxq9MTMsQAF0dsr2kbOJAeFWPFStqOSzpXHo054V9ob0jeN07YP51QtwvDcEVuxscBIbLFpBi2
IgR+f2KbDSoYImgv9L1qqIbIhb2rVtPvV5vpicAFE+qH5Ea2RiiezwvWyfv+nhNsYlJxoAZD7q8z
XBdomH4Cek2XZwmwQLL2bwNxTZw/hTn1/NeYG8/1RqL/drQRpvsUeaBDXCHQSm6jOkRwBfBqd/Tx
/Y05t9mr85cAD9fNqb71Ltbnwe9Ry8+M3F5Hdon6lQNJIp1qA++PQgbsJATUuFkOxZNVlXaIFCrL
cemtFsiau0Bl80/bn4/boyj9UkN4TzTT3sq9WY6TO8BmbIGjgbOeH61rqtG9Tk6yypY421C6JIfL
Bc9xLXbKNUWs3zI2vTzHj+Hx+dvej1869oG5eG3L2jeimKSjcm81dhcbh+wJ5eaBJNZnFy0nWFLU
bu7MGsj4WbLchVRM8Phu7Hnkv7NoNAUumgiPG5RHmSzC56Kmmruv+298f+7mIAg/kJ4bqLwx5Zao
k/dtilgzHy15GcVRnz2E5x9xyfd+WNiRSHFZ+1ARdOISzRnJQ55xRvJdwA/NM/pEMUNeBs1TreJk
eNwgPClT7oZ6RIKuIqT9Fp/pmPeHY6DFmr6GFES3f82oxEESgs6OIQVBOoeAJpitBpPbMRm1n4Yg
2vmlZaq7u0QN014AZ3krVFmWnyyDuOla0H+8wX7za3H+XNCM5tqqP8/IPmXbDIYlBoXNCTC0ngJd
50hNdzw7Z2CpZLXNXRwhCXa+JEXFyDhO853aLLi1/AW1hgWqtWB3G0/djaZW/1qiS6UNO1ggZN5F
WlbD7aTwZnMonARZg41DeT/INHZeGBd9KqKKyj8FGW9HXkJmHyFuZ3SCZzkMzf6qwVXWuxjFGXb5
vxQmATtn6166nV4sHltes2dXvSMtF1w3BxYv8GeBeChep7FZ3xjauN9zJ8O028wxnK+PDhCKs/3O
rTPyGFZrHqYH7xgx1zCBkVIMKVRPv44OG1pgqxhLJByGiccRX3u9EbzzxAWIhZ61tpbGs8pSO/IN
LtQykCKpVIx7gD6AS6nkgiRgzz+3wx4oeigQ+QqYIGHVpjxlGuznnPuE1TIflhkyogYToJ4A/2dY
oHLSpGArX278yVkqLP5+KudWMt8VccfT3kwaPX7kVXBaBnDNdX1ySclRL9NCzuwevABJ+1NgkyUN
ihkwtSlCHiBXefU/o2YIYugBlB7lyJjEVJP1e0vccJoygyYK5AeQNDLbU4w9jH5Zel//c9GWkw5K
fc0rzkNR+0xuQCZOkknhfLEfLpq8qtiUZnG8Sk2XHzxWMARvngkNoy/OdiRey+fjFYKNbxRwHstv
z5GKWCEtssI222CUqd2NDWWTClC14j68p+Tjcjt3EsbCUcqK5j0MdnWYwvI4CucfJmXguUMtZBGL
5KpWQ0i3Y0hMDBowd/EB8qBV1FG44f6S47cPIf+PYZMOIJRbxuVdNXOmFBQipWY1/KyncW5qyKJd
7O55/+HEA8lEwmy/PQCegz6zBo7TuJmy80cj7LsPTgIk2Cn+Z7AfSyIctJEtcCRsr6MgBgfOpkSf
WSEvQBh0MNbaTk/I7dC0nsh1hGPhgdjLY8hLo/RiBdnQ5k1OKPI4Peb2mlvo24sU+DebvL4he1uP
PX3JbObUtMyirpFqKEykVevHtslOQLOMTr0FLysv5tFOBiXdWT62SjIio85bSQj6Wzya50NCuZnS
41XzS3aeZaI/5Zo8Q1v9d4JJvynkc3893ZPdSU2xrnhyNN1XdTvcej/9V6Kb2gOSqZ2c4/NWaO3u
N1jM7aO5NcrB/CdSglGj38LrZS+faT9T1DgHwpLcRfjWBCmauzNgFdFseuhz0FdFa0CHdqGdkYUm
kxjWqIlhpdoHuOeHEaTkl9DJpXzyHT69lWxzcohTjvkY9+eVkjFL3on60Y2z8prsesteXblQgGUw
iRhtIIOe9aTuw+SxKgzkjrMSU2WsGAE3uWPV/a14fdYMji4ps+DS39p2Pawx/RIybW8xXnrsToWI
VeTYbGcrqzwVvnZz5aFAY/FQlrAQrlbt8MC6m425ebcqEYXvLn3xfgNGuALnSszxdz8t8kPWquae
TUeVaGZRFO8PFCEdbg73bS+ThGHvDP0xGRymwze0eghtGSrWL0f0SIJJOTSNFwtTBZ8n7wMYxkcP
lmzr05uYFG6D3O9jXupt5LaetHq0CdQaxTWinu426nbUkOwC0X41cczTrdIF7JS63svGoOEH3kFX
DMDUsHF3eJgDx1kXatnE6UAMmGKjqPe0UCuhPDKqHUvFqe1999g7H86hmz88xKrK3M004JCuYeyj
9ZaV2PWqWjmUdGs3ZlUGd/zs0apMUfZBXe3YjmlN15L/0S400qcgn4JTMncF7X4YRavwPUt6Pyom
b2Abu3T72ZmUtSothK71bhXKd5civ2SlfYBMJWBhBcggTYmTS6lcdUJguTCbTAuzPRqvBWjRVydh
waDGnixszpvKnXzjkGrCkOywYbL6yMmy7/KUjxz4XNhTd8VsqTy4dptTjWllA455HMT6hET7opBI
DQObuaQHPtjeZdW+Jh+rQQpDwFdXiviOpwz6AXY2fRjBsQ8OJAYwvs/M+Fgyv/usNYU+GT2fKwtI
JVCSsLoq4j45i5FR/65FMEUYn5//HYwg9sJY4DJe+GNCgjuF83wyY7F3mECnc9e88dGGe2YwZnVk
AToS7sbzvSC9icg+83TImlO8hquMAnfmxDG7sKBO4aRSLhGQnfKYHkfEG9fGcT3aE5LzZ/LfPEVL
d3WBdltM9YQhRlltl7f8uVjJjLHoJNxtX5XjGiCXwwzpLinL3fqpAqQIlAyOccvPq/5dnm3xHmVB
WQX8iraPwrZE6iLP3BJUykVbcppnKVQJX8HgdkQhMdJ3VULsPzfv9baD0Y/Jc1611BFcvp0qyIyx
igbV23BxpNhgkkXVhA27SbWpWKpQ5jx1p5MDwo6aBgQWFsanBrknoqATQWsZ9kjxk+7spk9x6VoD
9riTqH3JWQ7gKP4eeHbX4oBPDmtFxmHTvP19oR1wU+s5KJQYDq0NRNsoDnfukT1Lj2ROfKdvsdTT
h+2QBh14nmhiTl7gXdaK3dkkXL8oo8JjDLQN1F45UBpa01XuG5dgioBQmsdAphAo7BkLl3T7FH7t
y6y8ufr6Z0kknjnCKtYwVdtBsHZ0b50CfnZ2Ftg+i/CnBsg330jx+39d7YLXkj3LVH4f7HaWKabv
9a5D0bSHJjN/b41iUJSFEu4r3lgbsa2vLcJghu2d5vyvlIsnE+qIBYcwkxIBSfWzhBKvkdHvTbPL
uHLaHk1dE2hOJsivnjKxYvYirfMxVG7b9Ne6armRn/ifTLfzj8Q9GIGPH7q9wFi4gg0ksIun0Qw6
1e2eOg/+Nl/FrE217vwScxl8CEH7xqPtxSSmfAQT31L/LOofBL3w6ypZF0Qsnr989tunxNYr1iY4
LL/5WbIoUksIsTp5KKbp7uLgWo9b8h4bkhUjH1RbhtI7b2pRwrzP8/sl3TMEyqyjf5g2qcqwUrZ2
PeH9TrEiPedFDQZ/+Xr5pybVzjWZfSWq1evWshvbrlJXd46ab7k687HBl7T9YLXlXIyeOhpDktx6
pz3vTnZYvs4iPVLzfvzxbN/Do/pLeI0Ksp7kd1YFo1IKfZNPdPaXxEPfrdxm5GyQoO898hvKMCPN
L1tEsQSmCSfDlZFYhS/z4O35Alb3QOWRXVgcXbNby2hLQPY9LEXuOCKwd61gIjsOPKuR5hFG7KQS
ZA6Wr95YGp9DcMhppxNxY9a90Qq8zosCrgw/sCWOIc48jjMZONJJ6OQgZShF+8UyTLz4lHFedd0B
LTZUF64K6hx+gbljU3QsQg7QDk2FvGmsmQILKa7LCsghr2zf6wp4UYmNgS2UUjghT6qzw9j9Yt2w
sDRNcHpdRiC6R2y2lK0zOqxbeVrzYsOYg67PC33uHEZb3kX9SFb7clfpuZSXcLSIduTKLW1JxEUb
3yxEC/yToVWcUQZ5P2kf2ZknAOZarzpEMQjEqsGH5N3u4BQn9Cc+oLAnJQRXuGFlpZ4Cak3iXNKo
QM49tUVDUe6fzMhAjTa7wWMVsbz6gwx8xoDYuyjiWFsB8z+y+K11UUDzbOJyTFmZDTTM9UzzIWls
D39tnFnrLrTSxlmFB1AzVRTHAsuiarP3TcNmdT0WCXeugmxc/FvXXQt209ozmSrtJLQmp4DxicCD
YFKwohSVPwudqXjoRzWoPz95Aehd1QGk3KWEhAdsoNf4AxGuYgqqD8ARRCfIXDNeLvOJi2O8eFnT
j9jNuY6TcYMf4fQRi2j+Nv45FHZGfoz8GdWWYqX1qsP24XtbOLxED+UbGSyiXcab7P3V4dBTwo8g
NMfwms9YdKst2nkVdOxX0Rmyh6GbJ2fEFuEbRXQx47IXndiR27xTnjAGjpggsuVnFuTke1714SOv
ggPZZke38Z0QODGhMS4iIYfgAQmKMiAwVnmdrHVYHSuYYDvBqVKRXYBoKXvSeFsfA6LVkcGjyPdl
n8mOPTRbO8QlWtSoaYn4D+ZrXXTc2ali2jUkGKsrPWWwf4N7x+teHrBr0eyrnBJK4uV/aibniJc7
zkaBAkZ3GB7cR5Y+Se6Sg4fKVAFzAEOpqm8pzx25gZil4olYVif3QdXmxM41KiEqinc3mbtsJBCx
dnwCw4MrKMIRJbvK0CVnY/kOBT451sLzW96qQhvIdakSuPeQtlBAtwPljvm4JBsYn2D7ZS+dJPWu
LSiSYBF5+ID0RqA9RJWvErxg0YQ6GasDMQwIN2gR5mGhWw6JoAGHHYbK456ShtJZLA++hZnLQYak
Yc5AlTcp234bxtTGODD0s1qpyCCsvcTPC6o6rcBwkIJZ7cBAsKb2nW+/01sGmOkmx4VVYfK0gOvP
5ae8zbbH/o8agC2YOWLQNTh1+iE/giz2LxsihAfnvEytioAKZ+8p/yqrWMe2D9cmZL/J6khLmfvJ
/WiyOJfp06Y7cJQLyqa3QBVJ94iNXIj8HWdmZICsJ4eRFz/TTqDciJ2Gh+HbU4jKDw8gbViNjYTs
KEVe/+2hN5ElJxEO1kH64/kW0kpCkb3160gS/aCxFhxkf7NrGpO5eJs4jVmBrHwO/zfU3lihmgVH
6C2giUquwgV9jBgAWL0WbVnQcsS47gDNgmbNenaEm4WLp+IvJmD3EBom0Z71QUM2YCbvNBHKwtUu
OkWMZMtOEeQfp2aKumeVjLlmhn4fOwAisBXpLUkfWRAOwTSABV5f9twR3gR6pjvQzvK6CvakPWPr
M+Cn6twFPmh+Px9t0S5s6+LRttXV57QqgMUghl9+xtMXqBI7dvZw+J7cuMwvk7tYtNoBL/UJefkt
8C58/qwuFLZGNj4uGhBtjwjLOgurJ3QuiC5dJMwUSurdbl85UekEDTlrPWzc4FLcCzKzGKmpjoOq
lxC8KeR9KgpzRvpCy7hDn1MtPB1yydMEWNRD6Xxp8Ed1EdzEv7lkCCcfqYCAFeTULlqxTWd5D1Mw
iqxDP1RU5Csj9evfxqYX0XG0roNRzyqLm2bSAGV4gIg/qQoexsyKTkgncaZq5d8zwU+LzapG6CCR
FnxsEYIpORPQj2UDCnzQMSfznohZzvRcZG66MgU3I3MqP1gScBdiz57hNXiZ6XjvcsHrbRHJe9TF
HCXsiSgSSs5pyPTrX4/S9fUmyCPtP7OCAvB4bqKYXKaDyQSO40JavblD6BenFE6f4GIFRe6kNpC1
U0ZGEwfK7ZB/ekIzzu1n29gjcq5jyrzehVOyfboP4hVz5WtQeBab8wcJkmx1F4zCnojaPzrMLNkW
Tu+CMuMTS9e3weMAAyl+RTj2RFXlbyfQkvG4UhQIGI06jhpE7uoxm65hlpuy8VD9ifSlek+S8AKm
RN6Fcnn9OlYO9mYVuQdzowJOAeH5Ne+j4LQL/7AyFHqFzuVT734IbkBc7rFz9JPjMUE7MZk41Ncd
BB/FhkE9sI8X1RG9gsZy4BK9teF8U6RpScgUVXMeac6QdQVHYT74NImjTSeZx2bpdNpvKQW+eGgH
US++cO1N/MiqtUWVEf46IuqJEsBuedOeEDF7Nwfq+GTPiHzqmlvOAUo5KvL4hQ2dF73bGAZH6JiU
V5V9y+QOLIVVc09cCI8Qa1Yf0HseaKoLRulBFH15TUwkwstZvCMDBfSnbHFYrDeLcawFyScg/IT4
CTbjn5iSNuu4qHcF2nUt84vRZ6xcGZ+8+OotQH4qw8W72Su0JUH10lquV8QIUVrK9ajcPsEPhvzE
46TjXzHdN0/+3f+uR1Z9LE7SXfwxmfUvzCZ4UHfq1pI73xSrycTwkhOdGR9heTYbGfkhSThwTblL
qYPc0kswgEa+UkX+IX5hyyVlEOYrW+G1f3frS7yltBDlg5oW7edsOHniBzTIh2W3ktsX2vYdZIzm
zscT/iKEi8eNChhJto9PxQ4MXKDAgRpqQQccbSUj7A/dwyLFYaO4qQDyZkUT2pfqeRdoQQX8RfVj
w9LRX9Xk3dwfUvMpP+n5oDfUEeSIO0CWCd2JUJ4UdnaEW4cP7NwOrhw3kBMBqeVeyIwdIxSfq4Mg
WOPSfsdgfMMycukGoolvb24QmZ3dZiXjO+xe6ktn0C/tIINusBHaRxpzVYH4JjF93r7EyxMvFNqX
qLFRap2+mjkfYA1NKepRxZUZfOSS8VoU2p/eVUKG0IE7H90P9xOTTJsOBnCW1l2vWW1gfS5ug5Cd
wqma7mOuKaDFrlnmPcrH55YoAxYvlLlnoedwtWltaGouJq1SqK3VHtHNu13QCoUu+BV9BWT3WHbW
YroOw77qvKuwpU9IThwX4rVG7HMX12wvgPXHcTqeY5pvCFik6OGi1enX8Xn7oW3hlfK0oHNG105e
O8a8E5F8r02iNSYN3DsC++O3QfvXst4U+MuGPQWHsrYzm5Z8sZ/73vIvG0CwOjs92SRhc1Lg06zm
IQIHjfZu+IfNUhE+sUgmtRc25gWfUdKrJVacoDV4DSUNdnQbz2/fJ1k3TikiR+W7LxDFuBRwnVL/
jfPKMC6qtd/nDHfH1aCygIdCS3IenrykEMwSdTNDgbHI5U+FjGArs5XUoEfGuFM83z31fJCAd2Dv
aKe7yFhjA/0I51snjWMwATvadBH8lN2JGaNM7XKvHKKmI4xAkbGFm13LcmBbPDaBP8TGMrIm2yAJ
fQrvWEBRLKudTVxxp20CGQWfxsbANCdnPeIY6UGHxzurg9gwEkjt8G9UupNg70/koGGYnskJCYwx
4rkead0+cgtrS86lJ7c+ZKTfoEq8DgdyXKXclrlK7osNpN3P90az4vjP67vKgRjsfq2jMD87R2zE
+LlMjd/799Wt8qrdPmoHgDuh2/yAUIUdHo8Qthgs1VImOT8Fd90z9FdbHTdTiaZ8hvOLlUBDrpgs
TvBZH1fXEy93YrTqn5c9zLAGY+pNkRYGOSct3C1jai660aZgYHtF4XXK3wce4iPIEDI8mon1Y/7E
cOoC6RCprVXycrdMk5tG7Tgh2kcp5/e82gJKLMZqjwkew5sHqrL/ypPHHJ1MGH6hDeN3vWRFKp3n
NdtwNAsuGRIXGhiicEKc1TAFO7nzfR7NO1cMDrg8VJMTDEBgugDrKUE4erXubS8En6lc99kjUWAS
wOICnCZM0XEMWPDQgufWjgFRrTLNn2S2iRVx/R8rMB8BnVgjPiNIfA2eIlKLO9tPFLwNSQypMlj1
LPuHK9GAltErow+LaJBcliBSsc1zBlqGl5e8gJviZxGCPD0HNTWenZgEo/jIaf21BspkMRZM8br8
ufDBcZdXiyB1CYeNnEuXH4mvjUXi5H3dGfXLMxe5bSAyEfbCqaj9kSCPJsz7OCLa1tKPHs2LEPb+
twJmhLztyHli66j2qmDQYLLH5BAJFSrLMHmzrroEYeYceBYy6Og/EMcYUdwg4ZRSKDCSZ6bFjNsa
n4dUBPSeodKxjNwagFnh3ajHbbCVtr6oQH/9oQlgH+jZ5lqemA8XyzASMjOBH6Tpzj4fA2kOs+kr
bwWVgxk7+BEQcsAz/C1UFQoSQDUXTDrDkiJiME5T/Y5cGmjahHh+eDzh9gcjTtkG2UvmDptS22s/
o0I9dCntbm2mX4M45zgqxQDm+HFYVe/OXJ/RcGG/0JUQifLk1F8+cy91EbwdRhGKe12GsWVYnHYL
etn6DdvSHADWir9bHQeRlNQ5CHpBmoRz18YTVaAZM9kUOj/w75PJ2IMn20tfpKyR4T9UTvnQ44PX
72OuWC634HJkyTMx37obFQ6tWSFqTC3CL9zFqtdkd/3mjRaaCAk5EpB8OvHECDMCPuXUlWwVU+HW
MHnzQUTIK6kmgFR2vLpgivTGMprNIq6t5iXX28sMglbIbcjquUZ3Fr7nSkiavYy4p+tYDXcyeb4L
RyXGjfOqJ036Qdx8PAkosn1K1zG9GX859b+fEF6yTrpsjSUZJ3tsUJf32vBl5/+VSQUUaquh6NS5
8XMLd+9bSkTI2FSuYCpDOidwRIELhxOnYHpX8p7KH1t4bC1KM2VfYxmcZomwmkmisN4PDhVb0YJS
iCTSl7dr666Ha3NUvKeYeCJhN0laxJCQWB5X/d6hy61upb9/r0vI3u95n4FhfXfnKzN7gJTejERD
8fJbUBEIgtoItnXNrXUZfPtVQsAZqERs8GPjgFew6czrF+7Zvief9UjK9ICWjQvYr6vgi97orRHv
b39jJYQXj2eF4J95opIaERhMXvuggWSCIK35PzyuYI1UaDmPsH9Q5RFXaSj5pBoHRXBzbdcsdhOF
iDDJeUga0j7FOPH2PsU0KX6/IYjewzFrikbQZ8i1mAP0zFQLAb0zdGmVsxgXv67bslnAodwpycWo
PRYAXIvI99BWU8wraBqA2fR9lUZv9uuQrQ0/U2qzDuzKc6fx1KMvrEImnK2DwLAb+ayvpa3nOGpt
yLBHWGy/GkyUTx3dfbHHk5s+eRcb1scXIcbz9K2dKxa8t8toRiJ4QgEW2E71+c1HlPzA/CgyLArH
5WnqysLfx5JfBncwTn29kP+03RycQniZB7/Swze5RIaJjBKOPTU3oz8uHXDA/NFP4XmZMx7QssaV
UHEqd7yXGnQkUNDAWMIBmSyOl+28rHkr6LePd+Btmywk0IyXTi9bunp6E1cBVWMDkG07VuVk7vCs
NlpV6WAc49t7YUWaXzy1/D1atni1fWlpWsoEKxEEYB81opISekHlqo9gLJU0NqGS/ObPY0u+kZx7
q9Mr/CZom2x9eUxDZbDZiqehdU6KGyE4rMGb5KPhXDxH8jyqa7exb19yP9QHTjw1wlt9mWIYcoHk
P3Jpjn2cGj5SAIVB2aBNL+9SjjvpPrQIAUpxwvcGrDdG76ySuiw3VAtNgfK13r9oTDJ3/kZuqmbn
vYNQ1FUoN6aUXNOXgldn/UCkF62YL1Rl7gFXFJJlzWVTp0xFySuDGLpdu5+zrUj2oFsflnC2Jhfb
vitn6GGByqNj545Q3+RNYX1OUFmmHMCPwI6pmH7EljtQWXLOrymc1kTY8hcjSONJ8JgIGOJN5XWY
u6gD0c4VVDxEHb4rhVsXuuGGFPPBcwy3DQnUNQ8a0hSlq2H0olINr974bAqxKroOM6L1K8xbQpfz
bpnA5SBKKZzaLmcUPO/C5ci6KkyTKAKnkX2R6urUUURoBDEACFk3mhNxS8X7vtEzAwusaUnEMWys
wRRaYnZR1GyT+FpxzvN1BfLm9C3XOwofuOjtxBHbA9EQOvyIHXCxeqs9nR6uTCqv8dfO0EdJp1ut
TG2souSEVtl9K1BvJXx2F4WPPgIdh1ZTkVoog46JIk9kLG2hHBO7zw/EJkgxpaJMRHQUGZpNXVrg
3NqAmpUikP7cKCzvf0p9uk6LuNfCtSvSzmb1M/XpnmbDTE7n88hizMNhp7Kkkqt+jABgtu93rBOw
04l3GVVyJ/zKhOEq9A6pI4epND2aj0TaOJP+m3qe8yrqawDP6atycCYfLcrdOmO6PvlCgOnrB13/
2GvT9auWwv0/BEU0J8yS9VP/FhNr8FDyw4qHWtSwVDrwkGz1rDNFMax/co1oIwSICUG0ILe7onbr
JmE1+QigAN2v9/N1AQ3cJD2sqAkKfZucSEckD9xMvxZQRIUnQprNt1gOf8GoBaVg7looq4OWTPuc
nTk8ERHGx3rlEWNqnCtDIlgjRsnzHf5DENENgJi6k7IssKmZUQPmh4Vn1gWANeKgnWfTjIdoBU9j
iJ2Nj451ZHEweqkRvuiYAdxJiwUnnWOj+p64DFq+yo32EyYbF9GJ5RW6cwyqb8QvBmswRhB391e8
xgc7WF7Vu9i/v4u4c1WL9rI0sr9ZOSe8wZxtd9X399xyTrqfR6VOd9eQWRkr5l3OvAH/zI9569Rd
GT1/Ctc3oSz4lzv4aXlJOcpGvYhYQmMYpGcw5O1OC0xj9ssVDMhN/i2spCrI/F2qzCsZtuif8XP8
iP+YQohwQQwkyx2yKBXsFXyaerLCdMEdD1YanXs1Z80XyDX0PzCUChK57ZaKzVKuTUzyx/NcyOYR
JopsAOAXwk5MEsm6sQPJTh8t28T14zXFsQdSPnGJZaGsNTGuJLXc8gfkAcao/V7MPq2h5xt3Sit4
u2fJdAE8OLzIqwmK+SgMoErKD2AM77ixGYlzsvXzjlrAnYK69hp+atkQdjeBE2IBnKff5qE2TL/M
7cEyeTyvB9TzEmzChLEZqaJmWJitGSKecq2R9F7VmqFOD3SjAotwnRQxslMz6oiANuszjpJP8z7I
0OiLAh7FraLGDZf0ILXjmwVhj5SZXsmUxyUNKgRlIgPKNif9LBkikHr8Bbd1pKthx4a+qsd+gCRo
SGYlPXb0SGCoaVMH6fl+xRNx5+i/lfXQ5qkB00IJPPN6jYFBfBmpSr9HT4HPRw8LGfcWKJpRUCjT
Zbv3YEOXx6vca4wkfICELrHT0cVQMx3KRJZfBRmsWsCrEyORtoQNAAEychm0cys0jYUUrJutm1t0
CtajZiRp/td8XojbCbqiXFv/RpT7W6CmSKKT2i6ODcRpw75p1giwIEyrKl8gTsqa4nwMeg06EEf3
CWxiA654gbFleDT4Sv1ymvPNf6y0TujYPGHOOe0+11TlzvMJlBly2aLsYzCCCyKkjQq9wDxGOwSq
bRTdXYXPpjXIskpedd4+tuDq8a36+oBvi+73gTUhWIGqq/vfCcHddgYIL5XZuK0y9iIuMnKM2nxU
KCBgdjvbr8qOG3aXVtJ5r4x1pquRnQ3RPjbCbjcty61s67btJAi47uGZJnULnNsG6kkhh9n7eIA4
a3/6rtwJLhfFgqtAi3TAs7QF122mI82Z+GHMkNzDCMsstdvDGjcWYPKFf9nPTrIbOgHHxTtnfiR2
0i0K7kvwh/3HdU8jK8d/iL+SCUpSyY4etiaXBxyQFuzUcC1axD5VGTMvH1HA51uXj0jkFFPzy01P
EMjIOe+MGJeNRgtmzPGKWGRSW/1USYn/vINw+OsuCuLamn0Qe8HBz7hx1Sidpq6NvT6jW64UUajU
bE2xBbdXCBIPqtqm+YwzXDxZ8RXwfksoAdgDLOl7dN6jevXCbZ11JJqresp4jEr9teZtlDI9DAlu
7WIi1nC5dzkx0jadQ4kBs9qhjpJ10AWvpXGiEKbAjW8urjZtwE4j1c4qWz3t2EiYAfXDiUgsp4MO
lqUVyksheVKSLhntAc/k6cgM2QMDPdM1cMP5vREbfmXe+CYz//dDkL+/7YFtvcZg//QyQJfo8hKt
iIKWkMgAddsn6sTz2hue3OMy9nLkXvhUndpl6i84yo2xt49jGzbLerbB3pD+B3O2OKTrDJ08PgyM
hovLUw5gqjU6BL/uy2eqzF6I/5t+0T8t0e5yidOMlXXtsg3XnHbgpnE7QCwqHfrfAO0QAIOdeWws
EBL9yVr4Sxdgjuq9aujcUnLpJEY1IrduENt7V3aGl8aguRPtH4He8++3EoRIQf2bgXMu40SeZ5Zw
VdcgboAh+gWjF53T5qcbR21h/CFswft+7sIP3nMKJBbDrk8W/ydmJGoU2hcaNCfKBGfX9e4rczFL
5QN7iWk0WhDY61SexZbPZJ2Zzo0Z2mAcmXLSpUWHIBvmBmnPHyOjpmA1ebcBILstwIVvOE9Uxuqh
hC+2Sgz/3Zkf8+VgYRe6wKdAdf/cVCoM04AXSSuxtV6xLlHCaq6e5Zk2S1HKCku9yCP4Ru7DUXMC
YjK40CHATdfGp3L94R90nh43kAiDifgVgZe6o9OTHQmcA/I6mK6/qC2wD+7CODacxGYV6SymL0II
f6YvkggPr7bPGTNMmcCDGpCwacU0AzU6nh4rdVV4O69GK1gxDhbANUA9wbrXVpBbb7mu1r99OpbX
nwF56rAHF2lBnpxBgbrebA5lFRYJoTfVzCRYgFGvjcS7r4KDIHv2QbqGDevtbGTdOexi+ApgfO6d
w0/BC4quaqLkVqAz+ZDCdsZQvfZHpgKxZ5qNE0yJEDz9Z0UHEeEA0PnHxOEgT/i8BUVbgP4RGiNc
WqxfNrXrgSiy2sIo29SgDg04eV0U1RHObftj3iQm2kuudfzp2s4wB7UsWhIAr1slXQL3IzoBK/US
suVvXfxaXLZmKv0KlK6Hbij7vSgPre7Q69kJxlmZeMIu9WxYcfZQYU+ge5ceuwVLGg5s6SZRpHuB
XKkqYZxFC+j1c7gPZd5OxGFS5erMelNTpWbFfb9+7iR2wDI4M/c73HDkKAzOhOdJrpbfGTEddpDS
TwnYqJ9/MgDSz1rrvkxfk0AX4OJHCKXCXPqiapfm4wTiFwK9KKg9N3mHRWllPlWl9+j6M10IIV+Z
01BVU/Ds2H51TaA0Bly7w8IHrwO04lx6lAfOVn2Bhbq0ke7DX5J9xvLo+gx8HZQH9yB3Y2M0KKBs
O0gr7KJqIS0K2Ezr+U3hrgsiBsaHbTYMJzMCKVeon8oj5+iR+Bc7kM33egC91JFyR3gjPCKapS/l
jy2X9jKr1rY0sqL0P2fBYANiM9dkiKhZdeE2RiO4pfW0PfqOhzPjnnDXlHmmpWHdnZEcUDqQzvZ3
73ZVPAnwaSSrjTX0UbAr+knKt73tiKJ6D+dPZngCroeN0FmEnaY+O5M1W8QZvUfkZ8cgdUMupYDc
W+FlMvKN7dms2kWPPcI+ElAf4W0OG1pbUZnEM93rYtBiuo7tHbmc3bxBXUO4ay7Xql6sELlFluBm
PnyNPMWMSTmJgO4RCsDOyjEJCQVAZcD4t8fA5/nhGlJcN6dEDA4QXtH3DkAZejMxw17kwwpnboIj
NEgYRbW4mkGy64f9CsJyFXWCdvtIeUiLdNzI9+oNba9hh8nN4NAawQJS+4DhXLPeZAR42wiedb9J
4cYH2/an4t5/P0cgdBbMFFuTOCgdxY95WdHExSPj5z0KKVY5iUM1nDJgWdPrYbIZ8Dux51unWLqV
0NhwIlhCaHZWmA5RIN8hQ3lExXOim7xJZdcj1873hu+bfBm5CJ5Pm7iHJX/bxdq8G61CqtS6EYQ1
P6U5cJ1A5f1NE33EAE5NpStJD0CjgRn6VUK8O7O8Gyq4WTrRoHItmN6QSLvqSeQMYzLzFJqcxXJu
cs9qqw3uB0z5OMV/9pY36Gg1ENlSI16HIgal93hZYjDnoEP46rQV2wibjjs/+2lZmK71RZByVoQU
TVSDAwsT48fLbjJUH2VQBj+bgzrVCWZixfoW15L6PJVy8OAMP9npnkfjYoXK6lsEEEIvQqtIU/Mn
PZMV60ZqO+9sQKR8fR5YZuldAkNLx9+hYw6HQTC9uQPYJRxCMk/0BzMMQsYz5/TWy4UfwYa95c9L
Qo6NTZnUdijgQ8Lrd9HwgZssMK7b46gTe2cJzZGqZinzDDZyPDOqGYxjeU7+LpbX6A5pA9EADNip
hbVix6pK5cm0zL++3HAoz1Npq7GdoJYK8suACpZzC8S+4hsi0Pvnzi/5XxVGBz0FHzCOFWwJKp5D
s5oPfqVBDXyLRY20sjcyXkq65Gza2sfPxJIvU14wl21LfN/+O1Ly5ulR2oDFTns+G/5oyUrqMPFV
pGz6It8CrPCr6e6HrVy+ujAkCZmNdK6L+J5Xp+ZHGYaI810asDugDoGXj9wRvpwlNttsrakYcibh
Sb4yMnjnXUBU0ngva6lX38tcXBOWKaffWm+x3boyn9EyOdr8geXN4h8REP3Xs+igtLMStUpvVC15
3I7JVj19IzTXgDBsufBwPv+UDSEcIlJPr+FvoqWcHTwnpf6go//JrpIoIjoUfs5SnIg6qdoMRK5C
mzNBFs496ztVGSprnSt7V/P5kgLaLCxNUMnaEPM+RxYzkZGjL4nX+TYHfsnasNrEOcXBD8q7d8ku
QsRQU0elI9ShH8x03kpsUj1rrk0yTf6nsL6iHzU5tNJx5A6Ax1QHsYjT8UvOiQ3Y+Cq0Aef+sOYs
74uO4y5vsTtD85BRB0xld21TGTFKjHQRTGIE64h0kcwSohv+h04B1jY8bpOTsVGBmH/nqxSRsx11
VwSbM3mViL0sEgJ31pdiuQ2bTxsWP4ooIO5J/0RBkSE7pj11zjDoTQNGGXrDk3lSJEOvyAX94QTo
GreWEodiE21MRvGf6qnhsSdx318F+nSztvldT5PcCHN5daQ0EV2Xc8shHN0K1zvYWbxe09ef6CFg
H0TO3+Q2qEXEvs4257yvk7mK45SGqNOg36egMgdlJnMcLXm7ZLwynH3bhZV4JQCQd2rVASYoDutI
SHeb4xV3josqG1DHe6MB8sdIkQXVLMlt0pu2gm8aX6M2JjWNIoMCUpkz2anov4E3JsDA1JBzkNJG
Y54lsMkMQE21mNKZoWBqjYQlP7s4bdEak1a3P92b9vEJk9dqKnUjOjVRQoyQFzgKKl/vihpZ5Zre
pjJ32CMkcq6QGSLtlWXJsMrkT/TtOX+e/lUF40zDmp4t2AuJ51XsJncYzMuGOO6AGbzH8Tjrw6Ip
EiamQe1UWrgWcELISwYyS5mVNp3Q7WQNS8ETCcz0oxk9wkKx7lL1jyEcR990Prz8NoCnk3h74MBv
6SN02TSe27OgVCIL4F/8AHUSood1HFA2kJJ1UYPBVfKN70DqP1V5XUNRpiXLH/pJ0tm6yyEQQWYJ
DeYb/aLKRKM8mxkJrdp2C0B55wqSVnq1h+GyBxtPagyeNh6jn1mn44QL/r21tJ8wQwNXHz00PLSP
gVh6E4dLET0+uC/mogCi8eELb9gm5QO9lMngAILXt23A99bhvnhq/o6Icsi7c+1XlDbTL/DCJs4v
33SQrR+jGw76f0/4ZwuMvjjAz/0nEXFWEtsd1J6RD5w9gjIfSgKp09wEcPT4DAA8bnby711zJ/Um
NJZ1fK4gGvpq2yv5ClqTr1eulbiQ/cqoDb+9JHFSgsWf/vZrk0+1A7nBULQAHBzWL3FwBGcnFLeG
KxzSUwLQGGDPIFdAplxi1ybAkK0zcFlBRDIzYSdKuF/okL0uBztHRdwcRHRkHjaBtm3bUsHLSPEn
SYrPT0cNbbzmSkADdpT8TW9Nbz446j6234j/KeIfYGzA1PHKEUBpOBGbvjHhQGnYW/48zzR5Mt8N
KVuAbyzHS/OgJj5rWC8kPn7qbTnoFotR+tgFBMCyaN/ZIP9RKIqaowLXii1533jVO+F9thsOzYx9
FIUrlvXSQbDOjIzZDa3bUKrFfhC2mTD3G9XckkVtBk/t04BeOpVOX0eRio/cR8xLDUimmNCTPTWP
OIBZI9rWm4cLmYDcf1JYRp4q9rmuDM6qtYq8U0E+wbS418xV6TZl0n5B/1ZpM9QmcUOdd7Kxy8Hw
s9AU3adngGTcbVIMrdkUZLjuzg8sMcLdmKZuMB8oGoe36W1Nu3jljk3esVCBJWNzRk8J7czc5hBL
i2WDgv2u2jOtd/CtGC7WfKkEOlBkw6lb2FuSZgk60haPC5ocuAmc7pyknTvXP1j0hSXXweQvakOk
2goeB4CW2Syhzzjnxw8bVCVWkJ3jDCvSVsTPQMTEAb2skhwo04JrQdFWIWSnLwsE/uq+LR0cAA7/
PiB62nq7rbw0pjmMZWtKQvRHhxj3vovEaAHEI0+vIROoiO+98hok7gWrDVDoD0EDg9QOnQPK3+/1
hczbpM2Do5F83MuX8ph+DyUSRdxbUjoNByp3LJTA1ATZQbMIhE4Z9e4Z4H1TGCCBGjHAq5PVRTDo
/l2deMc/6P0zAIXTpzdtCnpNqoxOj5NW13GU9N7e81lpweyhx1JgEkfef/69tauWmAD5eVcHp+wf
402B1HHr7GQixF++o0qb9Ei8afDekIjWVKj1MMNPIH92+fyqHJRjShl88Epcvt+P9L6CNfs0dMZX
dKUUkbczyFTf8302xCa82vyTdM2LE3/LanLJsjG8NWZKEVn7Tc/wvn6kqEr7nPedxb+/ztUbOf7x
B31xaGMY0EumgaLTTUg0BwH9NRFhZDFJNnm0sgokIZTYbGpHiT3OWLe51HyW/IH3IQHyUTxO+8m5
2aiT0dWpDQqYybaghS9WgBitvp6NVupSyTaNm3pTCe9R+jGLTEhtJaE92giAyAjd2MkPFL+Xmdtt
RKIYf+IfFPM0bafxR1uyVsrydgAF/IMPvUkWda4GgTVpv/GLqHZMcR1ECCMlYYFhg4dERh+hc2aB
MMk3SFnWXxohfIpU80sLS/hJfT2I1YlEefeQRZ2NJV4rweyrp6gDkGODY7a8h2CA50IiWEUYld3O
xHTxEQ8gAerUH/2CgRDeY1kU0PyP6Udg81UIjc2msJKs5ImwylbvNdrY2JUfLCSOQ1j8cUfu+XRN
n4u+3Ns47huT2hQhtOBUdE4seQFu1wPhXuLLN+oSYkFpUmiUnCj6fISsIjJeuWpQEyVLbMC99JAC
IoZf9mYrxB+k26sJyyR0YMRA/wawhAIj2jEJHa5BPxXWjiwb0N1AEWdgQn5ZW9Obo65SOBmIzsP1
y6Fry/uB1dobVBuiMZRwMBlROFUfGHTqYKIDCoYPpcesPyDFUlX/EL1tS4QrD8D3fx/YnPAlM2KF
fo1dCzDenBfKUT1DPQruY9gaA1rI+0i+SpzXIv5Qm/ZtgxOY5uU4VFvZyS+SRLwzrLMpRwAgMdrF
IXNwrG2OOPJZDN0oDqdWkfHEXN7SLIr0SrCqX/08Sl3tcLkg2kk73G0yMIPV0t6qsI04V/Pg11ku
8DV4ezc2kt+fMP55X3B3K2lv4+NhVttOaKeQMqcg5YrayjUr760wYFRwWuddIwJh/P9WwFElSdVk
9xFTUC9AciKOY6yM/GfNcHXt+af4aGc72BdKToALB/PJfFVwOpMbWObLAdHcx5ulQRYKRLXVV0IS
CSgB76/CeqhhKMVMte4zUrpFRk0zmRc9Va57DBIMEJiWNV4T6bnjLf6TMl47OvPjifYyy67MMdr7
j2KECXIgjnlJ6RyW/3yZTYSuXl8mnVK4DYrVPMPWYnOCF56ylgpKUOKAWoDWzVoRO7U+oyZP+/lz
V7l/D29f1XS5yhhn+P3u1TBWGAt70YOL7fKmE9jh2U+OQtH2rtYLJ2GjgYz2B2XruPBzmzBhJOBm
pJX0hxCx9WBl6njKxdk9dh58aHsKo2KmqObk4aZcyHR07zn0u+w1d9F8dmIFCLPAWoyKUtcL/lMz
7C/oMTblH00kWczjkRr9CYGsz/VfzgCvVUQf2d2P1sAc/rso3cJD9QGZky93eI1mLymsButb5My3
yPEighfnX9xbcqah0C2SgGZlTlJ/wzRLOqbRDPTg5HdXPA899Oqd7c4ORq5DjFKrzQYLBGCpcTIS
j3C3NDCN3VqXmLYQNMaXOi4dVaowW33UuOAGxY8wd0vypfJVpHzIZ6TDQNV0j1tyDeotIRDg6XxW
L0jCngMHuFvCvuTEoczcE2qW8hd3wpf32ZuyxWs742xHHqSgGTEFN6YiFBmHJRN50S1USH1Vld5Q
HsvNByCImzHKSoFt2dPgX7OVSj3gp+gkSw2Z2upY5AJ/8hRMvilGj9rocgc1+kUtB4a+yIB4UjNM
rAgotwcQal7W0uXEvbj4I2Esv+kVGMuMxqZEQE56DSodRgvJTDZnOrQGpka81cQ7wJCcyqx2W4R9
YCpuc5wXF3gHhLmlZlN3Q1imZdAulCdyybfuaLg1CJhk1p/Jv9GijcR7zoBpig8Bh2+zFo60F8R4
lkSuiWptxumo4Q5JwX4pWeKs6D/ZLfelyKGK4TeSxu7cfivwwZZIbiYornZ30jqrpAQebi7fAPsu
/4LrOA4RHGlvqZuXv9c/IP/xt5R0FggQu9y5GyO9l4sm80y/1Jxk3NeWxtSysDiidM0iduK4Sp4o
4YLvjroFeFOvik80rTXqX9B0oyFa8JLbe2NNpKrR8xp+Xbk4Dzb3bOgr3HE6G31v9/cGJO7rnKxh
JvCkSW/M+chbt+JJ41+XE4fzIES50wdpBx3wGBWUMFZ355CpufKmRuBXuNhKZGqrGvGR7biKzGr4
PWIymk8djsiMb5Z8eBdiTCe4qZFu5fIpMHFPi//BmAvVbFZwUkQkNjnDW6ljdK2Xc27DWB3Rx2fa
rOT2t1cCeI7sxcbtaDYDBygfzVw5vRlCc5eYQA+WGQaN8qENuxwlOuDpR1Ex2D1nFGierPFw9yze
atyEWQwksx1h2QksSwUYLXHw3cyBiPygDP/WVDfSmBKPLSgPvgwiVINcxG1DDvb5LZPtAvuabZUR
K0yW40HVIqXliumPIBk9ew1NdBh0WCZYZ2wVjngRdnFogvsCtih077Vy6CnGqzaOYHLMJiInspWP
zfA1PvJ1kb4qXHyM4Mcm+59aVchhHbEohEYcjnAIbePxw1gtFwqKB8rTBS5lChfRANhc7aQ/pjMI
c2ZTfrqPZKQDGDnDbFPzlaiVe06NGQcOoHssL6cihuuxMygx2VvxxVgctnl/hTe6G6z/LmrZuGJS
pybY3okGv7spOrb/yGLszvLcB+Nsru5/Z/i7RKd+ylFCFzv7Rjrq2I21EVkPrZYh68YHQPt45HPP
6H/vq1yiS7CLQip7e7w9vxnLepCza1lOJWIRKWg9WgAWbRyYpXzzL4u2aNnLyNlPWTAGGkjYEqhq
Cp6vwZoxgT0cToMOA639VfecsNTGJk2gUaQaB/lzfgupBKRwyEbbNCBLIibQRuOlysQk2tifiyhW
qKHqL2QL78jRkC3HZXlfAxushKLNJpJ4cLeIpIIGdyUH/i7N1/j3QbRCyM0Hy4sXjFnM2cLJNk/e
oI0VabzKqtndrlwjmsweissNvstcj7nHNHlin/3/5fyCIAN0QGN3nXMQIXd3WxLdRllXsXTx40Vc
TuTRjRKUkgs6SfHQwQwphALNdIfUM23rHvfrIKoJhoK7i1T3cGJzSNZ+ca6ASGA1dZkCnAcMYbdY
wrldcoWDKBWhL7kXFE9q4mIA9vhQlScb1t/pLbZ2cvbpbkapba4dzW8bwQ8TnrXBG5bth+d3Qag6
Jh9u7BVbhBMc2UBFZgBX/T3J36NDZPo3PtE8SAFsm8RZscIILbc5c+6FUtOg5fNMNIf6xxMiC3wj
3zh/9MAVBMELvbg9+4rXymbG9ipNhzFxFlHPgIMJleEYbJswf0Y1qSbE71zLVBYPpuXiPp4pblI/
wPVSDqAtDwSSzf7tkG6EhpeGZOjuw604kD+Rl+ePZu78KZYGqnVxk8KZAUqAJBYcr+3t1OUqNCjT
0E7Junw2RbkCdM15KpPPx0pqTKJf3qfiv89X/027KyVz86MLbNQqUZbSygUaFoiamuvsfBMePR91
Pq/pHB9tzLwtN/zgSjKN9WT4yxkGJeZeR+W9QmErDQnAtXlLxsi0wrBhu1X7yPrxD4BpvoWf5LRF
OlPKvkwtY8Z943bgXd6dRKHxLk/v22b7oY/car3ybDx12NKi3S0fdSBMJBVT/6aW6EadXz/VWstQ
kdNBSj4iNwVypyte4wzAkKrMof8SdWwB81ivHgwUxzoJO4GJL0CKSK0acG2YQ37ebJ0JqoucQXgs
2jozvEtfhTfgr8lgdDSZvcSPE10ppd1B2hVimxfd9aAwANaW0iofNr9Lw4qKIMfJDKtCkHdCD+X8
TOyARKb3U94Nb8McTy5eSJkjg1ztHMHXJ3TEvNbzOOTPEWWBdGYm7jR9HDu2b40OUpn/2X5WcgNd
tGe6Deb662S9L2VBSoeG+Yi/85jDpd8Gil3dj85Ns649s4gr1GIVQOIIb5yzH1z8GhivtVp01N8z
9hzf+iArYFUz4jmkryo0GBYqvEoloB7nQVrhc+2SX9NirPvTpMLLf9G6tnfvKvqJq4ukbGcZoQfM
ZoPSOIO6FjCtaOgh5+wh3KLt1gncFr9AFwti/CN+iXX6lwCLiD2ZNwZR4pFoZzdtcABPASCJn1l7
CSnXbm+fPRicAX960uaAbSdT37lxDQSYO7+Ty8/+P98v4JtveeQjdb8BGI3uE1zmWAhjQGcQOtHe
yDuU6T5+/aOpyvfeAVlciOucavTckh8wqz1Hp2nQCmd3TDiwrAiApm5Nuwjss/pEBxNn4iwedZ+O
i0I8WYiReCs/lNVSFfYKSZF9ajSbfr1ubJdmjOGTeSaR+2JAkwefZkckiOz3Q/i6dTOaZOTSvB7o
W0IOPP6yOyVxvJFUORpdCvbYw/h0hpy3PpNsGEvDehumX1O33gdij91o5bPexZlxEyfhnPNynDli
qtrGReA31S2zyG4DaCN9t9pPpQGe4pMaCONjQ8ctT0orjc9rvHM4hMTWjqVDdGhwcv14hupN3xE9
HuDdG0QhYENYJ+ZyfOrNXGsD5f/Ed2XLeJA5l5lGpLKl4QWlu7z90RzMf6FDzh759rZQWBolp60a
6+ZboSeOx7/7hi5hfhslwroKTtgBGMyETzpqaW1IcBkqSYH4nENkEpkVK1jIJ2uA1brzZhPBRLkT
xjBDb18wkTLEpI+OSg7cglBm1DbBUkfBanmuKey68aBwyvbhKn8eYUFbmdiesvgpaEYNuV9rgX1s
DrkO1bQ0YYwr0SnXSxuxKq0mMExveryr/MxRrwcTgHi2r2VkQVOmzkFWRAL3UrvMvi0eKw5KQ2KZ
yohwjyuvCXNvPMLAO2KvSweR6LUtGDh537kq86hfnprL6XmNuj1qgiRCE4GsFGkqD22+AxR5tVsa
SK3KJrZeV25oZFDEaTeMsLmHdKCLUXFKZny08uNf9mVM8TDd4d4m4EUrE1c4lmu+QaivTDyWUQ2A
TFTLGUh5d2CkWC+A1v7bvc8CN25y4NIAonxQC8IXtmNd7nCbR/PaR2fs1ytyhBSkUObvwv5T6C7i
+DQYLE2OlB9JQOjMtemK76dEUSwkuDTIMfMuUmNG7R5ZLrlkDQ4WVIASHoy8R4tt9/tmeT3ak7uH
aqr9a9BRwziNk4bS/LdVrqzgTeHcOAyWaGd8CJzOkGfQIfvbBwl7oqCojvh9o3ygVk1nHX5Irr1w
bTr+NhqVhETMtquLXUgnfVmxvSJw/aJy7h1DCcbCIcXgwVB+nnaSNBOtS57uSoI8RD8RbtzELunq
jnh0Ona1QIRWQcEmwrNe/TRYwUdJ0FSdWslQFH5q+KrZW1Qs4WYYhnXlDRQQwbT9/HaHENtGsIUK
TH+efV2nli3AcCm7SYPK9ZUdbQ5ratB4Bi+uqUuisYUADBRyCXXVnOob+ANV5u+QMoH7hAgHWgQ2
Z4lqJqyxeSyKKTz66z7aOF8Bw3tquOO3UYM0DNOiW66hYOVrl0FoYaLOvZ3mVhSj+VqS7M7FiQwR
0UyGmzx33x4b5KmQYgtxP6c0DzIpewJ4nbE02pYbY2BKPHAscZXN/mjppwpyjcRYRkmSdrkcQLQF
JoK+CyvW9DAo2/yAuU5AAXknLpiZ6UQFRGBKey0lBDA/Gf2X94ozxByCq2/zvBN7zOVoATlZROQQ
cH7/oAmz3rKuFX4RNpRar11Rssw0lFw3KBeapiPv5ywnRFXTsr4u2UKMbkKt/Wtn5+13vqx6AFDE
G1MoFv9TNBeY4Yeyrg7LziBmOsZ8b9KxqHHc90mZOk7yfk/lkEmL2Mg7RNRXeWwP+W2AF3IBnEco
6OaPDbTeSytGMO+93uxhn2c4GldBXa4UNLsaxoLRstprrg0+syPwKgbrdVLT5EKQdqjFFEfRDImu
mGz0JEZfgECGaOH2lGicekYK9fYYONTelPp+h3632Bz0CC5IKkE7XChFt4q9LszE5ZO7/tpDnkQL
S6pYCP8wU5b+pG15BwwjSDsoP3qwBRAVO8Ri86Ae5JaPmAT+3L4TEHwpP28t3dAXZV16iRaAkx4e
s/N46UkvCkzfYDrGhem58KLMhtAJxA7LnQjyfMiJBTrT0OwAjF7vkuMERs1UCqTOjOdhHh4S7DVP
Na1GWgkPyFGfMz78f+lx+m7MLqn4cbzTJ57Dpb4rDy/fPkfoMTLr7GxrdAzsn2BXDvILq4An62rC
r/gW8B4LwnTFGnt+D4IXXb2vbWec3LoWoJHfjIw+IV/zuQgZTzSklWV37+H0CRLNcVhq0PTrF9aj
ta0cN2enTnJBal06rvWcT024KYRW4vlnvbI+NSzz+/jltf4DyTjVQirqwY1cvNSWlWl0ZXvHmfgo
yqvbsggfjANFD2mTeRszAkZAZJrLoFrbRGFTovcS0N8l2nwx3VMkYWlwrhjOEIlDkKEw3ArCw8LC
smPpUDgP3TwUUu8/RMbkr4dMekucL5ocvR0HnBSrUxH+MPED2y7zqd6hEqMDHfWO20L9QI70VfUl
mxEc3j0Oz0Z1elI9mVgYq7bWhxC0Pj5dvyQgvFonsRnKwnPQs7hqacGlCgaq9JgpdAhm/41IkGxv
Ti2gDHqkd3CMGBqEtesAQ+dTT703SEdmvaCU0uPbqHOO2IOKtfCBoct+ReorXAqEO/oqoS32szpM
79ipN0+9K5DcYak2CHiyWai4Ei887bX6ojYBGOs+hn0X9x3BeimBQvQZgKFc77b5Qwvb89lDzFCy
KWOPYDTdJ5lwMTaYQ0e6gN1ONwlukU3/FJnys/niKS2OkT7e+VZD6Ml5PkZDou7bvNXM1hp9aglf
TDgdcLQc+vl3/wk/7WCTJm6ybkcVnIFZqyqLu84rW3h3wRUkFXiK/5LkdTV2AhYEmmjymEhb1POf
ZCHlmPthEolCs+G+9JPFHfUKOLs257MGWSj2JejBg9iBT5jXcXjFdgc4XiW9lv7HFj3lnxy+Ii+j
GmnWp9AZaUE0nGNwJ1hx0RkxxVuN7Vc+iNTe2nw5QKJdTqYTmKooFGB6Z6vp9FLZ8Pr6kT+btjB/
6TV1h2UIwyslwBW47Uh4oAek6BWD8FUw/R9INcO3n9Em/YQgssGpwSqq6CGEf4HSxOhsTZOVUOeF
cQPR9CzqNfbom9t2D/iEvTGmOg5mhzT+HpVhrFPwqYPYKqMD78ryqf1yZ2z5jWnEe20MT3nFUEFn
M5tZRkrVLFOCuPasjMzysGZmM4TPJDFsS9rw8xIdfKeJaTYSeM1VwWzSXUhGQHgCvU9WfZ9Nvg2Z
fGMBgOqA7F0BtoaFB6TgA+/dPhyDp+thxq/l4o7FebPj0lIprYVOb2AfMGv1HDYugTzGNxXHP6bd
0nVJBZgDh8DYCdte6TIo7G9ZEarcsaW4iFx3PtfmRyjUO9NBHAAgTLucllhz0DlWr6Ni7vsA87wr
bnw75vWxjpM9mySeTdb2wP2LXgua8LzJ7MqHOvuXLGFUOIYNCI5V23NMf15paH5A6YMRwkk28MHD
JDaekqgsS2gLf4SPlw44lzLwC7V3+zOKFQxp0oVyCKch7nauBnfy5V60iU7Z5wZUFvV+no1+eXHu
rDZxAx3pAs7kggSIUoD4hO3lGD1wRKIaZdtCyb9JBZaQk+t8nueVbBauMiGFOdo6Dzm3d4qDXdXo
cahl6c6cCulJ4LhBGIgD+0+iYz6rjp1+aLRse7CQhbNUdvoRTzdlvK7LLnXnku4xCHdcX8o2Q/sr
VoglCDH2VXIHtLWM7HfUHIRgXy2tbith5xkxjtC8Y4waV2YKdbZCrEgIWzcGK6MAfyJ9kKBKbGp4
VEppoSESCAzSExjJJCPUkG22IC/zTqcZvCu4Ve4kRP/vcQDv5JdTeYkDoVmA8WP1a87gz90dpRCB
Y0fE8tbwXDwwLdZORd5sWiAUE4BfQuEizU5gS7O4MOYpw/DWT+/+ACUqFaIKA5A+gEt8XQdWn+nk
+GauH5SYxPNG4t1aWGEU1IUd6BtHIQE8BH2iP/oNIRiNaW7UXYqqZhSoxiY7XRQcb/I9PeKpdONI
n9+seb7eiZlrVgrE0PxFDot0MNTyd1f+pR9MuJmqddHJtVis6HqhAiLV82XBvtL6J0eg2OEv1Vgd
M9JH2lDb9eLwczqoZMzwdztkYNJRwVbIs0ErT9Wid4Hfh6vqQiU8hUdDL2CczUHcUVBCfnbMoIYQ
2o51jdlsdhX++ys9eKgEy62GYBBIeok9j/1Tpou1trfXKeM3TYwrBUVuOrlwTwwl0iQf0SDstpT2
+57TE0FZnGTp/MAaPE1QDMCvvh0RUitJIPRz51oxXK3nnxsrvy6n4vZ+GtMlB+lb72VZidtCREFW
4kOJDlu8WHHzFL/pgs1N4sQoGcgdVPFTJlf3vduYLifMHZWfl3LeqfZryva/U/qqjr19zsxaCRex
TaUvyVl1Mxd/6lrLfi2H/MLtOq9zplv0w0Xoi7PlAsK73C3P5SH1dY8WxWlgo3OW1OXDiDE0rBx/
eD7aBGLZDdE3uDyGm63GpifrLfKc32XL5QxUiQTqOEaVeYfaCxJQZGS1by97OQ4e+tfRR6D6dzOf
FJJNiJtZSbb/77wvxMXn3iu9G19eA0t+3Kxev4cIY4nW2oNGCzzJ/96Zqj8VzW42fK+vSOKNP3a5
ptbV4MWyNBvds64dDe12pIbcw2nHL6/r2ZLSsuPip/BSknUe98uzllLFVr5EQc9MTtVA7NNd23FV
TafciZ2GwowUHm4Uhd4iDqxk3nqywYiJ+ILD8MMj2lXd7py+WviLre20dv05eIjQ+hnsMDAk8C6l
HykBGVUOUFLXD2iRqwrEdgCzU0Z3WCV/aKFf0mfjLPVxhKQLQ0sd6d1qQ8nOkP2yIfg7+73YsLKk
yFKV0O0qQ6QSzXYDbO8v2pZSD8P5ZhvEyvhKPiyIvM8w6+odv9Dkmooz6biAhMmNNaPb13iGRTlz
4zV7ccGdZ1hfEcbFulbIahZYvpmfK2BsnXBg7QralDvVKqN2mY7HarDovFdzEQ/mkN7ssMZ8tyOr
jwS0cX8/q9IHbQ7moQAb0gf0Kyojasi4omqjjWhI/AgJZUWg/HHo2rALzl9vfTq5aahxAYnMhmpU
V87Xwb1ZOk2DRHQdvIEsbXomlixmwmPwoSV8NCNm6StkgWx1Zx5oiNQa9tgDaTAt1jB/5peE3IBj
/IyEdTdliMwPY4vcRATLCTRgckABIU1Tk/cG+Wi2sY3LgDVtpnufssP6B9ThO0cYCqyQPc7rmeo6
PKNhgjiygbmb8XUx7bOVDcQUpGUc+/qN7NcqIIH6hwPq6Xf60PlhH9JFJ8/QZ78h6Z9+g7hkwrWf
q7BjibZb7flKJglhiJRRR90wcC6ParAfiOlqQoSAZKoeXt7zSj5bNuZMacpodd2LZuD87vIAEqmv
vEf3mCfgwHJ+KFwz7RM+rcirDrzAvzdvfZNuoZ4QdV6hcINy5rb10vNIf6ExPagwLTnItWUI07gk
SN3KjMfmajk1giWBqvF6hGmZ/RmMS4szNg7Y3yDpKEIq/uwCsaQIo/vTAkgsF2FEc3r+imK5Vlbd
RH7oaZ6RxfyYMKlzs9DMdLiYJWfldotxyQk6JN8OZQBD1KcPVozGWlR/b3ntd82UZ3Web4nl29Z0
iRDqgkwgrRoDmEJiOFwpfsEQ0ssaErTyelWXI3Pawd6JyeZoQk/wFpOaHVQBfbnjFo19HeHYS9Dx
QUiRn0AwohBIYjv7HG7r6bdTyU5vqJsoSVjnP/hF2cKg70JE8yLjHvCQ01AJBkhYTk22Zf6Ispl1
NNG67dA0k4ewXotsZ9QKvMafEnUYdyLXY64ovh8Mmol5bb9APyZ1bnc/mKpaWONWbfjpTjwGBpnX
tebU8p/wXxu7BP6inU8esP5C767PyDeoIezd/y1O7kHJneISh3G+VxAgWdxPo5xsOLkXGx3GtS9s
vgWKQGc8FNCsXSqny5r+0ckEvj8x3ZoQup6rhmiBPjzpHNYDBkQNsBK2w7UTXNaofU7gitwcc/Ul
7qm1T3VlCYipwfo4+1cgYSWfoXBzF9+hp0sy1KUSjPiUPu6J/qm8I7ZB1BEWGOjKDKSg5qTyHyVa
3E6NR8bZztO/yxvCzV/GKYWAEoGmE+BqngcRt8JU1/fcSuEfjRIsTwnBu2/bwKNd8sgsfjLbrAiS
QRniuM3Bl335fcN5+uuTiIYr7w+PTDF5ZHJbREkLN4CDFzFGUnUdy1qgaHWzKN/PHfro1i4pm75G
Xd2WIXyJ1YskIoSTV0MxHOm6x6lCD+BjMLnpKxsb0lfzvvZpKpBGFLHFnbNA0miC9PxX9X2vlC6+
X6iE79TUHdoLEwLuqkTJHYSdojAFZCEC+/YM+FFEZ5/Bv0FbwEmvwjRUfW3J/00m7VksafPJ9iZm
qNrB+T6yqj/CjZZY6ZUwCdGjoluosZ7q0FN1B2ajBlaJlL+PqN85V7KpmsYhcCwEre0t48LTg9xH
ZxUEb35b4ruFYfSshfB35ooakoE1b0IunsIfumDWSCjDlLYo6YGjeToEcOiZFG4Z38wOxmxjWUTf
NeDHAmZi0IoxPGxo2iwYpN4ul+Qs7Ta5WxJhPxR13/QrJ8fKI9KtILMjxilkM5l0+HfQQP/BNPKg
LQqVvf/uX/pXlVnfU2ZeT5iomYBVW9Wh9dqUf6UN3AMPJ4GSkYGuK8Nizu+C8oK4XNzUOG9lrOv3
DeO0L07PUqSSOLPD8tysx1ekOS9S/8UGYdlFtkWFNEqnVlHC5W5rnsk7rbRmVviYq8jV8/GfQnwh
1029CYVGaqQizxXbpoeOy0MOWC/aUVPKTWG7RciavbRw3Zjv5HmbHICqSiRKAD2pbjoLclvKW3TC
Ake8Cf4N0FRxR4hIjQX0kTFB61oN0KJe9z23J94MCzqLVv8iYf9zjlRgMNtI7su1Sa0aHwoYjvha
WahfWSLEpVq6KIheBOtSHKEULF5I4gRzw8H13Pt2aSvcWrQQgDz/13b09kzDhFL6sj0j54IUV5ig
Vd66mF4Us/OiuZXx0vuVqGhTPH/wFmdSN0J4yiuSkOvbdrDbxRTDhPv47jsbOoDaJA54VT0Hb5xO
+m2lJSwawfsNGaVLOQlI+jynCee87ojrOUe89pcVtzGoSCE8Cauwc5y5jYz3sS2r7mBw9NlCPD4L
F0vgAf5m682AQdTL5E0zIvhHB21KAb0TbezjfFNnOFg3R2oyPph2ThHsha+tqns4TKjzG+tgkkAx
1Ln8JV4ESNZobdPj/jxKUjZIJvpwRjqNTtl0gFFXGMEEF8iI8Uw0KuJQTjBu8cpheKqor0KtfpJE
OHIep3JDHofnYCuDqDTA4FlrUOdxINVMZWTcYqtlstNc6EI5JIyI7YX+1PJdn3QFt+L+7w5L8EhZ
wSMSEhvOjpcQsPMbpvW8hj7uYg7lgssADePIwd41beFpFuuee5kNN5BbhNwAg2AkDp4ocJ7y66YP
Ep+YHEArTzDzKTHvHG95pZOdAkHTBhh2HmR1ySIt6vSnB3M/ycxSbRcB0iMEJvexYiZ1c6LEqCEE
eHSyTUm9jWVG/+pVVn78YwTabRBanhBcofFDmCWluUGsDemcT5ORsXCZrmtd+fvNjYzu+LxASslY
pUg2lz9nIURFYhW+YS5Ls/As1Sbb3DNN4P+sfpFzZR7nDAKDuqBKwG7KZ/tzTT+KuFegE96mxoFi
9aY6+72V+hDG7R0tbb9cJ6f/+knxVdoLg2sw3/VlLXS4J0QDsGxZPFSDNMigkMzDPyvXWGq1PKTo
xNf9NMINcvLP8CdAdvO4Nr8VusvYBNwcdB0GXcMKkXyHlVc65xMsurQbzMi8SbK8AE+gFvbSRUxx
bIFYHOBUtfoPidh7PEyVE1QSUcLOxYH6zaBjwhHVZGY8d5Ues+gGEW59qUuEu6YciK029VHCpEAz
OoO5k376AN6BbJ/OfXcW+qmBh0YUWjZlVzm8lgWzNP/hj2sM6s/g4mx4dJzUGZIVoCaZyPfj50sm
6bA8jAWo8zntat/2qQJgHu+DSR2P8u2vbthcKKvcltVdpnlASg8Ccb8lJfb0CnaKINxkrr+fnbgu
UTKBIE282kZSuMIFILmBrqcPdCgT7Ld4EWid9ejG//Axa7Ugop0cAMceMYoBmz1NRBvVH7yLPHJN
uO6JwAvnELkG70+F4N6aIoHxB6sM9R4S6DtNLZ2YHC8c7hU/uNXzcr8NzACugN209MGVLXvsqNsI
EaaU2xyNkEP0aMT9sguS8RDD2BViSGbucB+b50uGH52gB2wfXZYaMjds4p4iWPNZ8Nm8DOsqiH1o
SklJvGoT0O7m5ggRKG3MxfwOLsJRI2N+3jvYEzKRvgLYJlrmzAGrQjiiX4i6Pud9KtqYCPULZsOM
2j4l3I9r3v1yiy5CpdPXDV55VuVCDDMQG+yGkwQA0DaGG5N4A7saYoaFX7n4jhoTJ7mT60mkWpdo
UUpjoS9Ac9CdeSPn9UfqZAQxcWdCpVpGGXqTCYecdFV6BH1hMsOnrWqlc8GtdptrKSuTGivGMjZX
xJ6feW1W4dnQs16zEnuU0VIIXMGZT5hh833tcIUT1fuoWsTXDQhsMEwU319lj6m6OdiVx01SGbGu
6XVsGVB3cqujG7woeYLOTAduDYgvjKtUbztTbSjT/mI3RNHU1QcwtTDeASSezAZNnl791WCUTODt
5v3+6CvT+XtmDQx2mQ+SZCpTdPkTQTvZBWpY2ByjBWPT6huB8gTVtFDlzw9KQ+m8yqWumlDNqr4G
MbtXfYC0+8CU+Nv/QNZU8e2M0BkY707FEnhU43liHn40JWqWYC7dt9LKPl65bJK1/6iCWs+HXcs+
gcLlRj2CjTwt9b53kR9jfJx1fqG1h7SWUid1rwMkMgoedpwyrIDvLxww7O+cCOdivH1KDmBbxLkd
iLByid6J0/6t5HYhMKMA6p73S4/53rDspheY4NvxcIrNk4tWx4ajfwzQ5u5ZBgZ6QwqdNF87KGVY
IFIy6cEF1pNF/Wz8pQiz3A/AqDw6LGr7axLuDbtjhSDFLN9iEhbzBstG/bT3h2krLrYOfAdrD37K
o6Y/D1MRjdO1AtDW3AvwwsfBjHYOfN5+kSbrZpatbidHawFwn2ZljpXxk0KDIKDlaEYA660LGl+q
+yOP1oewqr8GZMIITHJUCK5G3ofbfQFUs8jJuNKsF0jpkwPp/Ze5f8kkBestBohHO7itevQ92axK
dw2lODjgoETc7Ggoy7dLc3o6ZEexeycyNXyKXh2k8R/WDq5pbVjPii7Iztn8+zWfmG1Q5RqyNmzW
dHrcNRB4Sz3qMnHEslWY2AUWtTm3LfV31cR/DXQHyp6AKXeNA+eKxE6EsXzjX54ZNTPj6rulNmnn
YrhO2w506GeAolI93bkoKjc8i0rNvWhGAcDH6ZFqJ2TrzUj7vx0CreAVHWsJSlwVo5P9zy/MZg40
eskN2rIgJw1gTvhUVI9Gxk49IiBiNcw+RixLtuyFidVq9lPq32fPQu3AEARoDS016bQdl7mN+tth
8V62Pu/XJrA4oKn2xU4oGjbCxzm8a9zFCog8qjBtacjn+kVrJ1CRqF3U0Oa2vHUuwU4S521w6G5j
jh4GMdxCB9R7K3D7hgvNW2Qyxldbax0VJWMNBIGPcu/LrFZ/n2z0PnrbBWkXBfHwPFHJJah1JTbK
bm40SyRwpHpz8KjShoIUd+2FS1Yw5/9yD3HtftAthSWmQgLP6WkiV7739h8gWGa4bDjM+WrVVc9S
OUWNVqnOlPG+nHRCm/AwF4wNGeXVPpOnyFn287/VAQLl4wyWzD7Y1xHleDQTpcjTlL8VAORgLEhC
Tg0ZnLbpo9HpoqhKP8PveHGoPf66pQqEQAQ+KI6TO3qie131EVyxSoIP/KWxWfHANTJYZo1Zidol
Pwzi/vZWGMshmL1ju5riRt4g+A79FBirAHyxGxQLsyrckt1h4eokXpDKgVmvk4AppDSTQQKTVLMF
xS+hKeioGggqQr/1CTyqqHsjoK1sicp49aEgtAR05sy2ADuzglsZSZX/LpvC3AVhZfHgJyBtiHLp
cLcqGAp837CnKStFskVRrkH6Dt5Vy/5GW6JkY66beQ4dGHcOzWlbriy1NZcXf3jYZXJT6JYxgLq4
ujFgA06Kc7zWTEydfEDCgvjc7X7FbDiRJOSS3CHJt1/wGOhorZFTWq1xBgoQrD8cELZy1w/hvdB7
CoodO/FrOEZ9nastsdo/4NyRKt04WmkBB5yyl3O3+0BAR0kB6vqfqzAOatAhajo0Oy6kttb6XUX3
hT04Qlihj0j8DAl4eDmjGd4jKxTpBgUjVw/nWp1P2hiahyWN5R3kc7oD53LBMsBFG2daaq7H/IjH
kWJ9sUruP2vZ/MJy2VeVA5Cozk/A1Mc+vBB6T1MG+SUxt/lBzK9s4ifGqS4tIZxtLbkmrCm1v/FT
D1xs2Nzman+KN/Jw9evUY/F49SiNT7gj5QF66Zm0gufJpxJzP/ieow/ioXT5rJxeHg3V9rcGj5lH
wYKHhAUTOAQmpVNnQzfAD//WvT0krE1IYeBu0O/J7cxmwz0/OJdb0/MN8z62KnOlHdOVc0wPi/tM
thkqysMNfm0sO6oTbtWtPTNZce45lkw4eriKQY91pmpQWzqOj4x1DjV2RKkyVCOnyal9ghj4MIGR
nnBrbFfD0mORUrSBPrDaXRIXjPL9rocJuKKQXuNcuaQXijBv9QXiAEDTu3DFkYq+66mkAvb93VT9
ZdigxBWMO0OrTYMkAlEbhICaX6sAMKu5LtQ+zzhAEIADnRsfLwFrCA8VlVoUYlShOW1mEIlihmXh
kyJ06VrX3BJiRgQkPnaegQwAZ+YHl0lJji20VD4cKQdVgaVGaC8FuHiERyiz+ES6FxoMcsdCCTbl
cHn/Oe6c8fb4gAOSl1SahE+CDqWxizFDd+MeScgoeZ3RXmJKNVmztDYKHHZd6+d9zLLc8OWwhgsk
djoY9S7HT2QRwM+E6JbTZfgacWlTJvU84Nnik62Jqw6vNdcjVaZSz2zFbF5zAqCw1B1U06ULql7x
6J0ah09IuOqJcqPGnu3dHQ0NFLyhubMURqVvGiQBYj3JU8o7bzjG3oVu1WICzlKoyUPmAAfJP2A8
4Pcd/Fdn5uaFD9wTHCDWIKSYVCXg5xTEIik6z4YV7gXRo+ER9X/aFIc2/Y+4KjcMYD73Ag8ALWgk
SBi0lGdFD2eD4L6TJXLwNavQfx7MMb03H607+IFMXlOT6XSch5WY1WWYjq1MLZPnZEFFztGIkjRR
QqmgyjgplHdUQ150lo79QBVs07Vddn+OP2/+cAU/oUb1cpZ/tD9+H1WYixcL0xKYDi0ajnXkPyUt
ffkyqjkl50p/OCeyfcGR7cD3MKfA2yFxkgXX2P+aWS4bZekYQNC3KMCQ+zGFuIJ/6gl3uWcUe6iK
s8FFfat3tMrsTHEYeaSi1W8tNKIq/8k2LXYTBx+sL+DhA4OaMEUqpF21SFgXAyCrmp9HnNkLmU4+
xsf6jU6FSGl1MdG6qatmnpKjdk5XeOyBGQY7zVtuojfS/+MlGxh4suhJUjtpZfwcIZHjLJ96/MOd
mxClJpveljL6r9KCL1Iezfu/rphmaYKAeGOBAlXRUTebKx/y3Po0OgOpM8iU1c2n6sK/MplUwfAS
YF+c9kOCH6jyd7ipEo8HtgWCSjsBP+T8h53/XH/gMus0JMgBZErGYKnbjq1AzFSs1DkieVl0Zs6g
waQ9MuVuXSGMH+D9KAdMYAxksqwAothcuRdfDrSVT5AK5C34ul+wHvGFeU8nEzh8Wc6kPoJsZuYP
/oz52UfxsaQgwOHg/XA1ghkqMOvMVNPkcCtE53OVbtMnXg2RbzIYv5DbX8LPKGKLIC62ugO2PEa0
Aj4Q7JTCU398rVtkGQXeFzn2OU0IKgOB43rG4RltIMClCJoAhGZJaoUbxlQV8g9bvMEZNwTUYLqO
NxIn+V7qwNwKEQtvNRCIY7Wh5e30g0DnP8kWWVcuU9SCl6TujnpqCItLFn7RlmDz8ZqYAV0GUBov
7L6nTx9KVBid+gVivz9B1PMx86iHYq7i6USgFG0Vm3C/jxp0CE0Z01ycAEsGBeRLWnl3rs4b45O2
IpNWwag4Zz68WtdF1TuFaX2FG84ScUG8kaT3W/TE4brLS7XjYw2ogK07x526gHvZd80HPdo13nAy
4JipZUq1LP2ZRKFtyjqwD/epm/5tJvlAnpU6P89Ehnm9vDf0GnLBBtYnYkAqgnj8AUQReecRZ6Y3
nGAnKHuAU8SF0Y6bvQB29OLQGnqFv56diYsw3hgYbZe9yRE3L2eeuU1TUJIhR8BDHQN3CzwwCyeR
zzFCGNt4o0RGc/B9A+lq43JIlSk0SqTb6kulyDtsAhGju8Xm/O+aCMValdyiRV/D7lJ5vzMBW/8T
292xMhkDlY2c2rjyGSWpMJg5BvLmBfaTO3W3JzINSjwxG5OkQWoNx4OGWyxydl4ZKzq05j+OxoyD
reGOJbl9lSN1W6K/7lFdl+/oRM8LlDdx0IEq/pDU3kf6jr6GtSbxkBxkkD6Dm9DMQQNpmMjPz4Wk
8CvmGe7ywYyPxW/8aWjnCXCZz8GRMYwAz0gcLxFbIRmXFOC5I+uUUFwQaRRZgbWVq6YVG4iUTuw2
ZQSiM5ZQclSpifDJ7Yjk8d3qUyz6OOHQpGvLLyK+cAwmWYTZmaQnpl9y1dkM+7g70+6IJXlnAg8+
tAuX7tPxBtGaelWIxBrYlgDkBZ8Ox0ymULD8ooz6EMyO1eTmZT7YKgjDp0vHByjIS1JIw5VVfwMl
tRqkRhHepRew6PtxGgO0YECCmH3cwtPHwA6xgoDq2vWYHFgdjMys/JF1kQf/9p1j+3uBVvALHQBF
sVPHKKQnL10djrjVTfksmiQ6CHwxWUnu39zD3uJb3Xy4jIxrDyJolnCPlN2Fcl3AeZnkJHO2ESFj
BArTR1yxSDZNzvzIEKIpoHLpzG3F54xh2no9+sQHtoTb0lVmEGKX606vySU6fy52asQN1aRx+Aqw
jsfW3SNAKrV3OaxXRzpSkXkTKeRqOxq/aHeHQa9KdEXDjD+piQ/GihjBWWrbi8EvZwRlrGlhZlK7
Em0qDwukRUoPAqMhQnFm6eWmpP8ibtt1mKlvsDS1XKgxJSl/ojeSnAQQ0AwZ3UGdECARa0XHR//Z
SQifrtRRshfDEuRhWB7GRAKQndW3F+sJLTs00z5VqB62T/7/WGigkFtK3bj/L03VY7n0u/fKqprY
YRfMJ53j/3EbCDLBanhwsJM+fjPaga0D3ZHIIaeJth7ixJHkSoIbBGq4HVJMnmKQO+AY/Vdu9dHq
kGaFdjvQ601f0LjGOL1mVvoeZTd+CzulFXSOymr7Rkf3NQXCkfQSQVewW7KlW9t6+S53d+JGE2ob
L1ko+l5Y6vd1iflabuwoNNIjlRF1ZIfdjmx9YvcrVnWqN0dGEN0zhaMlbAI/tjoWgalYOkQc+RI2
Tf//46qFWD6C39UKHfUuO7zeplwyHBr1PwC0OXthe3LT30PE/O0OkLSS+JqUV11rgeqi0hPgnIpm
u02tmC/cUWRy3f9Fl2ELpSQBwCs+lp1j+oj+KaQtAsl3ici4VGOGX0Eiy3m/2G/TKEhAxhPC5v/J
Lbt14jMfQWBFfAwMgIhihIzPKOFEX4ZBB6yFbbwhOqrlyiuU7QhHz57NiF9b8BfjuHLQJ4qZTh1Y
uHFQcXupISLZEyjxaTvKg5huFCZQjemslryYBNqDszWCTxBKQf8oM9aq/qnxwckVh13Py8tjKSK1
qgY/Orl/8fJ91+Ax052lD5UrRXndAZL1UjEtfI37l7pHPPhqrunjdAxb0aToqKMklftk2M1RiY9F
pi8pR9G3+puB99k41qLMBK7fDeWRrWtLn+CdLdSMHV7vfzQ8iqxaHvn6PUN0IOU8ROCH957GpjPU
UJm4qSIoXqv9Hoql5NA/QTNmV1Av/vXzYtqTgsIJd9YpOXYECYYxeb9aZcc98jcFYWwpyDmdReJU
uFGI3O9ChKO2lUoa/gLUD4jFX9u47FB635uF6a9m7uTPcXCExwFUcGZv7c3I4Wc0DJC9gN5b2IX8
OTUeiA5QhFLrWQNi8pVR/ET2+8BztXKQr3SZ9SEezn+eIlSa2t98wQxLYtKhCkOVdnnIiuOJ92og
Wr9JkoqIOBDkYibce0ILvLRMoZOkb15YuIBk4WDdEj/FHKZsXSsoa4XX3Fw/j/95GBmXJywQqsPP
way1ldccnint8p6B6IBNeYMrhBWMNp+MpRsGLNFStA71r8M3ZWeGF9acEqh259wIgJ4LzXBw/XjV
elQigapUZsPZjwdOpHbBuu5zySx51IOoK/v8o2T+k+pvCnfcZv12pFYkXuLm8ZBcWgoYqHciExQA
/laxd96/A1QRzbFTT/93k9Z3dQvzSx7vMO0Zhs9KJ2LQhQlLzYWMck/9HWe+6v8a37dTxeTbk8cu
0CFl5bYC8S8z8dBLyROy1uYjuK+fWMmQ5D833s5YuPdDr7W//v60KHL7yONx47TZ3pfBKRV9wD21
vaTLdBjotQYFo1EcuA+PPVBY2TjAaWZSIqr6RzEy61jB1D8X1Q4pvv0bIC4xkWEJexLVj/ld+WIJ
3eBGmZeW/vVT74to2Ti+cN5H4ZrRbint58GyqFq/HxQS+irn3ncksxjvRTr1eyvippqILZoH58s0
9Uq3RUotQrbauQulCA77HAUtbHolSZ9wc/aYx9jPBQbN01gj+taVi21QbUOXjyMl7+bo5slp7clt
EID2CjK1iTHNEsGpJ1fBUJR38sWo3rKVgiL+eOP3ZnBY2KyBN+HygKC0obiWKMpD8fXN3hxN/sw4
Vo3useAcsEnamXp3l42O+1ensHLhKH8qbS3W5lp1SnAHx4Mx9i1BAk6/CfhceFks/xJItg6ebOBO
gJgpcKYU6WHY+3EcBDMbkvDopqAMqoWLMu3dlv1ztgptQEES6p32ILG9vS+XiULrmgDZweR32OoO
zusgHmwGsSkWnfSQ86pqtKlNodS3VOnuc4Vl0jdknlwR7kpoYRvyScwDlLHgY7bDXUTRkA+XjQPO
ZvRU4sJfCCbUUT51G85jBSq0SFobfnBrOoyb0SMA4oAIDUI3gzuGw90VERCANm+lv6m0SSmwYt8V
x9dpNwtdPVHU9AIbtp5epxdBxdcGV77SAvXMlpITnVYjK2Ysj6l3TCXzv5hEb1lm2NbMLj2cjQHX
c5hMqMWGSYz6TBs0TnmhpXsBRhUjAYLs7+329Qw4s9efMXaaXMonoA2WZRQSfSiYml173iDkxc7u
PUV8N2qOBdw9tsP4znN6JVFrH29AvlTapxiOg47tVoqPhKQDUTNOABNcxFLPU3X0LBz70x7DAgKZ
87Uz9yaglSs2rungtafY7YCJOujWRZ+kQPpcTtj+RhLZEXiS9HD3p6JC7qO8KHCY10m1Q9LSCfHB
ls0wGGIemlDxyecYoa4UbwMITpYWgnFLoZtTw+efnxFfQaor41yH2ZCqb+Hhu+uUC14QeQuB4wmr
XjXtYQ3ZKDJr+DdN2YroFmwiruaOS8HJ+M0AldViuAua/1ZW/QRkfsrAZfWCuiav6Kr4LvlLtr9z
7bX5lclHGLs/K56ELKztcoc7/Lg3GRyPUxEU1NBnuxRS2wywDnwgkP1FtwbIjJMhVZ/hbP+xG9Ip
xz73qyQTS6nCc3rIYCjFv7uUWv4RbCvPvpPA8Q5ZjikHU3YyByy9Q5HpDszQ7cdSuItSYvq7RkR1
SQSVhQjKPzQakBGaIl+lEy7A5g/9+BVPGBJCvbipdOWEY+kt+zDwQvhh8Oo8COg8lWV8XiCvv4Xk
6pENWtJFKHXKTBzjYrsPxQbaceaTtm/4h6APFqiVb1iyiOCQ5Rsk0To2fAItahghdDH8MCrO3XgT
Rhqc62aIlRD4RSeMyh+jsa/GeqQx/s+KuiCvlYKuWleyqFF12lXORhMUAIo1JWCSafL1BI5wXt1z
VqQWFmsTzo8AhBcASFazunXCjPsNxWHFW29KigC1nEBDj4pS/7OiAxpob8BHMjCGxIeb954ZbC1k
7JHNzo42SEfYzVusSIjkA46brcqPvJptVhuRD4Rp390iRyUbVAYRy15oLO2RspYINjJSBgHGxyXN
LSx4dI4xNbC/AFjUG+DxCVxPKljSrT1jyuKsnafaHpfGg8qoW44pj+RKgrKGqXC2293JeiVIYwrT
qH7zUhutm/4VJVb1sUFzrmFvZEAreOuCKmCcv1SToK4Y8q8894MQD4Ppd0I7O7+1yV2zohk1EvPO
/9+XFRcfIfzTYrto+rNp9SGc9CP+GGUQwlenicD9E1x3DciraQYkFm7qQZc1t5vmuPp5Xxr6+XsU
UBrkZC21giXNpxKS/p9U/8opKYplFYCAWJ0xrE2VHGPRFLz8pbAaetZP8Z1/3Gd3CGEqFydblG/4
5FJj5Qu6GTBWW5+OngvnKybPY6HwQBYs7hOA+FgrRwqbDI5iXxEOcVk2AvRZaXGYi6z5hSnFn1TV
JM8Tqd1clRztjeevuHcYnqafy2k3pK/4GCHcFfxE94sworsbLIQiyAtYPA/RosAqEhwKa7mKTsMV
lHB3xhic/HcL+1DSauKC7upYNwgkZZgEv7cs7CEOZCdj5GjJ2Ackaq9C5KX3gYZiVzaRfLXSThA6
m0Fl+lPfjnOgCUmzrA/I3BC/Exaxg/Ae9enGguVieXoyNsuHMoth/YOX39kwTLAhSOeHgnb78+NW
xf7uL4vw2Uh8gXdWOB0V7pze1/Jyo8xdYJqm99I6UdHKY8Rw4v16EK2mdlAgOy/luk9gU8X91T5h
9pIVyktMFNTQQjqMjnOk98x5xDQs/4AAkMKe9m45uOMcZbkLvx0F6/wIdmW/Ogvlrx5S59njBRYc
141BJS5JuCO2FsT2htdyAYt1bShvkUJthFL4l7dnr1Ilciz3IgsD6m8KvWPEpRT1MS6I8pQBgXAN
wedoKucIWEl5X6ck7GBNonFMExdXszw9qQ+3W0hAkrI6GNS84eIy5klodXNKIB2g1BoaLeErPtHw
T2cLFTT22WoKV6ACihuzqXobEaeAxmwIZm/H63+N/HqnJT7vRJuHJG5Q8AWsEALEsL+vg2z3OC2g
Pw7UGGj4b8FP0zRzs8I8mJEfz4Hz4rXvkBcwWSlAAFv6T1UEiGqUxm92C6dveARGc4hiklnC0gPk
8Gp6wt8EoAptkOghJSYpgjF13XRqSxpmXdW+zu9jHmxBDL2pVCnuXBOXIp0uDY6E8zpWIT2cHSZT
oUX2UB5f1ejsi3pV/1Oi9qrOzbJ/8HO5GDppsSKTnVHX3+5GU64L2B8hZsSHz3W+RFPYHnK5J+5N
8p1e+lb+WJW93ddP6YWIYiF4z7BmeHEtvXDaYB8xfrri9Oe9HjBGdGtAG4yOTImIFgcD4YIXIHC0
y/q8L5sTRVEatTSYRDjgzf1TwHIHYs/Vhs3n3XRhqxkxGTHoNn6swIgWYUY9KKHgfwvR8x2AKyHz
S/hb7W41qSPvYUonrbko7HIFjGFuq7lr2cyHkUpr1Qqe2R6+HGPbUh7fkYQhpZmCYRBuZ2HWFrmm
cIgCr5bPbaRLLFAJSI0ZvBL8RYfp7nY8BdzRW7bkzaicyGmXUKZynw9hgS/z8ZTD0irrKDL5JSvS
10yPbTuTivt0Upu+Wig0RpdKplwrzBlXGPdq+6O1D54RxFaPExXsImKbTn2yT83hudaCpWNmpR3r
F+bhwcOVcxOUL+wkk4IAChXzWXXsBdfBvaXcD0XdDGSnIg523pKX40eyj3SsysW8K/4QM2NzUx2q
/EK7vDClvYn11xOOgJHkx+hj1sCz8mlucp5IQXZbRVZEruldZYOWajkhBCj2aJ2GCvTaZYpfaMW5
BpRE9a9X9pheCQlZUmCxj+4rAXh/wkw8HPFyT3hrsgJtXWPev59xUXEw9dH3bIiDOItWdkJds4YO
3EoT08rEpadGbBAbGK5Kb8C0yTbAZePTIVNZMCM+HlKjnSoLiebcu2VPYHDRCDqqJ4qvR6yiOyi5
IIkrzhNLDtoJV9U7y9UuftQ3QTDhto/GTMukSZ67+Pu9bj6HSxbQumwjK2CGcrpq2Cc/eNw0J1kn
wPY4gdQZhfie+aTvqfC6dpgNGGcvAe1urjstwpGkIjEbdGDXO/wtAHvpQuwH2rik65J1IqYrVC8H
I8OQJs6MynNbC9Q7PAMxnbwJ7SSfVc/tZUH6evZ4k9uQ4HtsWd83qwqVK+5yl0UAcSFGBfBYFG9J
utoCRGZSwmpFsL0Kiz1Y86fDeYgu+aYVzP8chs2JevAP7GpGILqwlh0fa9ix42Iy86HWHu0ijyxU
ruRjEYc+B7UfiMmNvdJVGtN/wOgHc6nhNRQymifPY2Jay9CtPWRVe7UB88MCzZQGgq3DTCV/f+2W
f6Go7cjW8F1yu8/xDW1esdN6FUCn6+FCvloItoAlkDpfGMr/BhraNFrdB/X8BSfgV8YQpjsaP5nM
FPZTDyf/xnd05g0KmAc8CiEnMO+bxt8BtdHO6yWSpcIJvgcQ0gkCIfinRQx+0wxjEqTAsVR7bKPy
DwnVwoP2S7zQLMCnMCE52iPMGcc7tKqrowAnfMiIsMK8dBWsrvUjsd1BAitocMoXkj70QDXTuokf
XoLcRPTNFrIvIgZgutrpkjDPmduDHLXYSjpRs1ztysHEPp0/bmQKrCkU9ubFcabIagWhaEhz3RSJ
lP1CjhlTsvf32N3AMf36Thoe6vCzefCeg8qlTCuYGiU079hzJHmo/GTCLJt7rM+AvJ8gXeC7Nrts
PN1OVrG3OsBwQLTR+GeBZLpqDZxlCQh7jJM+vw8gMaJw5RF1veeK2O1aNgU4yW3jW7ILPJhXyLVY
3/DGISS8E7J0Zx64FeROFgFQ6fn7pIY4cEVNWqH3azYQcX4fNcqHQo2Pn35Rzbs/qe4gHQLrGSeY
Z5o4637LcqSejmjZzdZxJsOeRxPGiYtT7fZ62QKiL2Ag1pJK6rnxjzpht2wI+AZxDy9MvGk5wqkY
azwTGyQGv9+4J6N0/WU275CG0cwDomLL91LIKvnwS+aIIVb41UWh9lfB8lftMuMSkVeesGjnHz9A
d3+9bOdvLni58tOl6mrufE8SHwrZsNWU+WKSutAsfhRDF04Gl1TufkmLbuqcH+BNFFpmmt2KmZ5u
Dyw9LoDwaCssDvnS2cO1TIkukp3P2UrSeYNQdMv99ORheyiTbTpuwkYkLBtkqwp0GtqI7GQw+t3E
dRCSaNkPR1h0ngY7WlASXjts5r6To7wgUeIVBvbSXOS3GjSVPGO+D2gF0mSg49q+sFyVUBTaAACc
PqaqaMwuxAW37whd9WPt4RpqADf4ZRDTOHzcIFHO+eRAOlKd6Qk0CW4u65yEI2MDiisTYRozjWHh
Lu5akJ0MCjdP3TlWL3i8zEsPlh4Xh9BjLflyD8CEwVhePCU1O5QHDHvImsXBKplBTmhqFJ/vaEOo
LdgBub6m+Nmp8yv/rPuFiDFsdghHIH92/aWHQvgZPMpD2tRGloKtUc8Xw22PHHvaHufUK0GmVylt
+XUO4RLbhWbaAtG1p38mzRFQrMobnNLQPgHugPDQTelYb02Uz0SQRFctz9WcwyGKZ45xLbeYWCPh
XhENVrjzZWBfKk2sUfkUoaC/qm8MZUMqgwejuWLNWW+m/mO79GVVMuMxqwjol4SQZjJLxhjWRcKS
WaJ6eKxTSpmFJBuW0dqdk7+fj8ikI0Fydk+zVuKggPsIJl2buoReEuuDSp/oHegil0HjaNI6cT5V
nolEYvg3yNSbwMb9TZT4gXh1fUCFEtS2miqKOzwE7z5HqUlCFIIA93YYT4LKVqmwmAqb7sP/qH+Q
lfZBs1U5igPlcva/11F2oH4iZDDZ0hycHW2gAVh4Si0x/KLvOf1IWx2nfJ1CAV7bLSvi0ynHL0Zn
L6ltgnNxjnqrLXRRttTkHeJCKBbTxYUlV52ZA8v0Czfijke3/XG5RIGO73YsejQ8IjKs0I+2piwt
VcWnpfblfeeUNd9lrR7JR8xzybcb+0/OffYdJ44WF0O5cald5ap18XaKHrf6WHMxtacRTrKxXPwO
nWgdOUptE7CrhcyvDUCP7EHl4enGrkIrGQ0YgZuyQOu9RI+d/wpZd2PmUr5No1RSA8roATGL5ad7
U5q2BQqZ042qhb0MgT+YON+wxD7HAwL5TdK4ECujpn0kE5+NC8Vsn0t1vCyLptJfvUrvvckWpQ03
SngvDJQiNGl90S139tDM4KvR4Vn+JGwS2VTORM97LgCqoJJyxkB3TEUEgt3QbyBqQDK8DaApzRbs
BwSfYCxWrANsYmS3cwniAz35/YGGTiN/b+CGqiJYo/lwwIEn8MjUhA/4btDGy0hamUR/AQKOa7oW
+IL83Vq77d9t7GcWNniwbYH3WL0pZe9gGBpw6wZvZC3Fifn7NmT82RkIOqKWR2mBNELWjW4AHbDY
EWonJkJYm4rnsYr8FxOH3+OMqNWKk2F5wu42hP/tpkLNgQBa8tmSKTsKPQdJopYekcYd1KaFphsy
8cdNyfVz4ZN5uOfznR6NPzX24nBsGf55DUaGsMwzm5dZ/A1qWw5DmOwFKflDG2rXpJSY3EVf5ReV
vkB59+3RWZPeLLs92xOFkPMGT5z1W9l8AO7H7dKRe9MsiJ5mISM9hNiohx8+A8G+yUczJXh6iJzN
Kwkop3T8teXQVjr5Bw36WRr/c7H4Oje9Yf6GQIdDJSVyqfwPMR08w30SDjXOKj+rDlVJRsqHShO2
xgJ40Sm7S2yAsBAt2lgainInEkZA5uB43cv7+UTB4WRkSFtj2j8PSSFf3KVJo2VC/wSp8uTuk+9R
F9jsf/d3o9IoxdTCvogNQ8rqZ4gvh4ddUKjnDPdb3iVUWe4s8WnWnUKmwh6lN9LfmWaEyWqh92Oi
wI3L+hMe5LVtw1ePUdJgAecP+hAlHf16LyDrpC7aeSjjPd81pYEA3iIUoCiGqnZ2s6AlZQQRkqzu
oxSTbLZwSDtffJdlU2biYyaaO3Ydx5fDsm2OWmDu9qMjShYHPW3858UqwLMXp3eAcPElMUaQhzvd
QrmDpe4LyFp4k4k2VTBnOD0Rkc0Vm7KlkEn9XKuiJ4K+utT1dvp3LeiItqNg1RBg4UfL+V5utDZv
de0ahZx/oZbWi4aqFB0VFzLRc7nWYHIJQMbVmYPw5MuOY8U3Mlmz23wuGsU9zp55ZQ4H0mITepWR
Xdadh3vzEBjLosuTLGkIbhVJ6A9iMYIlfWsm0JlxUyoq+5C7B8Zh6mduIWEjzFbr7y5QBpNDP7Hf
2C7T7dfyf7fr8mVt6XKxjnF0UqxerPECb0J/+4H5m12aqocfCytotcphxYZjCNfiRHVi0C8Twjys
kLWtL7Clps6hlvowSQGkceqNhep5vMFyCL8NfsvjeEaRp2azaK7TeRuqFTpVDlvL7K3JPxbfsWW0
D8gGiK0TLZd1WcLLmFAMYLNS+PJunqzNEUDpY2N6Ok2k0hEcJUcyyAyA301PQ5DQzeoHLX4W36Z9
Pp24zjDZD4+Ba7JP9rA3FTD9AIkobrs4DqqL/eqMyTSvforD7bwAFe3Q8PFalLxmoOoXCDKlqNeN
oLpmsywstZm/GBjeJF52Hxm8gRYIfpxmCPM8FvpVLJvYgKNEKA38k6CBI3F5xbw7f6MwmFz6NiuM
as+Sr4tzId5IkbNPjq8of1+lkqX6xBe254LSMcAvSfAXjO05LVEcOy5RZ+Yob5ZqkUzMT+vusnoW
CB/0DrKh4RPMttmqog98O/HOE6eTFIFrqmPXxlAHqQCwiINnmNOr/egcNdfL5U7nWmY8FV0xo3x3
5znfHtxk89MyNqRQ7X8o+74LK7ntkYrZjbbLh7R8DVQpf6NOTRdkwKcK1byAVzVecbGdc8poMeOy
e3+1erRZOUxIEIQnabeLq1a5+z5yrw8NGlV2snbNJKYSUdPq8t3hJYTJ+sXRYvWB4peRxhDCMJuW
jVj5K5jy94HR1MvOhmBhoyKzJcLOSEOgMsraqFb7cm4QHwbTR1jCuCLSBSejM2xZrkeeTsAeIt9x
GL8G/tqCU7NR+mv0aa20xLgzEd3KWCfU+0t1lGBC5h/tcEL9vtZULnlxYu7/80mK58JnShjTfaQ5
2YG7dOBvn2F9VvLEffjaKgNYsqQM5oXJt1BD2nHXIK8gsF+AiX3f694TjaOswT8Y6ghW1QMPHPX8
GVhtHZG4EPPZ32APMX5zbGAxD4i9FABcQd0rNscnBguVEB7LLxfrpxTR0SBsO1Nn0U5ce2P0ybkx
tPiNA7vVCMeZZ03AkZM+1JYwnnc3Xjf5ndyvQDF6QRvWz86mDGpxjdWQbGD2PKlSMKmQoLO0Nr8O
4L1OnaOPcyOlZEX0x6zKBhNrPjRW55t0rqdjIa7U2ATotzaOwJ9Zi07C4bN+1wbOOzqwg+0lqWYP
8diE4wPqwzGcgGZyhBL82NhZCQtU2pYGwvVL/n+aUomuc+Ht3L4g9XXs5YZvCHLvszVcclelxHh9
Deqb5FOyDh6Rtv5cL3zP/zzW2KGH8o4Y6A6fgvV8pvIf2rzpaFbuiSf9tjPqcuWxITyZJZTWQfiZ
rF4bm+J0c/CVJEmpEDvDXts8iTLoNWswxr4bE7mayhlcNcIx/xhatk97sLmfsrne8bW7Uv4JPWq2
i8wB3QpxsQN6v0tz6Y90z0YujLiosfE/Qi9swlqZQfa3rXlGkLHOVkZJcGLMOtqq0Ltp8rWIQR+p
t8/PsOSwcOzqVc4jpxf3QiXUug6xnP5SgHZErsYNqUz3K/vD2Kn87wqmFtjr4gOEWQLhbrOWd5fz
09tsCsNjXXKfvCV5BrYD/a5Ccb5uIqtvGZdUibpCnPKiwrkOFA==
%%% protect end_protected
