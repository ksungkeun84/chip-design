%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
oybZI7BGNUcb909lMvjrvyjfHciXMCLvhfWZfkL7E4wvECx/7hrrEEFvdVkjnDQNDh45VIR0qFHI
nUHz1+346VnrbtOkas6vWhSLNL2TIdFvgIGv2RdnOgvwDJJ0S3J5Q3kxTTwPO8hl/xr6EnXvGsIr
5XbHJqIgLP1Omq6az5vv504eGXv2DZScbFfQqJbOjU77g3M7L1WagWJr7ZlZgWNeTgE70RAK7NAO
gmM7P/d+A8INuBF2qwkHS6CZag9i2yI1I2xXkWzSZ3cDxSWwfvJLfDvRIMEjSpIHm4cUaf44L90y
FTd+hxedThp6xz3cOtXv3w7vxPz5ufNubyxVaA==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
6t/6Q3j9bRNr8N0pg9Xvf9SNYQymizo8tHyskvQQaM6uj18umhB5cpmElJSDS3HbZG8uDE9qhWe+
4m9XPIiMNApPbZuMoHY8hWIbwJfqn/ApabhnHx8M+Z4OcDJOfnawTfGycjCh1+UgiF5wWIIe71AX
tfTg9qEU+EtsrDbXy1k0rTJnAAG2gJc/HZuhGqg5diuGzxZwj3vtdNptPRc1AvpXlFMi8YJSXd3x
fJ1ZKUrXXDUca/opd/DUHmNI5xr5bEIChgulliMJWGCM9mRNHw8562SOfTIepF0/MtGrbevx/1xT
UZ4NKnqC2rO54TBd5yvTaXL0iXcb7s8IdHsZBjfo+Ra2MX4alxviG6ZkzMPi3O1Et8SPjyyoRKlg
lN2E8pI+ssl7H8s30jdmjUkgnJiaCq+S1PqvcFX+M7NGmBlwT/ajMuYsfqQ9RMVZsi4FWbm3h9Oq
3QwTnvMCpCgfOsC4btKOvmL9nHd+TZZdzUFWjuIv0k0NzaamrSNmeFLzZG/Plj+bV4WUkxVgz8cr
zOz8KXk/2Xk6YFtDj9yvH9IaH7pw9LrEGod1slPE6UjknS4HeK3SXVi+Q3k6zGdx6bPBY6zMBacq
A8yKpEP2c2w+iivY1/HwPfqkyIwVxlctdxQSjx8UySTAvPF6C8woRK8EdIxXUWINlR0w1XwNg9ZD
oVP9O6/HDx3GN9Rs/9iinySXUpEuJ+ejCQPng4+LBPeNO6p7VYTPlIhU1u5IKKxM3QaQZsjkmc+6
U8SRs+6TQoaP2KRWR3fxiaBDgn9faK1OIWmkNoVZGiOPSG2Si5JcOU57DVEz/vZvW/VM4XNVioXx
Cj3XJCTffRrFoUjL9t/+9TkoU8xC02QQ6GZ/o23GYJblicKiSOirqewT5QAB1cvSWGjI/h1iPGxp
ofRMY9HW5nmTyRewFfet0HPpzN5UaMcHBSYp5yVX8+ozRI6rXn4RpyMEuI7PJDSSB7wekYm517go
2rj845Qs9fnxjOmnuxWkbjTIK0pLlEGsROpuVwtWdfAZSeIoSkOHKHKHk8VJnqR8EtNFA5zrmOTQ
XxFmGqAcPadWixLHmjJ4ojflLB6Dgvfy7DP4kLHpscHe49du2vsspn2PdO91S495i05cf/f1h2Vs
tyR1ytmXx4l+Tc9T9wPmD9S+soDvbWVD7MQEGX1cAAh/av82pYXFEIfLYSstepIHTQ3co4fW78kx
g+7VuXvgYntqFHqXwVsTEnu2JsXf0VmTeKQIokY9n/4eUvRoBYtXZNS15Kk/LHUrQYJFbv4a8ZfW
anjKo5OgdEqw+6i9IdKQeBdHJZxAAfp/yjNN+Z26BOLtRiOmJzqfdiO/v8CVpnOtmklyQWyIIGwJ
UVgc5m/EcpFVBvzavgnjBfdvC76Hk26g/ei/ochp82ktFpUlxnMJ51LdsKh8a2c/Rdb01O2Phnkb
685CwSHZZyldFDn+gdlkrYQtkhWqI/fxwzfUk93pjRvRKj9h0h9e0gD4FgjrOdKk0CHinwklNYcV
gSR8ArkkBjIQEAHNvGib60ohD49gdmLoHrChN6wYdetNy/fB12cqxh1Dtb+IHq5GRoKMkcLld76t
H8UrOtQ5Z5Q0VUUAxlp3Jottw75ciItNc+axN17AeO6mDi0E/n4uKNVHpgzJAsTg21rZB9wj5W1o
uYbmmFignq5QqvZlqZXX5OY0NC9uNHezZ8/tDFwsryo88modLZkYCmlVLtP2EqAVF2GfIVp+g/DS
yOyHcbjECiVbvjeWBvi2jf1ocJLIm8sGXf+sYG5314sw85QIrzUnf2geBY5vggry39Mv4ENNS09P
Pczhkh8/UsbDtJfWqwWLlvbxlI9G4dFW6zI8XL+kPYVd1UcDd0OE0EJx3ecjjmAFmtysStF9CBfh
fpM0b34I8dUvGUd6JqoJ6C5hPuWCvfOI5I9m2NPgY5HQOmqDhnA1zr2zJ+Bo7XNussIRU3TLPDUI
ZzJkMkoi6dR3N6+ULF9dApGJWtNi73Mtai2RFJJMIzn6hRfn2l3moWs5PPs0/jWs5ppe9dK/qODV
QJXj03pnqb5CH4mTsdoLJY10ytrS/RR9mXWJQ+bPkn5PGbuCBItGIpLNCm9MS7/NjoJ7C/kI6Js1
OksfVp/JgckYi1W3QCU833gUiGRNxVzc6rbtkATL/e6eQyqC85bWDD9J4MiVeQhkSrCiOg8OzugK
3QflsOjzG6D/7YcdRAMO9FyPFoU8+5qLIuDkDSSPOzG6VKNCP3lbd1vI+WacykpRtd6/outqRGfx
pBl0v819SoJOCeCIwgruvA44u5AdvsC7ZI2gz74GA0S71H48WFGlPAGHrM2ecogGl3VpehMpYJMw
dG+AtI4uXWkYSauzPuQW4H+LWvymONagW9OySv4fTgmU+QGOAhvmtMYoHVYMBU7T2apP1YN6piWk
83MhBr2d6PiiKSheFAYgmGuNsxoAJ75sSUxYNX3ReWQ1/2Eaz4ypAjkDmPU6h+VfnmcBRVY9vaLa
XD6E1bU9G49Av9oEUd733g0GjqTTL/CHW4BNYDCdenvOp4skZkSDP98LB2yZZhVifiRuOGKKmDHr
zz4yHeB/gksl4slmGJ+F+AsH6TSxonp5WXjWoFEiAk21IeyQXej0b/yURHlJRaQrNT5qgfQNW8AC
2n60DYpXjxC+gM8ywXuuLACAHswfZ4v2gsYaTRn5q1PNbkbJLnBV+KW4qkonmq3RYq4PAgzhXKDg
Jgf6O6gcbO4iF3urzT4usMmnb5z7jsoZ4f5o02oKBC0pSMqCGinQon4YpVumHbpePRqhjDcS9rNJ
Hgs/NpLGn9PK1P5M5b2CyUrhoGoVBb0vy9WIC8chUlrbGlwXf3ydUxgtimCbNdO6S/KBA5O2vQTV
um9YdDCcGYiOkA8ior+/r8pW/R2zXzuS2TSAOSHbZkpZaxTo3gG/Q0rJol7rFmS/n2JQRP1wKNqN
CZSsfdfveRZ26oSEoxoO/mfNxDA4P7v5bkYm+c2WFScqIeNU1aB6adDihBYJiFQ97tKkgZDqMekP
8aiSDBAtXpWQH0gcpTlGsEf4W3PPwATL5YqXT3Q1t6qbffowS+5Q5veYkawVh61hRp4hfyAjUOkm
itkz/TfhoM6aZViv0Jz3d//WfwL7OGY/Yj7driWPsoDchOL4dsIhFE1cGtITq1exWb16cwntTk4a
xHDxYGXg35n2KcJ5b0AIh0njGuzEyURnFOy+Pd0LMOU4KCUl4wnOaQ3vIBSHjSTn8hTQWhezEkV/
Onq4cI9/GH7se9S/P3jE1W5n6DxHTbMpRlt+9RfmvCaYq1YRIseyL9ejL6QsMpC3ovfCWbSqwafv
M75iJznXVh8K/qdGtSjm7qU5IXBeZHyv/bEu6oFuOJXSFdbr4l1+F8DwM/P3X/LSLOktOB7tC699
fpOFktlKw/Bq906wtbaH48Qng8ztpeyMsR/UCzSCT6q/PX2lb+Z2zuh8Im05/URAZyS6pYC2t5TJ
mPyHBnnhODZ8Kl1T4TslT68H702XrIqtnReRuYP1YCbAf8PJYutYbxgmulp3LZp3+6xEK0YdZhkE
N+gRgXvKxphqEnR0IiZGQFG2GLcFDrqAaUhmZrLb4c4Xrndt5rhf5/4yMSvJJTFaKMK5TPnJCVT+
pEEjONDc/vNnizJjqW6w4+EqvES7ugy1IhIFm3bs+lNW/ummc+S0I0r7YJoWh6r+VWhWJYAsI/KE
I/ZREfmKGGwzY8JBK76DcXGC4z4J/OYCUVofbPzkjKoKWCvadtEwM9flsELm+Azpsdux8iAio+rF
NBbE7GAonzi50k6oBvBakvj/j/83wS/4klWroO9LcxlSL0fuGk+DOToUDGd7WYIOy5T0cEasrNUa
F0CGRno63zHikyYEnmNZuYupPJVIZshPwVLbgVJGneISB+Qx+DVh2KS5SgmrGNuFzXU1F0H6wRiE
7xDHS7ZcBKJZAh7ZfyFhEr+lkp+vO4LNbOZ7IELr985M/LxCTvJzZoFjpZwD4l9DHZ8VuU8Qtdc+
LLVM86jMIxWkA2LO4UKOeXfi8FMR+KTn55NLwMRZ+IeZzsGYIwPn+suJiHif+uRFu+cu0myWkWBH
VHJW3pvUrJ8yX10qJwDF+mPauRW8/ORl/Vq5jWDIlTBf9zhDoZ6sOKJnmEzDt63EfDH0YdmO+A6b
fPkf145WodjnvhvWc0EDTd22c7s7xgHI059I+aC8EBAilvls9c9vIb0dg4DI4I2129sYoGO7eCWO
FfuCLdebRsMFWgYlsaMgwte+IS6h9PfEmlm2rC9E4A9Fx269tuT68Y9937egEfd2dxc3yW2QwNVU
A1MZPppLRAOwjE/sTg8jz0P4VeYUtGMU07A6K2tRKot2W4FxcKKA4N9wPRfMB6J5C2oHqVSnINYn
C4gAOdmsKnRqs0HeUIhTBYNwp9CLfIZ3dQgrkilUeIxJHcxIP/oLHy1STjUDiXo3/8wOXrgkckcq
dyiuAgDf4dSmIRcRnB3p01+2yMRSJrlJUrFSCTiQTM8apzIaTVGqcUNXCyHtW36gxae023Lq1IY4
2A998/0IrduUwpP9uNP7nLqijnQ/sEgBcenG4SgVRlYs1ebT9ScKqIAkd3vcYb7oH9HWC3in4MVX
I8I/Gw+uSobCIbA3puoBQebXSdJCQ8jEFO8iN1GKpxAKe/a/Qi9+p+g+2hOu4qHKBtZ8hLl0n+Hd
eHR5GhZAk+MqJJa7dN01TCiArpegI0ugEzVjkZ5z8U2b/S0CEHuFiOSCcp3yFwjpQrF7Wpm5cqXB
E2Czf6tuLA8Q/3a2bsmnYn60v2JOZLylo2hUVeGMvpZTvugv7qvMocrOP087nuzbTxiLiZKAqeF/
LLUglUNZqdVH/fIGTa9B4NywG/HR09btNU0gpZlM0zP6MjJnNADzyu7+dPNC+mhyPom1zwcQvirS
0ODlawA/ha44FXAxEWTHUOFDH6To+Hyax6iglzR+by5DJxogG4hstm329eUWK2TXN32dsX4WGNQi
+vg4dQ+vXi7Ju10oDceo01p1G0alAxhYO7Z+K5qOJPDGxT8+0QzThpv2S+PkpvCgDTLe4/sGHek7
Uc2FXjCylnCLDyO3K/nsJDyaVQ4p/OQ6+lDT9uENyHoyPIAhT7+UndD5YdQwUWV0PLleBjR7/zAm
JD64drjskmGnNg+malb6COT30SYdlAUX/KUy5vcIjCYwEM8KuBUHGLMZpEoxPmSTPZJH0SmqvLQ2
27XcieippWbFKwlx1h/T7DMS/s8BkE5kjGRnAhdFIVzzemGr0WSpre86Jdci0Cj562N/30hCAEl2
agMFPR8rnhtEWhGHPVKk+w9VpOBxXDeyIVuhJgilon3M71QVTOMVmVlr1fb3GuUE9pb3EbpoT8kR
JFUTL7QSpUhO9OCaTHrR9IML3utztl5HnOCpdcDGGQcag7mwCVJG1TeOdUuY495lbyqzFRZda2sz
zD89zoNMlSgcjZT12YknDp2rY5RML+BFigkHZydNel3caji4FqlItCXqotdASBUg6cL6Nmm9o8cH
PK9j4NiuTyEifpiw405Q5g4YAsMwp0yWQpITl5KeXU+U6OzXGvJiwdIYH2xiQH0JDd5EpeUptUqt
V/ySW6dbMtA0DY7r7vHBO8DEaWRwaRW+vfQO+uDtOwUd0ndex+299UFdtDTDozR6v4KURdc+FDVE
pfi0WV29LJOwJUaxw908hL0hhRqPlaKAt/6B85atLqSyFSF+b3s+JMY5uhFj2W9fu/Jv7I3CLnu0
oDw//xraw7nrcZwz08OtwwS2rYvITeYRPJa2ncQsxYktOug34HO8FnmQyr31GSepr01tWBQBDskG
6wuOH92aq16k9FZJGRqPP2YWMbJ1EgB9QgG27m5BpK0lW9OQOYphGOnRLJz3ff/MFJTuHFEXwJ+t
QLj7eOgsehKJTpoQwGgkzTn7/4WGcxTrUBOXBFrdGdIqLQPplQhnd4Gmnsm7VAUyd+EELmq0ycSJ
l1y3JNcagCqPuWCK+KB0uhKC9mfv+eBleNTLyfiFyMQW9hoEbS1wItloOHBlBGLdmopPxNEjIZtT
LipxrXY5ufNBZPurmOrAGacp5t1zrR+cu64TnddtvS3oz7QHXigcj0cZ8dnoHoTjF1f/FDwycPmj
KJQN00gqfEbao3SOGND1tTZkrYvX0KTB9RQl/gh1JgXVnkpAGLUvMof9VVcmH8UuNH6gWUjG/xqO
/Gqz1L6o9L6Z4t7QOiCMHOhpR08Im4forBoJRxiIEk09o7itMsrRc3RJlM80AJHcVnAnPuc+wacp
D0rwxvNHXaTjXIKr3RQG7QWQWFtAMVKSoujE8oydPRR8bWwZcIzUhaX7ijZTmEX7t/C2/XvyxY4b
wSmqSVx1axG6l/6zyXc+paa6GLhj0liZkiYyn4jPwHxX+5z9bcp0O8ObQBUnmntFqviRkMKfxdcd
pmbeDlALaLikZcIMDZyNt6TFeC3pPt+l4QfZTe5/ij2xbA57FEKZojVqEN8xbu7ei+5sb05IELBV
+AdpnG9kyxR1iioCsIePW3NmlWD8KesdA2FYlegdWSL1Ay0O8/VtnoMYYDF5sd3dwu/9LSRxPp14
rKPXruHD8+yUu4ujjO/VIOC9OqrPNglZMw3ZJEcxVXe/E6vuGxgNqSn2vHi5x1L995sf3ZVH6oVg
H0liOwU0VaUvSQ3yXERSicUEs5RXOdGvtxMOIqcvGYJp95SekA1W+QgxNmyWPDMmOPfH9Zs40iAk
CIyNLzWaTjI7fYzuVRaZ6p2mWtL+Q/ajEvg79YTDHbUtKtcPIJDmB/OqyTEYts1ScdzygopVenDj
lJBdcseNSD9+pU0s7DRja68CregGDMBFh9F0bpYloqYRpba2nbbFhxo0MzyaN1AeLavmjnrE2FSZ
WXlyOzpw+p5O5h9XPAL1TTmlJGVa0oITwVdIFIiyiE/AN+qha7cEj+omc6kACXPqJD9t8Omc5CJ3
1UnNxABOag+DI+u9Bw096Ai3t2jlokohWVvXbkB8I9FFXhi6U4ijCQXM+R2p64bCXnN+cipqHQiV
qVmOn87W5V1qfn5QF7WGnHgIX02eW+v2oQJPw+wUGPX/k4o6mZa3Vd644VHxaT3H5Kiy2uke0eRX
iYd7ayyDPJ6TRG8SxkBkz1nhpSMwL+oF/zej6DgyOe/7Z1Ka8xzGAduE8O1AzvVK4ioW90vr0ewj
sU2ASUPrKHQgbve4uAgWGPez0r6l6KKKATpgfFEa1ib8vpEDrOEm4OucCspBEOgKnDOStuEXvN61
RRHF9U9pXKN5oO3c3ZhkZjC8jVgAQeBa5mo4urheKbx7yvZb+TyCNTtMgxERvcrjn/1/Wvh0rLnT
iwpxXQbHlfx9d4gV3bZRcvPszrXrmm85PAsjAF3hooPmPL1X86j34EDuXNgZ2jGuxiHpL4/3Xdex
7DXVqZ5DocuG+Ulp2/aTcD/oajY47RR5Msrhcaw0z8ryJpgux6j1llT5DC7v69RuLZadKE35kYnt
SC5pSuTptn02Mp2FPpnOow7aa1F7s2NVtBheF105jSR1st4awiBtjAG7ETQhebqJwhFK5ZwdkNeS
/xz7G8MEx//WXbJj2+BY2wqLaNRw3VvIp69VrQuIh2jo3Ot0vtulH7stJoJAwZPGTxEKExdTsPqK
kdK4QNqkHF3xFJSujlUiwUgI9QMR3NM8G8u+yq7LOyqEkt+EkiF/XGgMJWrvgZsSxIf+E5azsTe9
3oLvXggzQlcKo2iGZRMYf/uqAUv+ccBTF/A5hqNcNA9Atw2K1nDXvR4Nl2JpWyMN38aRkCwIEY1D
AqvOt4BctmqZLwQ7leALaCUwZvxqEcG9HYdtRVdJmVFl832XqZZzZgDyVO9Wk9qrOMs04sRe2IRl
aV4WsaaLnkJpMq80Q2waPgPRfPbBajli6XYHsnXCwOzIMW4ANsraRSmuvvafBlDn3Sjfj72iys6T
YglrWZiXzurmYQc6m2dmphl5pEbLI4/tIU1v/1JykKA2pmfOImUXSfrN9/4JJMXU7eV+Mw59I33/
lW4dpqhzzxiQNdN8erSzAu+ydaVWtiJtTYN+KpVRGdHMZwZH/jfuv2bS6LJ+wsjZDyJANZ4ae0fk
QMKT234ZRyZlJavkYNgD64f5diLlhew6MDMHswOdjpKOMpxKTIj9S+TmMqrIzL8t/0UtEXFauopK
Lz6JB80P8/dKqY9wktoHDkTGoih/Q2DpUOV2a7x6qGhRAUD7tGmti1cdY3Uufa9KZ0SH1kVJAU1e
MUKyaxWgX+tKMRKTinXrUxK5DEBs26gkuk9FzijxsUF7+RLkQPfdYrh8LPqoJy5wIOu5aoKhHwbN
3OphVjQ2jwCsctrd7XHPtpCupfci7DRrONQHZTbK5gXkME0gRTbRrvwRpvZRcQ6LfMPRWO6e2l9i
0VCiZWc82tj6VXUk0x5qWWNKfe1R/KLQuLUD8PZX/I/4MqwLZ7pANh6KrEZC2xly9ykkGnsYbED1
7e6CCVKE+qWGkPy750EatbZJ9iBG3pfVDGGDWv7wwqLq98TSHSKXuHVOD/34PHbAq83FqkmQAat9
V6ubejRtz3QVhZtcp3ysXrcNlZbvHh6S7zPN2ldYimTbPzN3SB5ubAABABCypYRRzaqdKUx30f0m
czfEkukLhHnHsrN0zA04ULL7K2DjRDrLXIP8kSO9dUvh4en3X06YHKk777/lEdp3PtutaNgyM2te
upJJgQsBAGLYlNnkWiccfq9zyrouNZG70vpeBOpVTqa+HBywjct3z2BStJ50fzeGbe4eynbuG7Yu
YE4VqUXHf6QP2oWVNkSPoC/rWh3ZzNiq570UEUXl+1fRJIJQQAFW7xgROppP6YJ+M+HX7cw82CdM
A+wo2BO+ZQIL7mQ7Tiv4O8MDjRg3H2VB0ZY8wGvUZkYm87iZiH5syonb88Oy9ZFkkOyyiIvogQ1L
JsrAs/GwQokt+wipwtHWPp7+YU86CxBYA4u6ajN76gITWI9CmvJ3pWe9h5YWNEisTutwUQAr4ek4
JlsHYDG56pytAxbOCj5GTrJl3Snf1RYR+6pJFYheioCcB+iWp2bhM0UZD0HEHSL54qe/o8DD0BeE
kG0IVpBRtN3V3ptr58sMNYzM9mUNY3b1a6Imf2jSK3/sKQDxs6rrBnnWFnEDEUBcCefXQEMsBp0c
ZUK7QUayMfs9VGRj4hwFsWnhqysbxnU4hlUBrhusVaPmsh0Aoh/Y7FRFaGLJ81D7HL8uhD7FyJ5r
DdKKmqsbx1uJOTYWNmaqCvEdS41VELJK2KOZ+ijZ6grHaeOAr6okH3Edo3vUMINPqsHzXtKYIG6d
kEHtMVgN8XR5GdCIn7z7Yi6ayxqGJ6szmfEeUJLeTUfq02jh+3/5XgTR/YY9UZsuG57b7HRPfD0/
GKwby763t7BlwEkb/kQ2umt++wKzHiEJz6gSknebuFKYs65x66Eh6HzyHrfQS1PqZP01eHUrDnf4
YLBZG6fo1OlReL2yvUNfw+MKGLAFlyxRFi0hSB7LKbCMIPQJYVAFxHBrCtEpAqCxpH4MEZuZWmpP
Sqi3gQj102gmt/qREBNGQ6DWT3V8ipH1oP5Nz15AIAifMctojfzELAtsHiN05BYgqARVceS1MvdM
r0lOzR27bniRqPU0xe3Jm+xUqwoyoc0SFvm/UFBiZHL5Wf9eVKA+gWEOm6f5rAtRiVYiJs6/JG+k
JqA1Pbkoffj8rvuwasHKtUuUDbp2Qlv4A+geWvxmv3SQ+jd+Fr9iYqnq4IXJNoM+k+Ye7tGk1QgY
cCK/4huUtACyTRqa70rhsca1csPTIVpNcMAfppU490PZEBlAM2WS8+139GW0hNr1NQOhh/60dTDj
x0znzDkJbGshwHjJAYPm5EbezcpRCtKnL+2OqDYebGRdehQlNkemQjtyu2bZ2LpDYo1Ail8Lp0am
SxNl4EjXq1oh57QWDLKjYJRyUSLdCrFfT3RS0L1V1HTIqyM0Rpb0l2lITYZT0yVsgJw9PZp1NOoh
m1/FyrKxtbSdCRBiMLds4Vh6y77TiP1txbEPFOxMkHwrnRMLaRYqnCKaPUXApyu9ogVUNEaVmZms
0hRbLw6X2qdglJwT08pvf6l1ySHSzv/pcBRuX3ikX8NxEjkGXlhY2i5Znpb97f5Wz2xPxBQqppTA
aDtWyP7zmR7K+Dqi9jgVJmDNa8GGrNdo8Ly6CHKkr021/w+S5Q6a5gwgp7jm7qDxxpcpMznZPdtx
4kML8eSecyd+wbOVtvfaCNn8drssysYNKUMbeZ2giqw5hcMKXlLeejhTPyAqipbYaikhxo46QWkG
dIcl+v0HSn90eBPNX5rsA+56OgF6J14ohtcZ+1/icEQN5if+jyT4XQ5n5Glyyk7HYGp257zrnzAm
Q12fxG7UHVsrBnKdWIUaathyAJdBn5EBEromn/nBHBvxeRdw4M3+ReqXXyXAQRxAp+Zo6bcJ+rr4
bHbfQnUwd0I+KPQzWERN6EUxc3pYx5j2cjNezrpBgl1UkbP0BQX05FLqpR2XmgrGUx0wCOvKTj1R
F0ZnObChP+DJ8F7mlOSR+IaWvcNtXeJrV5xDA3VWsI/1CMRi/+Hsn+eEfuVZBGAGeO1sBfSrcmpA
YA9V6BRTN0cAHPW6X6dpk2OKV6wmE4QZw+RBO5rgnbidsuBWk4rZODmwzGJDnsR7gF2z+7JEk45r
mVpP8wJunuaPbXVX6kwR3o8FtodEbVds9SCxT5o4ze9HDylRwDPin4BM+hOHygv4IFi0eji3U8mk
itZGVCBQTWp8XfcnUiFvpBa+Seqd7GYgnbajCapaCZLVms1u19bCaZNKocZLtsS5Lx1Yi3nIOktG
GF1F3PoUwX4z3gavFlC6UMfHVMD+cxbdaj7ta645SahPR4GLK9dnCAoNvxa+Ci5NBUYS1tZ7bEDP
ZRIpqOWGdm2CrDMLb+jl72TBnzbCrN9vh4i9xflRkujDtctMCt4Z+hW5vfTt/euTXHdrnRK3uzxU
xM4GF1DPgEKl0dxvz60MhRpKc5ZxjRgm9Nc9vvItWPKVdBKxS8SH8hQOLpg18TmWzW0lOLOj3ch5
bgXjwVDeV87wg46Ue7omX9DGe0m4HdXC0xsagM6dfasG6X/Cg/jtLeA05gqdECdteV4UrqoWPgsx
57q2EdZL4fegJLaNZZISu4PuudYSTlYSOXHYbj8982r9cYq6U1AEy6uVUfAvzA/N0gEdAXENZ9Ux
7uMwzhLtjvybRCnLg/eY8MURJY4OSRIKKgibuwDEuNPFRyELVm3xTIWcZCFLnWzA690CRH1O+P1f
R7niVL2xERE74eE6niNCntbKA86GtZu7mLcB9jVvnoEiG4mJ+PVlXEEQ8rgfo7KDrquuWN0X7ard
2IGCqiMRW+pF/UMT+cbRtw0uxj2gNQih5p25hnGWJeYCyVlTyjBwaWHLVnWSpv75e1rq27Kb+7KZ
ewRT3UXRm/OnKfDI4GVFHcyJliEb+uqp/Sk/uRhL9Bna/FTZS92+/hsD/xUaEgPknikV4tXZBvsG
xXUiJQYGppxupQHWngBWspo/sLkzumIsudwzuS+aJUmX4SPfNfNcKm2lkSzc8p1gfWO27gPTGZFM
K0qND05iSAUu66eoIScLcAKbqo7y69Mn/qMMZvP230iWdWj5C90bOaOuC8QqFQ67TzWJz66Djo7S
a1qbcljSov84JVc0UripPBCZfPpR21mZPgG7Lxbe8uPsroOMR7d+bcgEUfE97VlnCrhyfV/Cu4Nb
sZeI97hfivUHBVk4oB+bDdou1um1C84H0Nc69M6f6sGOn7DLpUHf+jRAtTvXOx/bsfJudIAWuCBM
9Tdyb+wfM58s5WFRGJ2H00n249EvIBaOR/ooRGV0qE8DQcu1qYgj+M6M43VzifssnPyhcPuRor5J
Giy2NMqVyn2x4zZLx6ZeQBWla+qIpTQLsS7+vCFUM4rExNLDQxCCpr68JJhDBAbL8Pb81TWfUQYY
010BUoXd8O66/W5iReEFInfNK4w90ZOHzr2JxXg1N6gfp6ALrGMHu1fMh0/Ez7eYRtPqtM3tMfyn
3xNKzkU2iuJsfzluWgGtivQEMqdb71G/S4hDkjoQntvS1TvApg0B5ngqT/YJw3Vxw3IlsX/fe6WP
bn5qBBl+ERiQwOgsJz0iykir7uamJRpXNtoEjR8DSVY3tWU9lLrMyXlX7ZaA562KWDZZ/ivTuUR8
jCHEzgMu/yJrUhnUo4NilK9Av9naOE8FOOUMECf22n/2AGHDEIUDLIrucyUxuFoIDz8TsjnJr9Q0
4LIzDq5TGYL0jUfnczkSMCRDpe+9xtt1aAxbZ0vKgRYx8xHY5x++U2RghxNTZ4ezgTM4QHd515B/
+KRU56MEgdy1ywMjNa1PnEwuK6iH056YAPHMR2Jo2wrsc0QY1LUWt/QDN1edRI3iA/mwL8gX8zBB
6bIKl1Lzog7KhkSov+zJz0mgimqv6Wxbmp0XMVDsz1hI7leZ/EYaB9dLEQdlTsdNPwgyl7CnGRRd
pWONOSYVM6FZ2P+B3TsBDZDFdnnU5VO9UyF6oAwF8aTTvQIq/iTIE/C7yhavG9AkNxpW9l7TyXYy
GOM8P6mUYV6LzljBEw+d+AM3T3osu7viwpjlShEOIzwSAaVEkw3MU6ecK7L6lEKXuMOsIcMdqtSH
lagLVJRpF+2BCX1SWslakoSpQpIYz/MvrhgV/eITV0xUtSs6w5cZgtcbltOvdt9FmBDZOdWMwiTC
A8aInXD/Sz6DIXv/WQyESRKmLa0SiDptgMEUi0O9U0/dWJjnVqk19/5/bgIwJM3VVSEmWlwKPlT4
+AadjZvtU7pLvzY+lCfK8x2/NMRUcX3PspNCUF6TyeP2k/J3Ax6Adi3H0Vn4zheLIbASQF35tONK
HwIRQ+9CgorpXAHSgfSX7TESCK5aZPnEpf/mlT74Ejm6Kd1h0+y6NUVzIHGW8coQ99vNQ0Onhmi2
+C0fkcSRRmXcB4pxW8lsWejeIFbbSb7MflSyjnHFXTfyx2k30FS7YAYEK/Yisi0y1xFUwTAkhgS3
GTr/4PVJ9l5pyaNG4j+vITCUyvuBpGEUMqtCXPcT18IxuHQ/SUAFKmbGpGQTTk8bfj+SvqFSJ7i2
VWTW8E9vJzSxEarEQ6M7oa30ns94M0CK+UKFAvzj7LmbbCQgb3lTnmMlAVtHTawhZwNhKmMgPutq
MqR5sTYEJKTizyfTn5J54y3s9EPMWmS6UNhtK4okOo8cYLisNlqeaWsabAJtie9AbZ6yBYjQFdnR
O3RwjVUK5QqDGGum281pXR3s/WBWaHcOQMgHlvPzJxGXmkWfejVmlNV0Z+oDF0FvfJS/HFdXYSMC
vd1qdTSrK85Viv3gXi27Ekaw2YrW317KW3jqzjKEXprFniDbtT2l3mvaYPkf3ru/Tb2BuMVBn1Kw
W7JTNxWZ1CI6thZYXr01/R9b05dYBhH/K7qBELNdaCvT1Kb6ZSTC3Li2qJpZemKx1kd2uzGp0iRT
eEQ8XE0pAw8YNx+JOGFCGrDYax7wrHnPG7hIbSj+fA8imLe7uXAL7Fjh67yHq9frgSqbHvLfjB6w
IaeJn5sEFGITaXbvBh/wFfJ9FZmu/12Aii4p/vT1qdxBZ+SaQXrUXDVHbcughkjWBgW/punXUnj9
+0LysXe6A1ocoI+UjXT7lsIJMBfFUjkZ5sGwh8nOzk49WUu3OCgh+zzyVIcKCHjz0VFZkLDEoPU2
T5uAg3B3nl2FAAdJ/vNIMQ+ZDdoJRIoWpQlyT8nm1/QcUwsAJCfXTnbi6DTSbSgJqLX8m/4INgdk
FOGM5xXgWbN/dNqnIHVQrrmlSalIG+Sdp9k738VCjRoqPx8roxks4Z0r5124OYWvt8YLC54Yh44s
Jugh5xCa5hUYu5tJ2x1O/3eh05Hq2VRXzK2jTVrVq7LhZuc7VEb6TwF7NSpqAbFlggfUAKVRJHlh
poXu+8BaU9feJeJyQaHevnmLlD7zUcy/Oz4gx3CLrSAQioPr3sygMJOEON9pWX/o3zJt6alyK/Tr
DycrfUGzz8d5qjy1ffgkphQHw3X3YDcX1XbPHmSeqg6MJe5VzfbxxuttgZwW6PHnfjkRjEAcwcel
L4RMnUl5tCYIF1lMa+9fbI4vXXihd1NgO4kk7ftuhJfCfeeq76Fu5IgBYq2Y3rlEmwg4B3XV8Yrz
2Q4/SvtMBgx13MURwAjNQQStHtuUGCOsAg/4BKSycYNG+Nnl/XOK8E9CGom/gK3btw0S5AWIUIwD
4oHSBi7bt1BtNPjfIb7wNAm30YKR/yip1fREhgL4GiChFHtZVdssvjasNOQdGMFoFWd2F9Bws3fS
oyAZXz2LWidMMLGy45UyS1IPo5vGVLiD70G9PUWZig1r7NM4wK5QV3L1+QNfOU8pivrSnKoESMLw
gqEYa5zeaMCDax5/t7qw/KsikpqUHCQD8P1HdewEWOPRxEbMfmJmXPZHmJMk6IwMNrABc3PnN9FE
BtyoHIBCFo4aA4gwX6H1UqmUp4KW94hL+pdb3mOP5jK3gaaz1PFdxLFBYy4U9NfGzPm3AqoY3niW
PGLptlst4tP9/5wdI1sPGAwh24gJBe8+RRAKaZOg+jfV4j1/X0DN92TCbcSnwxtSMga4OWlVQAyS
hMDxpkL3MZyiulSh6w/s54GjPRlRjBj/YpqhQVCSnwYp576RiYx7/ZURfynxot16u3btK54+Ity4
0pXoaN6jdFBP1suuLbyi6SHtYsCZo+xBG0ynyFdEAJfReWR3TIWuj5c397YX2v7dqzmCuVJp7EMN
gVuLWECL8NmFHA7J4OvTBZVpXXaOHxRpw0sXYj4EHYCGOk2QT91RHlJuW6sxQV885rqVCFwjmkjl
n56QO9giZkVJBug4hQvCDGma189zpucmgH9Q6+JG4s6vxTMHiqomxXjKGAbArM3bvnVm82flpu5D
sF4NULc4J9aE07y0ylzXwuD8QDNFefjt4B+VXPJE4eAMtdLZgM699tkVOVj/jkIsaHl+uvFGNIWf
uukzy660W1x7CU911sQkycweB7wMR3bC678/D6beR5OCHGKJPoVn3aKKVhl5/LKJ4Fi7o4Y/Iwmz
tv4hAkdy7UstKTBGWm2i1cnvcDU7E1qQTuI1cp4JJibDyv7TgxiNXpWak0xY2bnX9qTOtmlhCN6h
ZBfrkMNmFG+lRwdk3GVh+yQGO4D1v0jNlNznATkas34NFZSlAH8VeNyKy4qSanW25puZm859NhhS
b1AiHcYkn+o+vQ2gngtUnMGbQ+3o+h9Q7SKQFv/kTfUYq/aMAiET6T4QTtNR3kyPUMeJwqKKbZVp
vm4pErE6Y9X+NnTF3IGR0G2o2k9EUHtmunK7lvoRfCtC/rnhh2/9wXlpYqUuWtKuLhYrygMw9Y6J
Rl58CO8vyRtAFEFS7F1j/h4FSmemNVIf7aYOcePPMsYI4oQXXFKM0B4B8GHAiJ5mJARZQzkn3dAo
NWVdxlbF5PA5Zxj3Cugn8+7VIPsYNJ06G61TmFXJNpuZEHp7YjY6HrINu4l/X1yuyivYsTsS2NYi
WtLB4+KurVZwZCJBke8VCUzxoLLXaZ/FNAHNbZad3ZXkpGYBou4gNFbxN85bajqibiRbdpXP89W1
LePmb2fgA6e5Aq2JZOs0SqRZSvx2Vp+4KC3hg2iV9zll0pbhBvbq5Bmvqa1GVQ32beadAxAFbK/F
IaNgCxZqBlGIat2E1AAykDgVg2wOxCnB5tPrYSaJ/om0htuqHo2pgtc5J2GLJmzWt8vPGrX8Eq3A
wfcCOKusX63nnj/GvccFA9L81ECI6P0T4MqOfhW/ZJHARCkIqTLkbuoeI/QMN4m67kI+Ykq6cYbt
WBa5OGSDsJGsgsVjo3ZXJtYaAuyN5ai8gAmXSujeNmehFxmzMgPvYoU87h8P//eN34M6GzUmcv6D
imLpdGt/BXY0drFOh9Xt3i1ehLGlS9Wqilxyrs2XLUdWe3Gw+oZx+SS7YjA85IsOtAfHDyKHhz4R
O5Nxa+OjqSv/cMf/Ca9yaI3bhwGvJUcC+ZusubFbFvVvnRm9HDWrgk5cL/3MxSnhp27/YqiWdbnf
tXK4K8HolW7SsDezSRiQlgSEj3IKwiStFpSP3WhuQzG7TISQEu14nbxx3xyJI+VJXF1f++pHpJGJ
tNOeBlpDt8JwAXbmMSPY68E6+biXPr2QHHo6OfHm55bRVEKrYU/q0x3avt4oUd6WUciJE/wq/vhx
Ez6nz+2s5cqL5gI//NdjL28fjFgrMvU12zf5hy+TsT9lkDwmXF1cIawZ8TOrxu+TIpyosqZvi12w
S4Dl7aBbkQCTVO5frKouw7NzW46NRLLBN1YcjU4dYEP4SgKgTwwPXyYb2o6qFFm1b1ELSYqUV1V+
sHaTESIumrFx8gy9XoOufo7WniYVwwtoDsC88EdmSY8/dqHL5QrszG0vD7BBEXM8Y8tl6sZMnXdE
0oWCNh8RY9QW/sVOF5Tz4WAx1H8CPxSi8/3gcLr9NWsZCz32nPmxi3VPLZzDt122v2ndSgtqpY94
dkT4ZIxsI6laEZDaM4e5dUhioJt4sW/qHQJrY3TIX4FFYqel8YvKLJtsrcz/4nflE8yOswFTTRXm
cCPANuvTnAT0+xCo9jRpiYrSdiSC/ee+1X2LIke2CSzBr4zg1SzQ2T+lfjf2ICbmFUNH6oprFWi3
ipQJHSMxsRZXn3ZLEOUlw2ta9cFXIMx6k8c5g/f6dkmsfRPhljOoRbB+zZkIUEra2nyo8FTI9xZZ
X3AKaAB3q7+azaHYCV50wrO10H9ScT9FuZ5DsZoC8S2rfpgDqFQp53V5y43D7bPIQ5LquTlOvAS4
NkdgagJuynttL8cupQKD5G0fId0UQTT8JpPhnVu4nupvxN+r03Ln8IGRFlLF2X3h/4uQqoG/V/z3
VJ60e4l/6i3i4qZpnqsQT1X4R8t55jQFFwFwksW9wOLO6uEWPvnD5GQDMFvATof8BIv8FW4elFHR
rQNwvxzsVvgM2YXztWfRJgag/iar8IH3DL9A6AvcGFrLSKegxDnLkm+kRXSqRrsQrcoXFxkLg6SC
WT3lAo1mzywdtM0UZjohqfKfUioncrp3t3+hCEtkoZiOgZc1Jhga1U1nvuMmaP6IjoYpWZ45aNBv
+WglpnIhLnXwDIuoPev5j+ux1AeEP5+8nITu7VUtFg6wH983hDLNQ09tmPDInnuFJ120WyLJKJeo
QaWW/ceGcO1kEGlZCJGE4JmcRUFho5YD9bec4mcpkVecbLC4yc5guUDr9mKjjeMQ052exgtyoLh5
AN78VWOs5fGOtaW71sZdVDuFbgzxZvzA1KHPdqr6ujqT9SQ6G6Q3fpBKivt3Hclj5tocVyWdBMBq
99NL/MPZPNpaR4tHlbBqev7hkf+eN3WBXT6+cS2wGOZ7wm6Zb7cajAFKlYDMfN0Ksbhltw7hZBKC
mGzWsh7Vq+CjuHRYIHwXcqJJryi4NwUzTMgqsI/njcZFjLIbGTFxN4yOYmNholgUxr4Tzfg0SpVn
XOvL2F5U/SFbM39ml+wiyDHIJimKpvRiXXb0jxg5FIq3mAVRG4Mqz6XVpubGh26KfU1EYxv/4nU5
dcYhPcI1/SrD3ahHnPo9LVoXzGvQI0vrbOFvr/vxqrPCzaGVngTuNk1u60k0RBzjJPX9USMecYS1
/rrlvalLBP3y/7ShbN+uBdqj//46MWgSqA7XUlGpWwpA15HLSY4478p7cgLJlXHGGJmRS5Beffbw
V6cKmXMMBGvv0cKcz4LV2RzaHT07rQIFmUYk/FiaLJWrPnZcpmmdw7edUjqKvxld27gnzRYkA15A
kC/h2VSAJ0MrPyH85OfSPhehMuO7d9O4cgcC81t/QNncPWqd8I0CRdtQBdG8w7n+n15sm9HIBzWq
nFwEzVeEq4+l5+efM+an9fXHCdJxz/4+/BnCdR94CCeaTtF4MIqB916zysRw4Pbop4R+fw1DtzSz
P6o0IV3PFRK+9sVCdyVxnyelVWMY5nBZa1RPxyHA3vEw3/bUgJUjpG4xl74LJOKHqQefD6dYHRq/
DpmX1bpBcvXmb1e6kxQ3/2oOpXrMjq0iA7zkJq5WpQYeBTiA25Tsn/6/X+AUteh3vOW6E3mMNY74
ufQBrxpTSDGHE+emxrvrM50lL0RRoBsAwVnFay6hno3MFXNgVItcnK8wqpQfXqjlznSThNUmdlpN
jg1KeQhZC0sdgMUl4xPKAtnk6S2iL+9oZX3zwBT/PvvYZe0rhSSuI3pTg6rOaVUj7/xMqM7oYWe7
FOvrAik1wlCd63kIPxCKlWy5fY1nTS3XPWvLuZwZFg8pePNLz+PpPD/GFEfjeqFaotwWOuuEGJVK
w3Va593aAj0U04XMKW7lEQ4fU0T8dhozC6UpqiKzU9Sh7OU269G4F77YDBCerFJlZdj8+ZVtKgYq
fvGnNCsXDwncTxyS5brmmSbfn2am5ZJyrFdzCMTTjDSACFa5gkvj2Gbts1ZP1Hx/h/dMr0gkcdMI
fxdVu4D5ELxJh52PUBIM+ddHV/eaisstlLK4mYN77KFh46w3W/lDxJdj792izCJ7H3PRC6+WkrpF
BFaZNX1FHNWKowr5cYFnhWLkP6cIfy6nOVIZmXje6BiF6u3d26esobDdlJYkgWsiCz2uYkpEiVyR
WsyacZIvqeUgojxhSeVvl+H+1mr+79K746G49X3YQLnm15TPco8v50ACNz8YLiGoFZ3l7b5/XJVt
YFhXy3Qr9tjqZ6XRRHiSRJVMWjK3Zy9ov12j1HzxEZVE9dGZTyEbuy2g/6XR5ZDkA2CWGpkUZwsA
3N5DPlV49coiyWThujpCEU8EGbFENK4CSwe8iJMUeC1wFOye8qOjV6BuKJQx6v/pRFYXxW8b6c+L
Vu3yMzkEKMhjr26EB2CAg+etMTfAoDEvCMMTn2haGxxX2ZavVpqqvkaBqKN6BwqsHJKBPTv2OPRY
0whkEg797NS4B9VpFm/PCbjBdDYQ9JefxTZ9wnC52NGsf0VC5QztpwcTu4vL6Dz0aKMazZ/4iG9s
mSev15nwwspG80fAZ3Icd/NMZQKFh6hKaIcIk6t81BfJA0XArnMDm+me+Y4iKaMSjCUgGeT4HL45
tj2g93FNqATkgENqeDsPtINKTnTiM1crfYMKgWxAnLMbZlLWTEnWVcyD7NGHALNf7qtsvsaebdrA
jevUFnTTnXSIT55q2i7z6MfsSyhe4utodZwZ9t0CD2FG74/3k6wO8GrcNWxqJn5cc4LYvFx1e/py
sYH5Pw0rEz1AQLTO29P9rpu9foQdsNc+vbSwJ7R4nduPa2SJ1CwLlUJ956csXTkyxJeFB2MJdzYf
ibYCZW4Gb4ca9gORdC1/tjEtoJd8RKrFuzDeOWq4lavERJ7+MMn8nECftGeaJuuSFKd/oARLK6Bg
AVFO/dD42dkF/zFfj152o/Y8wTD9BqNLXPTHGfvzup2l29sQ40HdVOVprsXBy9rIO7gehnGHUnoX
KFBnUmyGIebv9HybvCFkMaPHVd0r+XSsKwA3NQqgeriKWpYHktb+Ej9kPy1qi/5ZG7JK5WRVUSfj
P+rR7JxZomqTnEelFuuQGK+YsA72DjPq8ae6ut/nmLnk1KvMDlL34egkb+OSR/k8q717Ti3HoWr4
guzbyfUtQYMQVqBTXUE0YhhGgzqEuK0NWSK1+O+/fIR8uT41o/PiIrH5siytIE/ObkGCE50DkDDP
Es4016EYzTePz9YzSen2WlLfDZ/0AbkxJoWqkHkbCQ6do7JQGdOyGfnJbEF1Vups6SxUrzrLWyi6
Be4geX+X3w3sgrrMVkzmGjqd8ra2cIBXt9rZXzRTn4Y5ajKpnIIvXAAWFGFfNc+Nr7O/R0dJQfZ5
/bd0JsdX+TBG+3HI8jD0Wc0IySNyolSS3+RWIqcmlkUSIKEWw/O4OYe8rc06jUtwg2l5Rv2n1Efu
LmINLeLLaE+6ocmNzOeAeKB0jrDxvbHdgcIUrgfAe6ls6gc+zICctRygPEYjlmY22eagunln3TOF
+/sHrS7Q4Z4u1qur2RBFIJOPD/jI5N5ifqAhbvWyWqAWeCwsABC9LVL6BdArFXp6tQTRcrJPi7B2
8JeB2Bd27MXLEr8TvZufG4nAMx9tFgwUKUISVy7dkhCFmh+CWm3OoEsgiHeelc/IJRj5nICcZj7F
pi9Bzvz4Ma/speMHug8VVSK5qK8r919Y72YVcPW5k4FqX6BoxMGgtiz8qnpdk4d6Xe18IcTx/uN6
+J+lYblNaAMAGJ5BTkZ+cbYQxvAeALEJhLKQXmpJ4EMyvywgmbgJAx7VFOxHqSYJRhIGR1bIIV61
cD05rphPTjV9GSqUR6JjNgFCWmX2iAurn1pa9VGD/TqyFPMjDNPHksQNhXtvzLhpRKIuq/2oab6c
zFKKYFwEsIRUSn85H9tkyEaK/TAs0kvndrtu9if4eyy6qlIxeTzr7Pd1NYas0NnuuIdB7Pv74Dw+
D2lPzDByg4mVYxESO/Qrn89CL2ZMKr/D5RaxPs7FaEpD2ZiCdyvbstV537LPQIWb79rkhRJz+9kh
KUeyqt693NSUzjDk8Bk3ovTDRXahWsK0qqOsZwBjDnwguQMj+w+J/QtQTwo4ycVRqdYOufdAD8Gm
c33mR7tlHBk3EX6Zj5RxiEdshdaCZkAGFjI43jc/9pyVcwy/d4LLBYdZKFPoJ9ZbKPfCWXwZDpMM
MA6mYSI1vMSiQBZY8Uqg+dNDVhc/1F2ulli8V8cOLzxtEatV2X4mBSlPfAAUUXVNwoHjmAwK8Xar
xFY05DW2l04s7vMM/Jd2CLvgeeCU3XuejXrXzk4f0PXB1gYh/kFzEp8y/A7vnygzwZXzl8wBXGIv
ZVd4y9n7PgCrcraWqdu1vRIkWPmIGTnnYQ5IpNNmWHLGX9uMQ653xkqI5S3jD0uiX0jbVe97YpBb
JceiSI4C+SZDAYyVJeZSzxL8iN5vKYChj9yxUmzq9c524OAzTQ8gFmQs2qPxf4crkEVK6qSdxqU1
flU+Hkn0GYrbApbq2Fntx7uUnnsYGCTfj4eHUP6Pl4IlK5qGeDFKvKl8q1SjWwdmkgwkuZp2yZh8
7usRU3tcsFLM7CPP6tRVeCC4WrNj8nUSDAqgPVwR/bepQUnGPNNyYcTJ7UOxkM5dNxsaA9rJGR9j
5+KjKfA74mxMu7zCdyZOy0wFar8oX5sM5w1JC1RPTwoQQUk7dyh1OaBMq+B7kaaKbTAJJJ6iKmhR
BdKLYGVDDKhleFqNHHBuwmxJwim6YhTDkwFgFhZ/j5b9vYTeNDLt75Aapp/syqK+qes1MGKWeNpr
TYpQMTAZdSNr5OHmpk7iqBMfHl7I3hLcnhl3AeOt7qxumv7LnLJfjxBEyWyvsrZh/kx7nl5LpnyG
Yd6liSyMgEAHcr80FBFC3pTQgg6ashEl0uJxe8Ds8sIkEDBHojv18Ikwyn/LrtjuZblIrshQbkwf
+lC2Tr40vAHdcyn44tBcdmal95yU9kErWnNzuvnVm9p7/eV4xw/ztCsx5w2f30GKozxbsiFAxVhk
kBcWjbgAfC0lzSEFCe6oQLL0Uxp4xcMmqCft7SSL2fCrQUbduJ4Qn3r44wOUC+UlwISfRhLbg4gH
6sbLPsEemWirkkPX7A+Na/C3Wp56vqS7CPUipGWrQE5ONDPCQ19bGuRxv3T7gRpycHorJdlzIbAh
VgESp3vV5YGlPpn2wFOXkbacumFlBGt3iXZf4jQGyAN3uJ8E0nVN6MRRkAe5a08VZHLLP5rB4hxy
cMAgS/6qv4YH9YXiPjapaCFy6/vLJmL3weCVfZ7rz5u4+TTbUfkzMyKQUhpNwfRDqxWIo650giIC
IgnW3kwC9mfdfXc9xFkOe7n4iIDsSKuHM3S1hwyfC6UpoikYAJ2s+2huf2XIQWGt2sz/tDwFi5Of
si3+sN9gYHWEzTTsT2lFOM3HBSaUDWOPnEw9baMESq5fDmwGSpDtJ7sgBHgAaciWkQmS/x+g/ZJg
F9oJqWV8termlhf/pjE5OYcLWEkO09wUKIp7q3uzazm4csYzjeb5304UuGDrpLN0b9IP+8X0sPXx
Mm1BrTSxE1JhqhVz0H5IoZTqu1/ecqOmb9v0CKTCPulWNxLO/eYQWuAb6AVM+2IbJSFgDmwIN8d8
sl2tIGrLNM73cdCKlYsIuuqO7WwZLIC1M1gIB+JOWIuHviILd2SyLNd8aGd9GnES5xhWES2tryZo
BJYxyVEPAAIx8/GDQyktfw6qNzMQ2THmRciCe2KPxD3rGQd3ilunfmsikjjTHEdU+dpPpnV2Uqg5
ZRe7ZarHAqyzzdnzfGP7YHSw/zx3apJwJvivLqrd6H0W4yWmE9nx6yLR0beeKU0VIwgBWtRdmf27
7dseSVXTRoVdGoTTj3Z6i6fN7GS26aZZ+IkP2URVRukpTpVbZ58JaihRLI2/qwhvKiDLN+dmZqhh
k7EtuaQSWCOchJft3bKxRrefnaq5UjzFXv5M/ECat1zPJDcT9UC1yjdj4PMf5sLZLq9s/5rMVbqv
9ngBhYQ8yCrZv99QTiS91Y9JMHOa4mvXebjHU941HfgGZFP9AbvpuLJGRFDEMs/TnlcwjNhS8MUD
Y7sjRwoH2L2TZQUKb4DKjHNUIrNVBxnH2FSjWPqeXevrrvhk7aUBNIaLLb8fqcW+ISWZuvq7QwGp
2OWDQMBYK4a2xSaXM9zn8gDePjN+RI82XT8FMal1qlR/clBsinmCJu/5K11xFfctpebeTcboV+EB
PGGot2auFkJJb2VYqmNKICNMx/eQhL950YJQzekRrsxnBc/keXcTo0/I8m3AK3h6fjq3d1j7BpDd
evYqe0jHK7kkNe1uINV4rEOy3bRLpE5zKzta3bmfWlTdZ3i7ncijuTz6e48muFjENCl2r8FyqfO0
S1e6odMFuy4CBh10Ot2y2yqQKlkxxN6IaLUmgI20C2znswVsxC1yuf82evgap5U/K2X4GYokiy61
AGngi7542YQrTzGLybrRxWOSyWBq/omsCULVatEP28Me7xDWhAo0k41HDyTd1QOO35h1gdCR9nAE
ve+CZw7IyYA5gTHYDo1MwaBhBy9aJHU0j9dhXVHtgvmm5HCqmpG5kJy7eSfLAoZMZxKja3iF4d23
tdi61j10UJ4HKdMJ/N6KhTPSVsM5lPoGsFqKy8Zp+5nLyopU4Nrr5/qBehfrrGDoQ4WLZ8mRDVXR
aNUlRwEAcd1GiEg6AO4+K+xYJ/ANCubeu+Ajpb3H+2bZiwe3M1c/FykmEap3v7HBXu6cJFYLAe5t
5unm8Tu482sqrtbM3Rr/463uFm895yWVDPtl5Rosz9qUhTFYxmBAanUwBqFO/hI/ETx7YX+dI+Ri
edCKJnZXGtVWE7VYGSGVBXD2rlL5YxayFQ1bl7COfMX9sGFpRL00PX7Wcnu0E11nCJmxvd1TuBBW
SybZNe4d+/MAK9cCJUrfLJrbKbrEDB2XzdtmfW7BghJ/SVOGB4yzkvNhJl3HoLkik/KNYujvYboZ
FZvMZzqmuZJuH4DD5MY3Br32rvvAvW5b8vQCsQpkEDI45AfADPJVb2m9bil+IKgm55YpahwmtSs1
1Ijmg5nMrf6jwTXm++tiQdH8pmYYI5W6urhZVuQMJ4hYC8BpPGHRoTOw4ouDM44iuiGgY0jkb6RF
7jPqYLB7GGBgBsBRZBhs9v8tfC/aRddkvRvzQ2r5b287fVGDuUy0jXMsIzrz/7+g+D0/+PLBTcfz
0urRtDLWLTdWEl6ENSey2ZxXQFb0RVVcNAM8IOCJQL8IJNEiKgco7Y3S9cYJw1fz45W6M1uObyQG
esU5Z90Ve7KZzk0hTpujhs1ZRDq6gXCiB2h0Yw/cpfLpOh3eX/N7ET6MXnsPrz4bgOH42iGpDy/x
WtwWclobD+yVsOm4RpE27WKU8JuWG3DOShBvsUu13ttQ4PGvsczk5L4l8lEMoSpOxQkzR7ypdHlv
vIOJQMtjxZzxys3KxOfpfERNx8+bCV8eTO2ct8HzZ1VCWFhLmIwKLNDAZr5svL4hZ5Ng96YV8s8e
Ee4YS2XROLraqGYGQDXpkCVA9PBWe9TftgKCrEeGU0JE41cqofuLFpcUqCw2yOMyAfE7BBNeIaT2
hRrs3u0MiYLOyMIgHdmNMtHT5dGYNWsxqFYGheWgTbPDGmWyKkP6kuTR/QbL9i8W/DkmuR4ky60O
TPXjUObDY5FS+wC0bAAdHj54aFcv21xvcvU+XgTcFIu3T/lduEYw6hvUmRnUDwzp5eKp63escg1q
KAr/aXmGA6WOyO/t2MK73BRjOgBOQQgzNBUaZzC54AuOdVem1PlH9Wuy+Sn6UxvpNQF0rUCqwOT9
z3OOZP81qIpd20LL5rCDTGtO2kpMrwfMPqO5amjHBR9ycpnzqmXIpINVEiSG60dFVq4R8yfqJs2r
X/lLtmQzt86JwZ9xIbxoEyBXywBfe1F47yCM108uyW9UtiEs03ko+/lDkmlucBhNehmvPoi0oxgA
oocFr5I8drG3AFdqNwXWwRd8oJgdwSgeZYGV3sePPLr4jTidvKJVCfvJIOT8/itFf8ARrqGlGbK7
5927WAUY7w0UM/iX9bSXcl61ssbl7HGACfN98BGI8HFjkCsrU6Q4HF5UaMh9YtYi1xHJkvb8NjX6
GxVXERcBYi66pC8Ggw6w0x1hGTmwTZGQ07xCKxDg5ae+Yv+q6tc3fOJuMaoin5E2YbaP1BxucmWw
gu8sD5HezQ8aXJNqDgiZ15tipoW2f8z9IZxvO0+aVR0LZ+n61q8859YxEfnvdb6qJajLWlpY+xp6
4rM3m3oGfj1e50z7shHcnoOWbVdQcckd7R5dEyPMYRA2HMiOMkntWd52OPwJBuqYGWeFXnmKoDcb
+wMh7XN32rk5LP0tPrbpCB2yO83p6EZxYY7GFUaV0GuUrTUoex8pr+m5kBWvs3Bks6lsYN8X35Eh
UHgVXiO2e/eU+MvklniNqAgauKFX0uH82SrJAmYyhlaKF2m0yLzTlUh7JyZSRx+RiYzQcAs5cz5X
VgxkyMMFFqjqGrESAqtVaoRey2kHJRh6eLWqBoyAP4I0UWwF9xZb43lNwFkEVGS9NaTBuaO6oHeJ
FqFRhcyRZT26j7TUgWe3MWb8Les7SIiXJuqK8v+QTyB1MY/y5yi88nRY6WwP6BcL/MyrgmVyIEqA
a42KSNWi08W9Wh1KPM8vsFPeZTV3p37cdV3Dj38XCnQ7p4eUZK+HJ9gSI1VcqHkkYk+s1XZHjFc7
cOzZXmzV5cTwtpdAsjjEoSqeEoZVEHOt/9N++gUwHhJa2QhgDW1Laeh0o/lGNbDAv3drS1FrGPId
mABxZJ5TO+dA1/D+eyO2c6oensWXZca9KQemID4YQc9TedNQBOTexlA5Wi8a7UTiVwFNSzFj/Kul
TOHSqBnJpkVZXjRjkQ7WBScO8zgjBeTbrOxjNqvw63qxFrDcDoJOdYMkXdF7CLVcHZJg/7uNJrfv
vSKTMmrHWbRQUB2krDUkEwxXnCpLRJ5wBRlJ7t6itRWDJlPBH1IVrnSXBnwqEIHvb65KBbddkPO2
puEDRcdVHM+jPYG7Ux/cLKK7nKUZD0DUME/3sGUZfuS6pXPDrRpQt1X6TN+IYf/asi6HE0TwMpNG
nrA8uMpJNifgpdmexOjX18wYv08Ln/wm8hdoyF6HuB7NAo+qsejDQIAdwyaexjiOUYHc3tAevXSd
mDGE3TSP7C1ZICjHQKsDsz2yDg/v9mcnjtGwQFGp1Rrpi1gv3sPqnPEtB0j1ubEgPyImdSXg7MkO
Aj9YA2HsZMLy5AkSmx3vS2W73RVUHeHlfBW6to6frljmUDiAXmQWltLCiFZ406aGuTxlafCuF+e/
ylxY9OAYGOiaitOCn4LEulXQpHQiYvDjwEwxHAMOCqQ7LKx8QnlsIn6/5FFerhAL4kLRhBcCuMM5
pS6hHlfU/Ps6QSW/W7s7tq0APAQmuRVAahbycSx/4rqfC2smubXPTX/m5XXL8TirWmF057yCUXXN
lHAr2s8CeEEiuHUUCHpKYjtDx0FOu2Fk3XIDUNCVkRBKxWSSN/ugLjDkPgMyX5Vdbi6Hn2ebMGzx
T/eTumj6Ek82BLo51kzNZ6pYolNTcKerq5kyK0CGynN8bLEydpav6uPlvoYdG+Voibbthg7cFFCi
j1B/O2R1MwerPT3ovs6DcvQWy/wi7t5JTaVYRwOGJrijW78GtWVF45hESrTnzx71vRTK+tG0cVFM
FoMM8WnHHc3i/ZavD+nXyyr0MNdm05YIN7KgnQ2lifPP9f5KrgPao5olzYDKANIwfsuAd/3dTfg5
WkSDbhSAs59xYQz9E94BN9G1wY2yJAF/rfewk7pR3M+FLVSU0r/OE/HWCDzkBLonKzLDBYeDDdbj
ldQb2bg9VluJ0QF1xvHOMplM/fyjrLgcfx4pnGh1ikbaNIT5s+UOuHlY4Y5jkVZjgYzyu3FP750/
VA4YhQXD+HbDKLBi2jIIvu6eaJNayD2zypajqfJHlZRIf/3uXDTnhy9LnRTERAR1Nn1558O40P5y
WtryqWRf6IicqmG8V0sIuDaBCE+6dNjReyAib16xJKlq7VilCI7c+4Hton3kMKro2Td5vkXlx+8R
7YcMHRLekr3ugl0xiIPpUoGAxhdAHC82+wWYnAQpUy+OX5FLtBtyXRlP6ywgg9wY3PRgvdCAwZlE
iueUIo3ljC9EJVmzaOc2WU1N0vb/Dklm5GPudaYANdiWWcqoGdnFHWeTU97e9LS8/pwFUQ/RMIOm
JAOFiBPzKcwD7ODo9WRI+NXhPiuj4AXs7T/LNQphWGwN/kA/E18T3kX5Xlt4r/32ka0BJC02H34F
UG+DVji/SE6F8DfddK7MbAAW6j205MNqyOWmalgKn76bUEyt33eO3R78ZuoHv4XBjORBGvWdjsas
W7tkZLqsoU0OE8hn7cBW4TI/O6VBVGljTUUP+wBMAya0EMlZipNHqTTAvOrLQC7mNKoDoYa/JE3Y
n+pXNVZF6R+YkAeenr0VmT4G7ORXcRJO347yj9WZmsYm7T5JwcC1/A6jTknMHcmFbgQi9mt6rm2y
KqSaEJnmqEOxbweD4XtHQpyQbxL1Na/xrJcqKMOnRjvBxqU61W4g2T7NqY1I7zOzBfhHtULzkHBz
MMMNQGgvir/m3JZLmBkX21FftTyD0VDarB4PuKHUdYNZTEafmdGRRgdz9tah4CIvztBY2HwK1Zce
83wTLarvFUOt34RvmYfbqSLAeNckZ31PCLG7//ugp1N2yh91TZ9bAIDHI2TzXn4CXFnql1pAWX1d
JYxRHfWUmS5gSItilaKT497aIlcvriA90fN7Mn3TcC1KyBGLly5ugVakDA9qbK92JRj0vXJKlB1O
EzTZcP+ShpXOEiJIa5TR9pvM8ACqe6OPiPiJHqD/6vwdYOusZ0CTzpDod1OnSMs8a5zq0sxBtemm
+yZ2aaYYlBqhPwkRizgcpiEL/MdHDui3e5u/HIGWd9+bU9BaQdIzakJibpTSACNexj/woAFo+56G
d6TOeikrUL+4Z5DMovw7TK/DPV3CMIvcMA0jCdDocMBWBA08d+XNNY7cHmzqXmcduAQP8PIq821f
CjxrrPfL4BecpLc5LQtiMI4GkpSIiwekYwqx/gA0b4dGhN5EF7O54qKb/Jm/BXAI/F5X8eOEumlw
fH5I9Te81KOOoiAanAkoO2vPm9kEz3QCIlwAd6S97uAmhWp1no70ALjNFOKr9NECbpLisYRUUC/j
YjxJvcYsklRkjtv38n5CSbbnuZQanPc+xu7HvXjMI2jQiZhBOd49wuqNRLV2vkpnt7TJOxcH2Nh8
76jB/+yBMpYaBiSE+cmrutVnYSOSx8lKnn3dYiLBNwJAeCvZII9UL3fbts8NGnRS9LEFMV07pHMP
T3H3ABP13769JredFTrV9UV/3cD9ypEEmQLlH9lNrEJhhxKkmtrritzYFvgqY/uApco7s43BTzqZ
Z8CFdaX8Qw09oD+hL1g7qzUJZKF4Qos3pVMPwrU8hLjePV7dENtfiWTU83qK924iS9M0c7huNc//
LL0peirF+o4RJ4xq2aHsbDduzgdmFRZrb+JTjlEfeN0m/6S6h5LxOVHv+alVZ7w8yhpcpSsx7ohy
fuTJfi2W98UFJIt0MpHC7uhbBVxKqagdigkONj50HNjFLGDKYxElJ7NzR7n2AEu+mvMLZ0pn9+Qk
Lq0b3Y+z8Kb3+nBCx9FTH0ogZlWyPPpUjPYIRKLxJMIBfB+k8gZ+W+pnZvfcq9+C3qCKmv6+lu/g
wJk0Pr0ojYF+gx/uGXgCSmOAv8tt1cYrB0jsuVOrkkxJ5tdu49SgJ9IhI1aTnn77CJkhwi46ZobA
i36cdr45r7kph6N+nFVphN2wf5sMggfxQ09kj+xPdPQ01wBEpWvA1zrF4sshOwc4J3l5C4vvrPgr
OPcT7VPTDhdqrgaGxK8SXm87oN6JjuCb3AZRpu6SPbmfs0Bb4PX7QMxxtOePZYOLmBqThps9fZXH
Ao6dhcOZUSMKFXl2rw8yCrGfZ3JkjDWdPUk39qnPT/PH22XSGTTDFJcqR7qwdl/uWkhRg2r7f/RW
q4UNQUhVlw8OD7YvcF913vH+e6NGNQ0Sd2ZfDe9xxQsnYAem4/05U4dH5ZRYI8nSmrxbdZPWZlNn
ErI9qdWK1ThurbSX9M1Z/fKIyvCetbv8ftGBFx+zGpoFKsxZAXJ2per7ChzhFKZQoJbra8VN/NqP
4ntL0dYXZYcdmgM2ZQSuVP3JRCysyPtjYJDHFqPsT2pJNKyRAskdr5YWDiD8D8lBCjao4+i1KQQB
9wB1IIREe16A6scmKdlTGhCdR9+vfW+cJXevBIxKhuaCPVULlY2TYINXr1QZgAQy8Au6utZlsy6r
cn4niovtucZ3s/Eqm24wOnUAeXrl9e5PncFufSIgW9iYJQgJUyq3KSuyVYbtVFDaTErhez9cOFgR
cDi8Q/tZtUpcvImUyrL7Ewqyonsek+2/IqAto0kJuP+venYGC8Zs/5+t5pYt6Nwe6cNaSDY+6mzc
aIDIkb6fUCrltqat7tAUO2eoxpLJtpYgGyuIlALiOFHyBYhCvDhHnSSUh1b86SDLqE/nHf0XEJzm
Hx0bw/Btc/MrKQJ8tp2IsqYGSWWvJ5U+T1w7a5VZCaRbcL/ML+jhlJMX9fq+fkXss/ulXztO6pOL
DKqk5qnpRy4LIwB0kfEf/4TliVTLPy5opqGSTLnUvMAg7fDfpOaY/7OLfvaQ/CEbYMOSD8oCbOxa
iLvs73Ijj4+9fm7JssYFY+vDLQheTW76BHCS1G3OJRbc7OsZZ9i/AKMHhkvv/8dIN+nMIuWj/qYO
rmE3cPrjom20hwfGpFsPt2LjU1i14GjAC1N12A5Tcp+aJn3QAOqWFkDce5xY3xY4hm6If5XmODG0
YNRsCowweFIC0JrpbT0BLY4IcDkH9b0DFqNOTSO76Rpesk7iI31umlG82WAQ4dW76cuR8bU10LGC
LR2LY2Vl9MftYokeaw9+SznnZA1E3YwMLFhVtzbjvIJi8wtqFiNKZebblwDmaPQbORH+JGzU5Byt
7O4LK3VpWeEq9DW55IO0k6PmeKIwNs+rJnYZFDl4hZ7x+LZfX7/Mh7Uvaw1h6CtLjVqDZDthzPP/
NFtuyecxURNLU316D7v0BhXjfv3b5JVNzEsmvVah9FN7KSQt6CmdUe+zo3S+zG9iaFUPtIRtMyrx
xsTxTweXjVMCSrtoshZwTu8WpvQYsO0UDZXc1MjdxDDxnFCsbNXJunGHFOxTllH2NkkwvCbViafB
oLvipYpPqP9s0AN1qS7GB8lF8QFlyorl3XjATGH/58rMUoI55gfyYmvPFvsIAxZQaQtkNCs2+0ba
o/+XeBL4Zp7b9xZdvAvAPxenues/sTolEsuDqSFscS8cJQpeDWMmpvUYNAjYVCmslQPfucQnf0Xc
88V3d6W8AUF8XzEIu50eRbl7tkftZOzJyui3ZWF4mYO4SIMNQEv7f9KXc9M6tDulgMVqnXCTHs0D
42F6dSHW4IkbeVAgZB6jgAFG15RRfTFoFrbBJgYnVlwkIXg+mZdHDoyBUA+RyzqRrwGwE1U+9Jeh
6+jh2cerxaX/hqH74obkX+v2Jc7dcaiPbl+qXfVo9xu0C+ILpe++MHm8kvU+G9yQ7Cqe2BxK1lvn
qXjmViJy0h/DJUovtG710Xado0vwL6ZHCqc9Bx5xxzlxpf8VYFwf3Cm+gvnjaJiEe/sQaVcI6w4x
REeJi05j/nOu3JiOtuxotXNtKgASGYSerFvL0X5GsGoSe6+bVJyGNWUTovOdXp/gGu3isu77xIOz
r8LkHXAqmCHc7ekT1rm5dOAHctq/MacUXQOT4/746ykrmHz1vaH7lyD5j6D3aPJF30wBk8PGbGGJ
tFw9Wx7LSbNDxaIXLxKsKQtHF1DvcYJxI8CJwGJsMZ96djNMNAHpwqcQzm8k/lHbI6RV8znQ30ku
6KvMtt+tVSQ+9dIrp5Y/M4hegqseCvmIYdTyX8vkG/zMwCTuUUqOjpGAE7tYgFK789vBemfgxp+2
3pxtfLAIiJeMVYvdHWVKhwb0jFq0m7siOYcMyHkISjvsSuzNHWEA/1hQ+vSe/SCI+t8BE8TaYL2a
sJAHaXQ5EtTSajAWI+UCGsnvoWtqXWuGjDX2suC4rtLbLHFnTe3GXk7yT31/SZDefl0rjcy/FrCN
p+xWMacdHOgJLqr91LAkScPDWTQghrtj2c9bCqnPB8A6s3DS/i9jk+ph9Qf2cqNjCVW68JiUnu2U
fe/Qbfjrh1DQ+UJzVVJrNzzhSUgJ4lQ1qyAsja7+ArALElyC1toDV0tNtIY4xrenDCZ+222AX2Jh
Qmn+GUr/ZgRFQUJ7W8yUrkkSRakZ2qVS0kkIFujcHo+Xn+pIhisUh3GiVWo44kyeynVi+0eX5LnB
mMCe9hFTXoZoUzK0iiKNRiJsC5isgiun2DSDtTVD0cbQS3vQJC/g8MpVd8SZPkJEME1xSqXIoKpv
ZNMUXqF7FbV+4cFs1s4EOrvY1SVB2WVa2HRXOWVCJS35v13lqm5JRFIqauUFXQ1f9LxcVDrBo11c
P9HC1hvKjWhCZhqVvZN9DnDIHbZUrUn0Eql9CDuqB3nynagCCABSxWMbDS1m7ZxvbElhILJj/rbT
RPgCv/+sIXvZefUIanKXw9wnq0yoIXCeR1XLt2D/AFzNZ0kYiiqLhjefdkXYR+l1OkBZ7/mF2EOq
ggcH2RaioPMfXkZsjtckt14B1HFinpK2cSyuimqua48TW0uq2OWSMTjYQW063RX2eiv4PEjAAZXk
spuUUMYNP32WtGITDJ5MmJHnyDusifoPP7AsFTGqhEKeiJepJcDXQ4OwlUku27ZgfBgawnbgussQ
I2HlZnNMAhaFK9HexYeQ2Ud7LO0ZIDPTVhf9b/KUQOfzzZELmV8OTiX0k2KeQgI2EY/Oi9+o9xMA
A92kvA8Owgmbk4jMkiFk/rk+kJcPmREwUwQKagvsi5Pw5DjzLHgGzcNplFmg7LRbgQYUs/sIMouC
WmOvmkootcWXyi0CLNHltr3QmG7xYdzLzha/5CBwTwFTk7+yMmElCZ7rvS0/zkViQfdwdY3GkGa3
jMD0qKqYqJPb1tSxpekmFifY+GdWo/5LVD09xcPkXxO2bgey2SRtBZvzqUSIrU9QUJEMYYPl/ODC
INDuj7dpy4M/WMDmfuj+eTT64O4QCPt0WG4DglryDeiA4+Et78OVVLjRFlncWlZTBlmPVyIrj3os
t5ir7qDaPmkTTDUZGBDiDUJuQ7FEJhVuSJfUMEmt1Rs5QbM7Aqy8Gyuu4yq9PsYXekwCS0Z1O03J
Zb7hPXYTy3wUAuBJIEYi7cXslLnSOYm7hiQvuY+sC06NIi7OEa+vpCBg61rzn/yIZjeoBSf7nIJe
ZlRXPhDnU4A3vbV+NPMMIJTQQZPGsibXclu9DjbptmFQbMYlWd8F2eOOPtFGu/SXEH+9ywq/tPWZ
O2++qbHZy7smC6YST2myj6yK7+zHdrYWaOdvH9C3H8wwLjL3h9DLQypa/KWCSnFDxI18N1ssNoPu
bGusOGxvh4LyihIGNOs+R0JINd3WR/v0ShgO0kH6eJ/Nu8ZPPiwHDCFA5JeupW5p44EmMHBTXsC2
iIZ740HTYcNwEdB31Z+jPTqvwR7wCnSwqe3UpiIR2fpxeGjajB0Q3eryL8h4qg8b83zF2ksyEaBx
pQj6NH7xrz5mgYFtyZbfGCxuPbMa9uoYNRTMhBGQx6e18cNarsCdBMxN6U0JXeIUqXgZAP3vev0w
eIgtbx9qyjFDbN8hle20RXm3AsKFGefXagVulOZ95sV+ZzJTbNrYawDCqel4G+l+WC6q8XlsLiuq
bYDqVKzGcrun+X95DTs/S0nXe6TwfE7fLVmwYMUq79rAt1BWfVPQNPBTT3GmZVbsIUUEiged8rlW
V8p+kuuiWkoui23YjMxl/3mItqgrpe7dLYFjxTeHwu880u2GXQB3y0ibxUEE/ST1wDM1HlG0AKdB
9IQqd03bkx5GjIjKJhw9lcqCEmfI8LXa1Oolk485iKxAlLMcoS3I+CLVaL3Gp6F6G0nReTBWai2B
DZl1w/odrv57xTRlGHwX4DJhvL7dXWLBqD7dVh87pxlG5wtglLrNgp3mSWyMYHYfBLhXNgF0jaBY
KkvB5G7vlto26plfh6DKlfg2ij4ElMaA3Yiee9trl/vturRU46bM01FZJbLv1YJDx3WDME+CQjN9
I1Mwr9Nv8edXS5rssoaVGQfx27DNQNrVYvS2lXKbcX4P04I7C5yhgOnZeDA8/SJcT9IVNQYZvAWW
vWUqnvSau99X4ZFuWnDhfNyVzD3BD0/1CRG2DMdERoeGG10lVddkds/q60VmSE7DBr5tZdGeyGE5
xVsvlM+koyC1S2aqo+sC4nSGZnl6keNA6gMqQB4hVF13KyXA1U1ZZTad9J3ho+lTNTjQAnthfyBZ
QIZ79BxBClQ8Q4/9eBr3qxm/KiHTkmi/sGgwp7MLL6VHziG4Njr2Di3yqBwlRu93z+a5hN2rD1Wj
inlvPTiVfTPVyG0yDWefYFCopodlHoZlW/AEX1Y6E49xNSi0MLEbrMp2LLG35l31izhuIMbMxt9r
HOdnA5keBK6L+JYGsfPYiKdbflhQ+uiObbltq7Djd59H3yOVvgacVJ+NL/oGDdKIUKlDlh9Kc5VC
y5EbEzgSk7TopWxF8idMaHetK5I4Nk8y6imD3wNww1+04KwqrK6HaMiC+/jAKzlzOha5wAHn30GZ
7f1xikfbGnZQs5KhyicawogqWnrDIstHasB0sZ5oU/tSVjenYzylIQTZAx2M1s+5OUaPKvr/ELow
CzoPdfk3VGuodYN6/rBPq448DHtbHBdmkP9sWc/mPXi3dEUkLmct6+UFvL5jdzdV87mXUVuuFXMe
Y4q3yLR6esxudtKcPeSljo+iTcU7GfRN9iN4LalfIeatstXoPjo79pRnhGhhsp5nv3lqYdlFBoRf
rMgSfqQIAhT4MRExmDadmTfdQw2386ImzZXGBAZZSJgLxRjZVMVAA1ppR0rSyEgVxOGd6RcS/B4w
Hu2wKkx/8a0c2PUFK4yurROJKrCtuyGpsA4yiEqsZd+OtkwCsAK8duh/QFIOHVQUrt+SXoqjJJuc
JcqnwdxsNJfrO9x62zVtyUtlhJdbn5x53234IfuSbzag6G379NMcUIfbUmfda1oq5X5SEC+l59G3
3LOmxvbfys4xaEUKhc6YiCTAuYETgievplNhr2g3uATquSr3tyZmdu9Gadfe7SLezOTSh0tpZyRR
AzVTOCk+YWgMkBRGMQVcJoDU3fw4xRhaLZ0a3S7kcu/9WnUHtUK3WBx2GE96S+1PeMdu7c9YL9Tb
6RsKIpDT+rzsPdOhYeApU+kgA9ww2Su9kOlIPIATGEdmSqXcclsL2LREJuoPjnDvfRqNTHGzPsvn
DFpe4HAHmLHi5RMvYktqwxlCZRp50gGDOjxugHDWAisZMiTfp0nItv7Nf2doExVoMKPqeS5Dv+L/
U4KWStkOJ/AzFVt3RsA5HzNhxgocmlnACqbszckVOodF2DM9ENJ44mQrosLNN8Zx3oYJ8uqX+XZR
Y2odX1gYT93Y9xmZKvyTW4f21Ek36w1AdmGCqxRfDX+gj01KqGVl8E+ScGbMnmpII5g+VxWWssi1
S76O1MCicfDr7S/3vYlltkBwuPoIBLADjZlplAlOVXF0zfqMRUv9nzgxeu1luXSovYKwA7KR8J9C
sqOW5bJrVWt7WCxnOW9ib3juUtFwteLOxIDEKwIdg6JiZdiNaHsfOaF76tHL4tCqSkm4YPGnDq2o
M9rQp/lGJcG91C+8ldaYkh+GTynmGSu/ypO5YpGHJQmo0kzxaVeBsQnX0o9xzuqvMf5eTbb8EcEk
lhI3r3JMmh/Kluq4zitjMHCP4xxz4wcleQ3ybitHa93fyDRZyTJffJMoBvx/B0oqdmiYtmX2Peeh
INAYQ2j7TYiu5wnUpp9gJPR9juvqg7TztIDcmR3x63Jefdr+xoXBHZlMknq29YmVNGFuktMNbJ68
WQdDvGl9d+QVfGghKjgKomJ96CNbwIsOxXapLOjLzipXkVlgtmRFApD/iPYbJtDN4dC5hWMzxHK2
ic79Ftgm9zQFItj8HfYnYzak73/P9K25adaw3Xynr6IjlEMaZqn/opa8ow5u9F50uRELeT2khZDM
JYfTxnNx8bqXVXw9LpWd+nYwFo3p7eNxumQnfZ1znASh03dKSEKgkAyBwQQmVmoa5R5tukCYSD7K
20Bx2fnei2shchZKcMgTQgIde4wxX3sl1DlKYzp6TdQGoBA/xvjmQCUIYWZgeGxISTdVSYggWX4X
GKKkaoCAAEbHdTqoDw+Pc9JTAji0aU7UE5JXISU1Xls1eUthCNn5IvKd2M1TEgnI07j9lGTqQlfL
VgBkBQ0Ot5x/koeDixh6imJH9S1CQtadOwPSbecE8RQYt34AZas4Gc4hfSTU3TZ+wU0X80wwHux2
Ul78a5cb1D2drJ/VLn7G2VROvxRUAtaacjQH7eiUHpiTbHW1VrXaFlHzY/9rRO/pfbgpaQ5/oJ93
EXB/lsEFJacKSLRtyPvdFeNaZzFD0UbH5D9r0rEgyvnE233Lzf0x+47V2kUBmr9dMuaszRJXbPV0
DHVyJmh6ErEvHdBNfsT+8l32ox3uuZ3OvjzwbbVBDzSB7mc/2QaJkALsd3zrrePYO7hswqH9HdPY
mTl9RQK/8bmSzf24d8/3TCZVcFYdpLpA3IPZVfZeKDcjFSlL4jQ4ctkqqjsHYPNG6R9isLOuurxp
boQSUf0mjvfoOQGevPu+KbJeC0xQexDDQI4YWWNKhe6A0aVmIg/3qKg+UGm3mNRDVLm6T4HUwX9y
iKZYkVBV8Z3YKRkeCl6ZN5ajnLmDAWKpiI/ppeF4uO9m43CRR/aXha3BuZ1XGlwB4Advrt2YB0Kr
ked+qi+64t/MrNpyixxxS51jNoGmAX9jiljcyJ6NAyjmwECWTgjSPZJrtmpTyfyMrYnV5CcZIGgV
HcAK8S5YpPSVu91ZPQFqgYLv4liGeg2HguSN7tdSSiK/VepLgE5eKhghM7bUfrd7NjdlgfLGv0t/
GggzU6DlQOj8VzW6ALVAZHuf23WVIdb9g4OKIDb51RmoolYoItbdFRdPTfphm1Esc8DkHcYS5Y3t
uTXm1a6CsGeacABp9JA5FYI0Ve+Jn26dn60LfZ1hpwOS6On/rHuCjciHw9csaKa2jfBwaHI/c34b
zU3UnQhh+arw9l3HwO7WuRFZog3dJUUegwqCrIhS6kuH0OXRzIMoz7Ti+MpvOV01ktidAiKg81Mg
9pU7712VVhdHk+/CWwYWE6f6Hn7swRPbmNguNth4vH/PhotjJkuRfw6qNLMt5t6vxUSeEJ8Mr89V
YsKkNKZeS130kJPSmUBYHH3FJga+Elp4hXJEQqjpSzQ0yh7Vcrxyn4uL2RLqOJfhhynYddvk2ex9
LtQDJ1znuCNfKtBlxDtXyBg8KhYqr6w1i+Qtah4SC2Ce1bAtn0aoJDHSH5b/ql5slHNjY+p2/QIX
dHAtXJa8Ga2ud4pTc25+8YMsukXIDvPW4GHLDfxZjnAP/jpOXaoaTZ4DER2E0x8eW/n5V5qPM+Vl
oh6lwukmQgJbyY7AOpxhoZ/HSbcDlfvxRz7YBK41s5A2EdjVTD1qZg7MMYwIhoGqzceoR3IzxdQ1
eA3F6yNBJPRr174kmBtWvaRoufRXvJNcrjcOXmeEf9g/GHiKrcdYBtEc16lR0G6xq7uImvrYroqQ
nqaj/YRnH8dO69VHR7x3Esl8c41Mrm1m6xjIA6+Kt8+yoHI/lzWKMyMgJFSCvCq+qTHt9LAhPv2s
iENrqgBP7EdSaQVuLTUYAvHp0RqxeZ1pXx5/4Hdnu5fLDeQGIq5pUxvY3bs2Psbvc2hIyViRT9+f
sQwYVM35OIQgkaH7bpfQY0NLPVmZrgToRX8DXQAHLxfdoInEk3oYC9piI/i/jJd1w6PtQOi9fSQL
WnRWL77JZ66otOdJyWFj5V9kWqZ6L+segyQAj2dnEDTTCwBHbysGDBCDCW76VMekFKQ04ndolOLD
BG7XZgNpZqLv3GUzqe7Oythhz1SzQulTOJzNoRH9g8b6pwunUI0l6sMUIqx+V6/BBsUbUMSTn8cb
vnFBogzXFiibnSXUyUbKMXS4dpZRyLFuem12BLbwZ6ePhvTR3O/3plzRdG41k+yxO/WhqIe6/fz3
1NwXOSSn2XvQhV5Jij922dYzQXYTlh3r8o/0xBMe6QKZvGSUmdlL5JLlinJm4U3gLW5hbSi7m1GG
QFdxQZ8PK8nEm9+kdd8Ob7dIdtT14ijP8k17duN+TFZBSQ/Wx4OJMdIrvevo3UxphBGxi/dKv+q+
2E311J7kVMSmUowoFjPEG1htJ01SebsHJWMbHHS6yM1Db0s6yMwfDkcNGscd6H7P64zKOjs+rXfb
9ENGgs0XnqMHPYiBpKBtlEVOl2736esEz3SfhxV6wCle4STdqdCzED05/cGtygq7EsCBUhweknLm
bHzmNWWllc3zK5ErrAD1t2N151mfVX2bK3mj7vvvXVSVP5ltY6iGQ5Weu7cMzyvMQp2Nlgz+dyr8
0e5YnsuPhlF2cEDNN4pcbwuYIB9t1pVEl5c1d6jt9jAPFd6WGgnTU/ZXQPvYdjnBX7H0RYLQJUPL
166nniHdQVn0Q2Q5WfuDXOEGKzAKTQygHpF1NVt3kY8hyBDkaJrikXkrCl5YiRGJlCu56IC7xv+4
OZRNnws7jZ84i2QUV8LFIt4d1oQrJVCaIlNSdm6SXi9AJyTRdpMjhOvFlwHzwxg7GDdbw/r/fuoW
z7FylJ8m3tAbisM8vgLgZcVeWu6pzRJbZ2cm4nAoyP8gdlHMm5ExIWZ1fQQENNW9iP0Jdg26rJb2
niQKbJ0BOoGdMRAcnQ+IxdBMhGVMUDQfnE76HhfQPjDW9D7cks+xuvuU+HLd77L/OJzpZDzXAqV6
G4OJYYz1monW1U/lYKaCjwoWxCYx2q/IKZm3sQ1yUcQQyezoM9EcmNRGCLURNESUaiUrUZsE7ZA+
RyfEpDayWAemALHzn+qkjKqFSB373YYRP9cy1VI6Y9R7SCUezs0odWYNoW8TVrIp63NvAoAk2TRj
kX10RA537BINfNFxMNT/uOBVSqSqVcY9B1ZRCJxr+Pm3BuoibVM5qgShEkWY0r5+b8flZC5Qkub3
NBKnJZDPLbB3owFJjGUbyu/dJQOALghnFoTheBa8DBeiM8fu5MMwroXBhqvFcXpImfAUraetaI79
nWj3iZzvfdAVnel2ZN7f/DMY4et3Y72PTJNtcEU9fvwKWhOAwugAdUMx7ggqBTLfs1/NMDO5yFbA
Rz8aN6mons6MSG+5Cqf9JmXyvBid2VXt+CyNyoiEc5vIJM0U35Lmo1Z/Lyvy/TVLsVW5J/7+nIG/
zuJEyMcmo+Rs7qHRvqUZ9LElrxWPSa43rbhOn/xF8lvPFEbojkdKcz16bxAdV7gqSlq84y7c6QFe
PTkzottnh/kUOqEt9fRp4XnXr31qdoXRBlqIRwkdYGaSXmGaHpJLxQWodWesn6i89VKvmgsXa/I0
KaFHQnNeKItWr7NbgPqriyiTFEh/YtNzXBqWD1GZseTNOI98PbEWdZW89l3zMR3dJU5S6HTBUDWH
F+Kc/HSxjkRpaSj4Gr9fHUFI5sjFTw+RzibiUjBcTNnb5EK8b3Kc5lUmAnTiqHepdRXt+TTa6fSw
e0StUJkbe1Er8tug0aaYXiu8hH4Ee6lr9mV9ppSCm0SgmWIAgeg0yRoAZTM65NvWYUFnwhgX+78Y
Xy5+dfu7r1nhWdzW8zkYPohfVP7fLFGOFlxoh0rwcyLSkFPrkC3KHlynYVZppVrU2KNhL1E0BoPz
M7HTBOalCZmN6wErSRRgeVAoCd2SnY1HBoo7X6gekHVX01SKUsYSpIdPTPNjAHR/JSRaPajdhO3k
NwvKKvSi9Or6P7w74Eq9hBxPvwitAAJeNvLcrjGsRyp4kEVQhhVegMreivhHZMoIuSTYC+ub/Xav
5brYZ2cyuTpAWdxo6D8LtIfsksijjM4SiOq73cBj6ekcuvCr+HTIsJOQ+dZpZRXb2rEuOPIAlsmV
AXSGL+hYGFGt8jzXxshG68ZTvJ/qDlnRRW6J5kMPfOnA7sEqRIvVmtFR0UkO+4AIMYo7WKtu3iL8
1RmzwvqniTkJvfwktLYV0f1xUVHAjWJn+hAb1AMnd90g9R1dE4xTtdq5NzpkijUVUQ94z8JeovTd
52WQS0dRsuqaOY6dhOasTmPScy2C/+7XaRPUDqm6WGfRFhM+NyZj/KA3WsO4Qz1LpTOKtum+zF1Y
GiDHuBduuMwE8Syv8N1GrfvwT8OFc3Ikdev74VPcnas4hlmkEko3rK9v/p+kOT3wtLp2jqIn6aVq
Txup6+lPJ7SvLYGiX7Nlmr4v3yPA2mgQHVlUZ9lKAJSVJHj9vllrT+aKtoRjIVvnrM2nFfpY8XT4
MKcWC4Ootgm/KZG7hcXLcxvvg5ODu4uvw5V7XAG1vzEqpINYTkzOLujqz6Z3GOmkWlVpvz2lnu0+
Cf2iacY3RKtA7FI3jjjyqUOtqF4/tEq9thpaI1xgDRIVlCsXjSmzOn02EVDZ2d9zaUW32rFy7MLV
lEkzM6q32Ujs4A808pikotzZJ3aKMB3OUfbTqxAtOum+4KQTvTQtOqJvdMQ+lZ2TwMczU3q9VD5/
VGl/SsIktYqloyI5Zi1zVA58vo4CexG946YH411gD8Mjag2IksNQs5+9SGbTeofaKe3DiLsgDXsQ
7mJacdpTI2MGiRt51Oow2/laGfWLr484jSUkaOfSl9bSDI163Djg6uyQdi3ukr18VQqfFkkiGm3Y
FJguDFDee5h2GQnfbg+PKsj+jQmyHHBpT/fnnPyyK/ot3M26sxbjiQuOwIjk9bU23hsI0F/bEzy4
g6B0/6m2f2S4COZJCXBx5oYc51njfk6bjAlsJ5UHUF5atO1RDuUY0qwHBa3w4pvy6QY5aGfIwJzA
V5yIzXOQeM7zMgJbFCgZhM9SaxdnJ9qbSiEt8JOTS9LUC1I2AmlB6gn12cuxrDsBRIEwHUTLRpF4
dbBcpaPZuyWKWu5ul6iTy8ovjd/igkCtbFSk+UeTw5OeCwPEvEr9uWE9kzwP3fi1FzPdbxBofjri
ZY3mieYnDBrcZoDvLH0v2luivmDxkfzaBbb5J1QHdVGxCAYWJVnuxdqk5V7hZT8/ZS+o3ixNrvDw
x8xVASMN+uCcrGjKAE+quSk56Hv4PIUbo26yah9nMoogkEOZ+CcSDQkne6R0GU6yQJxhkIbZCIxt
0LX47GID+TUer41kQF1XNHyfeYztYUw8xjUY/aN8+21VMgosC3olkYGkSFU552Y7lxb0k6FK2umx
7pWvGS3hnflOsNDq/C0XWsgoDN0+2VxDnULvxZj63wRLcV3kAdnCJq6WNpLD5sBjTT0I0Ih5ENkD
isAs58GBNelENh+vQuKMmSOfgtoS/C8Z1dl2F+EJVVOTO95O15suFDn3bZzOI+OKivkLVNxht4al
D4Up7R/qBzg/HckYw7CjpF19UMbJbCENx8G+fAuHAXQS2kCOjphTddQpYXx238iLy9Rf5mwmWP/D
LUDZup0NW22NHQLG3PF2R24snHBjfbXp2tBF/YhL89yMF1CRRsmdgjV9imLIAyctL3Q2XLpUnzk5
rQ3dtl7R1NSf8sakvJwf84Ir3bEl0TNmR1JzH7kIYSkllDv3KfLDPT5OHtHy7UhzGXW5LwZg4MTB
1F6bBrQhZHfvBT7LK7h1rAtc5XeTQLGJD7YA30bi/q4lJOJVVBpoqikzWT5K+VhaCjdsXdGYNlBA
fPlx/FpEBTG/qqgGAGZWbgOMrnZBec9/SCibKDQHdDNd63XUWpd4jNy8mKrRMcwWg5lGKgvROmvI
G4pL2IZ4vMgxCNYabiwckQTkutECBQIFyeTSFCRCq51yf5vhOl1r0as+kwrITQ2CaSgG2UjGrje2
+R8iUvRHqEWq6R7wteE/3HEb9CfeksHUNlLP4vA3Gzw51T8yP/nCPZQwNcLzP8O3ZlY08IyqODjU
21yd34WXAdgOqStS/ec2Sr72b4qYdcgRzZNcloCnnLc5AUW1TYC1JXGCG1iYn2b8VCHYkXr8pDab
TxAhpU8AKGgxQgH+X60SIax/Dbb0/k0xYYDyhEp4c9CsJCRRATxKO6LPeKT/5/plnja7cD+ggecn
AAMuyDy7zCYiYHjyZDhlAZUyBTQ5t21k2V5XNzDodJ0cG0X2blTYxko482kcrLQ1JifTFE6Lrj2s
u/KCSKasRp7ackaPtm0szNF6uwbJx9QWeJLCb8PCZ5zFqdbPQDiX8Bhmg9St/ryE2bN8csephdti
sWZERuVHdkShqle4STxE0F7x7kfee3GewEA2zj59j9w+e7rQUTi3rvRq1nNIA6fQxttv1ZhGpWJ8
vfuDGnzL8eCUuDXpSj3c83IzrWce2yjQnVskdDySU/AJDGH323rqct2MP0P6lHiWmQj3IZTb5lqC
4SW4s8q62m2HXENTuzXRYuEZlB2+4x5Cu8NCrEVQGTe1tn7eX7P+01adkd8qcW0QvA4OmrMoIJCU
z5QPHpwMw4loaz0+2t20YbsmppTUeJO9/u7N+SYhYTVlkOGZ3u20Q/tehVOnYFIh4SpWL99xNTxM
uXb/NE8cdC4P9Su2c/MkVa5mxZn5ItObx0fzlcsMOtN49xvdSFWATbNlSViUcOq//bfF+fSrJD/s
HvDZTY+jwI47vLkHx4siQWQS5eWWRxrM12523rvpTff3rHchnAME+O+S0xnPGS1TPs5TavyQfKmP
0enc5lfOJ7B2wAE4d6SwVRqEnpGaDgeg7o+LfodmNgbaYlFmIbcw47t9kjjalzGoaOTlbRBJvc4C
lqaF7yGrJF1raH6rvVT0xl2g2w7iK3W/2s9n/e1pA+ZbvF6ue6dXyO5pWRjZyMbl6IG1Si5g5hTo
h6jOge3JCXv3w/O68tNkFGHswNiX/Y79aZqe8u47nJNvVYqdwpL53hGzXqsMhXRw0QqL7hNvatBB
TmIeMTGtUR08G0eXIbvkT6Z/Wd2Xr4gQQD0bhtapffrxSnbqUbBLdg0cNkdvCKO0enEHXwoMmENN
4pTMCcxkQKFLzzxmPM9MhYHt4LDr8GaYhjWqEI5KctvpXLwSaRFZnsM5atRpzlu/sVJmbGo6O2/0
m7fq55RtsasR3AIdPQnoMpBqF/xfbRhwkBiO8+j+QAojhpc8jX5mMhHYwhFEiUvlI6iJkVp/cnQH
8ZiO7u1dMZwUr19WB0VbEAReHMglU3SYMJzpMsfpGpt5mHdlSp1k/tIJPWsT8nQV/BuSgY048vE/
j/pq3WP1Uai4Xs2QpiURrNwM+RKsGLugp/1V88A0qZJ/v/DIjZ+EfT/fC1UYbuBPsHFO0idoVWt3
hIosk7j+oV/oC2amKD8wdsTBCdUPZ2nF6LOoMXnJiGe1M9h9GhLlOml5UNlO/sJfRGEikxYT/k7m
Ym1kM1XX72eJ9ET9gUwrJSpgi87mxOgdf2Q+pCepkjaJpj92ebBEW/U5ipKpJxmoBfUlUEIDkjXq
eEl5JXQKk9EZvLSsH0RkoRBRtA9SzBK/bWLOrU1v10OTCGZlOf0cIEd7v4kOT0rdAMNFrJ/vHwyZ
wZPcAYHJQ3FYFF1j+sTEueapA8rkdKJjZQYTOTigwwmTuMRhLb6f8TsK8NQGSdS+lSGE5N8yj8Am
j3HA5DwNEn6VgcTvAYrT4pnBHQup/3h2XETrVUcKvJjZtktArFJK/IflkTCQ1oTD+Z9QThTnj+Qf
aBUtQoLNQYWExnyiD2tsxHQyWH938yOJl0ouUAb0nz3/bFPKVX/8eNAVpcV34r2ExsnLtJaU4HiV
e+4SCipHvD12b2/qmr6+WCkDX3XZbLLB7JIsmijwK9IzKh37gnt1Kr0ZiC5THwcNZOz/o7YazH56
p5FMjkHRSUhK3DsYGFkwFcI5CkjuG4rHzCd+CJxhSRr/judYYVT+up+fy930SU2CJKXifFriAqxT
2U1KHvdMXxikHSD4R130hYe2Go8ePkq6siKwb+KHfK7nAzOwMoQ5WymrVXBAte+R3UL2nMpYGX7J
Ppr0m1oUrfvf1EZ8i1mqPadUcC+oJ3lAF2fuw5xw5EF3LOKLR3KGT2LcgRWYOFeD8wQnL3euDI2C
BURNTpC4XlzIzPqv39OCE/yhDiLvZDZvR6tXKRf36ABp8pEJho8ir28vlLhdnhJ+1ZpKniBs5rB3
A5+USMEJcM87ELUHvUBXv+7tAwTpsqENLkLAiXyP9xQtVeIFqalT2fjJm82/euLEjnMdp7SFgGJF
TgrjoPYrl4GKDsMbxqr8/11pbLhiGgFGTHJJsc2m/uIMRcU4iHlfanONngEsAgrT80uOCsVnb3ve
VELbKv0clcS5G6rfMbMunh3WG490YB9M6gi8w1yqwYvcYxX3hvSmxFk5uwnWpAA51ozd1x91mtyb
QSvX9efjad6zypAIpiQ+ory/QTsbr1iyv+lmgXsedyaVyCsukPVTJBe9iFWwLqzhXMc2h7Q/QiK1
ULkZ6GCss4OcFsb8kejwBecxpWHLizerJf9olk+bbNYKGjd7ycleBw/g/pA1CF7kXZOq1rs+GF1I
Zm6Lh95NhMFYqLQ3n2CC8iXtgcvf0/JyoxhKpiUSTGIFvovhfrnGbyzoN15HiuvvIhpq01soSaMM
SV9bxrBssRR5nmBVYYMkG47gA9YmK007n41DmDO82FCVyuAUASQqNGJVl7OTWkUv5FaxMM4ivzMg
EzuKC4uAd+gMgf73qh2+4r4A+BeVmpv3AeuhYkLhjM/+gjbQDk7RbWOYzcR6frBLgb18L8g1Eybz
z/7JwA024Zvj+JAMsE61jZR2RE5vclCQRG1VmbmQyU4togX2re8dxjRbzEb88yBGICQu2lTXMWmx
ZqNBy3ThbB07KTAnO/Q6bM1Qn4hyUxXKfESvCSCfXIr5gAUh92zH1bF3DUMX34P3ERrJOkaIDL99
re4ug00R6GF3CPFzF+v4WR7rBZCs/Bc5+rhoGB8RQVTpcUMTO81lo1Dj5h+Ff9PJ8Z5EStqR+PfD
M9O3/hpC9MEoC25g93GMmZMVWuPrtX49AHdcb73Csmt8epNIPDctYU2Ni7D3yNmNS6D+J3U63/wA
TpAvLii3D8h7VW5bSiW0qgTQ/miYoyyUxszwS55bpA8T0VKfik7ylLf/tKO9YHwoufnYYKpzlbYe
s406VxqskzxoMj/FF46BhfObckKduC6DPqADwAnZjQ/RMIj3A7ucOpGJMsUUhQi1m1AGbGC58ECZ
IO5HeDgexgfP79EstMUWcWTQTQXLky08NlNPJGP+2lrT41C69NZWRULhe4OnfYh15sC8xY+x3aHU
DE0cUmiOM9wo+oro6y7lVTzBqcjTvPe9a3YIaGpHLQcl+vjzBXjr9JxZYmXlvOyYbAQB7cFZEXDH
TOAbWoPeRGmjeY+fLg/T8OGprE4pladOqz0VYRiM/wxxcg0RDnsnAGwvZgD2QJ+5M/3wcOfS/am4
DpUGx2UFmb65cpW/+i0Axy/lBHmoNr4YLz5vMHPov/NsBHC0m7TjUy4vffL02p5ur6fGi/AUTmtN
ddiEqx6Y4+Pc1ywzM0fsk0UeA3K8iJI/nyBD0ftdOzCGNWDvkXzyNwQSLtnIpbpqbUu+J9rBGvMe
2/UlJYD2VUUzpqgjq18PZLVbWeqUkQvxb/ajqYmv1sNcmqVPXBps5xNcV/afsna4wv06kbzAKpi6
jtQPH3Rd1RiKzS/uOcQPIPlcNF7kG8mXKzy7Dy097m9XFcjIZ1OhiYy+NWo3Tb0WOMeAvPADrgES
lyDZiFwSkucwFFZIWrU0vrg8xFw5IRrmMWsg+gbOLUjSZ0MTsJUL7S71rWwIHwQBhWsaYWpMt8iJ
4aj6BYTg3tqUn6u2tzq9EFnRwaZyA7jDcyVop7SxF4ZNtdkls87YwDhQE1uNg1tpQy2aRdg3ZDE9
mI1+Rx2VV4B+YN3l4Y/VeKIGyYpduIKc7eO5D6m5rdC8AUQs0BfK2lnN6ZseujrLV+mziAbq7Luq
gPD0lNNPf6o54w+I5KQHWNEkXHjf/iK+Z2sBjj8fuZIQ8ph4AX5wHa9z2VTecZcWfSue21w+IldH
LMSXkri5oP7AiEWf0wmFzCvO4Dt+uY5Bjz41OwCfm/nY1E8dkofLucP3ZEWuosZrfXYd8QIdygO4
r/ONuqMMdD8Q+hzDepRTntm8P6VIgwh7kwky0eco1ln4+ltd3wkk55bg7HbWa89SKvoVpP2vitaX
Y6s2hSqbinGWSvjqDniOJqMA+fQ7PzYlDmSTabI1RrLHVqvCAWrZ9gRHgzkKsUiuVlvzxIoo7f+B
pfLxAS56rnu8zUWJzBYHyOVijYWupnd1O55lYxeYSYPViyulLjqKaERAZ9QWI6lKN/syJasdkCi1
OK0OmvRMh8Gye+7xegf8rIDv/8Po31nEVSTtYLkhWhy4QHNwDNQfJTbz6iWQXHt7gIlgeAhw4ahF
9Yxbdh3AG5kmPBkx1aLkYfXT7MSrcsU0HuhRNphrNhtyrqcTKGaCyDO0e1W/uZRd+7NYIB/QCkVK
Wjuhshxzf1NQkNneFOptJbFXh8c8k7nM6vL4lrQkas5DUuxgJiZYspBaLu9+4e4UIXOImbve6+So
lkbzaPQiO5F6u0pVlvgZ42DxrbTVSNOkXPnQWFDbUGGepuX+iXB8jy/TWkFZSfvJrp0nAEvlRq3G
ZxzzWO6ZRHbuIJNDZAMH8gVgUAOutwjDrqi6BqMXWY8JKeZpynnZdT1ORS4/WvhofI6sFQUhinLG
gvyTGC1j+zv218NhLikIHDzeAixszUFxoAIlkz07JRRttgC9qkTYLkawWNMKvBxHXU9CpbvIUj3l
ZTd1WmWOyd2sayO/mNZqQWUGIa39q5jdb2BuCcMyANxydqnPY/2uj2F0rmAXeTe+TDrfjkIhvWTx
+JCpA7fvszPG8SU9VmEHkn3QRW0KvAHvbTb6RT9cWqi6AHGwgqcgQDafhEySmwq8/7HMCI+6V/Kp
7UHaX1YyYC8MwpOqv4UGHyzoeheVbBYF1kpw3K5X7DLTp5aRVg7DDxSawhU3RiPL5QZf8a9YsWD5
dYRFnQ7HCKEHYhUAezVjMjbFZW33mzLeLdDt/ujcymxGmIw+BCYGl6VS685YgQEQCK4zLZhPrf9x
7NHO7x25ERgI8S3w64o/j0dlmDjJc4kZlvYQyjWZ8OVHJUm+wb1xLPCFwJEZ5KCRlK1CHlNIWq5D
sZ7YTDBakqQYiknYuvxlAS0KhTntBEp8GtG68s4u3PerwEYdGEU3+l4UZabsGiWO2pwRp4WjXEe9
X2JLWLgQbN+REtXwauMVkRtpODbdH3eZujWEkpswEpvUC0GUWWZ73ogSFWOPf4/idWGLBM6LGUUB
i60c+6oNx0x67dwVvy228KkrRAkssYcy4boNCcL8xPVSvnsqM+587oH5m38R8gj7o/Sy4AvCk7HQ
YcDhZ46t98yZpxuxQ3QJjycEqWvEWFn21sj/S79sasMWEhGtrQOqHhjmuY9frifWtocJXr4ngXWX
tXr3eNzKe1vT9fwy8oqXcb9Qat/hq3kAhuNSsI5hCfIa/AwR0aN96rQdmhl5fYFKRJqBMFfThnJ4
qYmbu+/83+B2hPxj80HUYY2JrkhsdrJGnh/QC1a+5MTEMRXHsTbS76UhoVbRhfDJXIZ7b2+fKNWP
lt0pK/67DhDI5QvNlpnyd1Jai41fiUKC2/SnQMYKmqF/pz+wXZegFgA7xFKt8RB/2YWY51LuI1A+
RS608ABtUAgjnfF/wbYKwumEjus78NuRr7QIlV8Kyr1pTHn9i6/XeFakxT9kEDtI6Att1KAlW66+
gvHo7ayJbD3xIc4DOmMEK4u/O/ezMEAaVcDwKe9wCNJBAHQ5AunmLgsdSnZV2+GgKn1rJCbzgp4I
XqbDDDsAyJBKrUcGIq12krYIqLXZgqY0nhzi29ni5V5Cx/nbP6fI83WwFeq6xLlyGeefvvLmFr6S
xDSQwVswZNX5stxPMuAdWLwrp6Q5efOYXDQmZNOjVwUARDOG9tU65La6+B7wOJqCT3VTgWjQztcp
XvX/GrTmd+xJv8fRaCFSXvWdPgF1SyRmgDn4WxIQ0Ly2+Jd3sMxhFxKl4I5w4TUKMF8/UDAzsYs/
3lyd1sLKzsBJK/e4LNQuMUIhc3jkiqpiQfdqgaWLnJgK9D+u1ZepZwAH7F9NHoZ6CJ39Lhtak5x9
7r38YPrQNoqXwYgm6NUXdD+S+HL0fxxO6c/UpO+G8Suyhs9hloduJtViYlOANIgKVfPQux1ugfs1
DOm64BJaP1gl+lpck4YxM3AGTpHjrpGf1XmdAGFIeiFjnznVO2fi19eGTlyemegELlaXEeYPPQXd
oE4Q/EelijoGEoWTbtWhBHvMiIZFFEEvz171acLrvc1LqJexEjUCt4vc+9Vyew6AiffKzfAtGUut
nWmqiHDCrCZESXgCK57/q8FKrkgdgk0F0ke4t42KgLSMLov/BWsV36QGaQn0EOv094wFjrjfatHf
DAOQo/ANSqEMiCsgGZLMcMc58QCQGNXq+ioE5wsvttqUY903Rprs7BSJ10/367AVP0klAOho29GT
ypEcfxSzwC8X3cvctKZAXmKG5o5tv3Sr4rcPqoweB5YncS51sZyoTIjIyYw/2Y5gqqtx+eJxVpa8
G0YL9Hhx4KaZQY5dwRZM3pR8B4VPFpma8qsCQ5rltiH9P1cR4v9sUyZjLpINZ87afsh1qfbxiPs1
F8cQTr7wFX1u7DWGQOI1jxC6/kgfUJbdN2T5vwNcpwRBti7G9qRoEK18aj/Y65w6U+0yfKuF1HIw
Y3gaAWDCtD/SBsS9wRl81OUqMqeMaH93A1jG5F7hp6AeheAQEP/FSEXszt9mkU8/ImSw3hLEUHQB
9iXndhf/4kmZlkqAbeAaG4XPxAbzNDJ1FiqTYwlyxzmvGWvxXExH82m19Oewf9mHknvpxpvFvIku
7CTTK32HnBZO0tfw1O9uIh7GmvhwaWekVp5N1uYEO7X5NwJkFym5bzJGRcaiFXhVsSVdiTlw2EMM
UTergEZiVQ5msfPVg7b6+ud1UgeUHh7boBkdBZsC06eTiwezobwQdrkcjconm2KEQQEZuzpOGCHd
CadtNeoGCbn+sprOhWSFRRy2cUFNtGr/xEW4JN7c/j95zP2UclYW2LTb3E1P0/5Gv7pblWf+S3KB
rmDt/8yWHav81is9rOJzlZ1WhBaPszws5eKf+6hTpvWJZDFUTLayZe5XLX4I5Ub5P1fH3BXDhuZT
GoX50JA2CeWyWS1OZfqX6XtF86qlgpsRsdm9+QrG8jlnSlHsn9ZuNUjyWKK1CaBKaAtphomPuTTn
Fexi09IUWcloe9TvXmiP4nGa9C6qjyYM0ewN+5+gPyUlv+IxNbjxTnWNPwh8zADdoGw+z2Hnm2t6
uVwI4QF1DrrECw/4P5lXkYRlhHqddVrY5wtKC0fsNFcap+WnvW4rj+azilub9jIyU5cQ/w8HlfwN
EcHVWdRR9u4L8t+Qb4wmDMh2n5alTCx2WtQKgelE3HDwiMtrFbhPS5YHBJFuqNjHe6O0Db0Kue+c
JTDXFt3TLnmp7cAQd20oh3W3p0vuRYPWuLqHp+8YFqlaUpNYSruhX/vT1fw+E/iGpr/5O4YnEp+O
ip2qan/ZVUAeBRZ2PYOFPf8IDuo8sWIwTaITYgFD2ppWnYrxLBLy2OHhn4rpsovQI78NCqxTQi58
/PCPl+tiaxZcHrAMi/8GIohfO4MxQfdkxKhfwOY7wzQmureELNpWMuyadeBWzuOHm6fACAEBLo87
2iaKGQAIQVvCOTEwEHU8ZHDHurTDEeYvWXQtocybud8ooK7GAdrM68b8t6QKoPEv1VDtT07xzjfF
f3Ct4x12WGbkAvOg9E+F7tIk+W7fy5ChfiERIvcEp9DOyRNvqDCLPQ5WfuNV5+QpqMEXwWQeDZlV
3y6q9tlISnsefFICteicsXJZllpEBaPLhvkXMnW2vCcyai0FdqKu52Q3bWRBT0XPlvvXq0CcqA33
d0iXFTbxz3oeqeu635KUqkm8pGHwMRcPcfi0cPs5ntltEQbM31a4WC5SJYL3gyRwo7gISufdMZgW
1/fov1Sq++fjxjpy5F0kNdBkx+5EFCBmD141o+/VeYZs2ko8SBIWwfe9H/2MQa6UjAZEl5GMx32K
6g5dBYBD60qIkK3FWi606Piq6+WMYSoBU5f/07ARs8lqjDagQBqFFGUrApWV1JTMdv4535kK9/HX
L4Yo1VK1NJBEnKvM8+3bTWGHThEwTEkPhTM0eKmxP2W9BQMItELn0C/+OZA+WQv3rxRSKPFWg6lR
gSesQ2cNRq6xpWwyu9TZ+8U6qac3K3/t5zEww7mcuZ8YNh0nqQ8cNdaViwmpAGVR3W1ritqJaIQI
YF09h5ii2VjqN5fuTD1DkMvl21lHP/ahkhEoc4UKgODnDQA5OUfFDdLKT9hwCiLd550qhcKHyF6S
HCZGGl/aNE/is4kftKYeZF/FTUURw7S60XYtdYncQOaTJy0EgbjYB+npajuAreRmWqA6TTz2mPLB
8+ElnAseNCAXg4bN/nWWw8FvT/7ZRX8ymfHBp9eQgrfZvNUqDLqJnSevaTWFLXp/jb7bF+Z2dISX
ZC2kwtHScdjZwV7PJu9RKW2NLs+Lfc1YJvpuUP0l9A+A7Q5rCAYJwj/oIYl3beOxMePjUqHjcFZK
K3W6u2+tgtl3sYFSKJTJoU7RPildupsgr8WwJtuV/7Ih6RAycOpSuAD2WiuOq0P8yTmi2LcMpR1F
JMEqQwl35H3IZgeqUuftyCxCY+7t5Xh+/g9RUaeuMeuyTXO/MJZeRDo7PoaZulxp5pfkmA/qVV2W
I5gI1xs5ssvFnD5OCtpa/a8d87fbglEhPUAIG2+Zx/vz0fK4Ulr5bCBoi9tmKokpQY8xlEy2vmKV
E8DB3wMbhwxAE2KijmaYJztCJEVRD90iFAIW6oA4eewDHWS2HwP2xr5RMJzBBcJoalatUo8VDiaR
y8JdBP2Cx5m10eEDaiPXIOgKwwW4Iq5ZN7o7S7aFv2v44STYvZKVoPoAN7MjDP+BgCVe0ddrXSL3
ae/D3AdSFI3/x/qT2lwXp0WQJjG0ycuWqeLNWobqn2htRBwTrSRLV393T3806YThn3aBqiBNy5MN
fvX08Wp06VsxCioeByd8/bvE6XL6MiHHxDU5ma84L2gh7t4S2wjczxlMqyXNbx4Sgl4iOsW4TmMs
pAqwBWNyOVOX2T7GDTsOl09mu7kPLb7X8HO/Qj4BFZY6R1kLDXKDac2FZWmHZiEtOaS4iAse8h/2
nPk95ATxlIo3jM3dvAXChiq8BAVRpd784gb+HrOhPzfKGk8eADpwGxAmNcr3WgLqClLyKygwf9ss
xDzAHjXz+HAOI+8bWzhAEl//DhQLzKvijQ9e3zRPCCbj7ONqlChVU39I8e45z38MmurCdDMAvk7f
LYMQgbiTcvUKaMoCo4s0dHZzz6ZdtCf3GsDX5T9pBQ1DTC+YlY4Dj95a0PLz33n7OpnSdcm9wIb8
ej/hk6NyKNbj7syfndOkleLYr7PUcqoIVH4S7aTX2QUgtu4AHh44ddKbvAxiZkAhZ27aGlsXqMGH
+43x/GiuTk7qIns9x7/iceLity6TXliX3AygDurJpab+BUKCSi1iQrv9nQQcRbGivRi22wC//NkP
ouOkvykZ7DCV8an8BFZ5fWNnNFFhms4V/v+zq0uKZguS9piG/V9r8s0PUJBKvBvn4njEJfZ7iR5G
6E7hGrAKlWV0FnFichAs+29SQq37E/CiPo+mogZJoMWKzjtRT0QIXnK7J05BPTFO63BH10/IZYfn
BX5ZOTQ5KN9VDI1hZGuGaJSDJlFbouK0uFcard3HF8/99NUy3ehghnMjdRTLhpyPMSSl6orzxJR8
fWpmbjFzaeXhmuC+jeHw53e0IlXAuXo12vUVCSQRRNCIOb1knZZFeQ1LbG7flZ8/XnBZOfQVIFzP
mrldhtSSZVcjwZqajCI2trKHyyH6nTPYY6oyTl/8TvluDWxxEGZtr/R6IGg9BG07m8QI/cQpm0sM
Aevj0E1hi5yfsvk7UvDV2mIpXml7Hi1Cpe1imcicMppFEzybMrLAm01e84sky+PUWo/6aoKpWRyf
Jhr+lEV3X6lbaZA+C1U9CtY1/s9gqNtpXQW2f2Tmp9ulpeKhvndeduA+udslxv9BRG3rULgWw1CU
7Zyxcb2KQAR6v/pwzAGbtVvzQRzwFdKNJDnI6+wZ4PerXzz4zKEUUyF1P30y6M0qT8Y0HVpzESFd
aFTa2HA+UrqIOs2XLQ6yPOs1bzxllbdc3Vy/ryxjVDGhxQWZDK2eVzN2nW56A4UB2h9/FrBptXsN
fD1rmZ+ZYWE7WHg1uX/1q+Q8OWZ7UMXPB43iw5mCF0Zc3h888fuuRoB8VpTBvMueL/gLaQdV2fK+
AVPdYZh59Vwlq2a7cS4UUzM9TxOrSx2eVindSQ9DmCg2XHr86bI/wpKo63lqQeA3DPBClNF9drDj
wwEZL+qZP9UPoUTWmx1shgpoT3GWiQWE40i49mwxVqd5zOKO3yHuofqUs0KHCY6PiLKTtP7FEcy8
5UggCFDW1H6wrt4/9EISi0PNae+DRMGqdOuVt/ngm8pHTbCjM4NmXa0oRVKPrede8bYOvFzUONi8
nO7DmheOuHP9V1B06buDePlNB2e1hI7JkuZmL9JMQH66Lr0HK1VUO0eXd9C4ZcNbY11Bs2k4mSxQ
Cga1/Cl5hk53xSMy783Yq+2+lJbxRNE333GHQj1E2KXYtoIKvAT03oGqddlzjRLnfH6rRmvbpUrE
GeulAz6AWsiTjLSgUTtDCQSIWSfJCp5JpByWWUd5S6s4sDFIx2jmnFQDSgaXfo3ogccsdBysqsF/
sd9o/bS9nXcnO0tGERQU8noFMnF18mZ8K8/P0MKYcFQG+YnZKqscIPcghNol9PQQFU7fWnqmGioj
82om4iiPx89ol/ZRNG79OSMQKky1u4QgYoSCT4eDwvq7KXRaxIGqN12ZiRikgxvukZer9h0t0NDJ
N8ZA5ndijgSvrQoN6JqZcuI/EkbHLO8T8lxr8WXpGVQ70T/o++tgt7qPA3SmiN5Pk9jKc0+n+FDH
alJAuNzmI9Ci4jLp7vclMeKirAFrtPHrGEKgl2OzvEOCufZVyxNYrWpmxx1QXmNLWXWKkCPyeXb5
BKrcj99/ow0jGtFEqFMB/Pq4BijhQLj0f7LBPHkG+GlFxUUFPdHOpdL3fXGIuBmWorAc4Qd5vj0G
pvthdtS4b2+uuuoLWisY/ANh663nl6M07pR/8+PGe7LA3MVo9LX+wnWm2m2dKgOB5FwEiXEEbX9P
sbjKcgwuTXhtX6pGlLnCiSRgicXE5uw9JX4A88PBsi+Oib/hpl2LzgvAjjSCaPCx/VrN2zibDHIW
bccOWlJsxQLtgsUPPPHx91TQ0ciXVRmvjiLz4hBtzlZ73uS50+pke7dceRHYZkgw0Q/fSrfbJeDU
s/Go8c0q6EB2ANynBiEibYXHxNEei5hc2VulMQW114fDjWO6YQrioyLodbMp9QK8a/cCnLo5sXUd
QtGF3DMJPXEweEKB6gh7uLqsUPjqpJW7hxuLgPp37CucCv0e0ZX+Qccf++0RjATU1lA6UllMTt86
0t50vyrOce50Dw7+KIVF8iM0OifEzuWr+1mfmKAB7ImxJXFV37moy23dteYuF8Mz/bGZ/NEp3T1W
psRtXyXb08YWGnbRAfGrhKPL34uH0E1K4RuWUhSxdUR7eIboEGbQ1S6z7uAS0YWB5Q0q/DdnGYTR
SuG8pU62eX47VHoZwBjYx1+HOk1QiIDzc2Em4opuRYE0IEWIrLHG+I3sA9f/kBG7P7ls3TYFdQgF
KcfmwTnAO0xGR90Of04XPwGGUiularDABf5qp2Swai3gMiH4gH8OWABANyvem25ankkIXGqMfsj8
mffsY9SP4d3vC9rQgnxwyQYAKNp8opDy31KjJL2oCMUjew0vsNL6/GkTjdE9sn1aHIPuPqVHkaaI
P/yx8EqLk8KRSBXw0nOVxfitqRno9+RtM4k73cGh0SVowDYJO5sx2vMiyDxqpdhrcfrBstWUXq9a
pG5WVvNqGS+Eh8I1hYfgg6O+qN3DimSfNVT9QSc9++xsKE8bK6HbyYKwVpnLnKgWxsxEeDC1b+5q
3aCWTElpbnLcccXc+8AwmRpltzqBiqIcihkAtTFQn3jZE8unG432a5jcAJM8t1ngVtnSh/+pmc/R
6t5qQCB6MfQMBsVLHrru0wsfWJQ0Tj/jksFNyEgcvXHsp8p8y9zW9poH87c7fB7ePy2chrNB7oSz
WUePfQhRFMm2H5r9YwXHss3Jv66++xFZs9Zg9IVd1GNoQ5gNR994vMvSvZgJwFxd++0OhjcLIE2b
6vfm8S0K4WbFt2rVH2ceKHdnAWLYTnmBk07t3OWBYDXAXwAdKR0Q9vYsJBeMXiCaLtZz3LHGgaQe
tPZeBj4h5/tn3oxRUNGUEL04oRyggVkoHYNq3VydPryS3Gu4lxl4GTClZCpapZWhVNimIFgRxHLE
fiWsl3g+CAX3bYW/Ce8UA3HE+tNGG5Nas3LopnBI0witV93/CB2OZPjFk+ihQXZEgdBIpgPr0MH1
tbwqTR3gN/VOAi+Fbrz29RYuEv88Nvbv0Rh/lh+eF5XFVuj15JtpSEkZo8G8nHHqj3b9rN5MuKlh
X4cVGYHDdsHONxkKmHm/pc3nL3jV8g7x2snlthKecYANkiRBxvobH29B/ugpC/ZhsmGipqA+gZot
BzTGz6KucEYTIH+ifAWESkCfOYKK/boI3h1xU3EnyGmp94qd9EMIhJ+XoJoiKKGPy5WJPmrUOgG+
h2qf7CzuyFV02isa9Vnvy0Uf0THv6BZq4vjU37zeNlXVfMkSAJ3A3n3KeFKFhtuXw0NL/ZLZ8OxK
5ChQf9Uoc5davDlUzg11t8RZrLnXyAiu4BS+X+ucOvEgL3XhSKLOh46B+2TDQuSAHWpkDLxnToJM
ZhwQosSDEGgy+VOcK89jkW62BqbfzHhTELw1k1oOLDpnmsMdMlGBBtCF0hMJxLnd3T6Qz+UeNk1d
Ifw2bMFfLPUp24qqFipYrJigbO+BrjfdvqcP/xdlK776ctDuA36/XWVq3w+3vnbYW2sVQ4vtR0cV
38g2QDjnqBN0N9RoxeYf4s0kAkj8QdG+As8Zwft5NldBYu0Qmc80M5uNZJ6XmLeZIp7pZBU1S1UO
rXKYrFSA45Y847ftRaDK3AWn79/PRfGWbNw7XpoFgrKnTq4XybX7dAGfKLeMjGhfX6u01PeEkZwY
/Nk/NstMQXz64dFcMk3+25QolhKCQMVC8h2ory3vlsqy4NSKS+9BcEr3yKj+1VNzODGFv+LkTDN/
vWbyEcFZkD61p7nDvQ04nHq140rkTVvCVP5/6L40cIzuEOeXEvNRfzJstWNUFCmjz31PJMPZkyMY
KdReJKPwUaRqJPIGSAqAItjk3hf4evuciAqO7i2/4mfV1vMyGi4aKfeYWaeiX+ozkH0B0Pjbt2kX
/e8IDMueqy7ndGatY0fk1gNAM0ze/bTUe68sTSoHzy6JlbGUh+Y/VMRfjwcCQW/bbXOp9loIotOf
0FBzx+rJg5EjZWSRP9ZKHPt5W6gP76NxPk1FAEtGow8LJlhh88nO/vz/qQAApR6fsBY6GrPIZPWC
90t6jdbisjj0WiM2wMPrrryloC2IOofNhoVzJmG5n/0R1tZ+9jPavJISLC1KuLIrLvb5jxnfYf5W
4V23y1oYEyge/z22O6iUCi+UaNm+pC0etdrIRvgu/FlBxZ5n/i7JM/d+3fjXRXEdRhdcVdXwcdsZ
AaHeNS1tDJySZj3Ro4gANCJ4+GdjC7QorWa4Xq2l0tfweHU4p2s7aRVp5QPyFR3ofsva/74TSJJw
22O0Ev0SdrTg6UxG1GvbQ9DKXc1MQry3ZAkTBrqTmumkntMTv2uoNtvCPN/cd6TiFXDYjD5TcPFC
lMRw29d0Cw+ICHjAPw/z69f7OyvIpOu7EAeHYyKorzc5qv3haqlv9hgrxcsf5RwbahCIyID3wnV7
ohY8FmZoygQsSWi/73qFEB2LV3JwLJlEkXZX64P0YJwIl2ZE8ZySd4QYEu5/iBXQ9r3kshtqITxO
eG/OqC5whPfugdNg6itmYNUPHQ3QZqSraUjCqae9aSmFDDJ9YFHCO1CxU0p4B+yZiRzpznFh9E9F
WBHkMtl8PruEqCJIiC701gotQpz1BpSHn6JCJ5e3PAS4kBu24UfmqxFOQ22wLXDWFY41HJGmqU3F
LbqqRc+HFZWbyRxr2grCeFArI2zYYE+7Vw44/9nSEpkkx5HwxXvIdUSsQgVzRnLSmW6RLUr1hdT1
Afh+AVcYXR+1G/hs0oCLUxJXhPynYnHP4uE6zgfajAqi1EKbotPCdzyxWc6hucrd396Y/x4rtfPt
qxvLadrYmCiu3NPu6kXcRlo8/a7mRI51npY7Er5X5S5/WDkWg8BDZvyWzaPWVB2yThaoyOQfar8q
3LNuaR6VRQmog2PPpoEDEsv0IpBy9oyFGMcPi2emkRdu8TtVYgHnacN/+FCEQvwJdrp5m1N75gsm
2Hzd08CUQo3hEusCXrBCzBdEdP9ze3Sp8BhKYo0UIZ2Xgr1jW8fvaYSO+J4o3L7iQBKtqPgrX74q
xDdAv+tYpP2Xn95xCKWWPkTIUs6SJER821EwM7aEyK7Zl1G8Gc4S2IFLTVA+0wquFw/kSyPvvGz7
43nc3LK/cadlB48qH2RhTvP+tVzb84F16IsqbubFIUFfa+JC4Zhax1NvUYei1+8Q8imcAr9w++1K
kj6hRAYaYboUOtBES0ROfI73n+PLagRA45uusZoDww1g7DuQvirriuGXqE64R2VvQDktU0NWKzyi
+wcaemUYfkdZpDlq9GIR+J9W5EQWHVPZPMJMFgvooqnUBJV2VnEMlnCT6qVt94wZyEbKiz9+2uXh
EV1jxjoxkxXnVrQDHSG0D67y4svcEXqE8bP0//Vi5Nqn9sCuIx/2md8eNLH5nfJFhwIviX29dls6
Ve4f0ccap7+ozZG+9BdqX5geWUGAnLIUqRy3eEdGqXgSC69dmdsDsA+buExakjUb1di2mCQwL6kX
xjE1b7YlezG0UvxPF98xBK9TL8+TM9iq8AAwh7KGaMuYl1mjCussgraZ6ALn8JNf8V2L/DZzLtCO
p/pA05G8v1AOqo5xJCpuB4enpGxExEaxsnHcVIrDG9PvyN0qPbqFiScIvQRy1ma0+UMj1+loKD3r
Q2Mv8UYjb7m8ErNpGND1OzxLKNO7fkdPJ0PQTbhhAOR5I4/P76F9+mKZbr1qKoQt97UP/8Mvde4B
DwBjdvaJpg21jRo616eGlXfFhrb2FQM8Js8euwLqDe0PiResFew7wse2XQJMSyBfsJFy6M2EAzAn
MWMQy5PJQF2z3xqIsEUENR4lrBD8E4CMhR8NrJ75v98t0bakzpd/jxtSvEUyuLNJ8Vp1QT30UCd4
Zcv+dRRGAld0zFJkDkZ1oop5CqG/UNPIRqCV3IuM2LMiBveFfA20spaagrAquXvthXaTvXIQcfT8
b1ESnlLZA42rpm4MG9oixeLKZ5R88bkRbO7YjPVbWt9eV1cGVGFOBDCSEzyU2vbr++ZIoHTpOwFF
7ixJJmQwoQTQP7pKcH/7RBCjF+rHB5TGLDlwxXkk2ZtQHJCXIAUP99qC5QucS/J79/9TiRvYEyxg
DE0ezkURjr0jXjTJJchRilUcS4czfH+bNtdTL142twLVP7oLu9Cy+CAmUa0A5VcLDmfRge/qACkg
S76VUIZLTe7atI9hVIs8ZoBEVvILkhenhIogk6dpMIn2w9WIGA1ywwEoZKUUiOEV/2QIQRBSqT7r
gtoQM+KGQqRZMzGQN02HTTah6SruNFuefvOlIjqgncj2oFQ7vofLUzl4mXitnDTJPc5M/jSN9JOx
lPPnlQGjKzYY9RkcT+VsJD5h8JUZNDVm63jXf6LJ1OP5FLn3FKmfIU5GWv0ZAEsnCCWTmpK5AIIj
IgwHNxAl3WCuLffWC1zMIhdX6LQQVCYYR3Z3ZrAjAlR9ZRsW1X0z8m6sHElVFPLBukeSnHnCD6E7
UMKd55UKJnhcVG2A84aWjYG55XH3xPc92Y6VBj9lcNLZxhsppx54Pw7MH37HCKtsPRW7w1/y67E0
iFGXE9qJB/vjAoOgRvcc3vbARm3f5sbxcE94eYCjcyRN9d3u6aB2qI/hyTSqxMPlyvkeiCOeQc5D
I5fQRUV0o1gSl2u8j3GbGdR6XnCp0P4i0RO20v1z0yHT+QasxxFQeiObOEB1y1/NDXMxL8/0IMKQ
948s4hVpt/N/qDgWB6phI7qrl4VRBThh+agS1tz9Z9REuvU+xbHLOsPHm85FhrVUwLHN7XdvLj1Y
kTikegljGIqBX0LlkhzzA2ZLxebELOr2KwYKHLdPvo/O7K1jfSTvXAXQcxVynSVnhp5/eCzrgnS2
QRwnJNBsiZjWLxAXYl20yC4NOuxRFyfefC3CS6Z8u/V3V60L3BY1/1KTnmcEqf/MeC+1tODgP33b
3fSyc7k9dW0mxlWs1UuTBoRHtxjfEqpJi7D4UYazGcxSNGxhQpgQFRrvGC4fRq/AVTR+e6Pjro5J
sfj4d7E/Fprv/BCcFT3nMdCT2JNipTlHpb09ofYyNwo8izM63/nlCwCUs1VJ6rnl55VUYrvvTt9N
jNhWGQ8+Lt7cAkWwMHKN3mgGvBI+GxbkV4HnyLOX5XZdEQC/6zm9S5WcI5dG8/jZOKtxAqYkxFKz
vVbhGFsCMdHd52e8/upTwryuT3ZMWP8J0hSomI2R+l6voa0iqP8fsHZHjLdADh3XsBg27TiCK9GE
emzSeJrGJczzDZF7zTEIqOgfTWCnm0iS07YAgMjytNMzIUaMZIpeaqrXLh/e7LIR1tsc/tKS3vn8
YGywBHfiblrIszl458ofIVkG67XQuAg3gbCR0TtGNPtGp5EW8XB5F4/I/Hl1efYBmLC126tVj0t3
5s8/Ph5w4SDGBrJwSpKQphmag5g7x48fyKv2v8HpZy83BdlznimRsXtHRfiXx39Iy/ZYtozXxHTb
Z3Yt3YPwKBaCAnxVcWxM3JGclCoRY2GwQw3TFK21tw2l1vL61EgLOchJdeOHt7UuJawn6JKewB9t
1EEDoSZrwTkhEl+U/tu9l/Tn0wVhc0zbaYfiQbt020XzeR5r9YnMga9WNooW2s8bgwfIdHTVOjx0
CNUIeL9HDSiLXv09Tdv4sMfBlH/CvXJHcAE6EFnehYVACuIGaXdn0vcW4QNPLj6tjRfbVxO9wXWX
7P2svx7ripdNq9vYfACWtUMcqP566y6uX1xymsThxA1YP708DHMuNFaqdKADGE+01M0Evv+E6y+y
Aphe+n1u1tyIlqvcSV682sqLrdbN976rqdIBsxU0M1+NnFmSfepylsp59tVPEd8RuUMIX8fotiME
fVR+3oKY3B5sEHe2eMZhk5nuT6QTSG+Wixc3aYgqnpHwbcoUFxpEJdRtiaxvz4m9PheS/dG940a7
vK2GksRxRop+XUTdGWJwIspwZsdAa+kpd6IxLW+Yb340bnbmddkeSDce6AD5Hb9EiiI1IpuGxVGT
qGkIeH6fPpI3+WEtmbHua+/qTpafvPekQ86692utjhn7EJYXqDOc/ZBlFguPArYuKahw81QeHhqa
tnmCfDHPX7H22efD4f0gb3Ke/Y2RYSa9ntyolgbRbS8OhGqIbPo/z0WNHvjqzim/j29XcerY7vyM
P8K/nkvb9RH+ZcFvMLSHeMq/hx9P6ImHdo6JnzlXmwKo0lK+IrWUSnoP67sh/5QrlNW4PD+957DD
t4vYhnOp1V9fBmPu3uFSoOvoWG9P4SQeTI/Q+QRSWMpKs1Tllw9pIGBtl3m8PPzWEok0NNd28ZtS
C/10o2k5/MiVE2VPsj3K0lXpUBJngVyrN9PmlZigjNHch7P4m41vFmAAXRp2RT3k0gBNyjWHGNk4
Vb+YRO1eKZ6iZG1F7cUTRrMJISyRSj20U/+etb8cfwfXs/GtzoA1PXpSmcJudN3I4SjhSOOcBMzF
K659Qp6o7XuVRIgBWYn3EKDtiPDhzcuMDchYuxgBUs3tFbjHQesbN/25ygn1F2YhvMqoFv96SAhX
XEzp0hn1yXfh0UGvNs52cBqmBSeU/qyC1+UtDLUPkrA9V65gZvi9Jb9TZemfjPVuCvM+yHO8j8OP
fL8LnoSaM85trCQl3omSx8I5ljeN6v/oGH6dqWzT5XnKOZs5dJDyjWA66j0OZvaYIPGJF3nUA1mU
Y7+IdmM091x4LZCjxJcKqOgguay1nBalqE11RHBBwwVg7vTEAP1m+EDl8lE18BZidPMJFooPeQCr
95frDf3Ht5xZ6eQXX9HhfMqR+cx3Dt57ssrsl3GGWAR8bP7RNo+slVVnrbfmmhKh5rt883yqgHBX
ZepFY7UXRWCHTslppEJOMhKkfAtHBxqbLOHtTLlfQX1GQxBBUA7iO/kdGDWhWjn+46kub+jUANuY
ZEl3zJiPMXBnX75rw0vpyNnN65eOvdjuhStTggUxNdITk6ft6JSVrw4v08OqvrFRY1eOY6iG1ycG
Vi0pde/CBtT3k6kKhcSLUZwcSEAM8sCR6dW9xXe7GWe4wqAESX4arAtLn8WDUdeCkZXZIthC15E1
vflrw3fcfouBwQY5HfgHsYBDLDJjbVqQf0GdqeWTrKk3uu+t12pPyGiD6MLxCexQGXF1eo2P6yIs
6Yp4Cb+4DfaDll88OEwNvG9Z0QWpltJySEcLuK4/cMGECC3ShqB4SJYavcREKqsri6e/xYDKFx6e
bHCOcrLzKIN5o8FV9BZ3RtzExt++0Ps8OunaBi8fRq2xYn3WxxM10Hxqrvs8saXmaZDqv2GHTC1F
UQUKB0PRojbNSZQO0zAW1Fjs+IcuDNovEJkP+DzIH+d4e4xfTdNk48p3Vx3Ud66i0w3rbTatFKIC
OVqv8uXdvT7FAdVxrz3O7r9SnvW7KReGyrOPkRnuJ7B5AELmmpBvn4sCok2zbAsHksxn7h8TIK3c
NlCXoeMBsIVwYfXtQohuYLtHT6xSVsQDz9f1GOggW7BGsVqo86AvgutNkWrucm84/U0LQWAYFJt+
T5cJmy8CGgp+ZDuCYwCLp/AEPhs1p2EYSToIkdoG9QFsStBw1ZtcWBfYpap2s4pHq8AfE8h5c6nk
Mlwl2zVeZLSAOXli7+/75ywvP5Bi602C+CPOdHhZlAy2kNl0m4Us2Soypjoq3rGyVDemideTFb5L
HJzjkVfB2UhsolWV+fx7m/PP5y3zuVXX23cktRSQipKTIX2Illde880RXkxKc9iPShfJp8QUB3TD
5ldWlvm52MGwbTo9R33T/bLsmHHG7ydhU5bNWiznQUWq0mAKu0BKC8NlVtAtATgjNRpyStrfNmHd
BvsHGwhYNFfKXcEI4241SzanMOj/AXPlHxN9FM7pODIknEKDsMJpSgrm5wuQiWCOWXfhfcMhldN5
/qK5cpSroHtsI1Ttjl1W23IX21uiX7wWue0I/u7Adj/bvbnRZi8MxpPpJo5I6q6d3y/j2SYW9tVj
31ENFUNF69ClkplXfmTgPMXzKjiqLWcf3TqBRDRek87no7NpiX0Dga+T/WZcBoEKqFNBdpgvzK47
AzTu3bG6fw434Fi8e6kv1DuEDn9jV5ZYcXUV8jCI8fOIaWpe0gmEUtgMl3EmWEIBGvcuMmX2mEqO
1PEeDUcpXUjYyiExGXKJw/82rgvzvtpSbWeThOIOUC877APAdNKrK07h6JVM8gsVeimgajayoKyZ
vYLN/ImIhKWwp6+rg/TZvqhddOayOJyM/nA6IVzkJAMtuRW44/InBTwkRwdbPpar5TEDlIBBtQfr
ZdWJ8PkT2iyhEH8B2ty4hB4i8ee3Stv9zilqmIqLTAGhPgp1G14iNgSIs9DihakowoNC+DPkX3Tg
X0aB98EZZHstA06CCRoCsYxKl7N1uu/8Mw4JTPCIC+xBPQ11vRUHC1Xj9pDFepjczJmJXJMtgT/B
aPHx0xTK7+y1eLH3MuJ9gm/OZpVZZDEWFmE0GKTIObQn8OQT04giliZYX0LN8QYityKetVUF47Mg
1oKCWWyDWOIhC3o0mMviniIjvXgOJpjDIuAr1itboXe9DSbHX5kh8f1RUkUm9bkWj6N8C7vzUwu9
XCS3eZ4Y8Xom4A69/aInFwMm1U4gNfzRFSquMPknw2oCT89mVUjHoRLauJ8y2EG5TQSahXJ9QY2M
HP66z9YlSfWsEImQIzlWb7VqhNMF2NGAPRe1u32Bh6R4JtD70yoJNvpDgizfMHm+DCb/0cUyQdU6
tgTyljzGptqXB/huLqRidYKat3P4m58+ky1DEJiu6UprYp3wwAczkN3QW++GxCOtmr/jk+9b57yR
uvCk1HAhys9yM5inPVRFbyPVw3Cjz/dVcP5JPpHaW6jbFGyd/GOW1DLBo5YUDweNGqXBM3dcSdZP
MhPCWUae67CHWs+RjT8++wnVV0SVcojY05z+1Arwvk160vU3zT96lYYx6JrpgX2XqphT/AktsCSu
oiSex2Z1eWeyyae4S6d/nhsShyJU4NBxZxZXxjYr1EqEPn9nlqp8Oos4UaQpAqAs62LFMEMWB/rl
iz1BnS30EbO6jZb6jF+OgDm/p3CNQAEDS/ApTEcRbWGPTdpSXAJrTDYzv4KMY23z+FYSISO5HJnH
8NZsmCm3prTwtSjZ+rWM7/q9LlTbouAu6w7x8FrMerLul8ePa3yooJ85hk34UbNJ4nqcSM+v9mdw
avJg+LtS8MCRWHj0PfM7ReXx1iVHwFquFNPHHjskVKAfSgwgPBfyV1oQrUwjo3EINOwgsxrunA5q
8pMOW3h97teG4NRGbfML0l5iAEk7H/CQ6QG+vNonZ8iirlXENQ6SgJHTcikQq9HUgxaOs/v+ApVQ
rB9u8OwZ9i+PlOSbHP+wc+6F6pSg352BoWabXG8ceHDH9UIwEqHsStbD+AUlhenAURIWFXmWIzjf
slU78GT7BhEQyEOSr12MZFVrzIl9ZnpsUGTOWnjaKSG9lHpibPK0OLSjLdajzt/NGtrKS5Pt7+/Q
Enje3XNRZflqKPUkp2RrZHnOppY1b8bOPTwlGP5iG2sl1HL77ORTSKkSwVpHQb2wsUFC4v5Rn235
qaKwdkTOaMa1fpdCQ9mGyGbSmLANP3119Tn62l+38XrIX71MWqpEw7lXOZrtahn17agaKrMYcTzs
/JiRvC4sr9isBJ6UoaHiLaj9q+MSCteIMePmytMpiKaKsF4F360S2oA5RQaoYK+QNWmtATB9UW+1
gnP3jNVwLB5czwVxlvSvkePDwY8L1hmKVJbgcsNvGe/Q1mlQ0RwTBJgX+9hXObAAa7m8cnk1+Qfb
nMKru/NnLemJgzJAJsVbLgUcrIUUH093AoDy1EAL+vWsWRoPNYQcEwfOrKRkNWnGF1GqZ8gH4TDb
5OHg5RJ8dDeI61iPYewelgyZiDHaG5gVJLl6TbEppdQXeY4VCaGJ5jW6jCpL4TeU0ceq2VwWLS10
km0H42gjFMxBZf2MBfDk4pOR48cJF1CdY9KlHGOlFrvJHhNNoh0YrKslAa7/y31EaMH7C22GgUen
mXOVwSqoBkJeulGWz0nnMHLxd22yWvLJ566U4ZIdY70S3cCVwefDodoeOtAy1aIwRHkyWLPy/52u
05Smcorw+9+ZVxzKz2Bz2FIbuevQBLPXeGIDZ+3e8rQX1wuR4/ODQexmqwDbrGzwl9pwYGKy5bI0
jfd9H4OQZg92TjdeSvjD/GARsgpdYqfFRFLbrJ/iYqEV3DayrQmcYemwRj0zVBryzTCItDz0kJdI
sP46jv2RftrPmVjV/BcnXA92X97K9wet/S05QMy48qBAk4oIVyhXKeApDrp/rPn3eAwVEhHZl0g9
IOaqIosYFSOzdRD0MYzGTuL7376PCVdQ/2CJgb2K1D/p2PZeYFteFk5CubLPVvsnH+rD0qa57ijv
JJnnozmM5myDw1mOkuS2C5EHrkuksPIV+73CunpqNVs1SK+IMdELKTix8bsDP6GjO/CKp1EN42c2
eMtbbm/l+o+/YrAh18fD79puqRH4+6xwULY1pFYJt8fImZsyiMApcw29pyUqKpWYib80t5SuWeXK
rEeEBUiDrTFfd+r3zge6oBwgY4jB8IAmxg/MxTqO1e2l6FYsGl/K3NYzEmnYUQUiCypls7YSXuFV
6SAw2ZyLkGhCJnGDYNSB6Ez8rxhCi3Ts7QrGF+T5XaSsiaOxvGqDKgJD6xIxYMHeW39PUi1116h5
apow9s8iAjCD1evWwOlyKzmfxuG45VLlsCE9XWAfm1oa+626BzwFHAtQuIrmA4EyXH9cgHbZlvT5
JHPxWrTTZjXOg39QkZPk6lEnKBpKvRTXvAbkuWPVzONoDhCsABOTlIGzy75FYzQ6jJd151tSYWU0
X4YoVsww1OUdOYbHARh5HewK2V04DR5z1CeGwilne6X8sR+AKW7pHTHSI6upSGHljGsMMDR6CCkG
/edYrNNQH1sga4KpLIug33EhBL/bhOVZmI0mmOjK4yNLsCFvFhkb8iy9QIsMJCFR+0iovzqzFxUE
ugV7sFyv9TG6+IiHG1mKjOAnCEJ3GQCOee7f/q/8NFB3iBaGpfqK4HgvyPh9SwcqRoIefRUkwSbv
R4sdFVLYmSY4mCoIErrWL03UpKXO50M3vv15fou0EZL+7OOlXExDF8b79St7o0pIlRrMEHWYBkXw
DeaCs0MTAxKmUwW18T3E0gghsNW650l5BHvEK/zCCR9V2NVefBYZ+XPYRhV4fa37IlNPoJs4kPs6
S34ZGTgHbxox1QH/ZvuWFiR+AyCY22OTEbAvXUc7b1bEYPBS8+OwMz9L9v+PIDgUzrT+DFzwLDOl
hjVACTPKazBZlfQUg+iODO/MkWEMflKIVAH4QzD88O9AF8dmU2dV0D2Mt9RYmNUhZGnzNU00Ycey
TqDHcmCiJQwouUM/XJPKM460NiyROhuXFPUIV9taJa1d/dRDX8wAvqwprwRb0qOylobamPqYmcRR
oILf2mlFdyp0eKn03hiYGJOJcPigULR3T/bCPrs0+X/MhE8xcHV+s/yiQ7myx58gQW2kGzOrHbPX
p3n63uYTBGcTGr7vrKzZlrwUNWDXEaUfEnvofD5TYzI/U83p07MfTOz70hLUPd1I4Dxc1v9UafmI
c2UnTWExkpO84tlE0TSbBcm9A26u6DSyQ5c8/6iUgW+a4bZERyV+q3fTdrlSIINkJUqp24fPMkCl
uJ5cJfV8Trrpfi6GZouYYDoINsDlWcZQwyRHEoPjpFp7kup3BE8seQKRRTsbZ/53tZc3Afvqt4j9
Fei9o+sasBhk0DN92G1oHfyy6mFVgePYnr/Py4KtFs3FyvdSQ/Z0e6kSjVGsF97zisbvAP3+qd0q
Vf8+elaToTatr32WFqXmQnF03BmdszY62bfl2eG1levCuHz8w66Gdjyu6rjpQCfGHpPKW58OFnsm
/+CvYH7aOtsHBwMi/Umy6GUq0lFuj+HlKtcSKrJQTutQ/l31y2OdM563RJOH3JRmSbv2CTdLrJl6
3LvU90ReseGsT8UdBrCnywq6ccWzWMqoaxnj75K/KEn3gVPW9Xxe+GyooBSJ7CfejYc+6t6Sxnd5
kbfPpXJIWNR7Mh13yZTMyNvlSLooTKQHxzKCfMjmnk1kwM9+dY0eXrYZRnl+2aePFhyG8siUOPWl
VyS8oPePsgIePS1bTRDbZB8wX9/txgyUsR/ZQV7htksnscBsdeZs3atDlfSkEO4FhSqGNqBnJGQa
iOMFVmUa4Hjmj3fG8eSabQwBiNaiG73ThtktKdCZ3fbkhxn61UviAIAvc9NElNLJnCvVs4NY8scw
6fIkXCRhPgcr7RM/RdA0JS+IfIyChd+x72lVCqqi8VcDU+pldzAmlMxuSEqYvBym+J7itVwNUk7K
LNXg74aW3sFNEsnzVtzQVVSt6/JVEJb12GoNUp8TnBRnkO5ikFhsXJXwTZ/Q+fn7/mtN75KqdlzQ
ehlG2/2Pz96Q77sD1PPDyU4fXl8MFAD5CvzOi+84Higij9c2EAZzoz2wjOGQr+g9OFprOv2S3Gw2
8Jr7vl3eWonzT9s2m2g/MX0mfOzJ+0myrjkqXdCOJHxGCUZf1NVd9qykQi5jvryL9J+n8JaW8bWN
7sKCdvI9zjU1y5vi0QDmWlNfVuXUjHNcPVP708UdyADIQMtlXeyDmBUOQzQQ7MaG3EtDf04WpW0L
pYxeAduwxCRVtJgfEENtZc5L5CG5qPrv75JZkmJtWD/I2O0EncfT/byAlI3E/ucrag20jEi5Fv+w
vUzsrVr1oKIUp78SbKQU+bo3SNuyUgmisIKQsg4pQ0vjCdTmo+o1veCa5zAlxAMzItNHDR3/xFJf
K8wqnWM3eA+3HVs9wbodIXiFCSPiqKGMWnSUt8YiPb/RuaogzDpIRYD1BdXNnGaSx5sKj24dIjZd
aUEe6NWT38IMxZYKrUMp0ebfEtZAQeVdgd14NU/WkSF/eOuk1xBm1PUupcoBGe8ZsM4iqLvc/fC/
/L5nUIIYXSpXDX5Tby2jO43Iv8i0spQZjSfHsaewYHI2trb2SYPsq/kCuCZfvpt8+91ST3dbnqeM
hpCO/A7NQa0tq/eGepRndQ/hcshbLTaaFZoCtHz8+j17Nx4JiH0X/+2miByvuYtuqJoSVXN67+5l
vZgj3yhOm8FLG+NCoOTj4QP8clctvgpzx3NpsfUwdSUqRoHCG24wK5OvnDYIGWHrPfnu0o6CwAlH
5KOBipG2S/3FCNzIwVYBV+obeoOLPEGHQqGaOfhanfMBWUdsyqPt47fEjFuD+mti3E7i2QiiNweI
LuGtW+tu/p44oONdDFky24oGHoNMfnDLwtach0rvSS6mXLYP3lJaEor+z2qxiZDK23SUJe2wMalx
IU0WdV8mmxQZTSXiaMjt7nF95MvcHc4j+PlHIQzlIiN1Ufe1agCqelqTR31k7hyQF7FD64fXNgXJ
4ot8QB9PzPmLGED1IGcP/04+OTQRVeFzd574tNWx1lQT5blqabgYc7XlEZf6FtTzCubf+4DFTuvO
Mqy2Xce7MNp9p6J2vUeAzZREell8DcMzAccXW5qKTg1/xMyY3W51j/i1PYLyx4bbKku6wj9Pj9TC
qxAKWQ9737McVDi9VUMWPh7doaxMBQUuBq1rCv8mejlNs5wRgYUA1ykoARp8Pwyq8WkReX7UzLar
oJ4rFjGQX87nnGhYFaGFMRRQCa2VVx+T++Okfchm62uD2DboZFhH8FeAx6hBHMPAvl65OKghgw1N
joufBZ8gp3IeTjlt9BCspF8cNfGocFbu/RDfF4QCI4Mrttw5zJSjZurgtVMGA3C9hiUy/Xpw00X7
InwMG/2efukDUn4eSowXxGYBC994qTysfWkj5+Cwak0g7sUeFzd4dxPrP7YKSRqnFb4G2XWGcu69
LyJlKyzl+5SQ2Bcxu7k7ro4g/5otrLCaHWKXYVOJEs98qB10YViM8YuttWnx93oCK6W4vbAj1sOh
295bR84gv8chsbWBvnxEGHrbvVGDgeHpKJ1ou2SdYdwNvBFtAwcgffWnt4AWTbzTDR4vvTAzpUWq
SMFTnseR9O5KE6yTEFNW0zCAMoGhf4N2RaBxYa0UBVn5YaDN4q0tly4pKXRK+8Dvjo96S/QYcBIF
mtQikMCPhrUvlRtdH5ND/o33GJ3m06zhvvo4KsM7Bw1dKh26Z5S77AIkB90baYr6GOBBF9Ah3eXz
KkjOwM3U8JogkM7lWfqTFC76qxfcCmYOaezT/E8NpaY8aDYqk9jZtG7bdZdJHHKZZCy/emO3Lbfx
W3H2RSzhDv/ASdZFocOvFe/HBoHeRFWSZrKwNjJcxYAqfTKdmYX2yZNcSNdQscioYEFkKjlNIPvP
MAL/Ad6BQH9UCwYmTyg3NlNeWTZFvKI0mhzmRvvQEEwvwV5UEidXpXYiFDfY739iNir1mgrohoFu
9DH1kUO73YPn5QjmBUMGL0kCqEi/QDAicn4etEtCScbBUrshfcF8KhJJ01UcxRHvv6xHlKmKq6GJ
HwjyH0aruGOsEuPEwhLizDPil7bB9Sp/9I3rL/Z0vWeaYlciKwY9bqxUrF9mdFkZ1xOwyK2UT3K0
IlF9+R836Ub9yb/GtDtwL2oppoZkJOi4f3PQ6tY2a7ke3mkkIcBUWkJJmGmnIMz3WOw8FvP576sq
AQxwAOI14cWgMmwFnw/Q1CKmwFbk1GaUuywJn2eQUeW34JkwQVBGZ+Oespha9HQIeahStgGs23DI
dq+H3KlqEg9kF/MnkKbpnk2gP5lqTxOTpUCSgyY7+Gh2VleVHUVm+dPqh94XQLsTv0cd+014KMge
QPZ1dBwhfm+J8YX4jBaY7a2z5Sl2hpcvpj8Y42/8aPvnajZ5upckEWYQ6Ibgk1dtJu6m5wVtSHhK
A2nHryHpfmbxSp2sGEngsMwSBDgy5SVtWJIvJeAXp4gKznYw3a7iMKh2Y0I5ELzNSRfN1/mpJ1W0
EQvjodOkY1RyON6husyXcmBhIIyIvtjcxFUhX0dbmsqu6TEcV5qFBLeinU5d5LXoScx8to3hRT9/
chZk+PG10PeP5AyGG+RL/Zi34Uxj0MNHPhTFcEliRdoPrWJBB48/nMRKZHAWMzTrwFSPIgGfYept
Jt90iCY/21bCqF/vawrinOHc+2J+DrsLrNkuTfx9YPMQWP/VO1oWxFpcJZS/Tpw5+xooR0IVOHlC
6JibDfu8xErcXIFkzAN+byDxpsG6E19RZk1Ew9jbw3ATKaEOX7t5vAgJpqyvMxYPzkpW9wW8srye
FvY2wgKQmqgnbN3OXLZANkzMXQqNDSndNvIaSPY6fn7pqVN0KHaR+wsjlj6NanaRJtP5zTn1K10n
6FEXvJcCbZSyLJM2rk3uHGwsrCs+VODAh4sIfGoIrjHuJaylMdLOYHBoYgJgi5yfHl9YenS5Pte2
OdnJsX4md7zc9URqwJtvMRWTXTxGDm4ftVnSXNgSeNSoyxPHA8Nv8vVDqfJrJl+3nZFBxOw/O4cy
cD2dr5C32Urtx9gw50gSMlHqIldXstGCCgjOdVFweynntZ55K6uBOxvlOPAiUgDlutYc4QjSWiwP
8eEKtxoOqKl6AMNvmFNpak7A0Awg/QH1xYf92rNkBY2Bec+c54+Ulk2c99lAHQXVRyFfLmBLOlOg
XzcbcNaJ9bA7oYeg98RklDNMHYNAU72OgwzuXn0hu9XO9LKNec8YqnQOb9PZC5nbIY67AH5rRw2e
Sb4Sn/uBTyRK2eCHgtgVydOsMaphikHAwMLuysEQR9urbdweckL73mZcVbvpViXsJj0hhC5mugA/
WfQQHbgT2r3NdHbehEkIlL9c3wlsyrraEFY8OLqKCcbzwXS9k91Vx33zpXeiE8qejM/TSk266cWK
SmuR3VXxH+MaxtrLbl12A8K/g+p5MZajK/Y6U/NM/Pn4s8lpuAUixSG9TXCdtjvzqT8VV4uBBpFP
8vutYS8O7P4j/u/OBxStYv8OGwWgqppQGM8f68B8vlJJb2NY7k4/FViMeuwv7olE6FCCTYlSk9r7
pmxzVb52yjuM7AQdcohIWgCjRmbmfr4i+aEroTUMkmNtxblaEhegk/t17D5sGUTFY7wOuVlLxEqY
lUJ4/muW9B2YGN1ujyiq5/In+fiK2TjkeXalas8AMjGdl+LF/NMuBVi1rNshPtPOamsNuq8nsVfx
Rr86+YA4lD2ar5UYZwycmPitz04ZCNIIKK0TdoAhx4xWtoTTptTvDiMTPDwyHylmP4NiYIHB8eNf
NT7TDK3YydUVPJkpNNmEf9JV5Q7xA7w1RTaC7ASofw30xeqqR5Rjr584ZhXKdrxR+Wiv5PtH+5JH
O3ZsN0PpsfK7g17ZlVbgUmt9p+p9eWGf1I3ZgG/hpGj+lfVyLWOph9s7aO+BmCh+fRkInKzghZtf
yMD9jB09ibtmZqcBuspiOtoFoqyJHEQVN/hbbMV0Hzm4a/4YBrD8NAS4sj4fXZlja2wT2jK706wn
zw27xkygYBpazAXkH+FW/zPFadxDu1mcGdhP3urkeejYwcMVeQ7tWk2rtEj3mxKwacVvgi+UyJjc
N1zIzrOZo8CRs/vWIbF+llIWm4O+LMSaPSR7UsMibKvBtxVcxRL6kCXMmpI+DQskH18csNvrW5T7
2sdLSpmAIzuHs3DsuZ1RUfaO58fzSUK5xfm0yf9Xsj3zliSpxsbVDhHCrbI4zhwyqv/YaaFm5kN1
S62NquNK8yo5z+zdM+D293nWyNeUF+AjXWuasOTV6megDnrXXP26oWtkk0l8naLjblJus+mO/UF0
PDsJCIJxQS0hj+AqAKC62jDTA+Mjl/TYkqfVtEsG+Zf60o1S7J8sTOPHbONzhKFoTgCZsE+p+lZh
/4FOye5pJuAE6nBYmsZ5BLWQNlNSqrU08K4UdEGo6nzMqpP2FBxU1Mpm8ZPcoUOOJhAvC2xnpLcm
bTHufeCvy47/mvBcCINA01Gzx40BVEtUrY1hDGoiQyJRt6Kv+tc7BduZgV4H+dyF0OHmWa5IDibS
UnjJO2aa4fd4cljtxJpJa9K7IRozn1MWkyCzokn/Y2qfuEjIUi49ujyRPWd5rV86MATGhVrS7GCX
tMs/Z8NoRuBTahijOe3XkpzcH5FT/vKXECYouiRGxtg721SZ5OuQotQoh+u3ZnkWQJSLt59ShQmH
aE8BQ/03+33KORuFXtrBzTqbU7UHBduD4tNWjgYaalqqlrIqKZbH7ZaBvqZ9jH6CgrneHRyrAR2T
luL+FxZSfG63QccLeEMT9B/OxwIkht4Dis6S+s2R/SbQ6gfx5bi8m04a78qCNumDUFeNYPHnYPvl
+I80bjn8YVxpCPNqVfxZaMKclMIiDJi8xMzpc+GwJ2AlOvriBTSWG1+f82K51OJikKCYiniEtaDQ
ctYjGXH2Gf9XQlgzjxWzFJROI82JjLJ+WH6VZqZ5bruJSqizYYlusyQx/vW2Rx7PTF+NdmjakAiK
7/q234fdZJ0dGrl73pazS3xU8EMF02IsrrP8Qv/kY+IGi/8tYqEDIgDiBiYqu0zOL3dmiY2yFiBK
8lDypKX6z7DSmBbslpNNV2QHFlIHQkhKpDDmBXCi6jg2wAr9MJPh4YIpSG0xb3WPVNFWwByG2Q/w
gvQUm9RfeRJHz4UL7SGdRbbJKyiWAWbnlEh+zbWY5brTqFinGdSk6AAu+N2PYx/Tv4Ro1a4/4UI3
8Hd120JFZc8EdmoBkGv+2Ynz6kMFuzQMwcrVDu7EAMklY7dZJlexXYIqcWNUUR3cVPAuZbjiz5P2
ST6CJW/2kT60o5kY1cdDB/sxHeTFzTTK4G5moDEua8I7p00P4XL6wX8FfgPPxktoviFGGqT5LzLq
RR8FIjMHJbZ9NHShn5QIQ1ceiOvWjJLidKoGMLRXEgaT3TTqoGBxYwgWHquaL13A1CWfhkBu7pgV
RgimM1wFQne/EtpVUkZ94J6DIF5BCUTNxpDvZRZ0U2gyr2Yulfgc74DZkhe9r81aSjY8fmcyCANA
/qE1nVemEwsHWlvDaqdfZ3Pox78TRyG8exaTp/R0KdG2Ie2upz3H2qeY6QX8MDIRGLAc9Y+Xqhgn
C5QVYTjGqxbEI1iOWNghPjjXWF5gbYghOvam6FozYMx4f6TIbJxlwbty5I2Ttyp2N4hW0rv4Jc0E
G9WZtGPh9B8WkRPve4GgXtzWHM96qGxNf4cV0pSK5rN+WdIWAudB76Wr0hz2zKsPEvin/7Hupg4N
mFsoggJnOZE3WoL9XnBxL20Yx/cTM7NhcFLG3sv0Ak6JIGrgVAmX1kwHSW6o1WJHE5mVxDEF23LG
XoYVqAgmJZnl5rMNy3A/XI486ldVI79rAsElt4M7rgVF0Uokt8tLmMBtDRadq/AdfDQfLAKDSvBL
H9ptD8FLawayPqYiMKfpD5xE/ZsGvivEU28cj+2xVOA1U77CDDu/ELJkL/vclOPi7ITloLv5oJMR
QAmstoJMK8e+fBIlGMMvBfYBNnV6JZ7NTY+Tj4qQR0yaKx3gL6BWcVwmDZK8+Y0zPhhrA/tso2FW
GEGvUzYVXWQvDjDtCZ+RxabLoUTnMKrEwsGSmRxXhicM20UvZhDf5X8ej+qiMiQRvZ9F1whJYKO/
CiofJGdN0ttiy1v9rnruMMWgLtjtXUKi1MYhEAcKNYRuEa9MHBaJz5MgsaUgXMjErJZyfuTPTwKL
lAjiNuWSI6JLSIMMdZeIibJmU1cfE1kQRK7dK0r29sYWm2dDGwO0tkyXWOT/XVywaUWVusJ/Drt7
0DCx8RMtkTEzahtYMwp7rtDBq+RuuEOeKQIN4fmO/xEHIkOgQn2G1eyPoXfK3l6eQqOtoPg92IeY
b/7pm24NG0fdvPhpvu70hsBqv/4xNnF9NzrPvA8bj3lMiUS3GFBVbErzvufN7nBLvzDwTSVMBzpI
k4dz8pnf+fbA6MhUShZj3yLMq3kYmlVmQedaS7QcRL2H54NQt/EK1xK+n3PenwtswCp9jKzQmFht
sLIneR15DtiWNeZRwdBia5dIgP+SYD69EbAl8r8crYYciknl7eH+s2Rd/zsHjqcYRj/rE7GlVaRs
LDFfxHGEuwt1cI33uLWhJkSF8Az2wJUuloa6MktKv0SV1Y6hP8e4E/Fp1B9vPgB6+R9dfarQ9t1H
45o6FG6hIyjDfXc25icQV9P42/ys6NVaX+miY1Zn/wdT8V1JOd2udPNnqSjjjZ8m+euXzOA+GaEL
LGmCk1B3CD/ws+cucC63uaWi5JF/eZg5W8q3XmCP/3/OG/boOfrm/1UK1/lz/+HTUZoQNpo3qZWn
XLWJq4rE49UvyjJgqVaXG2s5ShAS/bekQ/eS+lhxkV1MzMg9aSyxrsRvHhEsc3cH7yM4eGnoPAlt
YUV5D2mOBXQusF7qGQBUvG5LlRXxPP8DetlUipZf6d5xFKkIkfTHCjrTsbi2iQvpzfTAlN6hJ6BY
pEIzL/2hAD2/UfnVVL0DCphG0zfJ/zgRtNb/C9oGrafdXlnrgd6dkATsrzDGrjsctq2laU8lBaHI
FzjlcqQxbKFStDQeIjuGwlvVv+5GLKR0yONV97PGtedVVdI88mzk/NGqrGROt7PAD95k5PsV+SUH
63NncPrdQhgewg4wSELEwIyY0xpdAycWWZUmdVPxAAaKI85GM0e3g0+KS7h9wDaapMYNQ2Jj1bA0
l5eLObtcJPzv1wuehRiA1Ff70ovQcNWcf0pomN8F6l2sdrWbY+y1Sw7O2O3UNtj6RFSrx1IahY8a
m/FHBzUfKNObPPoAJMFtPhqz4VrE9lQMClXALQ5HcRAFniavSuMaa6gG/emFZGkt7cIMCjpIOPuo
Go+s8nnVJ+TlkOrrmyaQy/tlREsbUeHwu+3N58bflv2h3q4B0/jikGMNuP7VXYhHCGHDcFQNOoFZ
6BaXMSOFVAfVutqcGzVrLsgVrU7hYefqmWZaOx54hUVnhzK0t/uniolsE9D3GVHjYx1nrPF4LfE3
6W3dbh7Ugfl0xkQn/PcZn2OsfCHSKid2dQXSLVc8RFXsd73jnp7Ay3Qq/2ZCawk8y3hVaisiY+zK
eGTfRCYGEuCyw1FAkorThRF8IC/TCaWV+Xk8QId1vqRTXdZqfgMoyC3utkrMmmGnOKGltXtXK1YD
kFtJUWkr/LQEhEq/1FA/7e6yv86bP8+ItE9mJUt+jPH5BXwBuiXpeFimqrSp//hDU62VqtC8eFVY
q+weG3RNA3dFqDh9AGleyJHXLwSpv2m7C6vq9HHbv3/i3GucdfmcxaUh4Z9lnMOGDAH26u0eZar1
XNs5iCo2bEybe1TqycOoaraUyY+z3RqUFwohrWrOEDmMVjpadGbFGXNuAkOo9U8NY3vlTeHg6D/C
Pdrvmg+Q7LnsppCMXXVZ/mKLjqxtcdqXCjJfMiy8YJUvvaOl+mdKJ23EdQT6IaIe9jVf+ayqDyWw
f+5TYWRJT3PQPbqRn1maHXQjeU+7bMAfPUuNNfFMSgdllMzcP/cyfvqDxuqKFrVkynu2oUmuzz+r
6kxJhOp27v/Z3MZ54YiKi6M+DEhte7tGisEWfVhVH5eGermEi7cRqHjf9A3btei+Se9VnitPBFWD
gAXET5YK51s/C1Y6xdNqdSq8pJl5zyr7dX6XRffGkgXWE0D3a8XSdHiA1k50TgzmLMK5EiKYENjF
CueQCS+NuBOCnAM1FMVtjWIQgFvCDfTzY1gEb1BE3O0nN1vOaaxMbe8uFTKwBQdSWaHJKqgLIYPk
iNBLSF8EndFat+xTGH4Icc/u9d2M/SCMlhNBt7c3qErZSDRqrXx6lypsNHmyfwQtFJ+oDRngCELc
KvQ8TEaJ5m6VEuTdt9lvLf40mR9RdxSelJ15L1Nkg44jpXZ5ghd2QEuzd0JWsC9tZc5q+RsUKhgL
y3+ApQw5xGCKdcD19PsGvsIhnPeLiQLRmY0nxbigXbPszvlGV4hqptVjCYOh6AeFWyIccSZsPbdm
KSEgRO/+RZERan6A1cCNLqCe9QQMnEB15g9OQAj4Hc6+JeKJq3sORQAQD5bCQrQ/h8ZMe3qLe8ft
iICcUuFr857TFB3B9lA0algDWDa4eE6d5x1Mmu6Cv/i7s54zqtEajbLjzyQsRciBy3InUQGPeyOM
G6Gvt1mZEltW2OIVlb9/9e+a/HHboqoiIZJUmHqCm9i4cuMUBDYd1ALfJQWbNwRKZ46Oio5vofMS
/XfpJBRi1cRIU0j4LpzSwFPe74/Kb/qY0Xw0CN3chQF6SVZ4Y1nPnD1sX6RmSNOBj2P3Wj1DE0lR
OP98Z1HsSj8INNUTbD25eWaG9Ym2KvYxVSS7wJSP0xgLYk/8sdZl6zhEq+Ybi10LrA1fQ0gWSDg/
+1dycqwkoqX8riZKX/CI4QyBxJh3a1VxQjzCLbgt1fOX/pk2bZakAt+msq8Y/D6S3PWw4TL+PzWi
xTJPDMUN7Pm6CmJwnxz6D/OOd9iC056pi9JlMKIPt/7w5AobRQ46nI37YuvkXLQeCDYDUndDAJP3
yVFigLn9zfn+y4PKR0AUXBMkgwiS6tH5x+vButgHNb3PZRA9YuB8qMi2lHNamqDFgVpBFIgh3Kjw
o7e5KnF/UjeGfF15LaX6yXMlvTRyGrp953uS2tsNOIMk+HcEQ7mGE/3Tqb1CJx0nxAcPNbfYs/vC
Dq/cjvI8zF5SBXphAAYvEW///8XTM3pNoqslve7T3+eWW9p6xLTeiPqF2gwQADVPONRREded0Wwc
x//pfjEji2nXIG7ge8a6t43Y1QSYUURIurE5tuZ7H6rCpTayhPOjIe2svnpPkT9WNcNLI+cyGbyc
vNqNXGYG+BOxbyCP4lGYTXc5SgZMQjzg5zPj0X0JYN6DV0i2MqSky+4nmO50rmab7GTQiTARVM6/
QcMNUuj2MjFt0NRCAJ5Lu1qJ01OmDB+f0goRqtomhFWKJ6mSfp4DQP17LebX9mwmGzjVKwBVCp65
xdtLwZmySOH9kQ6LtXrOEFvunqBhmd06KiyVBzCUdEjKLZEtI6ivCCHDvdIqhwIG3H+dd94lmc3I
dH+NTbMmOiwy2pSh7zERZwsNP1SbouIB41o0h+x5dKPYQJkZozjuRUTuoPF5mVALy9hxvhFBVKnk
P3RdOKwdutnSn3j73Efw8cfkfeTrA3raMBgPofirQXhgg5cma7mXXnBvGSnUaA+Wq3gh/fV+3FiU
s5T/1LR+R9OgB8RkCsObDZc4Jvhs/QcYLCw1BIK8RduHTeSh7fAFyeCxhDwKHfy9p1KJFyfHQ8bO
vA3ZQQ8uXMe20Nt/pNacSMvnCTiXrtpGpeL8CxbE3iDragoKI4OUo+6AdwwJJv27cfS6l+R7BMQT
8O9IujIhplHrC7eh032c5KINC3sHaPG47cLzqXLxZF273xfieGujgWT3rToT48kn0Dfjb3fROrDP
EObuBibDtc0SiGZXkFsmun6kWYBYbuo4DzNHUo7rBzjY4VfziLZ1VCrMXCbwnbCkwk5SxnWwzwV7
neaqJLrE8O9JQboStW31Lp/sPJKUhPNMD8KDAky7V2D31Qfx8NnOWDibj4vQ3er0QImUgjYazqCp
v90OZ5s20aOjXdWtwHBsisWj5YIVZgeeO8ZRUFfcjUYft+OtnbPVh/vuxkcEORDdKkG7v3jOC/gF
GeOKHdPQUhjp2jRP1+Ji6G0trknXWIWoV8t+4H1tvWos6s6A+mRWi1GPAgmTTpGmmvO9UvW/Lg+u
CuEuqi3AYGk/l6oPizFMssomHzJKBfXbRn5s2t6L5wMBGj8W8Ru7bdiZxFLKghdEZ23MOb16llN8
UHCQioTEkZGQvl2zJ0PT8AFAK8wr+r4Gej1AzycNSBq5ioC++SvodEK1Xvu1BJmz4QehSAPhAaFm
dF0LmAGNQhewAYgFT7tzfkizVte3zvatSw1UfrT2/kcU4F6Fji6qX1eP17Miyd9AYJzMuhDKbeeF
suwIhLXpuy/oaBHZdwHut0z4XNYa8iVaICMrYWOMMvvORWgJQK+rg7F49pxvsu6cP1+INrrap08Y
etBJw+B3oVq3NWGDqC4v2RlBD9T6oy10FYP5NVcOKhejLgx/2VMtZGIKDZkJVlyzTXktU/dTg6O8
lD/TFe3dZjM6q4L0ws4yzpF8gXa/EvLYn/2FDVXRQcKYI4bLwr3BRTZf7VkUub6FMyCb5Skswh76
vvb7+QBAm8//WjjxfU8aAr6+/3F+TdrQXbSmABN6cum0eupOkYjBApm4MgSNcFUx25lAiy5wmg0B
tNKNrR5T+VDK4NvmfHSFNnQ/PnRlK0MNk+6PcizIbnPRHf3HLhFQm6Ox6XLKd6kNhqidLFbHX84x
zu58ZCug6Xm+tMT1zTAaqlz+g/4Kk1x67P9cAVDvEsETgYlzmkCFr1Lhk5pYUXfAxkgTfbPwr03s
9YXUyAD5al0u64bOZvDSpjEM1+7IhOyEM1IWFlDHvvf27epJHdxjxbNzndh2zgqR/yz8ARFxDr4n
PJkQZq4aue2pgTvmhJdlFvsQ1QhYUptXjb+Pgey2e2g5YEI2mm8GlXSV+6xjwtk7qaBNPwtjlK+n
f7ZCpciWw5e++rWPIWbxuhrjbPb3NhTNj6egq4WKI31Li783YZJoeRS1nEABzZetX+3lQJ8QQHT1
ncyNaDrFGdVwpha7iwIYS8eh4090JnjX3AuSJ1AE4Lxwg6pAbQjXAS403wiWgmsUmVuMay2s6zbw
6hy9Be1y5mIWpvt8srkSvJ+kz8G/X/Qbp2qY5gsm9a/MtVF8vTsKOOI+/d56tddDv0/DVRqD7Cxx
LaxNM4/UCw4WKTofc/ONNXiSzwHwQcjTgAywnHq3Uy+yTxFSezrZwGPM1YRLCZ5hyXwEHoreNvqa
Gt/9yX5gn94oClV1k27D2ccBKrBkAQoitd92TNUwEouSGoKo4R64AvLCm6wVZxA1ur0tta8EWRBy
jgnUins5OytSvb8eiHqsSaD88obAlKXlPVGZC3EEHWHx5+A0tyl9/Ajl2vyT57o7z0nTiM+tz2ua
n1730+hPXyFx1qmzz/bD40V0MD/w2/9jUVtU+DQCoOXa/kgr6Tc0il5y9Q4sVvIVPaIUK6GeRu2s
18FJV3akxAc0m+kfnupvXauK+5MbjmT5YolidYwI2vLvexjy3WEugcHER/5lmFylvlmAXGnwUy8F
UAvWEdZzrzXpTwkORksKRYQp/u0JmR4Gw4iO0nVG80HaqmrbtsghoyieyQ6kQRhPeY14PsrvvdI1
5BRwyS6bMWUAppC37sZ64VbjAeQqfyInHTmIjbA5J915xnWb9GfAV55wqJTH9OexWycPMvbeuMx6
tPEZbAdiqO6/M2PcgPdkAWDdPKNqoYjAjSQJry8W8V5MeUR0qYsloxTaE/M5ZD0xNhO6X53Sz+VX
AOqerZ+YLNhvQaiLoNemrOXN7cR7pE5h0+GwPycHMBkZLjCpFVJB5ucgko1O7VPokn3GTU7hw8R4
sFy6L4Vf3/bA/B24yb3ITcWfD6v1eyXZPbbder4OMW3Pmif2Fdc7BAj+XlA6k4XXaIyMAgS8AbX+
ckW6R+x/SKDcOLcVODn1TGMsdd70Gc8Zh1FuAgnQBDtfY5QMhy4AFTa5UdfTznBOF3fld5dDYMCo
q9Zi9UPSYN60u1QV0H1Fg4XCEcn0kcqOy8j5A0I70NEgGEwfOmFfjJEPUcY4aQ+qObbqbyDx4ZhK
YVK5LcnGRFIthTOawpLtkhVT6cUJW6Skklb41NGXHqMpog6BCK9dTBddfgfCR5cY3Svb3OfEA7EV
4Qb+AJckdrTO25M2b8LxQm9tZ71v/YWKrMga3e8sfXU3RLwrSUUcJ9NFv55gkfbBgQDXdWoUw+Ze
GOCMwqAqfi6nObYE8NYk0gd5AOecYJlsgWFOLM0660i+mC2vyBdkKW7n+yhkl4sMK9ubIZa7ZBRK
EVNWSh5Wvf136KkNY8AQkn0WBP+GywHJSJZciQir7RkUr2G/4yk9v4FWi6hOe9bhr2mlC5YyJEEV
c7A7MJKBDG/1gJHT+8qtv219D7jIymdtTAKlv0LNCLnVxrOmNSRZqDmk4AguXktwI0NvE3aVAS+L
d6BjkGvG1c5ZdX0izEdidvnT7RlLVUin6BfgDw8ay/zCBEFJvhqfaVlXaOWiok0kaNXCH8FkXkVX
JxBRatupIhOms5+trOlV73MncQ5CPhmJEUrPn2AA+OPhRzKINjbJ73cGlIlrGIN3yjTslon6jw3J
nvijEpxS9VFPXcfFJKEAsV0WJseQ38HY+aWD0dP/9uIK+gUTV3GpQvXIBAomqSWwXVz1c1mvVaTW
rlaytHzYQgDki0r9cdfRDENMdz+3AVrFeYRE/7x4PMDoH5m7hTel0u3nkH2ovdD0rHLZ9Wfl+zCf
HFElchVxrowGm8Kae408fncq2GqK1/wkfJroAsqTxfG31AtDsngvGdRy1rJrOYQ8yC2DePo+7BTo
4ig4R/ysXKyUD+v5BJHmfVELB0Aekaksetws0XPlW/UKDRR751zrKE+FjWi/Z0xHKBRUXtSCz3J2
plyIBCW5jNNcOqOrHTwDXY6+A3kX3qeDMiwsaW9y+zlngQPTZ3m3wS4g7vdEbAN6NLMyHhpgGDrZ
L/cwWgtXQaKR6gL4cL5BSc9IqOYgM5Rnmybyhbz2vqH03QGK6hc90nSewIo60M8UTaASnNgy+jE5
I9VDaZ6ATcrCIovl0GyLT5qbWJJxq7+epR2jpC1FVFetX5Q9bZM1xFY1zxDMXGZz1ElQz2rV5gY9
XleFhIn6H1iu5OpQaCPT89Uh0+T5ned4hnJe1ITapax6u+fCDmfMZIRCjx4CsmYxUeEYAuSyySJv
z1f3YOqOxCa/JJopnBkitzyEKnPENbSnjHHg49iyqq1T+jHd5DB5MHcwoEvBoARaQbh3+ijAQwYE
GqXePJjaRlsQPALeF+P34WzOnifuxKzqZKwvbWpMSH2t7yD1BIVOUUY+yMvyGNQxHWF2gfmZm5Hg
dRKSl8Ey8hiYHL8wtNI0C1Y+8SkdIA7oETjfa9TkXwf3ONq9CPRPbmkHTPoc/s6yk5JpRTPAa5/x
mLEhPjE6jCDnJ5NS31YG4iFQ/YzsDxBELMH64wSlpPl8MIg7oe3UBJ6UAalbqWFCTsznf8eT5Xkf
LDjI/RPtgyYp1NMJrMzzKX425AT1et0UZamfDEyWuP/Q1nO2LPKz2TL/nwO0GksVLuHlj6XGbfbm
+tPsSC+5h+ymYIRdCB3ivcCYQBGeqYFL7ZVBZqrWwy4eUH1y+66XylhWGfCSA4RfRu2HztEE4aDj
SfZ3/rnU8LqGBxnb9EaHERbiI55lmKr202zxncC+UGGau377VaBL6ZndAfwqYdMZw9GLg4icn+AM
Y6AtDWfI+iQqnCPzy9MjKQd8E+7BpM4ClOCduADcNqGbOeChOr6xSw9CH8ir++BsX8F6aJcY0HiP
61Xe1GqvrYuth2Pnge+gCliHoDwXgn7JtSi8CrQpMy2j2OTGs8JrMM8fRYPsqfwdrkDj6AkD123Q
ttmDk02ZD3qTJbywxa/BGLi4+k+NjNzbvIvyEe4LweYFcP8RByvzW+UqnPL3yqlFTxeygCf2uSpE
c1u8xD+MgrUb+VRiNEN4/oRhcAuyeAQxDvUOoFn7V89vI4MvM8DAG1BHJaaXCk9ekuziAqbP1b7G
0cGQJu02nkWMMkXuUKNKGq3UUj8aNYMFfUhHUWodCNdnoSWttEmOcso06LDFyiBQsUEylQulwi0Q
LfeW+4nnnUXXs2O2mFoK9gugPcXWPX3VUnUda3E/FMprGCmsJxVmyhn6zfblmPyTNDvsSnwksur9
vF6DEERslP+uP8VmWXF8QJhUDFMpoAyBaO2DC7OVHZGiFOi1c1V5eatiQSE7N3eR5Bvp7o2nqG5H
ku1N3zXBxnKSas7PelCLzCnR4XlPMYDM0BgBko5rRb+PaNTNjX1thULyuwFHrX7QYomUoiPaCRK/
kftYb4Fj6zsQkBN5impHo74AWxk62A0eKDgcEbV6/2wCfze3LV9hpxlefmrj6cY2z3tiNci5GbUa
gaZQ4uV3xS6xeY4IrEvqvayHEW0HEpW+Kn9B9gxdy43cBYh6+rgRngqCm2dQdT/N1tljKL02R3T1
d/p0y56aDPAQO5GUma0doGbQ7sFSgC6Azuho+YtJncSNfm9ZmnJh6d/w8mbF9Y7nvLdK598JNqN3
rw5jim/jM/zVh64rt04MjqG3yIBaF03BILmzPG1kQlqnqMp+m3KsLkrSD6JBAxBtX8ItQ0kkQnou
qgxZM/04QW0A4PEAiE76ntOabE4KIa2G49l0oqRHyA/2csgnEcq3nGeHgGq9XR6CpTDLv3xZ08CC
vn3ZcNotdYggOoyhVW35v+isqldQMNi5V8ncDK+AHa43YDAC0az9dVUePs+Kg0VhGvj5I5drxBO6
FPLipIpFKc7aZF8p6IRx++QRNyd72ikwDfAox+rmNOzQ3ar8uX5/X0h3jkEP6O4qoc+/4ManmiKf
QGabxMh7FU0MyJLs0xJ84IBx6IYPeSryjv+eeT8fGzwKQ3ms+iYGBp70qoRbOCjNyJkgQ9b1dOeQ
xJDuZUcuxUIk1BJSlD9bY9I9LVjfr3DsXvoqt4WJvLPTmEt63ib6c/GVLjahDOuukGZekJV50R48
qg0llFb6h8tFQdpRMSCpEkd+V6oNqbySlORqUwNVicIfLKmTnKucpwcsw3qUNCaDj0eo5s7Qq5Lt
Nfw83u9SfnQqXp+tcVCwLR3L2NWp1BSZ2EF4AdULVsF7aimDBE3JF6gc5fXn8bnjOiN/UY77EWi/
QQMPsk+Gb1qOPSaUkJX8aqv81Ed1UigtgAhRAsKH4f5/FUNCzC3D0LfzbITMSomFyccXbdOjXu+6
P5Neti90kfsQaMAWZlc+ZO5mz5QS1Lwljmix5uT54roO6VB2ORNZAY/9gmqGekrGPUwXtbQBmUDP
q+mfCF7M+SRYx26Gmzt78wQhg++I32D3G8mWBr/L9Jjb45sRzMMERtAyNqt62AOWz8EXdRvB8gTh
R/1ypGZdsFS8sU2MZ19yK9+HJVFD0o80j8zooHpgFLP1u6x1/6hEE8q0/b0LX8seACu3yYdsaDYy
VPx3AfrkOLEBrlFlTEOUJZ9bjZeD6xSaudCik+YXZ5PW/oc63OWLcNuS7OeD9r7E8wgu8Uf1/Jw7
5P4mondKvasfxfRukXn9TqfV2lvcCfyEqy3gBqD8zJfJtmBmrCyzdWeHDJYqgUwq4Op1xmKTeX4I
832sUFJvIlOTdweIYF5GQ3bQ3Y+cMDrj3ZMbVXu0GU113vNFDlQ2hxd8p2T+oRs7Paczyue1l7rn
Q2iVYz9kJbv5C+PkUItvyyW/GLa6Jd4Ev1N2EUbrfdevlx1pMw4GDQJp+Ztaob+wgR5RYK/cy+YS
+FKLc1c7YyUnl/e+Qgg5CYN1zuUnZdoO6Nj55+dyHo2z3XUP8Pn6zyr9/Lqt4ylnvbJakZYGhOqX
RMlvjBzodCPIjnf2ty7g0xiZBxianiXmQPOAz721ilehsMziKtePdJt0VeuTjEzoojHZsS1Q3u5E
ZKvp+NIZsfrPamp8fpGXCXtrZ9OYF7SoOG6cAmBB7f8q0nRpcdR6FW5FGWESNcWVWxm/L+sc70xZ
vlyTjFH+NiB0FJ/ob/kRTGsYu+FmEzK/kjd6hhSSEHeJ7sidLPUeGt7y/OrLUz8xtw0cgPx9LRVo
aXkX5rUkxNFZHrS7DNcduw0zG6xBjLiyiRWITfDZNcZoCiU5wDZRgmCgDV4z4tiWMx9WcdbMISsl
mdWf8bYl/QnR3plQhRVUjRzdfEQUZdwC1w5ui/3W/4L2nOqrouF3RfPr4g5xSXgZV7J56ZLXwkGu
6ZElzWA5LE/nkWb1FjbrdOcJMwvaMtdK+PiMCmvLjWH+rWO+fiXN6S8W3i3OkVFV1a9JzHZnw8P/
KuOObx39uX0/WZBB0QETB/NdUnDLt1cVhE7T2IjHb+ubSOwpSrrAtXSLvv2nn9Va3EClwSc6xTcV
LqnfWhcXO9sZnVHZnZQ1K2/IfEDStiYfnu9r7l+JzVa19+abj3Dl3hrSPPR1Ncfu5Pv7ICHyq2ZK
+72Uq16A2jZmBBqxgcWHL9emZfyblWUsByYqQgNJbPfXfMdlcOj7LbtXls0qOXp9QvaYAyZjNNcQ
H9J8DaDfJpGyn+/zKBe9h7tz+YXBz2BgQ4No/lzcx8/xeP5h3Nmkq6uAyzEdiNV0N9sP6xYR+VXk
c2ehhdufqv0lEEIem9UUfdGfOGaTvfHCINPIgnbU9AxkAzHkr0KsQ+UAqBr0+bszI6DuOezFa8d+
0X8zL8kX7UIZNtYqWrBCStm2hRISXkZTqtORDZ008s58UI7+rJopXeipjbhChJr8pSr1ddYZ66ap
pCRcKO/XOOQkcwlhzMNn5yAoX0rT+BuCL0STpPMO0O1NgnxBE066cqgT3q/NjftRd9gOVooYKe4Q
RpTPKO7x/qP7bvc1WIIi/PceMpL6HvNn8uzroeh9JBnHBmMdiMmsDkpzEkqJmBPEEj6vuxfMiU6j
fHFVQA4/8D/h0EjnZbQaIBkKlJJ8QpcFpmQC/7XBagHHNOdAjn+6qJOevbs0dHNCuqe/VkXH70gm
vSJ5WzB25kDxUnNjsioHP1gsAoXwdC0vssO5gtXAHXhV6XOs3+W64HKDDayuqK5jPvbSuWPi+JTO
BWRlKE0iLk0OJSMCavm1+iHJ1BZnk9pWVS5pj3uWHLgbmNwu3Pa+Zc5+axGbTSYspEewZT2T2kOy
C2LKRc62ZreyGWsHzcrqCZULGEElnRW/l1IU/XD1ECEpmHwLCboqLIT6UFUEMooBET3kHFXDpkNc
3pL9aP2dUmca4BMKNpsAYhxIKNLSE34jmALDCpjRHSw8SOgbQNTIS3kAxe5Tfv21+WHC1tfhk0Ad
JEylH0xA5H9+7YX+oMv29DxbI5VqsxzgzyxAd8PahqrIuNKLXCS/x6fsjI8ULBMsu1xRRpprcoJ+
tMkXRmUYqXQdDCNUMMsyZTGAsbKSi0syIoOUfaw85n9OsT/RdlGBMK09bKenGRQaFGsbsTKxb0BO
knGbn4kARrbMWKSxF62wbweYgDHHucpFpE/yhQ9AYk/uf6KBU/4fi+bGCiM+Bpv6K5hlEHFiWlDr
y4aYFqe60mD2qtuNTsmlGxj7J1SDEEsjSHhtKbp8+UhjLfen9Mput/+9AqmcpnYmCQjFdusFupIw
usZ1HVqOqwpBap6niS9BMOzlQcq7fL9jr4VintLNdkPOch7LEG1Qx6jQFTey8WmLliBrFH9n9qgB
owSW0/EyWDC9IqS/KZzsDQT+FcmbzQnsumNdFYdpg1XLUjw9xta2WnfDI/DVgjRnPLgUKRMthjNl
p5WMjDshbqsa9fTgv1Dcjyv7cLLnr66+BPhN+UKtI7MqzpGfCh0h9Ax0CCepcj7Clds9yspWFql2
C2pvlSVFzB9vc0uoUSWsnsrjM1tqN1LFL3cnaVnHOwODqhG2/7gYwYCx6jA9lV5RB73IdqXtsJP1
BR8qrJD4ztFdECu7r5DPZ1NWveGMdOPcyoYWTd00D1Tzr/C4YoIhSLx3cGGCFpG9BSb13eWs+GI2
eQGh4BE5AIvuhzGhMFbeQxUmC54z7Qp6kayI0N8DigP0ROVMTqf3mqdDm6ShhHspLh/ccdNJdvcg
dopiQ0F1zZAa2uQXLmIY7FYEl8CgtSxBzGnjACqaS3K2Rgaay9nd0Bvq9wY7r2us4kIYucUUAYYE
Gw8GR//sIdDA4iEImoq4HBK2DcYOEhm4UOBlJgPjlwy/Q6QULl5P0ecQzmf2QunTjmIkrryJs37v
NZuBuNx2p7GezPcYB4o8mjU9ewDch5Y1cKXD6eYuV5eAc65CM1ibzXeXAMYQ1hBVUPhswDm+JWjJ
4HsAkE5f2lmJsFHWEt4OzRi67FGKDLhUMyXkyhiawt7vitSxZ4H0SA4llqOw9sZ54IkGXBTMTw1D
2ohpX+ZoVQh11i41OYbnoz69eOyoVHJbyDfLlBTg6EeAzerH/jOF7FriL2LgPttav4kpcdf02/Ts
WCNdziYgkDFk+GYnJ9E7zXtFYoNnM1OtP6TRdw6xkhp9xTmUXVojnBlJvlmGdaX/8wC2WL8A0Sd6
5BQ7IDjVgeuEjI7W8KAuzjphyRq9v4OrizTEl4XsbftvM0Mp56JBzPcog2XDvNCxgwM/vXDiIjxt
OZqnJenNbJ9uPs08RnR1N/COXptEmszwvWCmctj+K83Kdkq9+sBtrxtI5WVwFMvjWApCHHifKtxR
+GuWd0LnnIBQCcHRCjTOdqXfTcR63v81ZNm7uf7altIQ2zZMxpvq7Y/A5yw2ZuzCnAzk7obsB+c5
2pl/PFYPaOwz0UfG/eGqVELFPKRZjFVtLORB4ryPszqJb7WQqISEkeI35k6Zkg7wT2UILMC7Xf2A
0RCJixevM6ZcN8ZV+ADTLM+tWVTGjbbob1fUzVb8a/W5089m0v5TKZqwKbCxlax+FEdu0EMxE+Fz
d6OvhQMCaMmf+1dQ1Pz2UoozBuAwLjvm5QoKPbqPZQLe3ZeQcvFQW6HqgxjKh7+s/NOJqJlI+qXU
TDx1an4pCoOfGHYOhtfo1cu6zsxQv6LhaO8MNRNdHsG2sMb/CZjahp7jvW4p9num/WQP3gzfBcpi
3NY9bPFahr2A6/11a8OMB23sAcYUu/a0VtsZ4jlBbC2EGuLR7fTi/gDC9hRRwtaZMxZmv+s/LnWB
Os7LMY0/FbWPMwDe72HcOjYaJ3EXPtYNcDpqdNDC/JHqvczk97nfxvZM3NKhR6aGuOjYwhPDDuRb
qMYOG/FJiJw3c4M76mGokAxHMwJ4H+zSI4nZHWfDZ5dXQfEMybirs1ekcRaTBHa/VZ5MEp4YflXw
P9QJOX1jqS3jFsxyPSZtOVQpubyhd+j3ex4XlLa6d8SmmqO3j/j7YsJDzRjS8mepvQ/nVzj+f+s8
D9ioHnE2dtqIecjeoZb164LbWFj/kUh6HBntEjJ8k63VvPN6D6Chh8vAAeFYgNzeTbxcAEqNuqRd
I1pzDcb6iJOcy85j22eTcht5Z0LkSjK9/zqR+0winevRhx88xc4Lu12cfr+bMcSGgVTS40uU2Tjb
dC3t+mDQNHmLOkWqJ/Qc1WRUU++ZCvqEZna+RgihNjwWYqwAL+/ItwL5THKJ+Q7quxcKy+CNzHWp
giDVmS16/hiyrFOo+ncBP5iVTXjMcIK85eikfweVHxm6NVyGUhM7+ViTQ2/ctRLBbjkS5t8A+glr
2MY6GhSCdgpZKMv4P4DZd1qBfoW29CudMt5m+ZmLAsID7lDgJTSDOVoLrFbVArmizTm+wk/nmHeu
Shlw2T8QyV7w90uHvBt23xAUbRCkUDDAWFkSKZ4i+FlqngeV/jTScG5GI2BYdpn3H2wgJJdmLYD+
wQSjhenGjn5i1a+dOJ0vnB9KDW2G5Hs4jGbECSZsQvX89+0T/l+Fl2l3KJxdOjtSrEfu6FjLj9d/
RJn2svknI4MDKNSKLQ7QFhR9U0lPVfx2xoaQT1UB1eXRgPPn7tZSPTqGaiRUxkWBHOMBlczaC86Z
Resft7z3mdPvpXT/YCYXuxHMT81PtlCv0ilXvvRbmkV564Xj151P9lCybYYrTviAU5SqmkIUeHMG
ncOD7w1PUMWNt2AkJt1V47hQ4Vvznm/lpVo0aB1wBWrY1ubl44K8qBQdrom+q/Xf69O7FrYf3JVL
vs5pLKNIHkTrYpYsNSh29x5NkW++PIZM2vDHQc8ejmHuTwQdNPt8xKjHAB6HYg23rNKxRjndZSZt
UrWWU0TXSH/KjF7I7ojuoswURI+nctlq3nC6LSmqWeKFx5FLxJgtXOuOTrSFUBsZOJvW+KkbCTmM
9H1j8urEZT06leqAFCoJm45KAXh1XC+/Z5lTmG3nKld+syHGub6qsqvpaupHjh9SkLVaYOfBl4G6
yRKw7cVDuRONOrsd29bbzfWH9ZfBYkTkAgWnYEJLsdp5dnHrDc/z/tkhU0qveXVymH/b1BtVYEV/
j/hZrUaRw8cBuqPUTiiItDdmTCZI8FUm/oCaf7OnGuzY4c6InhSf+JWAgIkePgSYtXWc6wLj1R+i
mkc88xwbCdj1Ehnei9q0xM86w4Wpl7E+yq+O3eoSaalBeMoOVSeHzh3oG/EmdvwZGWc2Uy5AZOJ2
xEDjak9peZbwF3Zn0frlbnJu15emp8lcJazDWTGx4hQZScbGHOOLhAdgCYIpCxl6sA/caT6kkmWQ
g8VnsEI4G0x89MgNjjxHqOsrzYaT+v2VzLdWBb+BXHpdrjezEgjfOb5+SlZYtrqUbkGHfbpK67bY
pZCw+ngM/IR8F7xWJMacGd1oaiTO0t3KU2jItH76p/3u60IqoKpae9Zgkr+ofNbb146E+auZif4c
JH5zkswzAUj+a6rVgBhJfl2rgga7OtVTVx3ZSj2xFN5sqpmYuvhi/dcE3VE2tPx2knLEXE+wnVms
O0jy+673fVgEZEdj8wtdoJct/SN5BvemOuog7/q8YAHzieJ81Q4AL69aXUGVbaHAIO6AYf/ug+qC
0GqRSPCl191Rrsbhf/VRF/EkaGXnJ4aIS9VxQVYEbBiCnUXS+p370C15a3hdDxJEl1emOvlqijbd
l9Jph/B0Jc75AKVPdcwACoTG86xECkOIsBbrBJd7oTn1FP7/MI1cWdTb30FPQo/sNdsePHU23nMk
hyYRFoR0Jv0fFU/Q9Iz+iVm9AQAgReUwCKYpgFeQZTt1XhN09UPY6cShLLiwzIgxP+Jqz6PXYBMW
G47oBHJ9s/WCGrjN1afLccBi9tSE9ESdpwKVwR76opt6abPAAft1fR3MIdTVa3fw8BR7ImNfYUn4
sKrQBKy5WF66VNXtKY/HsyWawEM4Cvl4t6ueS+ZwqgXE2ebiV8T/QLcbjbt1k3joH5NFlsIR7kpH
koWS3r2olnmrgg9PJW6K4cE8+aZyGbHsl6pZXbGT++eO3+tjBZctiiJfyiPGd24JjjO2x+VEjqd4
Raal3sc9cQk6F85TSs+QC3vwxZrQdpv7a6y24wvN2prp+H7w7Xm6r3OGbBvtz9b2R5aP/J9sczGc
rXcAchFV+FvhEBavXPOjKMb48qE6vrMG5rBL4iG085E+MdyMSM0xYeQmPmZh0ScR4sOZpYQGjSii
oAWBw5v6nkSlGzkU4nzBhU6I/XgYb+d7nEUB/QY4Y1C14+MZG/2/MT9Z4opM2gcZ6nvfZrEccePx
9x6pKW7WxR7IN13/kRgt9gtgGiF6skpZHjATHdEmla1TUYvuSa4ac18or6JgCOVxKFXE1CwLMrGJ
2oYNMDCW/mTacNhK4MU2lEEhiIXtL4K19spsRHzTFXlJJesNVFFn6EOduLoQjgAbOZ7XniC9fGXN
QoQGUT+lrKqDMifBbv33DlRw1eb1dSSPHZSjDOtYz7YAaRJP5fnam3JA6rnaHS1EdH8yE4GGGJKr
FN7ADwkWSx0fv7eezYBfxfRgOiAfD9dUBbX+pHMPvzqbaJpzszQWaexJNlQLFwusD8FkQCyLmqNM
+xZyp1E465xRPxsvAAwIaUNBYSKpomEMuI9vPxowac7yqOjFlUL78GfLMweAwSwKj0b64i1NrsED
q0GSaI8UbQEJq6Ov+PIWPHNCvVyC1LRivI+UgVTirQAJnS/ca0HIgP8hYVXCFfd1UoOP5hnH5v8T
SUwIMhapgKVtOkDV1U390xFgfSX8p2ra33+TLT1vYR2UUbJoSLq+GdbWc5NevhFTZ0Bq8Snn0tmk
GBRJiwpkdwzDm8QTLoqWdi/1piiFiBcgLyEVqoQlyNTMPs+A5Y8yys/px2zl3cJqq78gLbgdAY8A
awPHHhWydAZfdj88oPlvxJaVukBZHHnoWXJEIee4rv20ScmH4TefHdzLJ22IHt4YhQ6QSx2qd5AM
FxMFmhL22iYXFsgEL7h1mncoX9WjTeW2Ky3+5sVnVvAEJDZHOzGWHowwzVZKqM9HY8+1gX+SZVSA
wYJvbHmnN8v1mFNICTTKnLifCqvTIMmGMOzPRKF0eofnp1bYdXtU22FPgykpc6ALVXblSHO9Yp7j
CaRuk9perCnAa1RV+SDemJbEQSpRbSHccMNRkfKmjVqBTOcuWjyW3h1ewzAZe/ThheahyYb7qPTT
P0Ni2ly81foazhS7kf+JZRBuMN++9Gvo3DV8E7i2FzLKN3qQ9IsQ9TqTUTXeNdnQzxudotcGqEJT
1ThsO2G2+cUdyPHU4oJ7NbFDNuXze8jrkF35cPszNtGDn+uOrpQaj8fgibutbU0N/GDpLUeADNDQ
eOyVmlpFdnxz84LLpCgvnpeM4j/Ce/IOHZGkvLSUP3TH65hY4NA++M+oZ9lhEIzThVmal0C/4I7U
jbnsqTQ0q1x7an6cgZtpsyeZzN7fuq6AtG6PaiDpKpGkWx41fR07kBoW/1TeUrBJpf5Hc4VzXhYm
7gOTqNU/MvGYd2030PWFSo8xzPEZZpZiUfs9W/dg9LWUx8XwF51ylKkARMTyBzousVZFcrGdVngL
qwgjzwvAWTH7MTv4QVl8bPEuV+KzIaNb9jpS5mjzg2WYUHu6g9c4g3gz3mMqhNmneSDOmAl9FNEb
dLem7U5yTNq23jcC8niE7D6gsDZ2X810lSLN2VA1+TCtQ1iXRxqLG8FzCJXdYuifQR4WB7VXEZgi
voFs9g2sTuSOfGo2vk9//10AXaCspwLl34ING8qbTtECij8TXiVas653OGB9++ZaFT6GL9KfKjlH
utPZCk31JtQlP8SVv75hTSFuPj6lSJYZCfpZq0xC/Fb8FcRf2ZzHEB+H73DFxQGmM6cX2YWVQ5LK
nd5Kng5j3qjlSgUco++r5+XLGv49WbN5mfoHtyhl09BPOuej0AMs5W6wl9qNAW+1JbiEZc0sa2za
s0fXZLZ4cRLJBBrPZSOsOUXxLv+/tJOkxVVOamxI3LO+KgTDy6VH+RGSLZKB/5LPsKJnmMXq4Lar
uj+d7d6fgYy46psqsaRXpwjpo3k+mq/VQ6m7Yd6hb1KEriwOOtHZfv5iVRO84bIezKjIuBFIi+wy
iqUUuoH4HgsZDs5daxlthNNktVSFiX5V7NKmdlEtFqsmjUOS+K+XtVMN+r75p7lSEEK6jr0t+Fn4
KQV5Nd8uNA1Ip6EYkJt4BXaGcyo5tlPh9wRLBOOjb+qf0Gk0/H0uakqKqFIIlLnWvo2fb+CHKdLU
1i2KIRkEDf86IEQMdniJF3ecdHkZEySIetA405SuNYNK1hcMYDgzMoCS4YRLj39IfrpVkswCRDPX
elAkeHchBJ/QHHC/2L+kDLwB7Gy5zRXTdgbBBBKE8GGF35ZyPnygPNO+NcVzI54w4DBDmzKGZj+E
2K+dh39/MZoqms+oiqaQcTac4Qt2E8H+LU+dWj3SXG5v/zfpWdo0PTzgKCPi9v2tlXN9zLEoXx4/
Jxs0KMgi2CyPZBB30hu1LHhO99A04ck+t+jrjwiZ54TC8mb9z1GQKuo2hu6VKUxtCirXfLejFQWB
5w0L6odLFkLbk5konlFfGzifr0E8Ga3JN1pwnrwyp663L0XCQR1ulBAdcFFeh4fYRF6hBeSrNu6F
5VgFAdreJFCv9MByNIGheXPx+qPmirj4f79h2HTGeuyxiaqaIn33h//2HeotSjafXhiaB0OTbw48
220Ea2U482hx+a4IuYDOd9bZIS3v7g83zw8/C7UNxYcv0+6fC7VSpFNtFI6UQvl6PblTAPJNnt2a
L+zfqsYIiiQuE2fdLJdLNoWwcfb2nr2dtgtJXSAiPDxE8v7GjnTpxsRqHJsgiphD00F2pMTKDIGp
0J5IDwOrSmqpIHJCGCk0oU0CBsDqgFW4+Vg+Z94f8wVvOMUi8K+5XmYVs0sHfUIrEz3vvBX/Eo5t
WyTriRs6Z/4dpaP667jgjdbD2pVz7Am7jenjHdkku9zDFE9NMvBpPtGm0y7WNGDk8JFJCjvwWCH8
7McW/QNIySk6GKBFfr+VPc3iFmaDWv4CpVgr5cG16zGy0HL5Jz0OKSJg+aZ4II2R9I2s9vUOMAAj
ZChSdhQ09dVfuDRWkZavihAFrsREEqABeJLY7d4lFdRhOboLeKYw1X5U7QDl6If1NLaKIXre/y/G
RweiuArRR+w5843HhVqe3v250dhQ2cllblrVJii6WInsAAcSjN4Mda0sLi3v5MbBIcbnrr4HW7AL
q93H5izP/jKzAwegq748E79/EWpjU8dvynQ0OIVUIgxiU2+UavQzefeRiZw9m4p/pyg9SbS+vem0
5E4Ja4K+8q+/AceCw8ymaByighDU5NaZKxMTYFPvbu9KPfnCTAbrA50EU4GlqUpICytWp3QJHhRN
sHN+yMNB2gEG+AzuYHmG2gucp1JSl7JQWlnHiYUur6R9SjDWdjh68kxE8ga3qnUcimGoIchuoCK2
oIGhqlPlwrBSgevyvrly8rJ4KYGJ0Ox4b5AJX/Xu6X2Mtnvb4bwKOeqRYHotHn6NHc7pv6tt0vrZ
Ar7DCXPHgxOTAlRJ3WPqf4azRRvtv5TXwOzth77twJgkzMuRHtY5w8BQdp8OqJm22qTzzOURHrMy
XCKigesAnpYxCACs/Etyqf6ZqiwWPcISWV/LeBc9mfbCYFUf3lx2WZBiO8ZJClFw/oU4qeT4fmoA
GSI+hdlSRncqGTzEJ0Vq6c3pO3QaiakEj8j+Lkpkhwa+CJMu/jyX11/F6tdql1HRH09H+296qgZ0
2ER2ZPq5ALrlVyADNEBd9kwlXOqLnajs/TrZ/chcW8ijn8IPbfBSc1yPmrpb5sh8MnI7t663eKXU
GhtWIOCn5Wa7sKF1dgyExOYV/VRUHS0zCjFrHTuBTiEDXYoi9frpjNIYhiwoakZ7Xy4tSIaBVq78
BS6K1kYxgxnHaNZW1figEs4guEkoUILQgu9ZXstBPYQanokcvuFxRqUrjsWwEd3TOiJoWKDTy1UQ
kzjBi3KpeZf7+0zyzjAiBB3HASob957qI3FPAbYiZ1op0T1xV5h+RT1G/kMvFKWswG7yEHKRLg6X
k/JB5ehJCH/owboLH3TYuq0qOZeM0j596zSid/bJmyE7uoGu75pctKARkHkGqs9pJlMoKyadmm9S
JzPpM7bZTaAXfcdCH5+O29pVLw4Vxb1pCCcmHLncqzyn7mVNT9V7775521O+47ox2/5lCWzHLiDf
xVGZlcOwZ3aM1CHXUgKLeVpwwdpSXbPvYVi+LvXfuizfahGxGNL8ZEOz/iiD7EqiIjbbZz8HolEv
hwIkdUupKlzT2EouNQrkiFa5FnZwYjCr7QmvYshxTy7fuIFzL3B8Xe5OmT326EAOOdwGyi/WzNC3
rHgQ0woG3XmgG1Lx7WpExZgktxY5Tmb8ub+d5JmqOsWq7spx85KHJxOW4HhC2WRKtmFyieRhG4rM
VEwIq2DyYMCD/oC8/IXZmswPgYLrgVAY+3cWUpjS/mM9EgW34Imi9zqRqXLHa+a6gWn2Wb5yXFjS
lqks/2DzmRsSEveZNieoQFwmF4ETbRsSLJ2lUl8oDPtq96avZvAWwPzdf1bhmD9FSxwNR9YIr7sX
AV8vxiDsTbLzGrynWEqFfJTU9aGRUxsgQyYUXKjz/LYXKleKahe0ArG9+VcFbNgNK4RWuwNt9/xG
YEoZZxyvpW1cmwz+QCxyfMyfAShYK0LpCVTPd99nnZl8QMG5fiZ0dMi5/geN5WP43FKIBBZS8yOP
Gs2DNTalmB/XadraYnNtO4IGs1XPwBky2vawRin5J+mYIKuTtw/QofjXu78nIsJSbstcvBH6IBww
JE3FJ74oyxZJ/3CVzPO9bd4REMsRI3YWgTYzZpW1UqZU02ETqeEp+L87qy1vDTzKjyJWNT0AIN6Z
PoGRVxI6e3bELKois4ZkI6GQ7J3cgGH+JlQBTReeyxc9vZG75Nb6Ts5HwCOo0YnSxFcMVy/avGrU
PbFSFeOXTetUTNXbvuhpMWItwmQTrgiJg2amE9V7LJ46hJq0Cgxzk7H6xcwfBNFpxnmeT4p9vNl4
dJHKQ/WOvgDGzok2Z9FzAmI4fv6iZVskZX2CY66rDN8/jjJeVTgU6Rqv2gh+sw7/531fSYc0ihxQ
KOXVwDLkoozTxC4nMNfAbwbp8RlcDAdphYgpZw0jtGchp0SPfBkjk17kENbTM8e73dklntivJjFq
aj5AD80AMdBxGQz7mmNxgLy9PX1PJQUcbTTsUqg1y7G1aY7cg5VX+B+vAy2EKIMRn3Vsg3xRKOaR
dnoztnUgy8eAXdLFb0lLrTInYznQ+uCVSNlxAgOTr1Bj++QivrbwKUbw/S6R6qKOFeTlo3Ik7uHz
rMf09pHpvVZ1zYzIabuaIzejVHEzOIFe02u14ZNO0Etj9Nk6b7ELFDq3uAZOY0Wt1tCGkBG0szp5
kfKuLPMRwne9NSpjRfnSHv+9y3pGl9da7yh0RphNv2GhEbv+L2IqNc+bx4vi1R0JoAqRAFHPkhhO
E/jYs90bQLYDgwtZgYhaR680kTdoAzR2zk6BB+4lJ47RNvSpK8FftqV/eGKdxoY32Fw3UGhsMFCd
jVgLc0TyBX/129kmnMgbGo9gZ1GhAvfmH8fm+5rv8AjJBQjMmnHEIiA7bH0z34RTxMr3kskIZ3SA
kGm/76JMe/Xffent5LHF/pBhqZ4JsdkNEe9w1KPA06i8F01QsgSb7UXRXtz5rsIxqyb2fAYI0Ng0
yvCIkXL40leK3l2Oa5mcOwBeJ7HLZnbrj+AVxaLUde5f0gfoPZYqJCwEE0DT4PVcut8uPpmn2eBp
Uy5rFrSHghbm/quyQuu6jxU6j+LW+XbMcjaeutrhIY6OfVImXRlPwuzjn+9rWgdpt28Ktt6SNM5a
nMNPbOi01629bTzMQpt8eLfsTCrZvdUlSF14JTX+MOkbOVjaNHIwgL4IqPgsqTyo9aRoF4Wfggzv
YNzoFdx00QcXjFT4xkCFnBPV9VbTx2JdqvvTQMQscN+AHQLaPkUoQnrw1fNx95yOX+ucnlSIZCkV
gXpmPhjWTWUXbhdI4vKJmFPLCKI4oh9V+LVGeYbsfzZYifl+c+D4iHR5A1M9xNwen/zbifVYFjTz
M3lEK2WK/bVuP2Ks64G4xAXLhrKkWAA3rJx8TNKUa8KH/RDBQBMeGrR3OaUN7iFUjwZEIZdYrdxA
DaZtkjEba3sJhqps0xog9grDla5vJ2csqAHOzBzyCt+48DhXmC52i+WlC0+dLdzAU8SwLIEONvIu
wI09HrHbGqy8BKPci/xwKDjDzGWacIzPTvfRzewt6EavgKX3UbM5uh9s3D/8Xc9lIWibj8KawX13
fYlZVW0okqlo1b8RBSVGsiNPI3lelN49KlYDymZ/DYzDjo0bGsI0P3wjUgY/yHxwRDUwMJJKBzSQ
5Ux0xPhRuPZnee4o8ZHwJbfJs1c0zOtnjp8CBBn7ktCUKiwPIGq1oct+obhc1bJfWYe85AGH8W+v
OONlIzMG/qLZXbC8Iox33GAU1n+kjWhXaTv0W/kjrqEInMBK3dqKM2LvbvBhq2bUQQvk4Au1MXFx
aEkmefWKhyd8lfDmNPUUAvN9M61zSxdl2Lnr0FICmxVHWhMbgVVH1NstBVgDCeHgKjZN2SKNrCR+
Ik5O+CX2NnKqOU3G9l2iEqW6q+6z/aNwIx0vxHGx9IRd0/B5+kZrYTkFNG85Po3Zoq9VLC2YDnCj
vPnUsWS7H6brteErhKOdD5TwRgS+EhpKLj+izzOx1vEbTpRurtJE9W8c1NptdAkKYpiUj0rdTutA
PpQe4GK9vhHW8UoEPyDmxPZn/BbBqVXFccQ+Que5I7Yi0J63icq+kNDwp0zzIPh4jwzvufXoGuZc
212/ZkG/9BxFkEdSamdGgVmwmZEDZ2t7jkRWYU62ZnLo1ixZnM7uJ2sc1QhAKfWO166AcrFRBAv0
5hNwHirCq4pC5yhF7UW2oTqzwMGFgldbPNOsRaryR1Yb4tzl21bnhmuv/U565VB0A8v/VVW2XK0+
JqeSSCBl43pPohRFY1BlknqI0Byj4feyLA/RVEjkqitzsnZEABvimBfrXv9OMZNi/MYk+zk+p4By
zPEPKmJ2GCTZ6XgVJEZ+TNY2R8or48toeNme3nMHIbXGUf6p7klLDDT/chh5u2a87F8jLB8JgmKo
alV4FZBCaL/T+IJlGiiGnDpwpPVRdE2SJPUY/u+TjksT3FTO6J3csAhn2Wr6WLFl6nbaoc34NGNF
EHo6HmZ7beCWnhI7kdHXqzI8riY9Hm5/xr0fDxRB9TWfAPrVq7VORpxmVuY+vjI7+4Zx77UTY1bs
T71idmyaQ4WmVW7boIvIWVH4RKGhPJ8lIaedijrF7ZFjMCog8Fbrn3mAQruTnsF8/Dnq82/Nffz6
ZQEAbvjV+wcZKDSRKo1z+RGGAcWtQVGHDDdMQReyt+J5V+fqzJ7QN5rlU2A0dxkZWFO2+ufX71Io
1uqeF9OCrOd1ijiX66xdzdeZOXlyg6XbFhTLS18g15+w8MkuaZpoV7hQWNLiJhqnFgC+AnEGuLhT
7dlqiU87vq6GYpjnyaFdS1e/Bvjcs0eLwqxzWihSFyg/JaExTZZCMGKq/k/euYLLauVFF4ySTne2
ZfVXpsllgY9Qi7HuO8tkviOUHiOcY1OzOJ7s4jRQhVrXyKswfePsskrVGgH3kV95ermUmthOxVdk
QqzuGQJO8UABOQmrV6MdSVVfJOB9d+Sxch/NlpopdWWyhI6GRfM2ZrLrGI21e92CuNGc0AZ/Y1Bs
PVH3hxZAliELL2jDkuSCezvw5o/Q3bmLEz7fxblTpY142bNdwnoikZvpcfNpa4vUmG5zfhxmZAo2
E2Fxkr6f4DBw7wz4gzbLk9MNCAr4hs2FjQ+Zj+bI+YDb+m/wRYkcYQ1W/lnnLnxneNkvfTgYnfLB
k4oP5VopsiwmgMFn3l5Mkf+JxGyjIQmJCqKvJGVCvDX0hrcDINXGkMINOEfHN5LKwjeukT64p4u3
1DLQTi0F/I5yq2q4K6jXPqviY23+Vqg2mT5nU07kNdwt8o5D8FkjPZdFghFVLyf4zV6W9Stiw1kV
Dv1fY43NTDr2W2MN0/rrNNqtsa/RqDYNxeQSBSSEgWFbGQ3TuqQ+6iTIE2FEpuQ/Y9VspV9gW+ms
bnvE/BXekphzKHjWhmuaTZga1uqwJs7kXJfYE73PenWc+sjirrJxUc82Jk2KM0bV6mRMWnySS4yZ
BJaxrhFl/JV2HAi7GGl4wCPhvztLWmE3mqvihTWyN+u+iUQSvWi59jUo8ielKU+SbTX1/WQ85CFf
SSXPkn7JXIKZx4IqwV1K93v3P47akaT91WkADYBKtvpzu84q5P6KEE6KIt8YLOUMrS1BeN+Nh7lI
oIvb1yuEJDxJ69saBZjK3+RHaqhldlmRrFV6BQsPG0BTIBi6ud/yDHQG6gQcLEeCzikzT+oZHmPP
swzGF3Oz3iZ2vHmbgZO5wuTAR3zOeRcRfM5I6H43XEulwkSgLCNAWH4ZNhXdyrr4O+c0imna8Z/U
HZ0eJUq5jqKBXAK9bpojBUH1iLrC7rQm45EsJuB1CzZfqabaphmvOGRwDTCRsKfmW3SBKZFvxwA4
1fRoO3fRq2V7ZEXbheETm5k1WSNAEdkdbJE8+PuGscq8if1Z/dAgGAzw0zBVizUzOSEmGUSTJw9V
HisbrPladQ+LYsC8A5jrf86TPDpS5I+sXD5O67fnrWxMw6bOqkbOxT38Mb82yBEjkLVeCYiXyCxS
7dweCmu52CgTM4qHIpaxfkKkpovRbN9x3Ah7TygenP7Q75bgIGSQwpF1z9IStNAgDvW3mfraNeGS
F4wW/sm1JS6Mr3vygL2kRtW4tJdv1VrGVMTXUNN5vQfX6b71qM5QlWQd8KscznfD7MCLAW7YG1pA
iz0PKf26WkH52uhGfaAWvthckdR6VFPxaQ0oXYdeLodFD+wrMoXKaK5Nz8wC4bF7BUOpymDksXm+
VmufYKyus1tIMmvE4zhKKSAem7OIf15CDThp/8BTMzzvcxShrvq+OyV0MZV0TY2m3O8u0qUkjBMk
NFawdQr/GeEZScUi/nIVPw7efajV8QRtgAVBYQB3OodiQFDGk0e6qs0YK+QeVtOPTU3AGG0BAlv9
buJYv7+Wu4T/Nx6D47voEWZpFvfJxWsSd+TKBOSIsivXSKllKLbwCjSxjqWkG3MLsshFeDcx2wnb
yQxMFmqj80em7bbp5LQBi3scbLX7PnJBbJXizKmwZEY3RBigka7HMe54oE/rj9nTGDf8ZKrLI1oB
cAjMKYNFTsYhIsHz9p+G8e8gZ99f4MsaeMa2AWX0aq+uhJH2evOBpszAhzXqD+iK4N/K/iz483rg
31UiPTQDtHZfurweR2ib9QcbFwrbSYPRB4+lULfatbJQxgjUITWRBK86Of6bL5Zp9miYmr1BT3oI
OGonfHuiZmSkjgXQ44dxjgRtEmzCWQoKV9Uz3+ZY8G99KgTRu1v8pXv0uOZXkXAAU2JlCrZQvTwo
U97Askm2xdEM8OZsm1uO2KSsKX18pivFQxBhAZaZ4Ku1mfTmP7Koxf8BHpgvywuopHGnfOWE23wy
oFG6CuRDx+KJb+eF3LvKkhsYOV7nqQDKToOt3COQL6P9AvrceI50ZbzaDr/uDmdraxDF2wbsGyMV
D3ARDkNMwKy80/iVqld2boz0ZuHfKIvOkKFoftMs0sH7C+/1wYXMBascZ+3LZdVvmL7EEPbAnlqr
niQ+TH+ewO1ncsLvomDCzjUiPOpabJjW8xhsHp5jYIUeTM38gNL9ZSUOBk0LoLaWHuC4tnUBC9EQ
JCXV+Hm888Ld2o07/01ZncvmmerYJhacEAUzv/lC9BZUTbCCzV+LwXLpZ/g0ridV3qvniGUqaBEM
kfR7GcFiMiDnncpqJKriQg19RJshFf9G/Arzy1FAqb95PFmhRZMwD+PEPiVH3do9iuazC8Vh5Dtt
lm9RnJ9I9m5rdBJATF4nAe/keNfxdfCc+15auU2wFIWGovztXgt/10+OC3M91XVATAN5VIzG2X1N
e3IIyxf+3cRDjnTII33qgT0d2/ZaAqM/TVWzgGASva51cbDpPjZUqPjy8Cr3X+H/p7/8q9YDH3dA
1prL/zBna0KtRCRW1yJa/O9uYmBXWpVxO5DfpTlJtVrco/x0j6iGqQLvXHWNFA2DrILR7NErgOq+
Sv/UI/+a33Rg5JWesIM5SQrmkmAJs9OUQ2QbhLtjSnqBukmJUwP9ymymkrRuRhcg7iUP3r42H6dx
/ym4EUrg/Xe6QkVDFBWTCMmlHKcxDx2zEDjpwvQKpXaXSenBGayJP3CGHFmkKdcFoMvQnccEcEAv
/kC0oR8PGDPlJVe+No1SBzVkSlqNeOG10AsHfmq0aHGxX6fC8LWLklRJIxOPsJCQjjk0kGPgeBoL
/Aav84fFrvdpFMiOw2/xvKJsUiJRUVWrTJdGdm6dlOyM9BGtTocTWem6qCyjlTRv7GXC9xL4GhND
kw/aE7vvxpeNKGIm1xrSTOpRJOXB7dba1jEQuWXSBPeHXYqKu7tH+qDZPUUp0QJha4wOIzb7V5dD
YEvJc9vv16WvNmQSggZeAnAR92Jx92xjrrw+4q2aiVnKxhJzOnCNgpTMIpvmfYv/K1kOEolpmRXc
kUViy0vg51wNyLJqZE29E01YoOtq7J/NPR+vV9QbpkXRnvMzXB95d0P7ZQB6kdtPAPfb62jSlecj
GWE2SfXHTHcaN4MaiKN8fpkik5Ourf5EZl0T1ReeOra021TsP0dZcNm9mSa0x1g7ds/Fc5T5B+4H
elbC9ChvVSKZmr2j8qBqjcGQqh/cxDlhUQGzn8BJVnfAy4ZBsU10nWHARzibM/VTa6yasln+Z5rJ
M/d28lAloHmd9uSHlFbC5y84QCByqMHo8/O+4mZacCdGuTvpyIJgosF4oyqNYQzJLCa4gJRCJyBK
x4D6rtjQlLE/vSQuqVRzX8CjzYnfKup5Uoktbj5I+iTnETxt/9+GqQYcUPLXE2pEIzIkwB0XZppj
kQKOR4poTEofTwaD+irfjQxPZVDLYVnReZBlTBOwrx8NpbGisjs1FLtMRIfpOhMzbNMeik+Mvso+
GCADElJ+Hh1vvWDmu4H3J/SPq+i6RCW6fAD+oWrhga7rT+4BsfSO04eM4YD3+lR1GHfWUmoD3h3R
Fl1OL8UP0HC3CgukCt6zcySXpZOhBm5WDopKAkQ5BE0+xDQuxgb19cWLkBDIUhda22PAACOR9ixe
pBi1bJWXAJbWPv4c3sifYHXkqmbisuE7Q6wLt1X1XjWztIMfU4hT8xkaaJUtVRZ7zRZVDVwIfeq2
yCqab2UgBzfUJdPa/j+HGrhGk7tlobwfC9RV1kEJcFfN93Qqw125qGNQ/yyk+LCF+cCoTh87PLMd
SR6rJyBdCg6TlO1qbvUa/frMgl6k43tNUUVRAFPGne4nKGmLan6M9SZMIZ6IHR5Nks8YIYVGiubd
QbwSFbT/AMEyErIuyTvxoYckinZ/vda9qKvnlngaSGvxvXuJ8IYmfdWcCzsIb1TbJr8mb4llL7Xe
OFSb/fORBn4zsUWC+MYimHRmt1l61IAdv2mK2TR75p/Ksdds01/CCCRSQ2XXTYjlD4GB4zCg53ag
ZXoOYBacvzn5gv4DzBWEsLNf412/16lMhuHBhsqGnE3+Vrw9ycUSYVyAY+b9Tz2Dvo+GkzDFUF0u
bGtg5+cxvh4b3aDclz3DJF8n5KcYInh7ThPphXArJNL8/YlVcNOkHxYNCQnunk/8faiFSZEyXp9D
HnMOHCMKagBYDDzKJgiiYkA+povNzYR8LOX347O4K1SqMX5P1hsbcQ+EqyMfm5KkYL17OR3yAq6E
cwtVkaKGd0VZijykpme1QVEe01EPKqNVHz7B/k7ka7J4gUU/C/Bki+q57oK6gysjsmGoEnl56YWv
UN5wyYEeE66Ylq8lquLMimBxW33oAd59uADMI8gqaeZv5blO4xXbAAOyNFQ50861HgpZurFPMeb2
ZAIOsElWEBWJmhXcKi2oZlAC1dwdkxWPLdcs0jQ+LX1WyBVejIgCC2T95veOkEmBkqc3o9l4zNOX
dNhl5kK5CKXv+gPyzgpmgNXrKtjIwp/eL0oZkzs1AoXtfxZNdQMwcWKgdWhdWhDdsXKmx0UzL4Os
j7NuCbPg+qulF73US4yMNGl+InFqVI2kJYl4KodGu32ybh+TzwZUjwli7paynu6/5/wZyBxRy82T
sfGvUHzlhw5eZGTph7P+uE2New+BrP/RSelu/a3fJFgHZW5B3aBDIBQrUGx38T/qkmk0TmYgEl3b
Nfvu9RSyeImrrpt5tp8LorxEwygifYRhi4QOtHbLthzhD34OG8fl/FIC8UrrY3/fLUj13Ir9A9jD
TxQawr1s6EOggCkPk19QAwjmZusl6nrQB+KsnWZvGPuVFyg4FUcQOcbKjhhscqP5SpdPIQKzn1jX
/RQOjxul19/DnymNvk6N/pyLkJTX/lOWiD/vHzAqTRq9/VR09zAfawL1jnR1SpS5p/KvVdHmjrfJ
YvYWSA1IjJLS8jABSa7cZCV525l9c2VrvPPTqT20MHcq6GnFfLTYI/L8j98QzSQD0kL82bTzcIQq
+MpTHpFbztpY+DJgDlV40YYzCVJbtod/qs9yzT2J2lve5OzyB4Oh1H6R+jhm8VJ9+aaFN5BeGpms
qLcex8gLmnEzvyvqYklcX2XlAwGmV2uGmUm9Pd9kQYlEuJKEZYY1DHtyXiKzZV1TLJV4ibtS8wl+
0G5Iy+igm1IZ3mkY9Y1F+Ct/7OwiKu7rg+zELyiGBU7IC4XJ8931k3ztOdjmwe9JVxZTREiVXH60
1pZQ7fW4pHvxBzoPfz9UwhHQv3TbE38in4i5JfGXvHovFOzbOxJmh6sFrlUBirAhRsReyeTKfr0d
Z0XM3jqXcGw1cJrNaGnCeuANyCImKGLm8vTMUr4Jr8KrFsIpASx7R0DTdI+ukz2t6T+MSSjSzpY2
Mk6gdn5gG2+RNW8r1uQ2tpcPIsBgdmn2LP53MpC+DoFC3oOcgcer5kcv/bGry3OHKCbb9PndbGQn
N96LJXAx6lgwBixA9U140J/ek/EYEqZhZHA+5xwfDNps2opRN5kRRetsYnhDyj/rR8UyUV5pvpNn
YY1S96AZRy/p9viVcH54X542UoCkkQcPRlWAVEUPsASC+9zilHF9kqGDldEeb0Czdpohy99UBHyH
vjtBuE+pgid6m8YAqvOdvZUkVZnJFvjJEyGuTOdZKC8p6g2YVu3vXVmDVSuJDHtfCpT8ROh463WE
m8lRL0ZiRMWdqYUbkucrd/V3fjmjUasKzzd05xmb90huDayqVqnuZqM7HbhEJ2ddDiGe8dkvE5GB
NVQXGr3qktvg6ycTU5GTxusqii2EQmtwo6GIdZPSJk1LFkAAIFrgsRv2YUyh6x2YCqeB+de+tw1N
Frg7/FhehXbFa9mZljHvgsEHpbIZZjYJsVl3qHhWzjIy36+ItuPCg8wucXc2Av2InljpSch6Dehb
MyICBOJGHQmb5fpaBxtIzYxYuVK+/mklGMBSlbzxCubM58Du54e2StlpAjpeoPHJ0Q4DXYh2d/9a
pscvLbqs5z6W7O9EHC9xM7C5L+pOcDCHVjov6vV5/aUP5+c5WMV6VDEsWFNtZqmJYYkwQdmhjVyH
v0Jq9oo69gsJoirunNnYCt4ky9v3XMTbZJDmuHiHASBEa09/tWjPoSKBFjwlWE/1j8EJk3hPVAq0
qKbL9FlGwEaJ3DcPPAal2Ds9/GKpGg0Sk/oY+oIFCfvUCktYnD6I7Dkx4UdZ6QNf5+GCYuJVrv7P
LNWTrtLrlTIltWVeIJI2qb1n6/HfPkawMY6UVni30ktvBJQfgKy8/OIlKna55cirXcOz6Nh8UpuL
QifEohAta8/L/1Tm99kpNPqFSBSRYtHwB5Ru8sagd5wwYvYjj/XEk00ilyFyneTMHuDVpj1Wuoli
3yLp2osSkweqEmNaW7LKZYUzC5sSRsHII3CzNvx0P40eKnKyN7tnVmdj9XrBjuCJeb829G0z+K7X
Bkg6abjAOzYbYR0hPr7D7kY2+Z/6ZKeS/4Bg0EFEIoeRv5Vn+oUDSMsVeMgqaQvf/ht5NKM/va9Y
hTZ1gmBP8WU+AIKZmXhhY6eJXGODWOp544/aNCSlz7txNXXtoaYgbK+lDJJ1+h2U0NDPuDXyWEz9
dJBTwcZy10oonysZ6+eZ5f4GZvEW+sAqFXX0QS3w4fJ2Wz6wUXjWMUqL7X4YbdDpvTJJSlS5Ci0t
8PvqCVGMyyCmUErOpguk2xfpD2TZgpaj7gT14g6LFN1FI9AsbMkNbiaduYVWKHo1tCLFvnlTc5dU
YtFrew0ma8LZiVkLt/DzK39BDlQFSx8PhngzkQ/rSICil9Ts3FPDE/UGyfDqURUGhEsFJRCFgQlr
/ChIa/fIYzEdDzcakP0QRbrCOgqDI3mHGEIewoEyZw4muqxa8HLb7VPq+RSBndrsipz8k8tESgDq
WIxxPGquJ6nBZD3QOL1hjW4F7RvamMQpu3rwxn4N/nd0dFsuTEKsZIba4mX8l/um1FuvGp8L1Aje
EpP+3Hhhk3SbuS6/LHhbcGU5oT29ER1L9GbQUMFD2mBiWdRlclGh1ZdfOGLVWo+8ZuYBiMylsd66
GfctdXU2Uj+bGq7VKIYhjqijta+y/vG+Ejlr2bsBVi8M2DuWkWQjJnJ1L9SNXJnbzg7B5g/8kvDD
mknof7digMWhAwOmU30sYnBA1pmzMz6oNUzhSzFGskghVG9k0A4jvRcsAolBdaCV6kmVB4cojxKX
BFI8eCgNgD7+G+xDLSVvJOKi4xDavrJBQGamm4Hiru2S4JvRC6kYQL8IovnRcmzm0bE+nsNsl7/3
kNj36HAS7noDSOfP+jLpYsx/hWWVwHQTjssHPp/CH310O7AFPvwFmStvLRXjFiueflOtVmgh1vRX
4OKrvAxwDlyFr7b4XGVFUBaSXoD+MPXFow/wbcXJa2Kwa4nl61TcX03Np0pnka3qrou8KaO43C+K
NTmQ1SeJjMVEY0XPR0mF4n9Ym9LoA/dH2Zq6OtL/kOTY9YpO7hTq/kR90bKI7SzQMLe3BKIWt+0m
Oxv0wTJgn2kgBieKvQMi5/b9TXR/7EFG1nvFykRgV3EHZPQyfkOmsWPLeUqqyBEEVxY95F6DwRDr
/1M1YMj9ZzN0mHgX+PGRbBvQ/1I+n+4ZLKXZXq75SeUspZNK6rfaoDAHhAYJ4bpr015h9VL5pVB9
H2+aX1qdpS/TaB1UtaXAEGO0eWWGXSgJqAoTct2QtP3fqYU4x7JV+d0WYa8FSZv9T/YqyRmyk40L
EkiPTCsx4o5bT1xFsDHY6Kyg0aV7Ea9egNDyUMBZbHhbeijYQaxGFR/qFuQRqZzVk0G+Y4Bcbq2x
Jud7Q+uDR3EqnfdxIOZes5JxiVP0pdP+LEWCSFMFpCpgTqJDri7oX1TvhH1H8ZPofMtRdxnQ5Mvo
KO8hxN/n58SbLtJ9F8rt19o8mZyOXxMGX2At+343oBpiBPDJSwfT95/69h24oMkP6sRbAY3MwgCD
NW3xTCVkXGTDRqHNEH/e1JmjM/Ub/PUfk9KTkk/9iF0VxS5smfRfRoAMntojQcshXsqdKck0bXXa
8VmwLFdLpSySnsmONrtMLh5xtzlAuREuV6/xODpAu4j6HUsN22KGCFWnlhhgEB1WlxxRdWqNvMFI
7vQz6AGv+WkFHq1sLZkHAT5OauBtc8B16yTLlxzG7k7Ge9TI6z0VdjvuZZQ6GmZRMnp7gBb3VFPk
d7D0cXohlWRVU6DrIoAopQT5U3KGF7z1UAN0zRGwVzyi/e2N7/1LBa7zN6X4AHMF8w2nlm5Uaim5
fRV6Ph5IZXE0ad/jMrXyqq3OS2OJzMS9jXCFspK6333u0GDCYeLrvOn7I2wxhvo7hqZv1LoRv9Bz
pEU7DHFAYP0ozgbvn8TDCrhZmAEpo6eOEmpTyVQR7H9GJhNgx46FK9gUPGS+XtI5KFLkeOChrq4I
9wvz0p6SGO1ArFHSE4HUGIXny21PXbcIfpWgzq81k/BzvKPTkhLLorqQpUUkczyrPO905037800w
F7Qy++wCvas3rVvu6ibYLkmQ/09gKh2NOCyvABHZuyfsa57dGox8odaD6RlvtPK8aR6oViUh6Kyf
9Jrq+Ljf5Tp/g7rs6rrwMOfAon7q3y0h26jBH/D0FmPU1RSC9RwDFx3D3FvwhOF+Cwb4HgjskIrZ
dxM7PQY7+pdr2FdnF/dL1f+YmY2fHYYjDvmNa8WkoeR6oSNpsP1q8x3g2CI1hEhJ7GvRQcIftFm4
Yo4Ga756SGN58hacUIozqR+J5E2wVRjDDzVjLfSJ/xrz0pAMV7kETDA1L5Pmals1k0SEraeYDpNb
jnDTAgJd1IHV0s5xNG1Y47c/QIoYgXmetI9Krwzloj30yDXr3QLgU1mFvlS3mplbNadLVMKk7sWb
t9NeUDN5kuHbfK9iE77IqrECJ4oDi1P56ZJRhzKhB03D85qwZZIupfyNXOFBPGqL8dzPYX/FfpOe
T1jqd/GgLcxHckGygUSXMLHqUQGVgzAGcIbESs+4PMQT3MYE0JInbCxwHhmF0K9NMifhFjJg4wzz
oSnH9E83l5XygugVJ7VCxMP/TBXqsrf3hE8uGK4hIVPo9BhLwxBD0YIbCT3x3D7l3XlqCqBbYh3R
D2TxKZq7UDqvCjDamKe09hwYk7AgB1F1Uxv7faS/M/ZC9aFgFj+bwf7v9l2/JuZh1k3YWpqFtzSM
fDBTfG0ZqRvUZjvIVHfXo087dNpgfOHrl6YBDokiv538fBJpk1TIqEjpZtnMUwMcY4CwBHXLUmQ4
Ed+tvSTb1ZNivV6Ffgv3NM82q9q+ttOb+T2neetlaMfLpX/0YMuWJOAWVp2luvt8fLePngUC4XUX
z8JBHRAEthTt2HI2VWduWuxK6lYkvHcI2MHlp9DJN8DWqn7rA2yEhGB6IIKSjg3Lf8Co9rNs4L3M
6issSnLNWAHNhA7ryApHPT2JS9BTS3o0n20KOFMCogIZSxQWO4CvVygyrYY4cBHbscx+mb92Bt+J
+yVStkZWc2RCPahoc16uFYC4abCSSTIox3+5XHYWkB4F8t5ZTDoSM0v8UHV75mdPNbCL6ljoD6Ej
cdSyyTs8RNW7prEzW79kZOVdG4AU0CexY/HkJzmHxwcmFmly1PWaHRHrP+YEH+SshQlkI1kYPi30
/VgZfck9HA/DFh4xWCJBVsTYDo5S3S+1yjPoNvl2zO6ZsBQeFlLWFT0YnkxbWiI5py4x+mi7MSVL
ARflnj3KJXjd/8XWBq51HBDjy6a32TfH9LneBNBvRQJkA2pY5FRI13DKQEW60YmKcILUoGfKE5UD
aw2s1g9tc6CEgmFDJPK9HsrQV3t/O3UsXXBA1UrqxQyVtXLmYEPC1rX9V9IT8V6VQENE7EGF9Jir
Y+TuMjyvhUK5TB3Pxl8cNLg44InU+LJMGflvj18qvBKCTgW4EJrBZGZ6pvOG3acBS8OQkCI2Tg0v
/wWjooCvJxNmI69/SbWRJrqrmB+gETsPXY+Tw0NOPSM6chnQ5Rf4HMkQiqvWMV8DeUzR3a3wCZjW
//ZWSEGpzWCaF+8tfa9h+GgCykhi/fa662ERCNqd0G7Nfps+hbkyi8/ILNH7c3OTbQ1mK+cZSpax
3Ou6q8/m9yN46tQLhzYr+OepIRFeBu4/PA3F7xDrN7sx9h5l+B2sd0MD86S5Mc1sCjcrH7ne2hdX
Qx5czViCK10qeAiq2kRrG3OBJOO5tLE9DLr8NHGaFya2dpGKLHf807aJkZrvZ330nWEmSb342dWv
ymE6+sF3ZV7+3gHino1P44W5gi1XnerYqb+N13lyHiQpvHu8lIGZFTK9TrnVnf9oak2zsIbzs6qJ
dBH3b10kE0iK9rGomlnYDLL2cS5x6RJkz5dMJ4+QJl8nA1XPrj2cFKNEN4OQI9gvXwymkAHy/CIg
TqvkFkMV700YXcgV5tYywTS60XNzTokIB7b0Ota6eR37Rl6ijh4HU5VSPdN+SgRz3PsTmtsne1ov
iRwzDXtamhJm0BV3WzJ3SAdWjlaIKHwltkk0+MRs4bdtHIM9vW9/wGkONdBVFef982dCOLhbZ38t
PKG1v9kOQStA1eYPrNa8a5OD8X6peop+FpcCeDL2VdeOko0yiECY74oceioyREwCmGc7c29D5Pd1
TspjPqwMJeV05nJviwLe6LiA7y3br6mxpFTsofTLkKaeDtgNLTXoeTWhUjjPjM4DbjKiymELUzI2
vdLlsEOvEJ7sywqgmMALqjVhW8opmHIK+6GnePlWPehMGL3a8Km0Kj5j016a3R2xiuS1XtBQAtL0
rtLfboNPlZxCIeH1Q/458loZxua0g5mdTtlW1aZaURUb/RRBEJlP8yXS4cjzpu28im905u0EGwAk
fPGEtgpMLNDTZqzzfUSN0a7s6oSHMW69UGe7wcNLl7oBRZw+SEc97xDOs5Jbcmu5Ehtu1iOj91LT
XX22G74WgSkbflOrKGcoEw4nLR1+nvxu12DeLH78ceCkFrZouDtH4OCN0wI3BKgcLT1hgF39KNvz
gkp5wNISzFBheF0MdFzlcLCgLKB+BHuZOPxJvooTA8fx/drYMBKImCW3CxuvYuGBRUBifRIxR30i
HGiK2j972s3f8uGE86JKIsKWkdNZzszDBKfL45VWbJ2qfB5x4r9kCn/wibx1j2uAhCncSNRU3OLA
sd6cFiQuPMnDZMtDxk8yJR4sMVE/3bff2PTJ/PR9pA7eg+H9scLkjsI08Za0py8cRKiYo4fElkEQ
r94atSCGNSU+WcTcoln7Mc6gM5NKTWZIt0rIDu1lWQDofsMsnYIZ5dA2Dbtv+Q/J3b/EgHaLRwvr
ZqzZJSrK6NhDChmj+QJg2lGGEYhKB/TzbgFLWcvr5M0LmxBM9S50oxAWlVsK1J9cfDD2MCjIK/eH
SQcmggxgAgJSrd5etpAuHJhiU0k7BfxijpFyjNw75EiRt1MTNxkgpZReU4fOJTpPAnEpwhAWOPJr
AxNKgylsphhq2aW/rpIRRw7AD2qEm7uiC4PksjmprV37+Lwej5N/V8N5egFlxxt7hK+YHZSuAgm4
KeY7gwa1RjnBDUVPT1dkgh8U1H8fQeiLM8sYhdQ1Zwmc3jnv1TebJkY5wJQwnvIDyTPJR0gg6lc2
RKGs5Nu4XDqqyi3tkz7vUsRwtjW8zbeKtZQGBTWkglRhyxvCpqPCrrT/7p4nlntVJp2Z3VDgaydL
pYf7ZMMJEmb//dzhIgCiqfOFqp+I4dyz6jn5wtmw5dl/LqMF4QHWhYP6HBsPLmgrIdt4+3DAUAq3
yhnr+kppCDy4fPH1z8QZ5vFab+UDEJzQp6e84wtUZopPN0EYeVRUjmgyzUfsKsM2aX3BLnifX2Hs
2aLIxJFw/y6Nb6iWGWOeiPfibGrJKT85r9AECMhxa8Dwb74qKikgMnAmMNGLYEaYauUnk0hTzmca
usiZ2c6UEvbXClZgPCMdyGMH9zHg09muvaoakXtTLSdDhnNkBxpXd+p9lCbbDLDbObkFJYyJ785/
we0Gulu7kmTiacoU5JsTkYN6hLfQ1c4cz3KYqeShChTzb9pgeY5zoeyDDwgsNReGwpRqIyvPpp5T
jybIvB4tMVZ+xh43rSv54CjjBwbNu/Kg95I7F8uHbrbEfFgYfSRL6vRkECSKL6ExsiemUjhAalan
NTTa+lBINOwAnrWGg+OliVkapqVTpkcH39TpRtbPn45bEQ3GTjj7SeOmw+zbA5xtDrPx8MRocNIS
CJool2BFESVik7xNJ6B/1JUDS91oeHBqF1S7hm+2yCZXtpu6u2eFZAaGkVSjKOPZvZ1G+9u9JDTC
s/amM8zHq97sDz8UICLVEDC0wy+HfVrQ2I11+49LRBKOPy4W5WfkCIUY5lsl5p1g+b6czRBEoY4p
1RL3gGtp1bb72B6qLDXObpOtT3O6FM5IRimSisAoTDTsz+0La8nTLrsr5P6qy3yShf7nIkNPFEuP
SFnGFkEapYhKVWTega6K1rt2959WHUT6MgDSRM/LO0W0fG5q6Yt0BLElhTihN6KeTd0Mc8MvsmPB
7SwmVETo8BqzTHjHR48wIynXjJQXZrgy9fuE5YWAzMv1xOB3ZnFOeW+yu2FZhyt1tKslF00zRSVG
937zEd06sqPq1+pDhBuH+c+5Nw1Zku1+oi6ieZjkl+wnuX3Hr33btzfesRfDSjIl/bmw2L+6xufJ
kk0iMGs4xCXRwvJW6yr0ogC/xk1xJ6OIdDwqHpw4lYPlP1ynuYhBWVrWKibr5W56O1adQ1aEbMPe
qMYwYjcs7ciC/I/6kgkSbYIS4A1j/MmqpQcyY90h8prmipyEfHPXh3XrYoxEPh0BkrTX6gfjB+jD
34oF8SQ71rDSG+iaMdFNAlKAeO+I6D7gWdJIUFo6AYrzzmf3yk5Roo672fMwfI66eXd4pjetAjPf
KqFZm2XAJmQIb8WtlOUif9BS+iZW1Ax/d9b1irazM2iUBYeKo8hmnYyYGAP4ZJaDpjsMtD1FkzzJ
nHdVcpK2HYdRUqFM0/aNA9Ys+mnUr0iBd3x1nCwREoFU81vydXSNOYomP8TSEEXSnJfYKgqXT/aw
HdfXT/f6vpIYw7OG4b/JaZj/6U31KOIpDkgikFm3qewlJBbg27EgmNsuzGP6M4eraatfu1xiKydE
8umY26JX32Hd7AqQfkx9saujBG/+YEPdltHGyD8ECn1im/X5xSPWYymo3/2JcAE+hpq3br+RGX8s
ltZMgiDb8fwOpUGwPvV4uXSjOBPi5Z8cCCuxWbBrmwpVLpry74S5o2xEJZd7VZnj8jLXvOF3Q0BZ
b7okjVaa9zF1zbTuwUpQPiVa74cU/UfUOn0bLPo3GsFkO7hrkBE0B6SCheAhSLE3HkTfkOKYhgSA
P4Ov8n1cd3wyKTu1PNhCiG+4glsh2fcHphXIk6t7pTeaaEbauGytlC4OgepfeX3QYnTY6rA0YYH5
9lE2604wvKewUfKe/BLoZZNaWNGCPqhJg70E0/QosBPv9hvYwtGY8td+lQ/U6S3jmICv0cyQZP9V
MsYysdyzsqS936Cg2RyzKoZN/QDIkw7bdJx+3mNCb/YW2aD4x/IN/bOFacp7ncY++jxErO8Fkt82
aNizdceKUCG3dJYdApYm0XVLrwtxYzpo876WspOPXYWKRdOnfPdwwnFCLwH2wndp8A1kDzglCc7L
XqftEKvZ/kAhWLAD76KHy1yssxGzwGDaeFTX/8havT2UichX4HLniVgo0LWZD/LWz+tpghAcMUsX
gtb1D5nyFVNjQjIT+uB2lbM46eXeORdTqY+OpGbpD857LTv0Ac+j0/Cy3Gf06Iu0Bv0/9eRd2cxC
Uy4UGx2jAoQUINcf/t+J9MsyoavdqWKkWTq5GbOGUh7bSlPZnSaHl7s/XtX8I+eE4RInwep5K8AN
+dIzXEEQHqJdzygA5HjSDjNzWTf/Zh1skyfNqbjiJ6KPVYGFenpz4K7/Lu2QKxPggTYqo8Ljlz86
0mTM2ndX/mMwnwTyyUEW9jEZD8wb/YN/38rfec+KY2Bf7bY6mz63tzXAvdtZukNf+wyaNPDSyPLl
DbBTx4boM9n8CDrijpG3vBrsML73joaDLBlUGpn6TLJJ2ECV6XNNqLa5DXqgzoMAsniP+fGfobnw
3bdTNEJFnyYHmxy0lMIRnfWt/ucDe3dGY68bJDpe2XOncvWWxYWMbKV3x2MTd4qAzUEEUryJ1B+3
+SuCGfQd+Pxy6ECZsUyjflZIZ1FFs1+YJw/llq13l/CW0VQTQxnXJPGRGLGRLCDZoluvWT7sltTd
NYaiMJfZmmsXODhcOhPEX1fBSy+47pT1mFX5luGpySfGEc/FKmB6U8is+MgfqwtkHgmxjt6NP2hH
ff9rdx9c3XKkXK/hC8ZxzaIeHJijnbS+ntGsF7zHHGQfWg7Ta5eztD4EKZ6eVXaNS2tIBWex0Ldm
DHntJ76fzh0pe2ixNIkc6G9g2b7J3vX0xoPx1uXanSSi0PJAZEVe5xOFtCj+94vryvenP3kWrmbD
vS3LGHBZI419XPtfyRCl51Vm/REjBgSnj/06iM91JxCFS9EM0P8DFJQJDAJlZ9m2DXV5c3xKRtj6
W0CtzvOlbZHr5+BxlGirwCus9ppnyavIDWfAisaWJTO2Qq94o2LFgsn65mUVSob7ARV48iLAcGhf
s2Fj7h0ol2+3kJFrUvYc7lK//9dVwXAvu2tdken0sVH1JVouOs7pGinaO0WBDRCpKjPhdMCbvm6F
tmBwpXzum1fYXXEn6bx8noMhQeYsoyA0zWZu4dchSSB5dQftQu1EF5vG4EiyDlmbGtEMBOesSWkQ
calzyxOhvGxyxknMLQmoBcaFlPg+CZhVja9Scxy23kE4VCOoC8wTqPEJiecAWQ5obl6PEL2dfmmb
aDObgZQnjxLdcm8u15XHA+uw96vwWP7MVG4rfEhg5t9xOzr8ADeg/jg3xmTU52wsq5yDwUd6mZQR
JReVe9EwyDIsr1zVXcaZ/CIQOpAJaQS2In5FyGJlOHvoYqNINMl245oWvGDYkdJQKiRodYc3qbXh
ySMuCvsJpFdFH0O9qzH85SHkB4CfbLFYMXblmjcVTvauuHw8JavvMhn9357uLVwR7KnkhbgvGeRa
/oJ0qQ+le22XZaPJRYTNBFKtZC/NbKf2RyMZPfhjY2sdQs1tfNo4v9A5cmIIl3WLiZ72Hf4Y4g+N
T5KMp6lXulVArlLCZDCX1g7VX4qcRLRgCwYa68I9LNV5KDQ2FgyeKQYIEDVzjIEiIZjgkumhI7qQ
vjQjO2Q9ggn0r0/gKcsf1aUmFC2H3pgCI/lSl7dhyu4yivIxAHa3y4eIpn/E3HtrsTVwdKGZS6df
pg/U8PKjP8qjJTL+/ldy35B5mULRWUSFKU/jsM/iLi8IvcSbZkJ010/1KqO61hbSyUGPN3d8MO5P
XX1CyUeBxypwkRoX8M4v/3SJ+5Z0UDzUraK33RooADCX2jY83Anpie5HVUnT3G7egCiPX9uOZDa0
9SZ6PGG8n9PwiRIQwUQS5G1tmmOU5s3nxghGi1oiqWOgMp/sOwW6bJnZ/HDKrGdwkBYXbDHagJkH
S+d8wFrGJfiJhsflrMd+NiFWVedO0aTG1cnPaQM3+UUT28WLFiTC3mecMY2Wyk9ZPfvpI4pPkdNP
mWep/j1+40UJfEjZ0EVlPyzN03xyfvAS/FGV+7Gv+uz/1aO8sPAFsLvbqDbkwDDPu1CFxAZSmpR/
kjHiJLVDuf9Vcae8jMsnxAApJEy0mb9uPdURnwVjpd33t1K2UH2ZbUXjl+iQfS3vOWbIOyfzTq9F
ZPDdH//4FaEdQ6spb/0UW2SPk2/c8kLCObsDz4zHWYihmMeDzhNbNlFoLb4KPWIR3ZmGrXh5eD57
kyrzJK5w0Dou9FsfcUKg4qA1fUsKlQjm6b0+sUzMnkqrP6bIDEPasN41e6CyATKpmWEKz7oxeUG5
lLyHvU/+N206ys2Fy34ZbJukOE0AZ+LWRM7GlrktlVbudkDtQe5KEuEyh0EGTBsMI4pVvyd+L8xc
5adFX+ao8iorZxbXk135S9iT/dHs2eRMujX0043JXV6ZQHHMDv8nHwana1voVJtYue2NLNWr8BfC
O8pSWY/eAUYP6siovKIVZAKFw6F46jSvuBlimJeMXMFSgKxXmRF0Q492Mr13HNUDQt1rEeOXUyNC
sSC27H/SA1Wzye+HUbgMX3Ryt0AMuwjLFUsh+O+x+IyCsAwUHTvBXOpzkFshTIrv1bfk3bgOI6Q0
+efiWhWbKrkeQ5YKJKsU2AYIM5YWZ15Z7yJBZRNjYnS88Ak9Fmlz8jkajL/bXSbskRVgwM/yqa/g
Ldp714yoAPjKQVO8EaC1ZwZcQAe4vv5d3pzziwCVF6JbMNGKymPVFlaEdO+R7OAZdZD3dIhJh40r
+EaOt7ddyd1iehifL9xQ/hAkQoiZPhD8ckebHMkwa9YJT6bsLNFMkuNYHZqc6yZLBzOAJtrPjPWj
sWx/CdZmPxhCLdB8Cwa3y8bNsu6vKC/c0Icgw0uCXANeQwcyCMRMquSBHLP+glpKrq0Pn1oQUoG4
awJwUfujGchgkulv0Twax5oiRjDSjbfOIp8D001X2ARJDBleJfwqepQjmkCbNwyZ1u6GQky55SYC
yIX2tok6cbEoeuUkimfbQgutrahDIXn0sBkHUJfY1PUiu8Yzw9bki+9iSzYHTy6eUjdwqfMiUvYR
VQAit+qgttuSurTvDJpvTXYSPJmVpZ3H3d6PxizzOLsAmzgAdyBJRDbspjNuW5rDe/MQNGOUrcap
bw4hq9LdAKSJiPwpIQStDltIbfEIQE03Ti4E4d7U/WWuMrs23JVgrWbMo2JsRiIb36D8hDL31Eek
Vcua8D3oILZnrqYFWc1KLl8yalJBlYjrWyxEQtwrvFB0ZJ93VST0Mi2UcSrpBatIHbQtD4TVIPKg
8GqP7hkLjM6o3pyczWDpuExWC8B2byN5Wz8uMrSLm+bg9/Z5ZCTRf6EA9JKxZNkUPM8guCe8Yivk
EueksyKN6+O3uyf3X9m+3ZT8BddSr/hYQgV1haa8tehdK7wSfY0dU4R6yH2d2uoRlTNzAn83FtV/
NqPrfB+nInWQqU8J/6QGgE36Tr9o4PW1H2NtQJ0z15zSo9U5HV2S+rDYqGUS872Z0wJ24pskjDp/
PyOotf615F1rq6+6Ht0BDyGhG1FV2dhKi7DBzYOK+CPeVtITiDNKDAPS/F/EMaq7Kq7wJfcgpT07
Xh7Sk59DEogvpyWQn9IqPTM9c5j2EH8Sz0ury9Fr4joWE+b53yUsGfGHb5G5rwjQDm3NjB4B86Hi
2Me1q1J8TDHpX7P8ML5+s0wc97LIShFFL+DdiLdwxJul+SVfkJKntz1Ip+ToEhoJU92b6LNwlx/K
pshMWZQZRntKHfdgcwuf1wxpjAJOnw2J4cmqd9GCoe94SuAKTccRlhcfXBIU1ALN+vA/C1c0AS+P
+q8Hbs0HvFdt3GqGfk/rCrqWRoQscFX9x/jcP5WE3Egmr4WzVchjda+a6L8CKTamCl6PrHr6OrO0
cTUh7+Sj+4dSKxE3IaG2WLKk9YRtyhXOmKIsqTRW1rHy+tI0nkOkz7/b/RUFrwUBTpNvlzs/pBqu
7K8e1/FlZu91wfWOWY6Quy4jKKkOQDA8pN6WtUQ4Re13dATsLRfSLXhEJlJQvcBHOx6rMZ+SmgzU
m6PgR6qzbKGsXL6e6p1CQTGBLwWM5cVWAtduTJLBOP4PVx6CyMF+BEMEGtpdSqh0U165KVeHVgPv
gDbb5DrjtSY+xV4pUrAaspbSWlRMC9s2q3M354QoQeDR1lvcEEqTMetEGZ46ga6FitMuePRLL3Fj
88b6/p9rQA2qdnc6m1vP0GBoQQ3q75JwH6JsnXoylEkdTzhriysk+H1vobdGOy/z+gnBo6OZIMwI
afdh/7JkIyCPKwLwyX6Dn6kJOcUUo7gLAHKpztd3/rv/euDHz/CyUjGr6eWrsfqJ/vQX8uTS8fTo
wnsb+wNH1/CWQAZ0P2N0h7VF11ydbh478a6bf1qCCvNbLqBWQrmDTtC1Qun9VHdbudBKChW1mUQE
EtrmiYCWgh2Yaq44K1TehkHmaWEDTlVB7EzB96EPbgPfeEpILv6S5PQGB83IsszsVxWsNzJQOJT0
Pz79TQt8YlPMxJ/nFUL8hcPxNDTolvkXxQRSt7ptniqPkDz3/TDzvQnq6Oghx3oR0XJmAL0O8twl
NCSGbPgzAPHgc/3SDH5utGP+GCaVMajWXdquM3fHMpZLSqNc/1Ewqzrv7/YTqfR4qY/R3j422/g7
ZbRP2Oy6LSiNYg8a0DvpZDPE5GKcLqF/YyzGm9Tr2zP+ae8Sd+IOKL/KjppMY/vyVBWikRDMBjiv
tlgCPP1y3h+3aLBmhB7Uo+FAiR6uu8eTMomxqaqdzh2NHRI78qSaIgsA42JfF5nM2YRCUDwYk0zs
Usu+G+3rXdv5h47ftvRs+XsBe/AmVWFVtYHR4iZYX0mZBdS+T1gbZr0G34pDIa0i0PIGs3mH7pip
6WNUMCeM4gNbF+Pxu16moxXAeo/paWX1SlW23PCtOblMsqZuIoxARd7hkclcKUtYltCTyILt5xEb
nPbP7KKq2WW4fgR/10+4IZH7l4SrF8DywAOJY8WuNLkQcbo5yK6qTeGZF20Rg6dlOyooLVvsmgkI
v3wfsyH1HPQTMNiG7xYCgbdx00mNHdAaIg6Gwai+X9nb2IkG1yiHoNEpeA9l5XgW7dqsdq5lM9Nf
ISGqpsX9R09Y9b8/WX1BXCWVWkf7K3mZllFW/rDkWZO8hidiIRl0agdxGaQ1azQM+i+aazx+F8Wn
pTdAUbR50fuMSmb+Ik0jFlzzP5fiqayDv9DBbciCssTL7JhArA1h5miAWbK4w+3dOqadhHGbQK7j
j0KvcWAi85Ca1F/GzzOsp0izJglhX6grWpdGVK07Pibc24QuDHDoi48v/XP7aea10132Dtpcn4Qq
aX5Cjx7PA5AdT2Qdpn6k4zhbtKo1V4f9di2mfxjnTxSUZCX90s7Kjo6uMvQutUN2vY07TA9BybJy
hNnz9wNNBTyheMzq2kX2wEpGTYaeeBQNPLCNlRI1BmgB5oOlMUMu1yn2ooTNk30qE0smEAMggah3
+tuMvauaIzckO4B2EMVPwbmP6gQcFDXEXaKD9Rbjw7ZHMVqlBtA65X2moMoUBAxAKtKAlxodg3Ve
b0uyYiOlPl7WvIGuk9qJ6qDgjaHtObwh6OFOFduCdReZVNHd9rgXJGAuJr0wIiPLmeQKYftFbbVv
FndIEB4itst/nHVJi/H5iCbfb4zQLwhCQ4zl+yOQs/USLOuVo7zYOwAkcQbsf8rSpS0d8ItF2ZK7
XFDG4pIOXnsXrzJaAiF+/wAa7D7Bt8K56jUXUj4DpU7WrnBEXEJ5ltXFK7Jm0TfdsBLXtbZvYYG5
9lU6h00vQWRimSKW2IVgN2Dy16XjrbaHSEdMLpwjEpQuII1Y5ol+hi3Pb7O5vfCSKFgekbHsDPGC
p3j8ZnNd05Jbuzq3t7wRafdQ8Lj9Ek8PbQwEL66ipjUGDD0aWrOx4ICyQJXxcQ0XJgzKBSBVDKc/
YvhXM+NsFD2fRNhPrGY68E2qGa43r0WgPVByc4PSdnR4cLgqVEaR+06hLS/Grf8P7QTSj7CoMIzY
VvRxix0ocW4Ux2nRE2x3NG3zmxV/8AsyspaPm4hYgEw0ZAPti6xskPZ9ATa3HZOwNqncesTLwby1
4UDJjdCWEYj+nn7Qf5hlkGDv6WdnsET3tZV5b24UedWtQzD2yUywtYY3ITFe9+i2v9gvK4kSzHxr
tACwsrOhfpRnr6btVx4ULGRzva+G2kXgIev1bLAezteOBeU3ZNe0OgOC3+6vdoQeT47Zb1+rP1bG
ffRPfSXxHai0WIoCdl7y86UPZHyi16YTGQoEqLkmhP2zJAmgj2DoW2Vtg0QAbjczwKkQFGftTTwq
IqHBRSBTvXy+QJff8vqvIn4E3IAEj0+ShhZJxgWzHrejx2mRGRc3VmRlHTxD3I0IIO7lh68yX4nn
OC95vCG/C+IwOxtO/sAjDKlm47MmOmWs6+ZoV0PiBqdBgdag4k8v9Je/fUGQowkmFitRStUgAMD3
pKUXckEpKRlTRMEB98tvLi+8YfTvY1DNVmM7fP4O7hofnnXPoaQTczMLQrpc8S1ACZuIAa0cHjC0
GLC1E5p2xcuUXGPYcOLln0xnmvM/jQCG8VjSnvFKD7uVoPggaenUjkz28ducPV1TVQSkAJ9nE9do
DEaZkrSHi188VGI1DUVcS914OwM9ee8rm8IEfK8CdjnsuMkWimuULcBUaOTo02obobI0mBn05VaV
IdP70Adop0f+MirwWnrwt/kItzCC4/DVeLBh4hBoexRoiQlPoSbmMLGfWCFCrPIDqgk/stS4IYFV
kgjTnI2gLl7reh7LbKghA4g5ATOQzQWqg/18IEWvYAN4D/YPCEhld01V1fED0qDKQRLiiSVyvmrD
+sBWMNtUpYCcc45/zdt57YQgqlaptXwi1VINKI+w1BIzzhzLBTEpypZFTMIn2xcP3tCWCfV756w/
JyBDFQoRT8maHQsYfLTboDiophWyRboY2CeRIyzcBoSfS59ZbwqmKhUxiZKS2eXVgvqMM+gzcVhS
rIqJMR8l/arMaqzmDShtf52Loz51XlNwrFOWJUlbJTpjubZ9mPtoclo4DdS2HspVHq14FdhUz5yy
Xu9oJRAenqMWmOM/V1nRUrEWqyz6uxz+5/RVpxhoRgNACUUCuL1ssWZkAMMTHSvwxddw079Ti+5w
M1REvECz8Y8bm9Ttj0apHrc0yQj2lckv3xiiIG2Btf8JDroBqHfA+4EMm0jGk/kitvLT8rb3I1+4
kTUstfUTEgkDZtLu8KBu4u1VXE03/KQ73vItP4UxgR4yxmIq2SNRxyrWJtZYwTtQVTXFBm4pj1R2
iCtFQOE2+I0nKY/Ohc/8L1sGTekdOkWBlxEvrZrmVJNEW7IwmFbAELaqQ4LTFIB49PrbezdB9fPy
+67daMyHKVVgfsUejQWSueyk3CJPoYufIU1gEs7McTrG1E//u4h/BaQ2HRI/2RslaNDxD0qSWbyD
emPuos9qPvHzs09vmCs/+NiabQFuMgBdOg/+100eI9UR5I5m1ZnOKpsf+rPW7jJAxOqiaDRebzWL
eD0BDlb8hmyx7K4LmS4bZ35YahMWAUAXq2utPuGTHpNmpPOPQbfx+kXZHGM2c4V+zvS36zKza0ef
Ilajw4ysHL+IGIBxoLri1z4CrXJf8waiwyNTl+LbqDcZ+aUUPySNM8r4o63s4Dzi2AePy4A0qOKk
uFJiAVzbyiXSg+hIjQFvutxe1atDdLEg9fsDa8+6aljEUOpbbzLjcAvBphaqLngIQyoot1zgx3F+
zSMhOVMCG2lApH7oFPai4arVaWXC/QvMyG+kzH3uY9BSYC3DZ5tGugf1GPw29ei/nQvYriA5DF3u
0tlfFAUIV8TGi8owr1hysad+l+bAMTyCNrqTATz5R8jshiQhtDGhGB8W+5B9a3OA5VN6lNEJRHR3
UBdQ77L040HT7pD5Soow80MoaomYusFEMZdgvNJe5kOzZ9LNNm7P26CCHhFf9Ni5EN0rxD2irZE8
uwoyxBXAd5HqrbSdgiLRx2DuCt50EFmOcDW/Fo+pR10S2xfMOFVG/twrDqikWQvxucZKK+xELvQi
nMHbiuHXQa8cwepwQs+5hLDqNibgVesVlSkkioRxmYTP3dap94GlnnO5xD2jO4Ro8hRvOKnwwtbJ
IJfONphMBCryO5unT0Jm5mACfCHJI9Qat235Nxf/0SuJcjK7nJglvJ3X7TrRTVTO8DbNkC3foTJb
bxYvYqlVUPb7c/EGc5pFu0dls5U1G487cgBqz11DerKXKZmTKs7xu7Bmb+Fq3gW69Cv2sWj1QVnw
z3RvXXmYVmagtH0Im+pkdeq8Li7jky7vRUJjqEOUG74AtkOI64FuI4ByshNOqFH2LiEqmkvatcrR
yREFyla4lh2D24WZ9OEJ8lx+Hnl+YwiDp2HY7nvdi43OGhl+PL8CRy+JV4B9Qy6lX7OAf7kvqYw2
qA6S4JwYzBeNi9Spn5jeGq1LGEKVTIhhlQTjMYExWNwwo7ZFhRLas7PiNQrtjlg3MrgKJeJwNmA/
0FwBr0RLIrJ3XcYyom3OnEd8t5K/fpi1J67T4rjVw4fOVnEvZfgRrORkOW7x1G86BxUkXC+Tn3Du
+rUyapCxdiw0SCZLNqzQiDUgtg/E6bvJ7ohmLeRVtUzOACwiH/FCvWsrwvNfKhB68qWhed/AkFad
F+Jgn6GbNrIyR6Ym2mlYZwj+eWOrOqyWUJuIynBHaY5YQOSSVw+E1frEITQ678kLDQgKRhodEghT
R7KxnfYax9K8X040htFx9N3CptYDaGTaYVYRp7jil1ODaYynAbQWC3uhBrwglf95td9668vr6bva
r+h/EasHOPp0TFCNAO/luzn1r24SRhIGa5Oa+10Gpb29ueEfC9YxcMmCCJ8knEBIzjYC3vIJU1al
MAodJ+HGyP8tj9iixMGNlQHoIbeeXyiXyPnvhqzxc1E5O5YEYoEs3/Jw9CJ8tbeFV4MdQk+O9/kP
DdSpihlRhk7b40HdRcXvDkybvfZCAwFiMRFFpmcYQK3gPdphuFSvyerRklFsJPMi81BdXBKzl+KP
qDg36UuKwAKMbAjZLy8JzKxWFkJiJ9J9zUx77R/JGo33trfiN98ySy60+SD2pbycbWzRHKGuK6Px
rNWdJGcMR47LAtUxg0KqFejL88Pa01GbtA/WNUIQqzJ/6rk18CSgoUV9alX1fIHEQCXuYJmWE9gA
eeoFX37u44RTv2viYEDKNv3oj90cL7LEoEZCtv0Fkm99Ggt6E+jY5vJ/0J0xm/bYQrnMq7xK1XSJ
teiiY74U5fRS5WchpuI9NP/+bcRYNYx5bFQxZOsv9FqBC8XuuNt10+3uOcbuj7n26Xbeu4KbXkSU
ngNsDDhaNVBx1bXn6cSgt6ICmBgukaZhI5B/WkWd//vVHxOcTtMsIeGC33L8twQOYchrV3ycbpq+
TBYwRs6MWVivyWn5OB/KFtpUl3VkW6zodKI0tG+FBzyri2HodrqBcNqWVi4xS/8vrWH6s34t4epm
7eACEewGLGKT9peURzvqK1nAI1YYcFYLqvGK4ykKj8YRZKapL2MzAVThXmzVzeLxUIF3RJqbcdAw
6ej/ZrrpVTtctMdPA4cRdWhWDy0QUgpWz84UNxVnJzT4Xr5cEdrj842us6q19gbupA5baxGx2YMu
wyaJpK5o10loslGJ0qnBA6DyhHykQEIgFyCGtCzzLjZZiFAIeAn+K8uBukCO6zwclHDSfzikiKqd
27CUMXf727xAe6kjUwLrpHqjsKLFqR/+qvSm0LJcT8871MzGqqPiXqejy0uWC5eCsZ6jL3pbLFoG
V60oYUoYyOnBF7v2tF/jCkpyClBd32fQ5iUEcKryvAFEuDEs/Fo6liHppiye1YsGKcM/odVHPOdr
VXEClUyQVIEKVS7hGP0eoaaPoXgOhYiukds+y+OZ1kXFGxRokmY9UxxAAJU+h1X5dB9LeD74VIyi
LbVAhc6/gXRc/h04BMLuooXq4qP39Php0JA51utk8E8rCaI5cpINQmEtZ8Do9UPpHBu2aIRZwotI
KRReQWChjuw127DyQieL+UU/X3uEjRz1baLNuvGJ1yTqZ04nGdqONF2QL9MeKRv6JtiH2een9IAB
lWwgWVW4E73TokSN1XJQThnTn600jn5HievpPFOvleKTJ7AdMISf9IJ6zONYEhzO3N/VQcJb4f8l
GS/QXXY28WfYt0vz0XXWzH6txKJDO04N/b3sdv2t5vyHa1sctFRAjeOPZiyR4Bl3Qqqoi5tm+p2Q
8iq9anJSnivchplOPkMMVjvAEi4+u3kOfZQ4SSBPMPV3o5/Kqd3/UB2OilXN5dibdp9lE+kDrWDA
NEVUySTVN6z2zBVyt38RmOqp0YEvzvTpmGiDFUHj1iYXHMja6jDHVyk2h2A0hujsnvBd7+KH68z/
8rdGV0edTGzXoMGKVVdruzRBzYU0U4NVhj4Gub3hImeUCrN9oFoSq/CkbuZjwlbuR6yTjMZW861+
s60xr3LQ7S/gJ3Ntbs+I5k5AK2JaK7Z5kV0X9bQo1YNPuQ79XeWl7MfZAeQvvy1U0UOgY2Jl6yIP
zyaPU+se9bA761Jngzahw/xDFwR390tgWSokGsFQQbgg+7ikWTabeqKQqbOXOG1pe2I29MV6OWdy
SYD0A4f/BcfjIBnHtGKaPblnCb/fuwrQnTSBrI3uEWrXTFxlT75yXJ4XlJNNDgNuWM4hi6vD81M5
+ceKSmpmb6eDB8/NPkEgR+nhwqNayvzCIHdKD3/cpfbsydsu5laOVgHurNF/0GFFikEYdsXvqIcu
tSFZzpxVEElp8BqZ71DEbigAlEK42nmS2PzxC3uEFwhzrqXxL4mt3H2BtGKBZ3zD+KBKQ4T7Q6Mq
c7HGe55v/GsHAR6AgElBqqcGaqmu5ApR2ZhbIHgY+LcumL3vWWfizNiS8e2o3adBpeBJAbQM8b/L
kJVHfjovuMPtGGBuR/aYAZRnGRPfkQsoVMOYsUDzej3xUyaFFr4HBpov18nkvJt7bpVGCrayhEjM
POOBRsTzSqfTOfk48ti8ZD08v0QVaunJwC1NSTLbWodOSNiTa2ZgGYizSKqIfwf5rjcFENXMdiy/
/Qm3T+EO1i0CpdrMpcMiDn5hTzqHzzl1XUt2RbVITYWonk/eiGgnrdkneV/Aaepu0WEzdrKPlWrG
hSIOgA26FGVuMamcm6r/jGzhGTXap4f3wKk7hKugPPcetpW4YjuceiNXS/7UfVKBOdz2j2IrBOCK
V9y6tqDDGrLacjBNlC3msdfa8XrarhN8Td4nm2ZIxTtoXQxJX7rnPeXYwaV6FcRcHPu+D1hWFxvS
JFhN0tpUC5BsFfR0IEcyNl1JATWrGTS3o79qKHkWcX0gnjhiJEBeSgoi2qrMwOGqKSlorrdr77mW
IkqvG2JNIy6gLjXE8YXtUQ/KrqN1fI1DvOr8L+ToaqOJqLDdatMntM95KbqQC9YD88V5hbLkYLMw
Ln0NWQ8VkArcbkhMmgQaruj1D+2dPZIia/dM3mlI8mCQvEPwMiIPdl/eOlwdba5BB/f7DbMmj9KH
QNkvVYavgPHQxF2yTFMesKy5zXIU2Yu4ECMwuZ4JWgOjlQd1Ju4LrdUEcbhJfFppSjp7pqZJi4G6
zjbhZGNjztWcdMakXPoz+YiT47ue8vXTFi1syQAtSLOpsO6YaZqEzcV5C5X2lBXT/fEHiFYhqeWb
NmY50asuh6wXaXa2zJFErqyX8r8Va9zKD0RT4yffzPadqdKxDadTc1fEyHAzN7NYdf30Hd1JhXjK
TgAdEN/m/0SHYp6Heao/pGAPfhb8IUiKrGAncZgyu3jCDm37a2cRl0EywVEDRQPTgovl4eaEuVLu
sZzYwWOa2rYom0hGuvA/y3rkYwldeqQdL0FOtgevh4BOpdUnYnh5BL+soHnU8/KpqKR1gu1i7vXY
yRPpd3Dpd9IP5d9727jbGBIRB7QALhzSF0bCEqAW2I7/ivDJd9SOFe+NpRvwUQx1u5OtOnpOuIRH
QsyVuEV5vaTWs9J/jtqn0zShIx/ubCLk5mehfrHIkV7/Pvu6EZXIgqRn6MLx9nrp1VLEi1vGAxGA
LhSl440YbY88Cj9VbxlkTCGoNTctYFAQAGUHoFiJpdDCU7YioIqV7JAmQ+zOgQajUCX4TatNhTA5
Gu96qcFM3fbqw2jpC9iwwA5oQ1YpGDIhAr5UpqFQ8iAUfHOlg+NBbXU/pNqOi5EITUZJNUZYHDOo
FWhLh7dDs43eKMhIF9uP1vA3ICmk/4bHi49QBu6O/8G8N6a4klcTQpWeR2ULYM0IRylRQtbIyuln
zDWqH50OSdmoSgVF191XnTljycAZjtNHNbp+adCPzLCjFjdFNLFEuYdD7nyhpq2e5A/HP20kX9xa
UT8jU2kdicqhiqomfQN1+r9uwoCS1/U7Yh5wNGQ1NHt91W4PrIe0LTSZCCg9odzy+nraI3IOtGRM
4TkBmop/VLK+sfIMLb0yq0MFYoKJR5dcNPBTVZAOsKEChPBa2fCgtTE45Ir3Gfq30IvxP2Yimy15
sDVMFlbu3hbUBRaV2HlkVOlRZ1JFYjdTb9sAfSCRGdVviFQBMbiwOfN2Y+nyuZhMeV68wZ5nIFsT
emaAs4NpR1Yoc3/5E+qRxqZXDKpy2bowcjnRsUM347bspRIZNedJkUiZaXl51dD67ONC1c9tSlGV
zKv3IhcoZ5J85dEQVcnJk5q/h+jZstkwRtbt8hoV8S8hlohxfGUacfahMVl7apWkRLzIJGxqHyYv
S9boUShS1HlX0OKQwDN/Zahum0xWQyalk6k3tH/3Rx7LZpC22LDKnYUAz0l2fNkzfA3N7i5/0qUM
Dqr5iJOBdWNuvgTeVgs6KBNM2OHxPurzTylgyIT2AB2p6QicLQ52gTGg0nSTWjuf8g0bas7NVdIx
Z47tKb41O3B1WaJTSdnK7xRvigkpob6hUTTNMC3OwBxK83taYYuZXuxtMiE9yERUDpmjIP4RDxT2
YJL1mfj4+IJ1o58c5YQ0gcMXHjRmHNVK5MZq2daKjo8OF6OdMpqofBEP0HVXXzReqkNYJp08d2un
mmBtSGpxDvPksHJfElJEscEw+UvynRb1shslZG3CS4MGOQeEzPO0ZueR7vAeDDgy+TisPIsbIhIg
Nt5eQ9/btSEHBhhtkY9F9CC3f+pJkDtUl+HtX/asFdRK/tB0GWRj3IBMzurOzDI4iJjfd9Vlxsb0
nkAiPcWVipxTbgw1kpHvc6AnQmBPZFH4PMz0/6eCPSplci41sQ89fb4gHgoTNoDvpm7MvXR7LmfR
smnPkPR69UAoU0O5LfgNFhct5n5OW/a3SHa4+tILxjO09zkgon/LMny1Kzx1YilZMEiYmp8Cmhz6
ctkLztomW7xvnMj9szzH5NEOBFWlhlGruIG+ofSZPCGYfZN8YKdmMPJQUyXDKQb0bP/istgY0FyP
/NJUM/w5RIpkvUujvZFQxgmQyCwI3EDB31OZ/miVeSUEluQBg8XkOTHV82RvV5vQ745Duv6EgN04
iXeosSYaF/KiYIr3YdAF4i/ASjCoGPIqzZkYRNsjNI5tZNX/pqvJLsIZ1E2/PwxcwJqFiJzfvfqZ
c2CkjvD7NOVAlAo2uJpJONhouzkKt3dWXD1OQHRgoBznxdHZREpV14/Q+2p1ubSBUG7uvxMkD6ql
yzz9ElwhGgmgnVh4Lzf4pvfqPECJGt1rHLz+PgjteIPQLaa3ogDNsfO5u+K4vZIO+Zjotsrp8FQv
VXHBE+R1UUHKJHsBca+5L3gHU+P/6JTXBAMab1270DXIGyP91so4cyHOvQU2kJ2aVdW5WhuPBbGq
aF4dDEQfjnqTnhsDZ27S25eZifYYl7NYiG1zUFcaMh8Pd9AFKKlByqZB0w8Q3U9onF2L+O0brmwG
aW1vck1+5V1Jc9L/H2I7s4nmtcZ/MB84R2xZonkrJxeIzz2JM2y4rrbdvwBUFZzEx0XzKva9jx6T
8lZ6X/YVQcI0YhGUK1h7Dx4GE8n8xFYguXIp9xwIyYUTlim/2JYfuPFF5f7T2vEldp7U49WLN5c7
VT2TETsGdhBYci+BTWW61EUbVFrcXfYrKpOlN3pUQFaD4XCdYjF8pd4fy+Xwm5eSWllxWdiTfDsX
tRQaRGZYcBhh1/7oa+WIx7u/W1RVymUoCF+SKHLsN7Bq2cfE7otmFkh7rdlv9pmMHULa/cE95aMj
xImE6ZR4d0HNVMVlIKnQM9fJQ6D5xDpI1flWOAUVgXOHTDofBDC88DA/igrIyvyq5sZpAdtK7ULn
CC4LqXU5dtLcN0clqZteRjJ0iyHqqY3H3yWDRkz+RShaOyoN0z6+v/r9AP79QzYlER2yPjwqGEgZ
7RMgC3R3KTHVXdtf6QMXBPMV7KBVxRYw4Nmc+2GmQYB/RV+kMAn7aHpmdy6dg7rvhCDVGknZCo/P
xrhZ4dX5gMEsGi6MLa8mQumRNQ5OCvIX2dYkMLx1vqoXQftlRS+G1VX6bG3u5iCCGBE9gKF2Qnwz
oTHbQW2qwnWk68LtJ6Rb2yj67Gc/WjERnV9OYnnTIIVeZmTbOOrlgV13PpyjXAo5C8DS9Hw/GswP
4HezRmtjxiK8XvvEudmW6e9Ir2uOtWITXVZrIMCvhhxRYEiEBDXU+PokMlBG3ZRcwxFe6Yoe/V3G
b6rYCtac8+CRm9pCPNDK2FnDmvv3HMO3Ttv+b16w4r1tjUw305/R7OrF/1KhERSfI6O77JQjonw1
2voQUNWM+7CjWvq7oj6n2lx+ME2RU6JfBHYCTfF2vdYgf8OAbx4NNwdyVC10+Rz216Cf9Wc1I6r0
x5y+ixiut8Akhjgo3tCUFG2yxvc9bo6lCZTTLzHmXE/Gm3tEdTRB9EcwV98romXww6ycqNFG754t
4nG2JHCpVq9CDnOo5dp2ZrdUbjhMXTTuiaayIY5NYwft+tJzV0DFBKBuBHJxymqhYuZWxtRwM5ii
HUXSMwdftPupjwQosWuvGSNWTjS+a715uhIrcQUgdp1Bi4dZ3Lm03m91+2G5j+XmdQKrZC5miInz
zAoOidrHEdt42UeqCvJQENwLXRWQzDBUzLvqoBJC3kZXcXarOrnu1yfujWYSHL9xa/FDf3AQXsEg
kLp/OHzAVaysmepMAEAYUuNAQuBC/bJ9aOTxZifXdwVNbNdyJEHk/jkeaQHxVYWQ/3yeEy1FuFxi
FQnsr/on+QIArcBv+cPWdtMeV+WALT936SiUO4BQRF/EKDETXkMlJS/MjBXP6IpjEALlT59SJP5x
HWh/liShGpNs/777zxbI2TY8mcOBLDW6oVZfUp1BYQ/zHKRk4khCgziQH9M3/Zx1WJTG1ms3sRTX
yqk29qodBCwGh3hy28mKyrc7nvCcNQjTBymlbC305BKqEahSnJrRd3fWMDC7ACdmYa2B/De86RXn
6mhg2GP5vr7Pas93eDSzjXAzFRnRAFeCatHrTWu38RP5lLnNMfC8DOS9DHoJjuuLxajM29r849XV
yDNO5Gcd1Gcfy03QKL7peMUPbwl2onPvYz4mxZJVr0IeLULa+g8kQkvaQ4r2AOL4+qeu1QR33fAQ
3W8Q4IQcu2bwP2OvEl0uO03rqGfmZ3dmjldKEZK1JbgYNYZGp1yFMxDyHAy2gw/6a7ldAw0j2TAd
zQNMO5I9/eeorf7Cn+R6YDJsEYPjUT2+detJgQdpUB/4H/jU+CcYYVCjqLr8Cibt+2i84FZA9WWA
otJwUShIQy1bjwJcK3lubCRgY9hdG283KtZlsYFPKUzbc+nCjJd/Yq9GovRJsc7aaMbIfWrk1rkU
Qmoa7Tg02FOyIhWvBeBS0rksYgygkbOv2VubQb8iL0vIt0pfL+3AQ6hNN2jsNeLW58vmZ6rw0thT
5nSxfBgxJRt4z5Kp2HIeDvYpX6d/VhSLhP1NncR62kmLgAXTpvRXj7PSuSBx29WDfVjhPNQftfoT
6EPYlSEAB/RBgKJI+umHM0D6m6r3K7F5Rn+oHYOjaDJEE+dH6ApNICzvyLtVN2QcrIiS+TEd5zCC
SKpDPkysAneaBx6XugSKaloW7FN+gLh01Pt1f2jX1zE6LcHGnodpuhhXqfQAvjHS06l9P3IQGqcz
aQfMLakGKSFTEODzffyvuGYtkkgbQlJr8ynv3vdamIZ6WtrljEAKNxvqkRiQ09hWCg8f0BMuCB/7
Foe3Xq8GGrpSv3+GkHlLuZlNxybPxXDvsEUxil9kZI586+tbkL2tqE8f+yVNazP3d8196KhPXpKf
UmqGdKcLy+4riNuW8HpYLyvlMkcJYe0VClHLIXXT1025b2FgFDEN+NZMNcx75cD05pide2L0b0X9
IIfO8JZSWESbe/U6+H/t5AWYETKBeUyOiZbzfnBd55ghrjZhmFK/R7/YhR2GGLxR6Xqoy+oFhLkv
KCxL4kym0BrV9fN1Q1KIwZ4WdgZyBwSp18Wy/7BpTzuNB9bw90tt5mwhmk8lXTJ9/YhFXpBQKjUw
hWKAXrBDaqgvJtdpu0zd2nN+IT7AU+Bdko6Uv9e+UkcVjhQFMpMtvZ8m19DIYeQz39B3xDKA2gRP
dlIoA9nmuuIgOIXZX7hl1BoxjCEJX5s/dWIOtFMDO7of2woBqV3CK6yGOxde3+1j+HeQiJGDRwhU
vbiXgo1dTEnaSzlKI+0OXBRRNrng9qMR54JzFz+FoBiwx/2UtAhFnPxtwlqAOXpe+f9ceM7801yd
w6P26mL6DIz5X+Ez7PY5XwgfICF/jQVT1Tc/155QLOrdUizGGnCp1BvS6LWOZ/HVkrW/1fmMJ/jb
sDUGkLpZKABxxsE1RBUkZeJH/45t6xqg4JoI72C8rNffstc5n9JXUuie/FjQmMcyqRB9X9f9cBix
VtCMl/6kJPytoEGClgDuhfAMm215+NCC1+e1s9eQ8dvhsOJHKR1GLr186TcCTniQI6vvorxl1zSt
82fi1nLJ8IkVEKi/aSTfKPJrORsO8jQtNEWZTwqWq6tvFSK/QDkyC0WNtlIpWegHdnw6cAcO3n8z
AT58BiAeX4+Z8+laa+NwCHkCJ4Lik2Y8S99mSgAuY2/6DAZi1kuQGspx5DpaGPwIrSjpGJJ1xVRM
FU2YaU3icmIJf/Kxg2eocptdihIoIyxQxNA8czkjWRePIizRm23Ier1OCY7ylH+bs8cZMknLb5SE
dFAoI9rvVbdPYbu4RsuKPTXkJU0m5PK61eVL7po0b9gvNkxeS9zBLvkBbcuzBk5deQpJlTc1Z71p
JGWodU8f19/M3R4UB262M3fg/wGR3q1m8l0w9RjaTGiLfHqX3V6d50dSAXPG9+UcbyGtcMUGS/PM
2JmenvM7MARMKBLdvv1r9tGTxqyxEEQg6VDzulSjsgZ+JgCHPXSSsL51g+Qv7KONFJR3CFPCCYDr
ALaxgD6qgCjXedCpvipMiNxQaCfqDUB9hVph0SQZJA7K+R3pKcXCGMzyS/egGJGNaNbDLifSgHKd
bG19yYCMfW+hVPDv04/UvOWteXj+b+K7KMXZhJySsaMsijuEJsankYq6VNI9oEbgCHUxI1L924p5
Pl8hcghpTrvuNya5wPmoVrH0buC/k5Zbrek2cAl7mNKitAnK28jkYzakEsVrCYEEes4fNHMW8OyU
jRj/kESNxppSKGbGM6swMykINM/0hm3XXaBd4AqDlVHFe4YB2ci+vdRtsJVSlTVPKTV0Ac3qPeBG
0M6PO2zC/huAH0KQgIZe4FA1+anvVhEfhPPl8YwtBILfhPOc9bVVDnaDWGlPldjlvR13ms2V+xe+
gg/EaRUOCSp8onMTeK7gO0oo/vJ7PwCplG31tqdCOKC3q4zzyEZuQR84eJMEuf/NxIup+umulJPT
/zN1x9wezdaekYNogeQt3ITAMllkwWtEwGSyvo/7Kek1vazr+zCbJ30CEw+CP50UfcVqBLv2QcVw
HB6qP1E4s/DeBbrk9WxPSm4pLkjefLoXoIwe+GmpxbosYki/hjY6knwtTGM/giK6GVKKtc0pautN
VqvGwIgArIn9oZTsPWey9IypYvkJO06AVMu9pU4iIopds7BqxSJ9e5p+ODsZaJnaaw0UgkNffm7K
g39hyfYLojCMXS+pWddds66y+d1JQ4MZsvpNICmEGV+0A5Zrjx48Y/Tut+6pydOC/gJjf34WgdSa
EFEW0GhuQEAYXepKwpjoGq6LUhOAVTczJQs/I1Q+sZ6NKWd+LfAfsZvwWJkHkUsX83ZIhv1lcQt4
Gg+APs1RCK3wR//24Uuc/0oeQ6ZHDbeApMLLXttJn6Afy3IPNoYG7Dqd7xxp8MI1ZpczRLT2yDUD
a4kA3N8wAAUId1+pbMVD06ERxPRDNPCZ1JrQ0x7EK0NcxCOMlxORkS9twT2kpg5kSYGMlZr3xwhz
qgdS7igHqG5F+ohIHUGvJASFqk6/zqQJGZ66GrG44BKWmCeKxJcQM+I/iDr/BmO6eO13ZDhH3Zdv
OBJ84WRbRuLQ3oB6EKK11ox/DUzkB6XaMgSBb2xQNwWl16Kmb6dXJklVfjmNWf2HaPsmAGjwhmIu
rG5U0gIq6qrCmsvPPNRTbm1YR+0mef/DWq/DRv6DBlU9tbKgKX3CxA0JzFMW6yNjTczy3D85C+0W
4lGP4/08hljxKaCsrYxdc//T+E3+9AFq+4n2a2DcCxSXfhqnn774f5OzmzxyWbDsj1GO69GDs8g1
+w+cujnEMXUTLuNb4fA47hYZT0s7d2qnksdlhItfUa5y9UG28hZH3U4NLT0XrHNuT7nc+ZQ5SMKI
sHksCXp+S7SSLG1Du1VxiWOiVUF2SJwFpuV0rd5GKd8/IBg+lP7oFtrUVJ7dgyMta1NpxcJ+WkXC
JWrLR/6lZVPr7TwO7skeU/ubi4riX3mudCAxBpPZhQIKwbqSiP3Y4S8NhrPxN9qhEkj3kClkyUCI
+bg3ESlDmt6wXlsGirOHy01mHJYcykAGrGV8Wi2hzCKuqQi+asfUM6eZ+ijddcL5d8T+NVFZYvYP
Rl/ige7YWp2b4bRLe4kMnSZdoyTcLLpYFaatZhOuESnMRSL1JBTif0zgIZhSVUsLxebJKZJW1+V+
WEDXDF300syiWgoN+gZXz6IHYxSUjPylWEEu8XidsVxfrhXNUM+gBz1L7CZzBdqxA0ZFfsQh2fAP
aq9kGpVDYGmIWcVMVhVRWQAZRyRBRn21n/DjZ02Lvzmecw1J2Cvzn2VDTbEtX5I+KMEKJbnrWcvj
IcuKb+1Y/O4o9mWx/ESzefRig2IC1ofzhloR9g8Ia13oY3h3gucsCxkZV71hbDD8xEWWJTLJn9/b
gIkxgcm0iyxPTt4CbAfxV1gC1gMhjqsAYATHtUxLt2Vgy342oemx6Cz1Puy0ydd/qFwkiRVIRM/h
bTsqpGgGPKRAPWdja04aVKRJbyZc54/9IWwx8SgC7q6eMu9FS0tMHcD/nS9g+zFiMLlEVFd9IUSP
P+EJJD8AdYitroawIIPBJIgRT0TfTCYw4CbbO+3A5ZJ/rXZpwSHTt5f1h8qyAXtj7IF9JpoHFCcy
TR+VqHBFBDgaPQ5xbLq1mrXdWkJHOy4dv/TnuU2zVThg+vGAsNd0IvrCETtKUWbfy1qrkDUFvJ62
E7XgRvtKCF2FeZoCV4+PdFmuBUWraxKJc8h4i075RXXg23tD7OO9lbAWynYm7mJMOW0zV7dS9Bio
J39o8diSZ2syI0DcRoVaS5wuFwrGrzfkIWys8COsMMhs6J9XjwUbsIvY+n5m3y6evEHMLg12jCsT
aI5WfbhdgqhdUonnMX4UfXt0Fiqu7NL8YlzL939OIHttrXvcb2Tyw+Tq0ACZgLsL4wprH6iwtLdY
XpG0yQDkHy/k2ee6F/4wv2SA0L408OKopg7KyqOsv2AUibL4OlUMHRdZXRtjRYV6bb9QB1LwGaGM
FFDCf1JzCJLimdEQGXdPrEY7Fj4Zu7OkY3E9te1XvS5GbLwoqgvWl+IttQm6p+fMekV2KmSpCsom
drfel5MBzJ2AlgLdqq5SFZSRPTpUn9E7Ih7aRTMsCfm6dgz0gLAVhIL2gHSs1qdn8c7FZOtHx9HK
rVRV5dwcmMGhHxxEi6jXP6ELv6P5+93QL6Tv6YZwyV4XK3zDSghJoB794XPPHbLRO0ZjpAQjANZi
AD92CFrSg5KoCjTnG/i0H0vnhTW8lsixyPBlRXkSKFTtt6SNLfI72lBYNQ49cxGa7l88tudsTpNm
6cVrQoqGGbhqXLr4f27BlFczvOQt8OPtZslg8RqzfaTkVJVGii20eVzMoAmRXkg3aXdQ0gArpiRW
ZjNmXphB+ZLOu78GGCB2GuiJbkFB5AKuZ0DLoBR6hWvxEZvBglGxeGeuU5I3/QMO1wgm8c1z2UwS
iZMrbaTNj7Sb8y0Lvmpymrc6220zUJmFgutK+5ALFKUCMObpHmYUSj2oCLE+Wp5N9Sudy+Vf4/wI
DXTfwtYu0LMZRLEvVrWYn5KohPla967jm0O89p2krY7y/tdoQxN9BOQacg0avXJ/9SA1a3udhpJO
21Zeizmufk93NHgl11/YfQLj/lgs4443Gxy9Y5eQ2hkCWPHyVvEQiibRAM+Wdzip5AJ2ev+2+T8/
kJDrGoUIgmnR86Bp+MrxdwWzq5bPvZlZRzCqmE0JDNIoapuK8Q7/phsi8Z+nPUlU3qmYur2C7wCk
/Hs54o23J4IaIRTtXx5svtju7XTokdt5vfCI1wWTqhWW86jJ7c+CjHEcU9GlQUZTBRuAuPpRGme2
yTiPXJAElXT2VuLyETCWh2xBCYYwbMTgJ6CxdbKOYNpxayVbmr4qM8NOjDTq/Iaz9EPSQZbEW102
b5VMnql1FYmp6Hc5r8bZYJTgQVu3WGJSuiGURDljAA5QLB31giF58oy/rMmUp6Nc5asx6Gz8sEtM
YFJwon6XEn6JYw0peA1xfxGYdFR0CcxpOZNp3B34emr8ajUH1KHBiLOZgMbt01f2AIQheY5q3Yru
nOBemZ6uiUKE80049ZDeOZcGnrJIPFnoNqO9aChwyiOuO+oTFz5b/gQrhZSM/QbgGlDsSWiQ1NCN
oDhFrLIbKBmdqhJmPmjr71WoPw1GWDqK/U1GGmVnnR5ppLgh6zFsrxKpVRs5mZXUG4pzK8ndmRQz
4eiAWz6fh43+R+uzXmrcHDG1+847hbb/sxaOrUJJCI5Nw0kDTvJl6GY6HFpAgX+OdqeEBP+I7/Ce
ntaDQ5ieEUs1QLMNX9th/7i3SzuAEZfWK4P2+5/XVgwvmgEqpv1pKehDqPXh4T26ALW1Sc1pUtpM
69Uxa1wDU8e1CQkhJ8LIvgon0JuRAKt65YSFNzSh0r/h1o4YTzGf7UcVqhn0oxo9z2TNGh6BMv8e
YF5I7woA5fXFbdLutrySboit0eCefvIeb+2satZ3bREHtDDEqLPCrDB++sxLV/yHpilXc5rGMQGK
8OEhJ69oYgxEqHE51FKEoLFnXsZd6akPNNsp+OpHSaSzpm68suGdJyS7zwL5HeGW9oq7lMjIsiDM
APyvYgWZGmfO8iW4ZOgKfigdQS/5gUSPwa3B0bYzSRbbQUCwyN7tCh3YrSXjSFBXLGBAkU0ra2Qa
s//hJyHKcqP5aseJ3Chg6t4ZqfEVbV3s5cVGKgnel1RHlXmn0lu++aT8mWen1M8mJjcDYO95K0EW
tCNXOdPuMUHZtPaWU8XxHMnqBVO4f7cfVojLRkoAC+fqlaCOEpgTdJ+nzM4uOh+A3GlAbst7DkjB
qva/BQ95TVxODYlv6eWqbR2WtQbcjyWj5H0Ch/AjC156+8Ft2TbUoWK5iTz5WQgZOgxo5AjLA3nI
UaMvwLgqrUlcutlcIpli0Z0qDxX8rJijuzSmkweNVEcKnK6kDfM9K3jWj/i85ouJL44QqwxZoDQg
GrCPsdPfC978QDYui/SrB8qXgOB/1dXrO0rXgn9BxAxSkLmTus57RmjhrOBYphWeu9i4P9XxDpYF
sBGNUCQBmq3z7uW7x/duy1kptEPHSwWMEl6Gb93BWGT8ptCzWJJQDWwNaBW3mMMuSGKk8C6IoO3l
+jOUMN2+csndo1WlQYs5ViEoqG7gotILFLFl/ieY2w2LDfQHMPZSRDX66Na60cr4nbp/hs3HP7sV
TKTW4VBiDsBImPBWlh0+AbL3z4NfgyF0wAsNBqQua2oZt842Pbrczx5biuO7jDcIDcAqSWHV4fUv
fZehTdTRrZZtfMVuOX666yoZPIaQKJiwOEKFkznnSkg/TOOICox0Fdo4T8+Ha3ia2XuS2q2q00oq
2RBxYYmtyaZFcojx+aXP8fvjup+G60edlIYvXqLTJPXM7Kkm3o1JkVX9aT+6mf6tR4akbtqIKQFt
mx54xeddqoBARd10VUwXFzLbBUDk9trDqi1g0Odeiq6V45qZ5uTBZZTALOFhYuVAIPDGqyU6oUmL
lk3PHIZtDd6RPzhmlsaZZa2D3EvX4fy7OIGKfbTlkOVyTuhHjhjWVDaVcEpfJH8dRFk3Yzl4PpDH
OIqP2h78Sp53xLU6QE6PcKlaiULr7YFb+6ooQ1LnOuld1s+76uTUIYcRCqdQ3i/CzA0ry2ax6+iJ
Zxs+BQGB1LNfpRUTVMcmQqfHB9jSXyYNJmtd1BMKDhFbG3VCNNQsaPjCJSGo23b/d1/UgERZDcWC
/5cw0d8DWLuM1C/86FmtA8eLKrkX4SOkb10Je7rYAtn+NeCYBCljUo84IVJLb/oSBlTjA4Z3T+O0
pOVD9YlurNDrEk6EUrYoBd9Mir1Qy8jQYo4EOYtEVp8qsPPQ84grXYTloIuCUHQUiT7Aoy5fTiu4
dnqyaimzoVkcyhgpVDcBkRUJa/w91idE56hiJfOyQ2GSlvcexYBBtkarqRz1+aIeL0OSrQRKihvb
1YixjUpPQruTCRkSYr6k1o2ezaS0GU2xmZxbANoJHk5gLnCQdG7douJBm9+FbSpe1CiM2o6dcZsF
93dlF881Zcqro6NTAy9mjh+de76DobQHjbCRIM+OyRWTJXmtBBPn4ILKnb4KlUxoKZTMp4X84gBE
4P0YXQOASathGivURLBHyARpSEzrHQp+AVbFVKdxh85rnVsxNVn9zY4yNapD8dvQn2FcRUECr3Pr
rhFCnPNftrdWgP/0mLpH3G9dq8EbWun/HjtSn80UNqN9ivphAWl45NaGRVy4sDlaCtifh3YE0zYP
JzsoGSPUWUFESb/ru76zk66GP2TZi2GI9wxwIgxn7ZRl/RiJlsU+cDFoCvpJB2MfOdPIXrxkdDa1
+BQJdQHCDBZKtJJnNSyHDzZTAlz0ktuvXKWpQk593A9dvoEAYETgYSj1Ga9OQiqZFd9OxdIrCM39
Cym4lfwDLJA7nHHpg/EgaMVCBwD1A3e0aCMsZhZgaVTmcjdNrcX27d7IHF9PtrWqRL/5bygb07KX
qr2KdL8MAmKX0jas/uz4QHj2UD3nK1W0BDw9OKe07jI6sYSqMNPqtDTOZxA2QZGKblccq/IK69bI
FEko8IoBGiRNkzruVv1ogrrNIdaLU3R0zbJhSOS9/2QzAmMVu1AWK0wQofQJw5CYRzartIpPipvr
q5sUMU2Nw3NLoT2ujjWqqij1kmmX5GfFmZKzMHia3p9FjrOPV3jRj0BwvYd4qUq7OomIeFcpjL5R
4m0MvIi/R3tbADPLQsHuxBTzYR7RCWCTCSdz3uDYqM4zidzZeC1O7QJPPAhDLabXceQRI5kF2rfo
Dvh9WSC3NxNMvmMQa07tN5m7pm3uDcoWzzOvLz9/OkSWwwSS9NYHpEel1iCvO/miZNt9nW8zTZoQ
vHlFQ2qqPtjExKqlhl3C0rXyYNafl6Yk33eSvjJVkTwmjhn6A/wU3rK6xkWzIt8lPJbhKizq5CsG
AzTf+cCTqw0BrReJcCj6KfwY0I3AfPo9E3UOF+BC85R9PcPobe0biVB1X+jVERgKioGYRd2h5k/e
NhkK84hqCWLFz7+75Z9Sl8Ie3K85OnJAgN2/Gt0uCC4d8YtF83JiozU3W4YKnVXtOSxOyaYqKPL3
jCCVelW6iD4jvwHvVV9m4XS09VC/1edvEFscvuQyO+V+46n4UcysVDdaosfpsvONmEoUuQn0Oy8T
U3bhYNc48w3pfcAIxlf6siJ/4/Udyk+k7e1cczKaZ9iyPVbwbQjuAjnZGc/0mJJxOsIls+hfckhu
w/taIqZuYWYHXHXpJW3b70p11zQGixvy2hE0/YpDYkUIGzBWNAyBYU/FHEyv2g471I0F1O/gBUK+
kv84mcHGMKX7Gn8o/92/PLSyoWmpAkfR6iesH35vrj9bvSUcc5PinQ4tTv1iRfWubh3OH2Jdgmqs
DysDiFx/fkL0enAwxe03BL2XJDW6SqRYnGLb9aqyBXqF6GGtcFzfeJxxCeo3yBFutqEcRyWQ37Zy
uTkf7I3TfKDahzEvneB9DXQVut4BbhTenvhXRqaHWq1fBAkyrmJLhLdh23J0YfMSVG0rdHcYFRww
ugIyFM0YJIkUZhhcZhuXh43Sy+6dLP+V4QZlsgemKYqkwg07VMQOzQ2PZvGuHmOJWqcwGkVev1Ee
UHKvH6K9yKrQSpOXVMQighvfCklBQW158EasX2DFk7G4IQWBNeWZOkbYxU7Iqx1kWxOFACpZWGii
GJtkeaOv75004GdwbktYSf7AZnOfM5PrhF8swM5MSA7DSJQRSoK9Cv//eTPakvrvUFVTcd+zpQQ7
9A8JJmZuoaKwDSfgNaE4z6ho+HGSqNT9EuMjozSKzURRRPJC9ReB5/jNV39az9b0+lrvdNL565O/
oPfBMPhtE6JlZowUd0W+fye+iFhW3jx6ZZIMxWNQ8U6EXV7TvY9YBMDNFsk5+DlvoCM4ukFbBHSc
aLNqUWW9/wfoIk95VbmqnVC0bB/YXK+z8+7FJ28kEKv5Guse0GAIzPxJjvR8swWj7RETWasmbbq4
a9jNzwZ8I0sRIAhWfKNceacSSLix8iPSXvgerMf9B9LYGJXvpG2CvnB0fjPwC8kUrqGp0pyVqwiD
Mp6dPvfRUQ92M4kij/0SM81bJ+UyooHhNsdlFS9qExydHrlck2j6B6uoUie92EYHNX7RjVlLmn/P
PgMdUW0ePj1Nb3ev+AwSy4aAqy1eu/0gnVoq4ViQpW+Ge885eXwT8RE23iyGTudrC5i2tfl6HgcA
emfJ194llKExOpYz/ASdbw/Rn9d93MV1D1o2bbTbv8FoSe6qfM5K1UwfX0D6oeC/1bxUaQIDkp0m
INyfCLCjw1oWExFN/CjpHOU/mO68x7uDcKLpXikHGwrqMv+V++n3775tnK/LgRSGPYRHzrQiIgBQ
Ajks5zPC8VaUXv+AYRBPWy+CywzkHqNfySrmszoMDfb4zUQnCyikDH7108k2Myp5Sv5fTYnNoqwg
KYJne6+rOKLFqqsMZZG7O31u+YD08zajdeBSuiR5WCg1mLAs5v1cNxaxvxzgKNy78fp9s0iZgBb9
lATFrgVfZnLQiKi8sJl+CSSso84aewm17jb+WL/zb3Pa8V6iEdVv0r4idj9EFe3pL1NUZbbKksWA
/CTBgBxNgCzttfSzX5mX9i5YU2q1gBVkvHiyA1OpZYfiPvtDmZF7ZFaJBtg0kvGTq+XvDygeXoRi
Xzh2+Mw67GQ4alaYVRRn+jCEm4eVgdnNT38zoE4Q0wr4cC+MFixWvkeVcn6Kg6PUf+HoVH7BYM7c
uYSIkyEnARjETYno+Ra/OrsJY9OqCjBOi8F8WypAmEHYScCGHUmuAUrh0wvC0UtkaUXjD9WQYouu
i/Tbo/2ekbY/agL0DGxAYtzURnrUbi9kmxxLQifpp1z7UVTv2k8MSENnckQphMVdDAwq0nk9/sSE
maQgBsKl8ZO8wXYLNlTzFP27E1oNVNGwzrk28jyCzH3jeOKLxoL/cTsFdPPMImIPtnDjr8Ee6msG
60ZJlfbJLhm5dHahuVQvdktcgsCt0jKmOxxsQCPQhU/AC21J1GN3Dihlh2kMIe3wOu9opLYOoUh0
chuCNEfo9TLd9JxNuNg2Oxnq9QoHIvVdO9pDyjPTu0mCzTpZLdwzE8bP3RbiRJG+Tg/TFhRe8soN
5GKolEZwmWYwj5laKb4fGhFrVLnRYHL09N0qmomjMZ9Mtmb8bZzGv+Iv32xSAlwBPAkRisSd2Ybs
RFrKGW8BcX970tbVCfbDqCAKZfL2gf6WY1XAyn5SOV29XJR1iLinxbrmalQ9359eeaP9xhgMJHKx
d3SBJlTQgF5I0eWy+ThtdCntG6pkn/lNe2+lU64/tVEvQTP1pMi4Yc1PIaFKK409gAKm1QYA00og
WpRR9yJA6BwyurFPf9Kk341IERuifzl8qVKNbYG/lHHVjtfBThXgG7Kwx9V1897JReuG9/Ea3msI
YDYyBt8erOoc1BYeIhHpqBrfbkDot/4/nMPJqXfj0SrHBMJwWA9GLJXjCmX5zCeuzkAUEZHQ3p1t
Ftd+SxGZy+rnr9wtPe+xIG0N/NJ3b02pwXDDRGZ9nFt2DgOCmg3YB63Aw7NDVI9Tdz377Hk70KCa
k9jN5I7cFYOUyvblKeSRQKfBJmEFL3A6tzRVmiMIBQznHqrfzp1CmhzDzMxvQ3uMcB3QycMKPO9Z
lPnrreh5C0KTBz4ODOVAZMWBMmpblYnZsENnmBzfKjDVYAuNPX4lh8u5vInpufsgrQ2ZR6hM5Gh+
DAb7Mr38SV+HlOoNBMx8g914gdxBqq/DzeYa3pZimI5XolB3psW2xIcfeXkSib8yvaUL3cKCZa+C
Je7H3hUoHKAs3aAzbWWCx41eqvrZhsaRfoB7Yj1AFHmlMl9ZUoQOrLJ+iPEldDcqU6MTgTCRHqRw
x1iB2QwMqzCNqkLDr+EbWPqNBkuem69E9gvS54CdgLF0ibV9DktXhWEmcZQJmENOV4qqs+MOMe5Y
9H+f8Coq5Un9eEw1pgyQaaSQa3yCOctDU79XStYutyHT5TqSzzPT/Evim9PnGS87qhpR3fqSGIR9
eEdeVrlT/be29T3o70bbb11mQZc6mwo5NK9DRSUzkcYhddA0TDcy587YYmQU+GCmRUB2CGAPRqug
SXdE3C2U70lGwP8+KhFnitilf61vQfxN3BzprZcpcxri3NlbS9Ct43S43QvXAHslmXs413hTyfGo
ZCBLOjrW6T1JvNEn2cp9cLZY6rB1zA8FVkzcKGSuS3NPmrHtEmzVRW2a9q/ROkjGmszS2mI656dR
QSJWVc3flTgUJRst4ZUgJlStgifLSM5vfY4K3soIqgATVC2336MXGCJEf1vw6ODMO45ayln7eZGY
F2PF+ze+ELWgVkNN6NmIQ3SOcAm8p44izW5hJ910zER/zAoRMFNUNsnSZswAUtbxK2QMlrcLNiHj
TAJy8droQg41M4NlfWmtlo5EE+nfEEiF2etxcR5FV50+R6GbXW171TIFv0tU7hzDX+IulR0S/N/u
uRDO3hdHRZGQ8N4UuSktJLQNS8Bqz/5CAHi3LOMImec61122t3aiH4IwRNQ7wtOs67oTK6qkeIHY
n7KVogrxLYpnQf/3Q005d1mBwj+nrNBJFfWrckRimvGW018+RYmBz6dQhakMCbc5HnLZoqrmwEAI
YCWtCNaVx2C7Y7RMhrXU4yKqcg1rr2oe7amiFaTcISk5cYimBHlBAVplbJgKR9rIv1MXOC0HJIIJ
6sHSdMq78zEppWrOROp3v8uaI7ioe2x0fc5vj9lnfpUp/AoDTActUbc0uKokGS534PqU4TkL/Tg/
uVp5zu+YKfdGl68TZ9HDSk+aN3rDkM+W6CNBKtgAOguH5irOb3cGhdF1hvJLGNFrzjTD6kk7QD9L
sSOBq+X0J3zKu4C1pPQA8OrH4c1XiSCgpAbDih/LpqY7k72Hl0IqqqVAf6a+5MbnoC1FG7FkUvAU
Iwwz8EHQOtCSaADSr20whQO79+twuSToyquqbVvTKZgjxke3pevNRBP75AcxyhJciQmnXNGTwXYJ
fD7SO05F5xwxvEn2s1//TvNBz2Vk7/7xA4bcQzeHd5izc2r2A8MtYs8KxcawdVrBeNcWaf0LlqlN
eDRcYTVpyJf+i1dCYHbnvTcRM8TzFgd10qaDYgg+dqJS33VLcHPyPBABMoQRLSOjizuet7RUV1TX
CQpit3WD4JvhcqKoAgF/BdcKfJJb8mPIsIzNlj3x3pwkX1in/7vWtM3XV8dq0rQLxtFnmgAo6iL8
ycxBragtxK0nuU30ckfv1bZmv6Yh1IjLkBZuPNNo6x4U3dBIoLfLOMcjJIXp3Nbwy1BYbgw5AzbK
PamreED2P9tpBA/mqiBKQmeirhe49XYRsoDOhoCnTyd2n3HfkhdRdBhVfOjeAAjcGpJBRKhWHPLn
Xh+7gAtFjGKmNMoBH0e7pWgpvNYK+lGZYqKG0Mqs3TgdEsva2nPmkvMzczpr67lheONANstYLb7d
fAgaH9y7OmLpsdxqb4grd9U09qZkqxtsZkVCEWZzt71Ese5yGz+vCBikv2hiB3X1q3uqA4XWSvV6
xwmQvpX2tHg0MvqGxVB2Xrl8IOW2VOPWyUyCoxzDMU6kLTb+ufdhWqlrt18eP75Ecwz3ka8gW4kT
p7MdVDabzx+kVYmRprX0fitsYGUz6+tz8SFTWFl2ElizBoqO9ws66jXUQmik6yudppLvfSa2ENuF
yTCBbHLI8G/QR3djETAS+v5ETUjtOBNpVboJJK7Zo7hn0h/oIzb7wGOwJvBoI0XeimCrKuTt4Im6
CkSDgGhuS6GnUlzV7lp0Nkpn7bJM/CjlfY2ffkx3rwqShoHeBNmmnyIlh+/UGqbJ0N2y7ZL1WBbT
HES01/cOLYfIy6iGpVBX5BCChoc8OLJGbHukB31KN1p2IGvMeyjouVcM2KeBZEn1yHDUrNbNXzyz
kVbry56KbQ39AH2SwYU1J+YUXEGFLjdW0bsNKjlgjFng85XjPSAArSfhJO1axvgDYcYoseub1kf6
Axac1xVzWgzInxrYu4Yrvl6bMrd+vjNodCiDiUAjws9q75xCZvMu2ZrqRpiO7ae/SgagNk7/SguS
GNKhKmWgfYXlOMoYh+Q7aEeD0oinDO28sc5/rxOLc0yvopFt0mTKcXOXAM573UxotFc17mOKIpUh
49QERdwTJEGUfVmzfmK6aJaxMrK9mP+KTDxI6eUoxN0VqrFd3tu5XNoU/ik9CkQtPHIcnaW8eUae
ahEtBGruNvEtVhKQ5h/gqIipzVJxLS1SuiMKrtDt6TwBWWySkL1b84mWFFbU5vdcyTrIldUnret5
LbJx/t5GPQtTTmE0EAdKeluIoN/KUX8wIpEMD98p1Qfzf1cTeUMUvs4bGvInS2zazBhMYNyTl+YG
NuXiVoSXY+e+fd5Nx31hjec9lgpU3l9IeK1+U1RRCP+EpQPMNKQ47HZ4jke7ODZkZDsGZ9YCfAFH
dsRGH/jdX9DE5DOst7U8+XrbnM8Aa+QAAKtI0SOtgqrRtTgEEYlzNna9n8WBmjchUtDxMdqB/aEh
SFuYwFSC9QbYLGCCvS/CD16n78GXNEGM6kcV4cB/iIEQqjB8LNihygXMihYAAF7QLA7iGCIDDRIi
7UmkQqFF5rdsWEPAxxRJyboEKFaeFFyF5pxC1zFSf3K7m0QuleEOExgEsHui0hxZKo/EWWlHmT4b
uL8sxD/D3Rbm0QtiE8bulH5XAQVjiRWnUgf9GrbTrQ+hgGp5fbzuI45aInkLJRtkoSJzwQNtTb/T
2WEFGMINTGuThr7EWpNEOV+3/7QVT0eb5f06uBd1xFAdGJTsnR4KC4xb2Soh6dwMoDqht0IwTcBJ
fkY1WuoQrz/ZqOiX30odpQMJKbQ+jOFT4msCND0SCHOc2c853VtYxVDlYL7bLuH5RAy3jlyACCBe
S3OxQHoy5W8ZMDsFJpIG5Mt5D0Rke3t4DuNC9VEnLdy48z2ytQ51snCBGI7TMWiViT5VyhOSyNSH
Z+wyPxJswvsda8VgYqk0XrO88a1h8qpRWokccUPYaToXpCP+b7qDTV3eKm7DhJsC6+f8w+nR9Q/h
/Kh5WLiPPm2mfE+QYjI45h/IWn+V57+IFR0v2/2yUKbn/bwOgt3zqNiZOe18UIlgIuar9DUrGm0Y
HTjBF1q1cflyUJYwMtoX1S4UAfU7nLcp/P8kj3Qc2ofNY4jTDA5S2c538WZS1R9n/N0iLtWqXoly
0U8QEu37r+Y/y4/oqGE5GDcP1tcbrcqsXXY8RP25gsuaiDHtGsytdl0QX9I0RtFMj1talGwnvV8H
5RdHrFV6UeC/PSLSVuwwEKre6X6hdO6N9Rb8zf966/Vreu6tvWjftR+lDD4WmAEn7mznCWJIXH86
6592uGwzztD4M3kwwka1cbY5K5gXaQYUqFk8xST9DcYcYrMSXJ6uLwP+tocjHjOc+zA8eedcEq7c
JK+k1GJ0e+8+jxM5IZpTwuFKSdrTLOiNSvXizjOVnfHbYjmjRR2bxrvLXOXqYSuYV1jK9kf4uJV4
UWaXYYeJCUtzH02jVEoG1PuqVuFpMzRFNGO35ua4kjfnBzDlawQbLfarNM8OKeICGIoRWTuGA+0g
mqNw5q4EYi3UOhAQniUuwMMHlfuqzYdxRUjaHp4kJRc3frTjjsy2qXItBhTbZKmLEWUOZy+K9Vmd
gcyHWE8ZhYwGtljwukyv+9rn3SSjQWq38LYIak97+7RgHivo8XK9ldqSpbF1nMR8vaZ65wQ4e8gh
/fUHdcNEPuUjbYqber4mbhDt5CkWvdvdYKclU0WhT6UwE+gYc8j4MPNLXJxF4CEV8dpRx5R87aMe
Q8YQW8X8qSdQ3PWAyp94QsyGqEkR3bCpb0YAhsa1+BdH5Ejafi2NSLbs2Rb0aZRbkWrfJO3D6IJD
yRjzti/lPbCX6TIJ9OBJDMW2V3NGlLNIoGrnNnzNm/Utubzn0+X1hk8JHh6Jb6Xh/roWv0/wkqfH
+Pr05VlKoK9AQ/V+vaJKJgp10bEcKizY8GeqLUjFFJn9nKkvG5v52Q+kM8MQCJLFzXyk+1bcHghT
uzjVAsglL9J6V/hRUN12CVgH8KGGIJrYItoWoiS8gzwu6NFGt+UgmVTTeFzU22teNQDFrnUuYYBT
HL9lm5iWCQ/XWGnQve69ILx+Z1oNjy4E00Fi6Oha9/QSbRkHavXuluJaovM7Lff09tlDOT8o63U1
jfGGBdV+USGlgeEpC1ls+J7gdJIOxXzb7pUqdiGAevgiBsCtYoDR6Efjua2LXyn551opO2vyiWQr
HFXJItJhxtLYg5hHAbD/+9Gro9cBEvo/x3Fic+ky3f3zJwlPd9aI91F4Jce7RdvRNqYGyXXyfsbc
KnLt/glHJ9wUEm0pkb1E+M/4v+qEvtNXBfGl1bYPqFRMMLJw2I21jmRvt+FavLUqHAyYkfkjHEPC
iHCh5MO50iMdMjlTxSuEvXNxe4gF876fSc9E6GZCuPnu5K/dnDmsaMS/rDwXjKwNQ7u8zI0RDZtZ
Z+sRtriHJK2rK3/ftZb7QegYzPU7oCxNVhxPeWXVY38LPhY0lT6T9R6kXMbqwOopvVHklZjr9LuL
VjFXHgPPU7jlmSDnf/hnWw/uYKX1u0KRQDfPjEG6f0N+eyIlGVurHk5X2Xd9gpSfMQp5NP3ITq1P
vm36LuvmZe5UPTHDkwk5XFCC/sHBf4+QLfjkGBKDy1Q/FxQdh7RDus5PRlHPhPMVcdzv2GRThGXm
AxFbI+pWpCak8MiQyFqy7GNqqhDVtXuL/EohVd27IZKYkGTEdS1kSBRAdnsAjlRIfwxSXBt/44+d
rdUNyCRzvETn3m8a1V6G/hSt4GoLcl3WyYGQUdtuX+MHt9gNnh6tl8+ZSHeu/8FLPoIYV7qPDPpP
GnlDKopN2ThFb/a3lV8bi9NlpiQSfTlsRYNMmgJry8yusEslHy+70FK2g4SwvaCGuO4zSzMX7kYm
+BmNl8iw6XMi85qaRzmSRfFm9w3zitps776bIgRhwq6ooGx7ijebpq4YBVVaKdcusK8QOzqTiaQj
BsR+SA4YlfUC7jdYhdfoTcz0KIB40LKqQWKP8eFKDhZ20+qanM08Aim39ZeW25eNSPn8EJnkLfTS
uqlqfXlbOfeFZsefhsP35QjtDLlIEXJ3fmGcAvrAjau8T1UIbrQTy+iVUt/T2cjUGRX/bTZu76Qb
NpnMIIuUdDyT0hOawk6tTSn+YgmnWw3f37fxZe17XsoLsDk5e02IVBVYuYIXoplTajT2dNNOYnxN
5HRVaauzyIFxJ9v6YtvTRM8EX4BjEmd8UfiCcRVXJ4L78/bH4i8pPrMEen+KOj/nfWm/tBTuh+oW
fzFtkWJwaWKzZO7Wl1CYzT/t+cQvI7zyJZyfqEBozjRAo8L+kHVfNdFEIckcjvVNAQlrfj8FB12I
ULsGVg4WDPfNZ/i3PNtPUp3Q1s/8kVCyMyH+h2PaQY089QP0NXPHhB2iGw0rYQQUkA7El7OIrGEz
w1mdjamFsqUFz2kVCp0SIrBz7yk+YkcGSMvGTj0qwOQDEeq8zOC9sDGxZRpZkcFTHui7F/8Qz6PH
oyDsx0HGXZ3C46hdwv95ntbJeXSd3HfFK437AqQDDzNBmukB/HeW4oyYX87J7M0ekF36sqk2eZTF
f5DbRotQiIuku3NuPM+WWTHvOndc5+TFekm1FEYJ5vzjVelPhr4i5Dm9QuHsBhQHVtxxdfsmPr1p
hDctrUzqmV5j9G6cQ/e1/XulhWbKdB10Q21fDrsrVhdiEQvqiXufi4NvD8tdojUCSyxVmv2Ye3fS
jvUr5oxVlvkpFAnKMpsr8Wkmn5zHqCgapo7m3cJol3+7c2wOjuBvXgnDuvycZDkdDmLF9V+7DO7g
+xDYExVXd7HRAXDWF3mP79ReSvzFK37fLcFP8Kg1muFiEmTuKkVWbKea0eG1XJnNE25lR5bF6OQ2
p4qnd8ysJ6XvwQDJbM2E2b3vKlcfULoGorwLTg4yp2ENsK8w4v/durHi/fS3CHxnfRVHfXsCdq1P
AG5Gg3BABs8s+SqNLEPHTJBLUJaSj3OAuJwfKv1equAtekX1UikBFswlzAp31gAHHTl05hNtWSmP
h1+1XLp6Rb3dXAWYCSUIsfFL8LWQHNHAYvPw3gNkuy9I4Zbjwc355qlqmJQLNcV7VCs8VKZE0PWL
qAKV8YqkdSW8e2odH36sn9eOoFhnjoYrOYqRbiLV5ibWd3n/QaHP8seb/hAMqPUZjx6G0J6lEDpL
12TN3UXn66kXhai20z9K8M/7mBL2mg1g5ecvlcNqd7+0iFhm4MMTxHDKstkweYDugp4taJY5cV6e
928Odx60E9uTQss4zIBPuveOgPMHeAFdqx3+XXYR8+C+B+G+8hpKbfjPnF2eGD2ytGE3Ez3Kd73w
yLJMbhiCHuEjs/3sXI8DZ7tRDWrZORiFUZprKUsvUSL96Vp8aLx+vmQ8ZbvAbSk2AQLikGR1k1RE
R8r9DdHqHWJULKOllEzIinvJV+D4gmm9y6cWUEMxnHrDIw3k+A4Ao5vVWUwsjHmJbKecx9mcki7I
mRTnlA84TNMJdJAp+o6ppaavMHCpgRNEFlA0JElk7AF2ShYS54fXWt60NOBCZ3Gg7MURD7Y7e+j7
+mzm2b8VcutmUj7O9QCx8WQ/hnPYj1Y5XLNM1j6JM94bd25KUsXmBzp9UOViA8KepaLjtavZ9/JF
FFuf9Yt0LGF7JFzbhanhu6WcL7JgRQlmaCykBJ+FAQNPYIQw4NW+SXyPIiD53Ql0TlKx8Ar27mNk
s4q0Lmb1FKcKq80WmGMvkRiK9uzmQXi983DIMqSjGQjlU5k572r2bOtJVEEgEoYDriilv16PTBoB
kOjkmgJKkdDuCUhohTUTannys9t/zqcgXHAx2vzlIm0jP6VKNo/elFIGaD6tuZpj1Q0PzY9pGKqq
k+Dd5a7JH7ELWHis6R4LD1iY2uJ0g7scVNruuAXici/n2lN9XYV4tNYOH8Wkmhj1x2oTdn5wkFwY
ymwBZ0NcVDEKaSB7n3+f4gH6qAZvfu7ESVpaHaq+p9A5703DWDXcFABLeZK6bA+0IZPVTYSPe6Fq
ePbLQ++hXnAeBRuLaoaGUrO81tkqiVNUxdhxD2FRt0LLOcE0DrkYVucBgcfAm+kx10dIZdzPJI0q
vVLOY2V+yyNV+kYpE8F7LfNRygg2pp8MkXJNXnRDrpQpNwFYqIBn0WdBCpdcyVQVP99sPibwrehS
UfYT6rHmQ7Pjvvplp7hM3zDYnR5mFExjOoDE5tM9T+Ti4xP0BcuLzu55Cbp0B3FocixkVRJ+MDi0
psyOSU67tom4KKb/vIAgkeuRI1XEkHNPlnxwuemKwa02wdgtlFadlZ8zBnUlnhtZ+El4tLMIZlVU
f03LIRURQ77ezznk3+yHJQjm82siQSDN6QbtfyI4OYCsXfHHeVtMe6fpNo9dFshn+tSABEKXHKNu
+6Nm029Ly18m2je9YsmT3D7cFD8VJ8irQCt/qOVo+/edj7yQI2we0r4dwFZHMPSuytY/MYou6SLr
TsY59AFKXpg5IagRIdJDyloD1KmR+2GbWMDVtVC5eD/gTuJ1/qVRsRwf9dqYXIv18SQwAXDKV0MQ
wjmvTpqFRFDWnaVh/PRE0cTkBEzZKAlUV7rbd131oJRitAfGCw8Z4L8TCYRpTPiMb2S0hzfU33qN
FCAGrdQ/X+m8/booRUD6Dph+XJBFXea3d0pKtyK7hu3er3VQdaP4G81buUyYjPnvetZK4YyDIBWf
uIjE/ixIbAsk/PBbvqz66NuckPVaaYsPBK3L8yNWmgte+9W4z9r5/cqfXEkXNPMHJGXOShTrhar8
rIEFge0e+BXHOuKygZ3lmOx61MzCQKPtZzQ8llliMqju9FXo0A0eb1ZBuDt5l+NmwLw8gQvsfLDu
WW9acmjiyDHECAk9YQBEEqng5nm9uk0E0L1T84v5AhBZZUm/3Ws9kY6w4OflHgweBGnnOqux5FAp
vJVfr3l4HF02I9HuH7bL30ZD+AHH6/H/AZQaRpjR9r0SuVofhgFfSCysJkbWsvvCGS5LKvIvWCUf
h4epNtAxA3nxYs8w76dY+vsK2ItyQBa7D9VfzV2zKus5DldpI2wdFWjpA3jkpQfeV52JfJ1SL37o
7JxHm4A9fAa6+qctkT495gdCZcCzdkaei1RbMpCJm1LqGPwHHeKbxJ16YhAWLzkC/ElJayZpiGj7
wsV8wN97z0oQeuFxR+rN0e2w8wjaYQrMitk12ijMMGpPMycOfch0hkbKO72UXjx4dsVLqnYoL4hm
oyPEGoPTR3PYqwD9J31xbFp4M22XpMyKbVjHm/i/agONxoXjlTVTzqr/MXxWdBavuW1ViqHQYj/Z
4xanxX+QIsDKV2htSuEDRlpvbiBk0WEAZwGubXxB5JIA/GP2JUCzgz5mrDGedf2CoFyBwhLSxo0O
JOiPRU6A/GymiMLGTNTSBRgzoHPEu9NtCMIxfHhJmXGhVWvukp97AgbWMhKAOIEF4F8uf7H1Qe8Y
18btu6u3/aKlI0zLgWPj9XIJdyde7BchjozGpU+hUfgbQJVXtQcC3VSvCRg+e/j+isbQceQGBhML
ANxlDDxd5cm1EWZS04tskKNcJvTYulc3R9tRv3tLZnZd0Qo2d2Cq17i23qQwuf1saYp0GFfc4X56
qR3GhzQ14YQo1IefUSXQ9nmehVaEdcQ3+3L+2XXEyWQ6QK/vseVQT2gjniN6kB9t7dcFb39gaN/m
9AhfTbKwbc4tQ7rCreEoLuYIMSPlB4LxHq3eL5vNSQaG10gqz6nvre8hykorheTBjmUAIVLqyeei
TNIOBg+hK8I29/8AT/d/1kzHv9Pmx8Q6GjBX6tPP7HVy5qp8HY1OX3UBu3lYigfkCS+g4zSYeihd
HRx/9Nm8u98ybWTkjwwLNQzTgjJXTRuzdspdrBtIQTHMbggmLQCdxFPCcXsRBnEismVNjrZvtGBU
D+Z4hZP5pQpYJtaTOfdsr5YptR+U06B3/LPkHu6QZP9IcktLGYJ3iU8a16NhGyVhOotGkJcCdQ3o
CZjGSu3AYjv4GlVWoZUlEx9tieL7CL0A7H9Vwchv5MJt62jfOONqj7zwlVPojaCcU7+nw4V3RHwx
2sWs8rSVCCreRGA0NbBMPNFD3N/g1g1X08CErdW8z5s+4r3RbdCFWS5mrO9y+W352qNVM/GTSzzo
thEhEIi7KYgwUfvj9ZBIenRUGuhVYR9cB6ViD6fWwTLe9ZLSzUSr14QHTfB7BpYLKnxDxq7Vtf+x
AUswaXfqnBKlUoAb8Dy55kc/RCv3vTQAxDU+7QCAb0xk55ivkbo0hJxN9bvDZKTtwR3ZxZ/1trUf
I6UkFfsA1U7UZw/SFLapFLkhMM/4OgUpI+iybtO+1oLvtH4G3DXkQsfELu+0+VUFwf9V3J/XzZC+
6rEGy50TKSRedUvVZhaum2R8+Hl7sn8UgLEbng04FQ+Wcxdy7J4iuGhaTKBMOU/tncFKPqZadSYi
NHbK7vrsofBACbYUVCDl7tlJ67geUdnWjxtwin7F3PeHRe5p3rGi99QkdZgqQEbh/8E7VLCYXuz5
CsQ6FR+ZGk7bJCA8iE4URC0vrnO3CtUHPihULXa9IKlPs0r5JAQrbUTM80q9dR3WSdm9w8AN9tA8
vFMNUqY+QNM0qolBjNTLVAydenppBhLg9ioqp5wuLaC4GnYLNY55Flb8C4Dnr5s+6bCKd0rUot4Y
BP+te1JFPh0j0XpkAFZ6dortjMntZp13jfKGAeOl6aLgDgmHEYXCa/s2n8/FZRo6qsK2vbNKPVP9
tsG8nrDyVCCnRJ+Jv6g2M5bh0EnOwXGILQyHAkJCif3EWsk+Z7Lta+s0O3NtO5B5F0R+nyFXqFI/
3jZw+0h8GBOqztpZpQxTaP4/Q6NYtC/hfzzhlaBrRxMMK7u+qlTJd08wOyA+jhexCquBmTYM8BEE
MDaVBYLsCFtW9ObJEJTXwb67qufQ3U4XHr0/wDDuLZFWW3K32rqgEYGA8on1uE8uadriktbVyms0
qUl4Cr2wPZtOQNRL+1S5tnTC9AXBa1TrSmYu8uYCR8LhB7vA2oZswTzgjWHpSrRzrMSq+HntRPui
22EtkYUAd/1BQcZajXy3VUMdSU7D5m6z6RUjj0/gyiszZf+DegG2jBocBuOtosssC90i9mhL2aLN
I5rjxrplzY6qDrgD2dYjqWtkZnGwgV1saJd4TEHrJIJ/MZeBWxg4wwvqz4WWAEEIpLrql8ypP94E
4TgAp56zDYR01H7M1jXzfr2A8sCdqyewnYgqXHQXvB19gyH5r52Ho2mwviI4WxSupdSYJ2JJdAgL
zB0lSo3eRv/S3awSO2agXd+trEBdWgFqZMaOj4NXq7Zo5LT9op2Dpncyyy7Imglm+wn9RNWeZHnL
C8VKAhRw9CmTupXJIb5nStG1boY9WLbB4XzF+gIVUZMmpaBPE0ZfrE1OHnQSlA2ekFdM1cXO4sTi
8fFG3+U2GoBh8OJtmycbIYvW/tJdlZkfCLpNpBAYd7XvfIRzv4UuDrkfEnxzfky//hckrukVSJvK
4sTgvzCpQ8L70APD8RQkscBynE8wkcCJ8L3uBBAaBgjJDM/GIexcGqqIdDM4TVU1ep2D2S8pvLH+
rGnP6R0rVqT+0sB13ItZ0rFs1TXCwO6so+EPouh+rRAb380Qa/J2dBPBxRgX9dlEzU4UFn1GDkst
OooNocCUdFH5Tf7ZWa8nPT5cxrPtEKr69r0GDxWLFZuNz3l/OqJvHZSy4lWLBkuCGgH5VscouNWJ
Yf8IQv/jPU7UexmuyHRfIMBQSfY4P6N+2ycPbTVyHPFtOwL0OhHcKLcWY3k+1bf6WWPM46i3Rbme
senHFWTVeav8K0xwv8Ai7CMDfiVYn3uJUvFts2E9KqTOSElQdqGyasHWs0/l58CFoAVzLAF7Bwsr
IEp1xtxDAmoCEtNVl2cddlUOwiDLpePVKJdH2LqZbIWTI6VHcUd/zxDOXQgFt66320x8WPUlaGXt
mM2Jt0FlCbMIClwjUZT6RTHUPyVjUw/vqFBhMSDCStsVYTiv3+vJIZvMO/bcGkrWlkVEaPTEUlcg
OWo0MCsGUX8KcGiLZq4+wop7FHPpiHg+MP5jFXnvI86EqJtJiRevKQn2yJSmH+UZMuveaDLQJrHq
Zqh+6+JnexhokJuUMa8XrHDU/VwaoJdymdpjUPqv/zxWIssGRK6ZWmmVz4vReS3MD62jlpOhdDRT
VB5nykYOv7H9yhTPHqPJ7p0XtsgUSVsOIa6xI4nABWKMMJMksKa9rudpb58VkzxZNO1WA+u6E9SF
/mtCgmSJuSP8RN7ws/zuJooUDC+P4N/W7LpDTvy0VZuWnh+n04DimgzQzMgMAnyhS/HFOXnuul+h
102JxvFHfHMJjPULUAOqVVUa4AGJmfqzpnRCVYcXTUftHwSnWVU2qHsnpm09gP/SgJ6bcothEk2Z
BgKLlPMIXCrYWCp5JFzD4hhsDasR437H859mbcB016KyFgBGmjUWfLpJwjUowAJdAkhQfzmWG2eP
e7/L0jTtKHTvHr1DaU9Ec9kJ2ReVx4doIQjH9iktRJ7ZUlXRwWXM9DPoXE4e8i4RnTrlo62czRzM
WnDvnyy4gbm2SO8kmYmXhQ5dcqZjL1D4gT0vLxxvES2OaXh01/783XpTJv+s7/ARv9woo2CoJnFe
ttxR7hFDNqjZfVXJ5mtT2jGNf6QyEynyRzCi6QI16Ilc1o2hy5fcnGeWkGakozOsv6R/lFJsR78Z
yW0avx0NLOtbHEznAcHW5GKjwwgpSojHGVHrOps6LpFRbcqO4Sy0CEV3yKMHvVPBsNRwCYPlgAXS
hzPy/+bfHQresVkhNqK8y0KAcwjXZ4ogogbGdaGe5FyUA4bVY0WX4Ydkxh4pghvN0f6vjUpMhue3
elY/Jw/F0E0Y5IYLqHcqpD3Wi+PmvBNIqCT5c4JXSAwTfRsvygvKlGSSe2axnRFLx3a82Fsbbufn
QQRTJFCuMGDKLiEHrE9OqU2eDnl3Rp1KKyiVZovA25v8HgFRNF00xU3ANYAoq+P+CcED5L2Qws2x
uKgcva8jzL0imwwpuI9yfBvnd0sYSVf3DLqd46qbMLvkO6uDv8bDE/m0B7Vg4nWwiZki2fuYVKgg
BAC+gaKzkAAAI/5Hu077Q5mDp8MCXOgtWJtzQAKh1w4Q4iIm+GQuTA2I4f3xIYTV18DlDNDq6jOS
WuH2H0ZQgQSyGZnbJQxfB7Yf8cC/CjrpeqwBNwsyvcSegoSSZOSQYNYbUEqmKeGAkjV+RassRo21
X+7pDFOs0pnq88lNQLdbUSs7/y3vcezNKdUT/I4hZQAmVghuRuSzc0/KHJf1qvIig+RpsLeLiBJB
6re4RKmDkcHT0nmu68/fVQ080Fj2uDOA3Szj8MYmuqcyvyteM3Jd8BY/2SPZrS65BwquDHSzwM+E
LdB9LclB0Ke3SMJeYMndcVhBqB/E+/LqcdzoBzcaJmodiD0vDuB6SO3qoinibznQCngoKwEuQPK0
9nkkqrX5rtqyDJh8jpMHliFMyjpiOG7lhto1KBvcwA6TSAAVSGf8e/YH5CcpX6Gh9tNQA4n/ZCk0
aJuGV+reEtZ4KypYfigYFDedFEvzepapax2ztzv+YrKVzANBw4kVYJay4tOuoVgHNNgEDMM9Br+V
ENpLEJD7Wa6ZYZsZzEVs3b0yzGooyicFOQRnEPG9Fs12FzgPIiIjkpcyrPGQkm1Agc1QQwVmCoxU
ASVv14N2hfztZy6dRDyi6WwMI75waIjc4oIp3t9pD84qSUDxkcukZq4q/rKdKnk5WEeN9i5yhsa7
zOXB2g6YWTscJl0+fwEEPhUU7b6t1loVUziCB6rl1/sjV8IaI7gw8q3ubZsev/lhno+WtAEoCfBv
u/WMAXyMVM9pZKWWfUk9GOTzCOZm7agQ56ddAMjq1MLL4T+KsPVlXAo5QZp1rvDKMpVWfd3nVymV
bq/uiSNsVIiNW7LhkG0vvI7kaO+vfu2Fsg5apQcoMsGwMxGmZw5T3u0AmK5hwZEImTFZeSEk6JIz
R4BzeySrlKsTdC0697tFPKpCLOW1SqXJNoBJMtMSNgbvJPbHh/UGoFNDN4AW2s49dn5XGTx0A73x
2km/wSyiUAf4t2KEik8PVxge6bH0dw9P8hJZUrh/f5nv0dTlB4nXJ10OLWIyTsSFLF0wEcdZcgk0
neVYaSdOAt2Y7pSm+s0/eX77EXWubtEJBGemNy0s4ELjsHimfc9yrWFgf/KPpfi/3vEOzbeSaFEd
tdQLorlkxNNLwVAJJrW4XNDRzFdarc+sf+bkO0p3kZZ6VYwgcjx22z0TwOPbdzPq4BvHOg0AIWGW
X5yxCqSp7yMzirYaUnk7tdycKHJwh+A4fQaii49EtPtgBSU2o6aZ01orG0CLpniX4gHM8//toOz0
MY/TRpLVevcC854W6xwAftFNyQUxsbi8twEFCHHM31c/JT7+N09kvmGUMOmyf5Yw7/WukNKLu1CX
0vNqGtB7ZIVpYZvq9ZOJwPOfcLPzQ8QgmszW5Ur4CkEWVjgrld/BgRNELI0PINwlaZqM7Q40DnV+
pu+ijKIBzr3vmJePz3KRpyJBQogoYSCp3ojoaUaRbevudnpY4apQLEW/dgMr4xkOORcxptmn/Il4
0EhaqpQY7Hvf+4+Pp5ZTCX1+rZf5zEnGCs5fYThwaI2iSPYBHWuYDI0VuAfaXYI/auShHTTNY/fR
3LxmxYj0u24zt+aPJU0XHczOpZOpPPiBAl9OGrRj8J5opSqj8MZ7BYwKWT1iDeBaMnYmUTkIFERt
9NabE6BCOoCzgNBMPLrDXtMNqwPqWc5ma9mR8w4jqHeJ278E0E16MzqoH7UcxIMB+M4AQdqxEQIs
kGYuAg9JQZOlopr1XvRHP+yEN6nvN3yv8Ks6Qo4/VOOMj5fbvzKfVDCxMG6ku6nV3IBOulZ0IjBP
igc4hFiBvcPRO7p93BpyD0fQosuyT7W6lym1wbaixQkmeGYTw3TXS3f1WXNfD8h9LRvP6wN5O45M
50ZrVqD+AEfpPFXPqpPn0eBJZftGgAYuzjQJD13g/DOon0gbXnebTbtXbEBpWyGVr7TBh38j9i7V
0PycDBR+/fMgKTt78NqDq9PhmjfAt6xPU4efcsCSwKJsoIrIu2IWzWaWVVbmV4C9wyPRR/7X08ol
r5/oRRogmVn9LoXowpn/Nk/JMHKOUUXOQQ10lIpgBiP2ITuzwSk8BH0uj7EIoq7bT7wQlP9dUTIy
CvHd5uVEnkQuQ+cgVHnbhdkBhhu4qnSYt2PByPNtTDWtK4AWRcIQGLr2nKMxaSpnG8YRogWzF6jT
F/wS2oh2IDj8nLTGhjajH6HcmVGr6UpkvjdAodVoc5h4vIuiGu8HF/YXm0j2USMaELTJLRorysbj
Nv8FJAXtDIV/fyjypcAtoO8v9L0PpgJZMgdvD6ZGPcn+g81V6vQFntl45AsY1fJ3K69D7KbU2b+i
xn8dgBYdHnHy5SIu+4PEsz0z8bHulaH/5Qzkhyn8KJclCB6VaUQSD6dL856bx6yYbI7JXk7/DXDj
UlEIGqGhC7+rhe6TokNgfTxlE9o/qSFnvOdPVT6RA91BP7cqC4cqAcw4QQLfAy2VKNii33KJybQ2
oEf+ZcSrFf3YllEcRVaN1HbvW40JxPWzMufLhZZd3KCnn+9lUmPcANiOO7ZlFJTB5BRZCzlDotqD
O8qaxqdkYtFvuFmrtiQ1QedtxYTkWYoEGasnUL8iLIAzemSTcQinVAywC8qmnh6TdLPP33fSl8Tb
FyCQqc70ao0/dkelOYxeXFxWtXdvi4aN4hVS/sBhCM3+kQFsQKMYRjQ0iKNnERXJwKINqVP+8B76
KB+HBZaJ81LAzJ+0+Ywr4/lu4a0NwanmY1L6Zy4WlSB0ui9N1QyhFSFfzjCJFD6p7azxp9Qs6L65
wsVthairwqhzjClXr6Fj5OV5iDEuZo1oekDrWF2M7EG5CjqCjs3GDgGWilUCFk+Kn9TysAQLyRp8
xM/gQmOaayIUpPuTw5n5AH8ijJGY9SubK+8SUmr36eiEPUfqnfECvN6wpdt5B2xKuF7WGOVlZCgM
kNv+b1Tm5MT/rMK8CsFxUX1rkZCn64A0QU4PxGo8SOou3U7i50lorP2ZGxImJemGkI3rscFVChvp
F9HWAE1vDkButfYfG24stbBdSXgSa3ZJVqO+kv+6ymQro87i0gFBQHkj+U/aKmu/WNSlUmQb9M0G
K8B+gQML1P0EmB94uaaik1yNHEQf6kEDVFRI0ac+c65h2ebS8bAcGEfitYdtmTrpS0eovDnKXOWG
8Q8dRri89wSZQT+D2IwuvoDMuDSOUMS233+bKaKdpuB4XLuOs4hvnm9C7y9FMfd/ejPI2pZiB0Xl
52oL5addPp/wADvDHmiCGmnTcZ2SCgTWiRAujE/UHUF6B9D1S9z4ovVysnq1YN53ObFE0kpXjjJw
uDmJQbpCMVoUacyGV+SniFC6qDyksFUDpw6f6o7lwmAMGv/6d5F1Rl/qaxShS9j7UWKcMJ0Omgad
ZymMBuO28dXo5MCyc21Zz5gQa8jOkpKkg0CRimVHYbnTzlaOCG3rfWVC0ggZeVTDYi7t+w/8we/g
I8Yfvq7r0RR0XNr0Tz18vTEF0q5RU6AbOKsv9U35Ycyd/sHvcEhqgZJIrrx/eUJ+XeQ7qrRwYIVd
ck2e3me/8WcmhhsZbOUzzNU+EpwADSDqzBq4Rhc4oSubRgvisIGlXtKSAI8kbwkS7R8w+41/wJBa
AUs3YIbNqXp+pwmCJb31rWw2Tu0p6mTvIdUFCmxaxeRUHu4PHAXKPB00p99eSmoRYZpf6AdY7wka
WfpkdiKihYsYKfpPDu/6Oiuw2+szEfSdbklLynDl2Hap/RmawQIg7f33IsKPaozF3R6T3gQYsj1U
wLteGvsEm5M+uUpJm6i8Vw8x1LhptJI6bTatmyJ9Yhrx0VLyzdDybl9G5WosczZMinAyf2llEx56
vZND5NR31BjrGdKxTMaZhiGVfE6620Ad5M6l83SAjKdmjje6zV3p4Yk18jjfNbu42UB5FZp9HCWf
S3thoQIRgpIvWINPw45i6Yuwn+A7aGA4GNwEM1oic/suVlZD3TBSGLBoRvWfRlISzqJP3AXUu/F3
0KppgHdWzb/IKnBK6/w7pD3GwwpBNESbN+Sy7R0Wm8xI2KKXbM8VjC4Zl9OuQPXfq/wcxj+UtOc2
iOHH5b9ulCIjc9N+SgnpbaTInrGbQrWqFNZ3omIbIxLLmwfTNFOfsevjyGa4f3T4IQem0JZ1kbcb
Qd4JCoeqizH0emtAsh6HC10i//pg2Ty92KzBW4gpbWvodq5lejFeVfIW4X/tpeCZUZLHDwixWjwW
qbv9QCWsFhoRTJBRoaSxZjEywJZJ2Xv/BkhUicPZDv8T1diozxfu2dZTo2Un5i8l5dxCtrvbfibF
Zozb3rTXXMl66O/l56GaEGpjpHPUNsxZmwj2+UhmfOqIbhG8hXNET8S9h/0b4yF1+hEkVGo/hX8K
PXE4y+GH5A0sw1lx1s+Ov5qmjS4smyW0nw0z+Gq3WfBZD0s+nbI1v5PM3UWam+ZUkDv8kDX9D4vj
L4Afa/iPcxfTNIg+KXXyzDcc6bvpc7ib92IBRePgQdvJWorXYBZs7xIJNrXKRktUNWwXNKdSycye
O8VMsWD/eAS0MMS+l19rb0VXJuRG3hgwyTrlr2o27MlMtXs3qsfalm6dBbjOoKDPMUxplRUy7vYR
Lo0a1GghrnbftkXeEH1u+VG3zHTMznNIOgdmA3AS4oy7D5phN8pJg58ZxqMhqsbZENBibdlWbvKU
fq57UxNR/2ejoYHSosWYUYYvQMBfh5Bxj4jPJEqycDtV5JAV5q31KWixMdaW7dug4bubXco/zQsW
FDUTZjWW13cCraNFc6M0l8j0luVsQkcFxvoRAmkAWI/AXf6hjaMRg9H6sxLgbBvafSWundUMMNGA
kpGegwaobwnv+5fAhr838sbqp442ZjVyRTgCYPNy4f9N7Pcgb0O9ls+oah8RSslcEEHb7uSlXQIR
dsKYTxvmwLA9ofEydBBycy329SFG3y275izZ2HqrYcz4lXKXjuHrWTbO9Pk1Y1t3yjo7/zNg31rb
ERRxzVNY6oV1FvAQDVG6sUVrgXcntccd8USl+DVnX1B9UQ28TkCQHtoiATzpRx8k88cAk5FXE/YH
xMGyYCTDa4Thv+ISg1A7p3p6CD68cLtkJVQ0iPojwXK/m15xLjR24mACz6wx+npPAEgycLWxLNcH
qbivq5bZGpL0pClpKQbJ/FCGRMvEB+KNEKFWrRjeUfrQojtEwuqYcKjwcwYXQ86490O/m4eg35p4
hMQxTQ9FaDDP/UlvcQBAshgh5HUylTiRzzE/4zxXUuWRbSGEtHwO4zwY/6f9vZqZs8pRw1ddxHZv
0LiudEmOHwmLHhoVtqRllWoxamejFS6D4iSTGs6hkLGlO7hTtjpUs4IFj1nLcqBXWKYqs0twsEyK
gE8CFbs2oHhdjxqUjLqQpYfy48wi3gArFwr/IDSVpwGIVQG9AhKOKnw5rdrJfBYKVxDyIZxq2Ww8
W6E5MWQKZuptS4Jam1M7Gs4gbzO4Rp9tOEMoF6fwRoEBCEm5wlL6LS6CQ/a55rCGWbLP7szNnY0D
BWIaNfYiyyIVhKr4YdEsQicskGhN5BLoR7V2vXD9smU47pyVUJd1NWr1HPWwa8xHSFH5gArgFuAS
4C4kt8lxpnaAAZm+E6AWlpit9DVbH3EPuXtXfQkvpMQjRG5voQsMpkNRsKYeb/P8KaGzMW68Ffp2
lq8+kZiBOdLIZ9g4YOKZ1F4er31drlFXK7Az6w8Q4vsSSrlgvXuIJgJAKwDmwzV8PqYBBGOLyPJs
slo9+RVpiUMVSZUpypPcZlbnEUYYvaobhSW0pKRrF70znG0Cbe5CGWoHFzNLnMEbS70PFP3GwJlD
baHovC7iefN8bDLFUR8l6w/FD/Xm5q5tK8pk19kBm7HORH89ivZOrIOUnnc4n4izBDw2dU67XJwA
3a4Uj/1OcFsSIsGLJzy/0MeDUcsebeu/E1vMhW/yPAMxPPTyw7uS09b8MVyYjWkq6tOB/SmQxhCN
gWL4z1tgOMru2311wIHZadDnpHzFBcK59NO3+bM+ChF+sxXIL+1vy1KgqyHNGGPrATP9slZqQlOL
MITUO2eq7HlA4rB0uHKNJTvKaT6Cm35uP2lsqvDpaK06oUHoTWyuykjpZRoYkarI3CIFCumgv9lP
fZLpNr3eUQJTEwbkvZtiKxuCNXaXwqoSDVTpJr2RoZZZhdGTeNON4YsT1yiSmmqDS9XDsVmq4k43
UVdsPP05qvVjHDeWp84SJp5S0V9t3gpA3SY1vKX5MG9GPizYtHsd2lGLOH//wVJ+rvPKbBkz6nSH
rXimsVDvnLRNxgKz5kZ6MHquhClK4mXa5WeU6MMjhtYhLXuwks9eCf10zx4qGt2Pq5KaHPrDs8U8
/nfBllWwZwOgs0jUE0QwuEn+ZA4GHmGmwJ7HM8bkhljFTXFm4+K15RT9QC3fE9g1MHrSYYjpj7iJ
T/U4211qpLz2cAdgFGwhi9ObWLl6F0f9phEGAmG386+xYsCmJGQ8GBM90r3k4U368PS/cJGGBMSY
3uIGJfnC+59DGKNgevOMdWcwj2jC8sFdgv5OzZpD0+uogJIi9g0Rornj7gBhHF/s9Ob40vhBR7IC
NCIqibQKRHSta85ALR3Y+VyG4HIPBBb0WxgwEZw8Duy9eAYPaGVRavQ6k0mFAtTuOxa98+jTDHZv
je36odt19L1KGPk48CQDKOkzJ/z/pagF1luDmVZB5WespqrbXP3uh3PNdLajfatLW8YbMiJ3SDqp
z8TzmK2Vo4uXfrunwZl8FPZAW1shhQdIAyesP1OurUwMbuad9xg4p0jJ01erLRX0Q7sD5xXB1KlY
FrxkNGnroQ1vBZHoLdAzMHGwesOPgbvVmv8Sk/TqyGuxZ6yp3LPOBHXu1vmuFYcSOmWyKxyGOxzf
SUz2cjMr3l3zQX0YuKTMV1h4CBth9PHjbzWDQWDmEbQNrYvkMbIDqnMg/uZ0D4q/+pMfZTXM9ri3
/pG+G98i2ze8VTJ7P0fkrxe6k/PqMt8c5D57EkdsrkSGFaI5mNjWCgXfN0TbTHHwp7RDYe/A1UJ/
HAmB2qV1i8CGUetvwik4W5XCx4VLSHIcgXLi5ohNsOD1Pd/M5PaIgFY21cODE2syjawOPuS9JLOf
OZ7dfsa6nEa+ie/kx6hcHF03eJBNEQ5FLdU2yiITFyLydz8GG+RNrUoQ4XYGrULXiF6F5CU48bds
NyLLbrwKYlgcvtGG6e3wX1DpEag3SUfQL0Nhptn/DayXbMupLhfuIpBEDPEPWXDeLma1kpqWc4jZ
5FnyjHRwOj8oX8CaKfYdk8I0C/CWGZAv4Cgn7RHzVOuRQXXl6TM/WHeZSvEPkO7PnJlTLGmCzJBh
V4gnW22XUQ7nMmMoZdNcA+il6mXWY1A/fQCCoidovl4MTwAxT/jK0PD7W0/cqWJMilEVXga50d7M
5ULBEHzIt/PqlvAtX9uOk6s1MliHu00Lcwxte7ky//Dzu5a90/aJy8ewW3m1Hndez7wmsGFHdFKX
AWF3t7ggjHSrBrKcgHoCqcyMvwiw0btUVKnjZ/8BVO/lfC/eyswBwLfMd0y6GliOXu6sHlOeh4ht
MzVNj9Cj49L3YOYtK+39QB9Cq3Bfz/4GTGonK7ukga7y9jNLcz0TJKtr4a0udvdwEEHLDnffrnz2
rlRmKxUtUlkYhXek6rQlmP6kplovd59ww2hmR8sri0PVOy604aZ7qcpbWI31ij1EadfwcgHeYeAt
hrKuxDjTDfLaLGrxQyZaS4KHHFqpp57P+RvPjuCJezBGoc2mdKaRXM4LdvcjKCih/I70nOVjhEYE
XWuiMU7EaEPh6K+s/wORjGTwC3qUGL1iHtJEdP9yrhlYdZbeyiwSKhRg+Th2ydlpj8ikcBUMj0vi
x9iam8PgdXQAetMNh5YFosrf8/+4HvXZJAcBy72YrJ+lj0dmtFgNKY+7Dgc/bPSlxrMJKTR2tFmR
DFO8kc8fy7+kV4osNdsPsuUmBX8P42vJJhv3pM+DOd6uAq1acK2BMK31x26K+3qFc5j7pxfN4WzX
1olWAKd/dxhxikmQMHFRz3axLYxwq7P6XddwKAMUKfzzYJ8gvNZ6uADoVISdB4OSwKWDSrsy7dVA
5+ym4Zsw04rfb/xFS+pIYkbutNblM7FxxoiG9eXD/o9mzhdLS3ZHghiUOkbiGi7nr0FtETtsCz1P
rGrsr/OhHqn5VJL5nPPLbUCdD17Eq7H9ukafLN9kH4WiP7x3RkGWSHnKlVIXwVDlgYgD6LQjcwpb
otjSkdVBnxTczeXabIZXKJFf0oRJwi5wR6utyenGPyc4zELp9oBX0Uy2PFj/eKtkgemJHDgDvyRe
mNCd4OSWMo6OizjK+rOc+84dEa1R0olKQZQQZb1UlipX/hQBlCKSG6eFlTJ8dIzU+RGVdI5piR2O
q61ufmnNNuS4ydaP/jNMj/7VedD0+M6pHI5SsO4TRWwlm+lNrZJL+nemOjXp0GF2Z1x4FEGqFaFM
m6SQtkPKoTYzDH17FxTdPeAGE0dk5xpQi8xb9IFMeqpWnSmiSkYbqeHNyNbF+2A/TkplhwNABUUb
Ozjh5hQvw0kb5NUz+PVuyWB20BGZZBHq60SLwNWhYmWenhz8dj7PtjMQbPrDu0MT8kPxFuxs9zMU
puyEZzVGSyHHz3iucF+zsJe5RzMdnTB7lgyONGVqdv0ZR4IXLMwv5Gu7hljmmtvCrsHZ9AKRPYxX
/oMVjPJvMWOGq2bgJ4qsOizzaekzGgCWCj8cu8DNZ+ss+srxekz6WKpCFYSsRLafskhynFge0sDS
gikrVeVLG6lsonUJ05/F9jIR7noND3inE1m76D6eemfqN8pcYtwnKOrPATRf5M8BryU7At3cIomV
Negr6NDK0YwSqflJkcxZI+RtwK4v1ToK/Mp/8J7m3nKwjE7WOS4DXKRnTz08BNoXy7qKVzETCRmM
W5bJRWq0ilygeFsjegtLI0TfvvH9/JcSL84AiiMcKURVnGZR5YjVRCsjG8PUWxHquFQ3yK0uTzFM
yRfeGnP6bwCoLHmuzwKa98+CVOpMakxmsuOopgVF2ijD4kt4LEr3Q2z1RwXOBugH8WgbjHk3KxAy
wkuZC6LdYbQx956W2OlV1MFfv+Cn+lWmbsQDtIw4GTdAQ2jB54LzBNAJCryrfS0MnsFCP+p25DNF
i63B2KpnAeHhBzj2rNEs3xrcnC3PFzFgAkh1HC3Ovvtwrg8OPZncdcZvyc6i5GB3L3XWT5jasGYC
w4KUEpqURr3TihsmNRvNADhEhLbdNLuU4B2nGivNKRez8U+sbA5YhrzifQd4DTeIHvJfgvz4XgsJ
9+LEN5akobarR4y6xDihZzG9bYAJxQgFG090Es2Fgr69P1tx+0RTDUr04vAFfTuO/bKilkj/qtnV
0hrP+2+Oy5Yeh483T5H9SjWM+vZTqKmpKBLbgMvtXCv9Zk6+TEfMuiViZR3NT0LcfcHVzNALtjJG
eHNr5iibfT6dC83n/EG2TwAwb+yU7xa4N2iJ8Hi1KwitI51fXDtF5LmmhanNTWdTRPmfGsstMfkV
u84zjwZDyCVjajW0vGMgJHt+v1uy/2Uq01G+OTytfz97izu7fJ1iAoUJjXzAld013TJq1wZzJwHP
tDaKRFFwP5GPdl31K3ftNb8kFd7IGpKVB0msy1kdvEa+NbtSW/N+e/BVU5aRfKc6BWzLwYVdC0NM
VL45UlzA9v/MtVrhf4NriFqSnDRZ2ZgK+emAApLEDpi+A3Q1s1g78Y1i3sQSXy3xo1FHElZ+n2t8
ZPd7Ebs9frGn/84pFKPRrqed58PqZ53xhA18wZ06PRZRneibo4kYXzwn4GlYX5CFAbhYveJ61P2J
/1v0Ibo3n1PlIdGrBYuMdb5Z9g97+m3NAZUUp7SeZqX63UVnxEzsS4eV2wh/kWi4QRLGl9VW4ydA
+lbP4tjWajRf86BEPB4oI/XgOwk5W2i5fjXGO/4r7/AvDtoLu/Ur/o34kgkhIcdIPqtAk5wpCPW8
fxf9bfZ2sJLQ1e3ZgOERkk58zJtLxYX6nRuXn23T0Przw0I7mtY8u/SzNf+fCMTpv+GRc58QueoI
w+i3QF/aiKwtOqwMYGyt/H68VmcGNCc/tkvrp2gGTeofsUmrBeEt+sJZ7mlRNL0iddkD+QdnByKK
nY5+oyhh0HjNTSw3Nym5nQSpBHiLMCBwm0/XIeNzDW7ZxZ8yLnwN5n2RF0a/HwLJqyuhREIf7mdv
IAN2bB35PopLlbkl9kO4FGfpCXo+Fju2vTlt1rFtaVfAsBMAu/SOdG/E/X3Ufdi9iTryKp8UvXfW
TBAAciPfFheRpKr+pDxuF4HGbusyn8S/1UqX/gFnm67/UNVM3YobvTEvzzVfUGu/5zEIQfrO6Eer
bQcC8PeJuRyeqeU1umy4HMSq/L62eQexUTq9Q1+BYwqd3CWuQdomSpA977PO6Q0pst8oElJ+epeV
V+Ry1EjSIMI03wcA9hfh6u16RUpeD6A6W9VwOAD2PqelMIVRar8OA9v5ai34IO3f/JGshsNqCZ/3
hPmKm1MaTG2CuUu/DCvHxcl/C7ttNSew0ffdyOq+YPa+RpPmEJlHTBiNYl7qFBWS8YfMdDOUIMyX
lmUhEfHOJ4IqRB27SZjnCg7ebsl8czILCjs/etVvLL9kqMcPPVx2zkCVRassykmbqsnNe5ONwrlG
p/8VdkeLy/Di6v6fclaM756ovS89My/AGMuSoj4lKWGToF4tfiHtkgeVAtVJVx83kbKHMDSus5Ck
naJdBo0bLUrjigVx63IajNA24b0h369XhlZxDt7BBBYHIl+K+9i72k8oQ2YhpUI5CS/QLGnvWFah
zjdvtazReqXHaonkk/4bbW0bn2pJj7IARs3RntHLjba2V7h4kM+Sloc2DZ2xpTTQgDnZH/1wwkmF
pt+M9uIh713QJyH5fIOpFBc5qEVeNG01+FiuRmktdj0WyRFoTRZrVovoMpD9cJTM1rqv0FQ2m8sz
MVCVMYWsJts8tlG4mMSFVK4OxT2XGlaq98koWnsIeED1HuLzxL1gvRksn+xKh9hB8P4vwbtnEoxo
fDe4SSjdSt39taeqez66rTfwAp8ZcaRbIPfTgFkEkjmcaayqfy+ZLzn13MeJyLZDHSrA+PR0EqJ7
zwPHwmasou5Fv7RtBzCVEDo3s5x7X8gvTbcaUNyOCx82Br/GcSJJeoLCId8491tyq/9/AR2cyMy4
I7sNJftnddFPNUSeKYL+UP3mPnXN7gxowf0LGUCuuJAWKe+EHBJr5EVLm1hhfYwS5EYDEWbwngnu
96wojOEExVANZ1lshheiDyybk26baHfZtwate1pSlchMmT1lnms9+UPr8/Qc5rea8TOQ/A35bFJx
j60Q1d5cL+1XJYIfefWz2zU4KFowjU8Xf9lSoQORp2iJPxYLoMoAUdzR0kskaxqCOoiScxsN95i/
08qa2cX+GiEnsc2I5v57oGAo6winsH/ADCTLxI1PuN/UClRp0hjAm/a2MGGTGq6wsXbWJg5nrzKp
FLEkUd0S3xkI5uDH3Vr2d0drba36M8svzwZYEKrDZ0+BFOMKaBobaiXuC5enud91OTs2+kzbOf/c
TuYlUDj6+y9QGqbyUyhgk3hWfkXNfRuPbaPrmA+7YnHTsOXhgoeaaNZ2LZPTNz8Pw3y4dnfdcqOg
WrrYj51FgDbeJ7eUY/VwuTvQLad6ru3nJpLO5zR2Y7Vt7q2X9nAJuWnRZamJ5jYe5vjM7i/cTQ+c
Re70hdn2yyA0vzSaQ3G+iROLG71OHHFyeeHhL/nU2C38j11kssFHhG4ZpdFidfOYMpKBr2h4XiKU
D7JHBc3RuycslWtvdhZVn+h3yVFKoJWabdheYU9+HmNjQcYJ8IW4XPorNhAZFJnllw9c3MBLrheS
W3HaU1c3y05gMpRNClqPY76jr2y91kGCRztXJPNCmImc96npo4xxht/q+79a9jUePLFgRPcAlt9K
xQ644Rz2wnVFRd7KIpwNyIUbOgkkcumHS4IUxhHs5ymdYpayp2t6/fLqQCk0BQW1jrap05VREaFP
V5Xg6LZEUXO/y0ayzU87I9EmFXdqd5CW45DOyCMfUZcfNgiM7bKYCQoTEXTh/Wo2vtR1DkjXRgH0
ZWNmMKUKtZ1i+9SVwkGC0Dx5N0ysi0qLlWFLK57hhu5Xjrc08x8TJeuPFHXZUPZm3D39ooO0s2Sf
hcwzUO3r4w9qDkTTqa4EtwcjwKd876nHXynnZ+rYGjK6yrBsCl+kQ8Ff6l5+xal05+PL5IkTR9/2
KbKIU2VYjCBq8xbr/ltcyE+/c6NytsFaN8eajwCOB1mI1akW+SgNVTTKFtWo/BLnX7GOd1obbmFw
QOMv1VC/PuX+qQ1YQjJCXRop4HZrW68mxHO62aueVpLoaifvYzFMINQn2pQpapCXZSigXmUTPkGS
7V3KNr514dhToNFHmXgVZ+i+JUdo82tPWWJkOCwLUXmaLbX0KgaEZQ9ZhmD5qAuFCfBpSBTBhVRn
/yHc5B9V7h3jCigFfui+fga4TZwA41Gy4LaTIIizuoQ/yAc7CkHy4dlCNEhoMStMp8pmUmnD0jXn
FgiI+ShFUvXH05Pn6+bKiO5A/N58hHF8Te4gHu421EyBAY6WJW4gzTwLThkXrKG1uUUZVdGHHP9s
dsuao90/OwWL9Q6s0x95UQholLrR9JHMKEfgpQjUBPNJ1UbaUVBTs7U2sp446glK8fumu8926w3E
AblzaPvK0FN4eek1jVoVJjWBgO0MCL6E2M9l7RF3nsIXAg6RbZV+2VBhpuNrT8VoueoQDr0I1WIm
wL1iZnYX7D9DE0Gt7a8mxMGIxGq86HFIUClPQBnWq46eHH2SrzR4YkGh/bInQjUQA0aE9PgITbUl
cLjO2ziCdwe9hxapUMkBMAlTw6/7z5wiMv40n1mZ5wt0dkVgvHzXUwWJ2EaR397BlbBJ+8L0Mv1U
LJh/K4d3Qv37SiGYd1c8y2SAQ0pdc6QKwr+GLEW1neEeJGSnESWwL4tC5dT2S2d2ERlWD03Z3URF
PKITPVmIBd9ybWag8UQOJzJDJvXlOw0T8mfwnFwce6cv/uHRStecBGFZz8fVWtwzpxlReCgN6aXA
aKhWI4TNoeoF5HWhhjxT6+y8M+QQShFDeIHud4mDoY1pXGwSfuJyJO69hBGRuWKce8K3iXLNQADA
vIJ9fNw7+LIPuBDL4W6DuydxH8OKIh/0nrxH3JlCicJtXJs7NEmFEgPs/TB9eLG/RI8vZBPlFOvJ
hbtwLiJ9Ya8UDdb/QbCW8zbRF0VFJX4vUa1Q0Z/TM6hXfCSLkEiN9EKXmOGMYJTYAdPNRQiyWulA
RqLorC5zz5A5VnlTZrAZCdLHwIATvlfEmtHfTnO9OrDpPjMdpiCWYLrOZxKelj3uS+zcApWkeSs/
qw/UopaGTRHGKue/NkdOdziX99KFa60tfi5zMF7/ZEyiMML5PZZH7cVaJD3OfJz4qYBgCpGvVb3e
9MH/N0IY/N7hU2/i7xNdXa7OhBd0vFnMCoAC+Ofmx0bGKSF7GDEslSSOvFV3EOcdZPKcwYo/C7NR
wWxwzqpD4uqY9czVUu/ZPEnpF8qDDMIkPrel7HjDdoLapDzJ5gy51nUJu4vDfB5oUL7AQGsvlKsb
j70Ute4h/A/JqgBuB+dK+fmVnRrIHqW+b5/m6gXJbnTyGulqnXExTu/2w7UIc9puW+bL/DVyxHrS
Q2tyMKRyrtT6ZzjlrfNELsEdkARKbJ0RPOKmJiUN+hwTAbrwW9TuHGq74DO5wDjtybtIgXzGIisr
OJdw5MPYKcdC5fyR1tGf9Qpnj+u3zHFugvSo77acULcrHQHoC9/8yLyJqaVd7R7LEUzvZO1d0F4H
OL+GuMdO2QnwBYmYz+88lKT8KDbMUEvDn2UDHwQwlTPou/VQx1XDK4VJUqdWm3ugKarP3XNZOrfJ
+KcN3V5V33ttamRSLUqY5SwHEbNeMkYcoKx3csCkgInuV9UdLcIlcWoYvrRZsRr0tPuH75BCqLxp
EVgBZoYJRpOQexWBCYSbUKTeHD+6pYHHHBmx9ReDAxDUb+0enYdkujnHROXP5SFq7J9lu7vFelLX
IeUaVyrvrbadDQb4LYxyq9nN74BhF0loMsyUSiIHKTtf0wyWjlpr8QzKV2vhOEdsJ7Au3xWFUljN
YlKl7J+zDHPJW91j+xc9kG05w1pyWc8Msj8+31hfWFJCCNZA5JH2qM3p3C3w07OrgFFyd6uKUGgx
iMS2OabGmG3ne8gdUcnKEMvNA+uoeFspnQu+dEi1IaljNa1oYJRQnMt2dHOseODiA5cGg+4LKlKn
UDmBRdeTTxeyJqQRIGqZENVn/vhW8qxYMXbE7/j+DRR6NRPx5qgBYyj1KRW8/0wKwUoLeYiiZsxH
vi0kjr2CxXmQe7rv8rQNWuxnQvj10SHUiwDcY7WVELwbein6E3A8/JeuR44K4qTOf5XEgzkTs8AN
1vx0oyXX/1p4CaCaTdGJ1RQc1qAyZ9fnxXLzN2zKkhRbX341geZQY09p23NrewlU7ror5PRyc88L
g0XviRdiEtFdu8sellQ/dMvmTYCtbYlGTiWqEJchelAW9C/J7Y1hhfvOmFri9KUyUx1LZkYgHv6a
7CO+khvPm2UvMgzVbYkJsQrjgZUE5NRPuLcVQdehYvKLbAaTNzUB4t+a6E8rkIe9xkbQUXm8LsVO
0owE/86CgaroCCbH8KN+WLpjCeytf9Wj+V3MlVJFkvbgoHjB1VrIdiqtAeFFtaltO8pYtnlP6Jld
bwdEN0Rezv7d6zVdnwzvTdG+v9y9Jw5nUDdoREE8Zmvb8PdJMoYTd7Iq3qYHAq9YiTFOBl4cAnHx
24Lph31w6QbipdwiBqh+VIIHfBI78UGjq0ApZv2VkS2mNjo/hnlXQikxdHhuLGIYTmoxdT89Edw5
Wxcoc3UlwBe5FFi/YXsRxU/J47osS8qQ3AcLJEHqnUKZ3Ut5k8CYFtSTb4kbZ/Ab84L2ZnYYRKSn
cr44OVsykM5yCsRjAKfi8h948/jykEWk7C96bpUD7lJJgBQYh5t6ubmFqO7+1E1c762gvYHSnOhH
DbIlMfoxAIqh5EoPeYrDVAeyHSUnXSfVmoDdGQkoYTEwshOVSxJxeSe3Fal1YJMduhiWM9hjADtY
Yv0MtrRffZgghVtkqKVw4RQYjHZZzDFE1I1792JFBv9cSUgTj5DiGgRiH5Wdjf9Rphn50YINlwws
czhvksWGhX8LByqmOrPXbQF3nr7avI8SKyFCrZ5RWvPZT/fb20lRc6aM4AWDz7V1yV8K0rqngmc3
WSMWXRxwO+tYNToA8s/45Kg1wPQf/icmMlamPIR+yXgq36VKEz8r8+r+ZXXOeKaiGC9GmOQcepzC
e37KvhsBR4rS7pcg6g3OlIeeArCepxNzFkMygwVoI2fN0k/bcyPt/i5sUuuv2KlpC9EKKqt7Sb0v
5QXowxS1KoMSUVVH7eVcfsLa1ecXGL3/3NxhOvpwCLH27NyGMiRdHGMDJDk/QCuDpRT0gt1Oi08C
Dxp048QM7uDNDgtrW23kvafb7IOMm7z4tFhMzWkhXWsTzJtsHapm6k8A1SoICIMb+KIms01a89vW
1metc3FmB6WxWClBOq6iUFKomttNhiGzdd9RRG/Cm3pYmQyvgzifOjbuVL7hqzlJDhOG6lvY4K1H
11Vi23x76gLXmTY28vp1DQXPZ7E6QNFDnXaqz64xCVJk42DcUa1jP6UEvSOkp60Fh4kN2msGb27v
B2vqsGle655B6hPWWtCurkziSS5CTgn5SEWz+mXfOf2RPIKXkgDttnFoUYpU6P60gZfOPw+FjdSu
WTi9PrqIS6mbTgaQKp54TUY3LwpAE5ijSlSmslW14UoM07jgsmLORcNlCcqkkoZJK5fcCkzA52f2
F8lzNse+yElFh50fnfrgVd+I7HtapUbFQuqB/b/UDuWglIcqTo7Vv91fyZghT2G3+VAujCJjOvtk
dnRFpxF6jOuYVPllslf7KLcFgbPRTDTm4+b7M0PYPjFe65NSCgGKSLEqKBPpWUuMzGC7BzTJCs9U
GYqfp1avidS414Go2ky27J16QNKosEKRuVlUy2EdgRFS8mPOQ8hM4fnqYQ1QgXaxPKISIB+Q08NW
wlReTaLBHT6WOoVaAeijNFoAS5Tw7MX/879AuR9qHJlyndIiEDTbVAcBLRRupEOOgsgbyOw4mENv
CNBy9Fz1vtMzGojuRPjAnLnaAqRFeSCl/NaK1ovSdU3LC0j+2jhaBbnVfr5YonuTIBnzkenzLwo3
rXVdYT4bu4FmbR2ukW+V6uOCRRELCbw8BPEYrQgC9Yq+PdXlRjeVd4851gzCLr4KxfM87PglhXwo
T1Hcj1kyyZjkzngvWR0idGHvEG8E2Cp/C+03CPSOfXPceBZ/H8ZrhNGwBaSIoVHWG8x1d5MKtClO
FgzIjpxdWAMahoaHy8bRB3nfD6ifwLDu0ajdIguwHqShCmDOeviYwzsMxM8ErxVL0/bY+f4mh9hs
NyOsyA+e3Dcw6qGa/WjNgLXA2fF9cl/a7rEUTAN4FhS+yKQ1jN11Y48o2RBBsAj6p9u7HnKe8Oek
3/5v3zQNyNnG8ToTdmdzT1G/1pMjcIhDp9KpW0Np3ONKf+J4NAfOZoygry6FCYOM72SoLXozyUT/
4SuTsSNkRYzpX3gDUDx0PBIUCMziUjp2OkD9kZkB2UVuSp+lD8cmxlixO6p/iFxhYVyGgeI57DdH
fyKwHKdPJxyIxYJcmQFlCGZnlAaKmErAI0BvgvoSTzQ1YzrG4RfybsIfE1jjd3D/KYcAz6WemiOG
pb87/xC7ThSVDtZwC6CQv7FmDNxKK7st6oAEUsCTOi8CCqGIvqyRfWBXE1gHJeJ78NlFwYY4xitb
X9Hb8x3SQIgAwW87xNg+cLSdtkjAl7B/5B2Vm0PP0UrsXCTb/oKVsTrYbnIWGEARD8LxjBITjHph
g8ZdsomLLcO9r/2M8bgEcAtsHoy+WrstFpoOAeM5wwz0jto7eRwcbLSzsNLzYLYtPjtsRZP6EwR3
pzd2dh6LTg4NyUN5ViqxNcZgwUV5CSDQGUyUSfUkcxk6lSxSEf4dsrpnvLq/v5x+PtsetqREt/6a
cT9bgaG1nBL4bp1c/YduOtTRtgjOSBtp5doH+2SH19X3NRqugY8DWp9U5lhq1BqswhewxMOwrnw+
09jLu2gX5vOp2smZV15t7Oa+SyRSchIAnRFe0CCpPMICvAzTTc9jnaoeZ8+GeOF/YorfrxjlhZuG
eVGUjWFEQbTrEAOso0Bx0L7X6CzRVxaD30FJuXLve3FmL6kJuwINxUTpS+3pV9XRmUWAapz+mqR7
Cc4qhn7ZACdjpcPCCmTFdl0gqiUHJU2t3hCPT47Bjx4kf50Xwnp86uNZLTwtkhRU5eEFHFJJ6IHv
+bQscl518fYvbcDgrL0NMF/SlTgb7Q5A/z2yvAX7Tvb1tqgWYI3EDN8rDzDmZjiCDZtMKI3e3r5v
syPADKZyOtvUwukREkUEWCR1x8pKc0zK4Y2JolgjHVPOw5qBPe3PzJFN3UuFTT0WWBnE5+a5m6Qo
gcRS0OqFt4sH9ZZMAiQez0J7O4W/2rsyGKnmDbTnTrh5ClJEKSUand28lOkjO5FP0xTyxQwJguXQ
dK9Ei1H7BCgxtD3U77khYBOg3mmPbF3YCTdxpvLVnX4xbz5pFUvsBNZuuGg9VV2BWXrpTHUvyvSs
kh8nFfXPkb5PsZjjtwAtDfUsKebqR7CW8TB0ONuqfV1wLeqXjRcr+P7yUlDIV2rmUB8EyEkQSMmY
ovPZ1d7eptnMR+Q2wQSFMRmqQaCcW+ACv2g21qWTB2DcsSNU1cvnohPwWAj0jyDcB5Z8bMg7225E
eJGr57b2J1xe3ICjtizVLEHK4oqcKXU/WZ5gcWyf9P8KhvehplSVX1Y/C6pSrn1urvFo7rh9QzIh
lr4nQPOmLf9GvTyGT/Teef9gGejf3D8K2AVebRH5f/4eykR1/DiP5Fj521psS/X69YbfA5KrGPNF
2fSRbu6A+3Se6uIj0rAU5wHOEQ3zkrHYd62ly+cXPWNTJ804XIR1GshNPmsFcNseX0rzBRO63obY
2YoBUhuUtdK8VbMT/wuo1qOZd9slN0uKv06GtkkpVQvHvUyjwi8MyAEgh0MTCvpKP3E+0+SbVSAj
5aZsiGdBhp47Ya+5dlA7PMiJI/ABW1O35wWS2DyPdH7un5dvy0rNuoJ3dIebLhMALVioxlruIobI
hSJvEsMd2pNDNIMa4ZuNEo+BlOb/zONG87PIhYaG1jyHqNeyXCRAqiydo02T3uEAlUnjRzJJ+14o
189rjDw04L22cXVfcDI5tzBbSCaJZapC+Olil6wxPlP6Gd3h/yMYAxUTPnMNgbF05c8ISIzhgQYT
3K8IixeACw0nqTw1zo27dKe/ZuSjHBVGWD8bjlwHBVWD6kiAuuFsVNZjmQoFyFjdiU9ltu/dtyiM
NcDNo08eM9z5yKr+g1UpWQwazswPcznLFePZtRzPL9cmvvHZxoXyeFR2DVyLfQRZOzwX+zhyBWqA
jg09pay1/x0906n3P/Lh5Upm2MUJZ2vfOTEIXUtPB2cGI2qgV/nNNAL34J8UOmgZOt3KMI9re1ri
RBFbI4D0ehGXVxpjS1sLg3a3LY2LU+920OY2SGfHur3mDYMNrZau/X+fOy8pgas0R1ruUSUa3lXg
BS4MyPVeT6ysWDgcxDGFK7U5xzrHu/UvDt0KmuerGh8luHnXlAElxEkHeF0KUM4gE0ARUmykz3fs
hqmzaC8LfdFdpV2ga5eO/S5vC6vHOLPH3+CjAuTL5ub7Ccoy9xsH8dtH6A/bO8oZwWh1y9b/UCt5
jtNBy+IE9OnWDdHJ4RX9uQhLmHH82SKuBlcBhALDf3Fo0nhAQNRZKwLjwvnfZFl0KWZAgydKyNVc
SFc5Lo86y3f9S4SlINRpfhUXsRIPvTydwUKbQxvjKoeYEK/pBBBYi4Q1siz4/oh39trCVJUmLT1o
eN4UBqcgC2mcvpgBIBG3VdK4e8+2lHRTDBkx8oDQZigdyfcFV4NCqN8rCsNtE8+41LSBAFadfhjY
zdbDV2e34TjIZzzVz1ZEAyRFSnakLaL9GxwQDGaTOY/FFOHf6kgr/o0nbiTXa+dKMhZR1mbVNvty
yUUx/rpoaHmVg4u+gv9JgTr4m+cwCfWrlVvJKHkVH2RXc2bcsX5VlSi2VA6gwmR08TmLE5BIWGJi
qaQToaSbQCc1rXwVbKVampK3bfFcU77Q6AM+pbFDJd52/Di34N+15QuR8qbu9Pw64wl6MadCvPbl
JPCz6SXeI504GY/6BlldabA+hkVTJkQqlVFRwE+aCykdnLwQuqOWNF3uZuJUC7JAHpgPWhhbHSSw
69ZPNFdkyC+4gGptgOjxJaGS/FmM7SQkfLxtw7vhkrc/Rm5MTQ3Uyx9cqxsbKLnpNlbhANiqaojl
JYPzRnMWWtwNoAhJgIKUgMuyOO685a1AZcnOgAaExuHGuf4I5a46C4dpw1kp1oe96sN3ofJcnTB1
DMnefDtDpDnwXAhASW47MkptRhzMkwByNs18nz8cm8r+vdeq5U52EmtbrI7hZYZGkQFk+h+fBnWV
sH0OgU7DPZRXjoQtqfZhBomnpBkA2qjTJutAklGHErJOOLVylLZNR33AbRGeFR6Dp8BvAiTI16e1
GlButhQkPII4+b0XBkD36aWEZV8Ec0eyU+35G4DMJtqB1nvlcoyP2EnWCMT1Z/2iEJmhWlqOvjup
V3ISCTeZkwcfP2xrcMKMlYd7+vZDMz5o8xY15dcc9LZaDJJtmXd+PyW8KymA9V0AuB08sSTgyq4N
jK3a7HLdCDKVi13LD5+4AVblhR2NuZjpxHy0FCXSqkWJwoldZRUrwjAaXtG+6tXQXS/MHE51UVO9
BgpraoBwrA4P9t0vqiGyGBnS5sQ7YLpftfQxLFHjrHb/wF03micAPvgztHIoG9W7bNDQyixB1Jw1
yk8a4jvF57JfREuE0oEczd0KixH6vXetCpW9JxD4MbyvPY4f9/X6Sbe/+JzniX+iWx+2NNpBGiE2
U1QZWN0SslMHaEg4R9jTlwfc4d/y2XEZKT/Qfaz17cElj2lVZaKzfRS+7NjbZAQNZ5261+++OjKc
mIIBhRgc3/iQVk1hGuxRllytKATikbFUZcvRBy6fiSsIdzQdrFPPfeUTSCwdiOrbTtQcr7tNmR4T
g+ZMVESI7W69unwMdelwrxi15wFNicv1f4BI1wwnwtecunr6xLk46pSVmDCIP84kEPKn6/jDa1nY
9gu3wn/yzix8FRXCoGfNEdBmSgJ6/6tHf5qXlcgIpiy73oTCRH5YnCNgrJiv3eNW8eE0DCy6WhR3
okSwmaohRZ547atqgQF2Mfi8j5n/mLPB3ZAmhlO9bqi1eoe2Qqm/EVpYmKp+8JSC3LM9qs+rR1w3
U+4gCEiSlMF3brBE+yp6p5BJuimpejUlGDnmHuWT9CadibLZxOezyo6MwCblGcHb/cWiNDescgir
IOFDIxPSloTvYIY/8liOPXBH+gc7i5ssa0y6VTlVfTAobDjvXYs5zGQdoXE2evVd8vpVyAg3Ahbt
pHkdx8O8lyVUFpozaAet6C9zAeAEEw03E6Me7SBcv2vhhnIgfQVQqKPJTAXMjRzm1gpJAutplEZ6
8EqYzfOpU4hR+6K+2UR58wx6KLqSaAuHHqUtLlpvW2iHeC12GI6fGb3YtvabFWjfLMvLRkAoy/bb
2LUb3QFsG2t25fbDpjlmxot6AcYzKB5mRs9rkCidg+qYQMWZftvQIVc8ovDd+3tuQsQGnbLpL8TJ
xR9+LRhS8j3ipscJZ5EH5Kd/KGwmSoQI0aCShn20e/jDF3tU7A9Nokfag7z5ZiFSV28kONe4ykJa
LfacajjiozVsxDWPI0tTvalO3veNqEsFvUqDObBpx4dN7jcfYrhaqajs9+JxujctLMKIy/QvJniC
nqL/dw5JyPJMc2l/RdmVfNCNGlpCnQetS4MAPd/VOCZSmTE5Ms4wXgoNiZUeLxZQaf7XS4VANWJO
kHY/37Xq4qJCXuyUWf+NflkQ/2+LHo/4r4OvY6KxdFFVPdZ2bkwPjVuwsOggOYFbVXWh8FvlV6sh
qsL2Nq2fokH/rDisoguOQGsXl5upzrtnnTVwB18GLyFvE3zxHeQHbbER7Sn1dCeNVUPpEVUCkbHw
FdpOmk/CkKrJtDHmlXG5f8a0Mid5fv543308zYUINekNP1HPsjRiJX0YsJQES/xjCXUrHmj1ogM1
VCuigP85RiEdVHabq5+kxFteC/ZMasfGTHqyoWdtOXLfmUikV1bH4jdGy+q+qaGqOv/tWPm2eR0+
3r3fZqQlPX04cDN6ox6htoiC444tz/NRtDBhpowj+1ykpEHHsTm/8ScFNds8V5oYhEZmC8RJKFdK
yS7lk5v0sVcKX0i6sgyO3a11oORDshC7ajxFJGTYak6Z2nHZNo3LuN88zzChp7df0AOdJUuwMLOD
PxS5PAIRoSN/QL0x/OvGOkNgGOtaNXE5VCESP5NopcBT9HG+C1Pm407YO2Vdc/3GPMttQ3ZGCxvk
1CHB8kNjaQiqnkcd5JAjt+gwA0iKNA99wWtIezf0CKS3IEYZjJa1SJM9cgWL+uTCxqE0LnD4FbeX
5xSja3wixMIBATk+9wuDtkZ/Mc7W8iTewYn7VUvanC4iel0QbGGiFiO+7SqoRKS9lPXru4SxmV3g
LYx9SzA4YmYBjFgiBiZUlGDn7VORDLFySZk+OkooTmkaUnzRxiD4kVz7iM+c6UsBjCEE9hhIaGNZ
VUetWLZgwYOXLHoMHlOAFXSJu66/jWix3fzUv3CcYx3eLJHrXlg8sxBkvGoK5t2ePoA3KIQMSP+1
9RbDgWvqJxBfe0VapGFIGy1S1QNLmvfa7bMPJW1yg6IQo+k7yQvoJqmFmbgbhN3cjT64WufzgRAe
ahBnyjJFrsKPT2EaLt7+nk1gfrcPab84ZytivSDjbWhOJL2dD75ocgNXuu8dvoe8vtHAO84xblu4
xsc6OoESlPRGcSEIz/KjMUdrtMvk1B7BZCPhD1mYYJuBbmdr1o00kx2jWly1AHkfLMrH/AG+DKYW
u457RbkdqopVAuuLGtvoQIDlm4ydBD/AuJgGh44OCAYaYYRkPZk9HwfCHHsXxFyqL8CgD9Isw+ZB
a4eD53rODBiiwRfz5gidhANQN4vqIKMK1hul0pln42drKNWGCpKvhQuoGEKuoWID8SCu4DNK+s4s
edjU/s3VR7PRztH203eve/e6Uvmj6EHICjMBltBvfeuqpPJOCjyFsnEcu0PFLBZW+GEdW6xvlBjQ
dZn/MGJ0Acg5O5lA/KaRFde/+uYOcHiQn93MNKuy4qeiQ4nnzt77Gz07unlMuk2DrpXnKITgHeIb
NyxTfbxrVJPY5S1K4Z6/y4nzVZ5QSj1yDQxJkt3kxKL23+mqwm4pzjs3a10fJ8yB/30LfOLN9XoG
i7nN18kEqc8ukdHgwwb0iZ1jI41tBjQl0/NpSrrv46gO2SdkbTBWDY6mUtyEIH7K9BqC4YJaPpzk
gIj41KGOqYJ+BpfAwUBhhHhWjbybAQeqL4bn+CxEsIU39qBYHk/r5V1C9Z0wQSYmROSgq/8bQLGl
dgymOxu95DN74UGz+rcQNVmflyYkykZh/s1fbFqlpTYK+qdtZxjxU+T1nf/oGOP1C6NJbOJeuG8B
CJRGjxLDMIFJx8MAZYiB8hvZ5Owv3Ay5GfsvphQD5/2p1H/6ds7aVONrWFZnsvtx+7Ed+PqPAdui
23HPIerPS1XIZizZtTf1msQhNT0Pivr1881h6QtuqALwoRg7IDqWnlgGRpAX+pCTRCEPfGnR5fKV
QX9z1uCcMoR7edrjYXHR8aglXD0wzTYPXXY8Q5NBksuGpWrTHJ9RKm50pHqlRt8ghC0Oh3XTtu2Y
IY2zqqmebbcVo/q7vUOm54xIA9YPVVDFrdKSzlpZDn+GdiBqL3mAg/6Sb5Gd50vAHWsMAbhjesi0
MBgxCv2zg917f58EFxPuupZaxiP4UuWQv0e36F2XWK1EtxUkjIMUGj5I/nsmKnR2kNN2kxxFE0cy
x+sFZdZUxZ95cGpRG5haJXYLvABJtTAEnUT+yZZB+eXxRIAfk5arpGYVWnqxB+WB1la7qvSzmFhk
U1NuI2z9vgX5PRHstZLgmy2Ikhm2FBEOlRk7bwJXIhOPWy4usrOmxT1P/6pKw34IldUF+3L4qd0H
BZtcczYP0uF+WhhTocRwyY/VlDNuRgV6sneXIlaCv6RhMNZW8vBxjjFIS0pJFQlwqhnYVf8o0x6J
Wwf2sRRS96JPRV91zg10uJdU9rbmwKpOVHwznrfyFVdF+RqjRh5z9KsJHU7WQuIEjpeFXSD3p+lD
su912e5ECx8/u6aFw4q6NF/TjmUknzeKhUqcwr423E4AKmWKribgQbEp0KUKFYr+veDtE1sWE9y0
PhwGkvme7tCR+wELDx4wl+I+YSZvK82NeqjjZ7QELf5WkHOP4AOJrKzTECVzDVbiLZOLlDxgMAbZ
vYAFeIpFGW3sIIDPmjKljBj52M9bVFbi6u8zlw6OR6Yy4bzn7+mHYg5orn5lpClt9TfHxasEKnG2
1cUNw2fAGqYTqtT3G0hrIlNRSVG1ffhwnOm5Ypo0Ujc1Bf+4VbJrgjiWlgmJk1L8RdalUslK+Mr6
6bpmMczCb6V1XA6gDLlQ6I8+nDt2PU0g0IruNNfxtFQVvQD9qzGQxbpG7oUiOxXmtLdYVkn3LiWH
zJ/RM07WfK6KTS57NsydwecXnrmf35JfxrtKoC3K+y4JfJ2d1ryhmwn/pAQMB+aM8wKKhyVpBY8d
f9LITGeTRRhB89/eL/SesAh+cYYHbAGp3f9H4kdx1qzGBclxQD88XOZi02Mckoyhq3I4i2/6T286
xv7CM4oPD9ke1xM8sNdDf4TBpmIwcruPb8dH5XHDZPlQ08zV0YFczYB7MhhO21TCtuCDPEeaXlOR
UMiXbG+z6L+T++NjBoH2MSibRz4YJIoOYsPthtY52sl1gz3jSTd1Rm7ZFgdyWRtGfot5BpzBjdnW
1NUdMkR0hbeY5MsjUVkdVrQ1ZZqc2gY5w65B9veL1SShWtuW6P28IjuNcN/stV4wFgzQGG7IrQe6
VwjU6sWSExMoFqf4IH0Wn0fJlRHTbQseqibVMRzg4LYJ9Zg4DdaEqr/PfISEVReEmiwLAg3LduKp
ruKx/0vPkblVsmuoCCG54NeNc8hBYM7NkOR+8rrF9w0wTkM58V8ppqUO5EVBlmMgs5Qig5balwZ8
zi0WwQvFSif/VAsYGbI/+3iAaYSiPmZ+N2sGs4jVgOmZ/na9JzKK+5v/9s7mbmUUdq6hnKvNnDDU
z6OeKcCg+ktIT5fHq/mnO3q+qHQVgz+i0o2CLbTMXlCAIK0Lv1cF3fPxeQY8Soy+bScK5vGuULWA
/Af/cvzitQptPHfnUygWUu5IPz9YtjDCwFawuzI26BJBRXpncVZkJiSwPJnbzx1z6pWdTsl0Tjv8
HhWUU+2WiMUh7vb+lxUzegkVGErcFlkm3yJdyNCWiwPUsENjVF1ipPn5/yISHK1RQRCJiG8K/dd0
Pv+Sjze1zfpAoEjTUND86lw3JVYa/fjSJp2+oK3VYcStswNT8sQqW6nNoVGY/rBhbMPFSNmeSnQy
31pNvv4hvkolOqtLNxBvYzeLdUZE4BPMz5r0fakBsugO94UQdWbdPo65DjXOBo8uqYK6/DPOqUdr
6S0Wotqur7fbtLiShXZGjI6zrnLLIIarCjnyzrPcS95gHswGg273VUvKW4+kcNoPutZ1D1zbUO6O
HTEyyMmEyYYPI96V15JRDxUO/SubfiqBdBu7OXzQkpQY5/65cXJsn3dPfobhoerKIdfWURtdJkuC
gEOQ2HOnA6m7TwAdVz3Q8MF2dLQrBKjgxSYVnWguD2ZVyaBwB/h1euMQpZCl4haW/Lqgs6Gy/Do2
GU3tk75I7HtcpA/qa8gzC7/lGkHNKcMRpWSZZXUmoctAEOM8zfsTSSNwANVQlhykmBUzQIcJsYY2
l18TWaeSttEfqB+YRHT83gNaoNg9JvIh80ozyIGBVjrlVZacnCwjTzuqgv2eqBggjX9y76FXwvDk
IyhYutTNVbnM7C2AAXl7oxnJArh81EcJD6YNPnXCpRD0b4skICmotTBc0/fAuXCJTwvReLNq5gYJ
v3msUFQnmjGfN5tH78S+oviLvC6OL3bQKPOMjfXjOTk5rMUVC/gBgjIwqAEKkkIsqzzIo1ouRnf8
E1qg3F4bhbrspuMSHYDpeSTy9lfOdDh8t3k1xhq8nZyO8VPJZPQGwjS0ErXf4LnGD3UBIAZTjcGJ
qj3PUihFuV2o5ooYEvPeMwPWSIWWBD45k0ed0Zs/n7mAy4rFcUVZMx2zrFe3eLad65b7D+fNqvus
dXZWTb+AzUaf21erJZkACJ6daGvfmGyzQCButRDFPX6cPfZ6mpXhl4oDFEBDcoclq2W6SWbA0Adg
g/bOuA3EmrFaRlHP8I/g8Hkb7/Z8aFdr2+ExFFoXWVMKXLtrRFARa2Q8+pEdew815Ya/EW2rleM4
YEXngiVMtrt7Gciu84XeWLJ0JOPZWtf5PnlWRH6aAhg9atsiYRuUSS7XJbdc8RtZDxdPSHyGY0b4
qsoGLIijQE7d1ht5ijnL1KfqguX3vLb+4xDw+6AypWdMXRCgEIDcYwxAeFRw1SXK27SHZlhMmqSd
4EEKEbyfE14rOFLKqYNF9CThFkd6Fj0pm9rYCUBS+3tUaLxwbZgNvRUiKVo9mKsYTGiVyLaAP5Uv
Q5r+JQyXpXJtv+CHOkLExXYL2HzkvBK6AdbEBDHRjwGX7jxjcagP5t/DDNRyJ1rfAfGoELegTcQ1
oA32J3aTmn37A1/J5CD0ZLemGLpOqPAUYRBpt6qj3Ji4ohsVwQ8w4TBnExw5bMFzamF4//TqwGY5
uu82QyhyDFAwmSfR+LkaDVIFNOQYqODdjG5AQH5hX29nZzlxSGjN2nQNvRI1bKRQVa2cKFAdLeA/
T71PHqYJ7Hs4M6DndfxONNDYF4+I4Oi/k9uNV7bNVna1s21psNXZDMbNxFI2dHmXRNGzrH258kUJ
qDoZGmOuBK3Hq0ybM0TrIGCpbAmaskN4CI5rHG1ZL6tjiKjUADtVCKSgn7iH1yiiCWH5Q+gpAQJv
RjcOyWYX+m2KMobiHeVt1jptx0/85kbUhggHHHB9CXjfVFVRACSw0w/K355EKlSCn5174K46rz0c
IiBNlqBH433B+fin7WeRdgyBGQWaOUtmhNWT80MJZX0OhSc+khI800OUJSILDNP7HAoIR3CLkqhu
yN2Sy5wIObdRLu2VgoVAbmvy4ChY6PoWuxegNR0T99ds6wWOHfXpHArbr/fznPqn53lxU7DYCWw/
9+Xw+fDere08p0g1yzqiRRBqsckVy8Ei9tWXW7tLJF4TVaRrCAVHtovIL0X97c25vbUZgHpLxQPg
qPYrJfBY58cheQB91OMrOPABSkIw20SMKo98RkSYW8ircVn7cT+Uff/nnrHBS/K15sT3FxrHtEJx
do3U9WRAq6CcNAPW7yRs00Ub4B8vQfDjoA446WScBorgDM8NsN3EbPCxjTrRiO/QuS+4FLhHP5WI
HrJJJ+kYKL7L7gD62TwfCVaSUXZD9F3qF9Vhof1kXshbRuD59Ck2bh7aIXvILz06hA+JsQvTZQUy
bsZ6aj7JtHEdfDjsoXT16udZwH2BWOQUZcUNtv3ITLQJgqPk5mlEH2IEsk0rI/nVB8FvXfzr9K4B
JkLxsBpfI39EwXRTQMWXxz6loamUV+vakP3xMA0qxfOEylwigR5N/6RBaEmnB3FpwZMeYsva3aWs
qtuWAibq8aGwJ9Td/5yMAKfaeQKFj40QZI2MZB9UdFsPsqzgpo8hgsn5VLdpGGXY5AI3wLPrSX2I
2R7x6BWM3AHoQgDOhbsj+N20tQq2GkHtKf00h/itmKP4IImGNI8JCBYbUJ5B6cffP63i8Kvfso02
qALd//VbqNxcGvTEQywX8DCIbxFKTJA3TPPoc7SFVELSEnX/z2p3KHqbVMsjyZCtqgDN/BAj9laM
MltB5v2av/c5hVdSHScQmB9BlqacmFX0BAi3xkBEgpT2kfYifSnhcfSgc+N1v4I4tNb0Nf+acFuz
IAOPVD2tXPj64Ju7o+u0ZZN1ZF04g0KzV+/JorIT4+Fk1Ci4LhURl8cSEUDzesJEhraJKWrb5sAV
GosQyFiL/5z+z8NMCdqn8zDGriEPKUtoGg1xLllKfspUYwvd6sfKObY1UcBN6p7YrQh1Ge8uoVlH
+j3Ky2l4Egn1giln/z9PF7HiNyGqY3BslUxWITav3EEcx1wQ3Wr7WIlMuj0E6RuvNA+ZoBSGdWT5
LBGH8tuZ7SuPyyCGysYG43o51vtwmVaDjkD7x9vBmsM8u4COGI6NU1a+dKCOnsR7TfLVw1T+vUao
YRVd3lHCY+oBiX8K1aHti2fnaYhNrWU7/bezAzf38gbalbR5S6YKN0w6wc0Rakgp+zCNwxvbYE7j
HQ48YKpuUjglj/r8m4q3jVSQhB94Bs53h82EHKPdUPpFOtqhyw4l2D/h8/ZtQJRyNzE+cDMKoBX+
KbFsNWm72tlzpIg1QRPxRK8BBAs1Y1GRnDM8FQo9FTdp1g4ZfHQPauyLu+q3owyBVJfAG8bNp+nK
v634tT2N8QcNosPQskuHwWPJIVHe04ZxYrp/sBzWX83dYwS5XJugo1R5DTPBbf5lbsBM4qiV3uXi
AscF0hK71yyACb2vl3md+3Pe2WH0kiN7DS2kjTiDBHdZ+xZ4JPJBydk1ovCQg9LCgQkD/bZRSGHb
pk0gwlmgMm98SS9XHDTT6BGr+j8tx0EN91MwdmR8QH3qlN0GHPSP+Jr3gU4DE2t9DaesUguqooVC
jLbhntaabkE6XoLpbL+Un+YfdzJBzjuJJIXkfDO+1nYRK1+28SEg3Y5IoMmqRdiXlVJbxqcTGrj1
aMFFJ5/tos1kbf7yySFOEMcMdH2vfTqYAQ+/Y0UairEdHb9Q1a1W/KMz59cswjXfT1dn9nSTSv5G
77m/pcpSd+Wcfxa/v3OYANpM3EEc9vJxkcpXSp1RCLQ6z/o+jipGP8t0hoM70MH9PYxaUEQi2CzG
zW/B7uKJOXmpPxCVK5EXI/QvuEP3UQenkHwuGHfGIlMuft5wj7QR78mFgn1w1Rj3/diEDrJ68M6q
icK2KnDRy4lML76Wy1dLr7d5Q0YeuWzf7jNkiesQCMEbeOuUMc5ZC9llUpoR1e1/vKPDVAGDnObq
5lTrUteGmdhQSVgmbCrcCz2x0Wh6eRD6AdI4ZtGD9BdPa/w6GKUV6awVbDjmihgdyFLxlovS5mqU
UcaH8DF3GtRNW4EOY6p3xMsridzpCJuyP2v4304pNVB7MRETH6BqlB7evSYm9r07U+IeEkJAuJt8
xZy1Y8KyzlOBoOE9kr1yPtjNIg8mHYULoYUb+huRefOsbvb3GMfS0XPP4KtOs3LHXqYpbid0SxAR
/PlNwhBp0o6AoGinRf3tFAb/X2SZA5YqsPd+vgeWoAlTuo29mNXIWGzC9rEceOerxykAM1XA8jmL
WWn4sh8ljLhpkzFmlA0f/IHcSzop2i+790voPxTLBEswMqxl4aDTMC43Lp7wN51H4ZnidFy/FE/U
zkkZVoECVufXWfOwNQNtrWq1wOCV5SoHAzA5erLZfxTWn6K5dW6R3riOlGQ5XvCbQIeOG5bPSWuH
Cn4jfA6lMwxNvFI15P/P+hCkeuEhvVUvNtULokwecdVeNCNCAZsAqfHL3TTx4t599qZ2dyWHDJk9
vO2ieuIOvKif8tElj/y676AfHoKEu/Q81t+RwSPqsZEPcAZUmwrFywwKiT7j8iKVSeAG0CuCG7/Q
9X8uFH3kdbh/eZKhbVCaP6gzLi/h+ZQdbeoQT9E9g61UBNEQ7goppgftobMr22XXWav7QquqvoNA
doaVENO7vb/RC9/NxvHbNXErukauuv8/hh+YRJXbqURimx5Q3EX/lVjdP83mgjXElgmmvPm6/DqP
3eyOeA5q3B6hw5g0zPAo38p8xSIfenMP2Xz0b0Vfb2SovrtGHr15m3Q+TrQlw4zcx1IXE8bw9E/U
mddKjDumTRAC+khVbuN5/tyylx0xeKIFpIwilorsRyxxBMXWMzPARLGNmUkZETPr+SFpYXswkSzR
+OJGPp3iRGupn9njkDVI9J14S7YiZ+Q36AAkcD1QZ6PXVlW7HAYYqt6PXOcctGoASPxsGgG653ni
n54nnYyHS/QNAv8ENqn7FTZ2dmMxXc6zAQfUU+P0R5W7pPTy3OASYcn3YyKAXUeuMCB3MNEiCRNu
QDcBOn1MVfqenKZ9iEfPJHQHEtSUVqGCc/JWitsbgRVi0yt9Mh5euxJiGGKKZHRXkpV3Lz1RVnJI
xL3KH3O7FkdD3nVwmsAtfQ2h+fl2QiSAnxaHS04/SAAMAMQkAFWM6phQnAOH3qmxnmyronYDJz2F
bJQRcO5COOXveE/15wF/zVfek7Q0a36xIpk/Z9QIsnIKrjRz6jHANNO/GzvCj1/oX61Znv0jADF1
7TEoCbC+g2byjNSZhsC0+r3nBBGdt1H5/Lo3NQgRGaVGYRpN0TLbRnvZDLfbGYwApRiwHjTxl+d2
2dM9bZaAzxrKe02ZBQeh5olpbC6mJxzSdNumDbqSbyQFTXQxINZgRMSVnM0SwxfzXLq6z9iTatKS
ELkWTvpFBnBiDyIQExjMX/RnC7jvll2B6U4MajhD/5b5aOqHejJNg5hVcEKxtOnzrgFsBQ2F9reg
X84JyHGJ6V58O3xRUd42ghtWmqBrow2Gu4KDuP0gS/VBspEnlXjTlUkL2kUSr6Fqo6cJnVdAM3mv
0KM0Dy+SXSKsUXf8Dv7o4K6X+C9VtwnzCKHfdeq9LbC7/Fs41CPlE0zLl1BYi75pIWOSBH5gwRUu
tgKb825SBCwb+IEtohDSui17TJht8EFYRaX9B7PMTkQBz75fNaNxJrRe4CFeDJu4Mox0iLAbf2vB
kamDbTuow0e4sGdIgrWlgf5FbmZpfu7IoNDbnTaQSg9+w+GZrsq6RS97uNAq6QylL3s9g6yKtu7V
QgBZvS7SWTPwm9UCyOH6tO5iadKsyh649oFb/LkbkPA54N3uQ9qfd2AI3eeV06Q/klfz/FKJTJ8k
QpfjzwZvo2Rsw7djfauX2oVjTiCLMu6CMdBsMzhsBJ11qCvk9D4lGp1ERoQ/pxHU7mGxEGfpkPbr
3Gic0P07EBehhILhb1I9sUdXSsWtm9bLHzRTGjT6pj7fBUQzH/ttZESQmSU95uaf38Gb1g/BTis4
ApKJ5fiAo0t6HuiiNfxXImwASGEDDZiqb1wBuw+TfVwqTcQ7Te0xtZ3Y5spCHE+cCqtIoTRkGv0g
aYTivwPBuVqt9BrNpnc1RlRrlAflA/Q1cZbIMzRKL7hLH3nmNuqX6HVj/ODqN2LnvXcXf5yB53oE
IGRqCGD/O6GZjJpUFf2nDdcUixN4BMbdS+Hfnta4E4itpsZ8Dzt16dvogpfUjZip9aJFNmdW5znQ
EoF+xF3pjkAZMXeTzZte2dLi5ySnPS8hDfXawREV8EHamtQ1uBbuLGj9yuCCvQMLMU1hOCHS5opf
lRVfAlAZZl0qsj0+TaL/7Jo0AX7CjgaOzjtdCDBH2AeSaTiZPgq/DZQO2lQ8cf3s9KgR/f0IPj/o
I3X5nisN70eCX987r/0w02PKVolL66XWTGyN/BYxtShZi/5w3/fBJ+GiA+VIxQYLtLn+CkVL+THC
SZK6ZgzrAECGOU/wFdlPpw6hNXdRv/g/Ujf8JZ+iJkyKuXiQuSIxtRwik4WPCKdCAQPgHQLwekRH
2PdmTh4Xeg6BIFymnCXSl7Mzh61wJ5Jc/UxwyI04r1Ox3ENtqFomyikRgTYPYXVtydmRUPrl51+E
e+5pSRnBdCKchwaF7tBMSlKVJKbIkz5EA6PSVLSF89AJs4Po4OOUaJREWBN/JGCS1EZPujivuQDk
UYr8Lp95E+n7qZkS5v5+WYqXAThYx5XeBO88DkHI4b7TjRkOhK8nJt5hAU9hxsUMPVNa1bvUGGJG
U49G1KmW277n15wwqQM31tegKHSkPENF8B1q68qGgIiMbETHAn0oHXJ4oFk+3pJ7Z9Y69GO8k2mX
Ac5AEov/bpSJ96cRUtxXovBjESdCCF1/OhT1uSiXyFtajg6i5Q5L+VcM5vSd8rmuVa9omnyVksi0
6xUlfI6KGLzi6OKr+UQwbJQkjotPKn+GLXRss8D6CdTUZ3Ysj471FxM0n0fL4XqK8sOpXZmHhTO2
Q5goJYMSGnwknTLzh0EKSiBXHiQOrTXn1ojVyahHXj2hx76mr99QHhI7af72e9Wu/XXgIZnIWFon
Ouw7t0L7PYiGVcgGd5HpPatBSQUDN7+9vf5zuBicYdZZFDljqaXh05eDzAzrNj0lSDLkA9FhmVRG
LVZtoLo7Z3kiCv6gBp08ZKxluqo5FrALOEg8zui/gUMUDjlNzQYune2MMchxgd64X9YN6skdsBvr
fE87eop5vR1fPlUAmIS0zn4pbs7/I3qQxBVejeZ3eGCb5l7Io0vIPDYIeDKAeN3kmnjVwbr6wEJz
2zQxLbPnPyUDZgfCC4R1KGbQT9likuQ3sMdc8LVy9MC/ri+rWaDP4/G1OjgBDniyUUDI/Re0S5yY
9JXYPyC+RchVj7vjX6/oAk+ecQBTYUD5k+e9+6QQ+8G0osBJHd8QHprlFeocbTjlMCLi+gfsv4b8
dbsNUoLUq2qpfM0P7CUOTwRdx2bc3y1uAXyR0IS83suAIvTsy4qj6+d0EftMoCjp4SdoaDuNNxL3
FLfs6Ue1IBwSMilFXUjMgeJzlW0mrj9sz8Cuc5qG53fGi3yo+7YS8WuLkvcY+5ZfeNfvsKBY80yK
eIS1qDGLXrfysJQ0wo3G4nLO3/Lqy4guFATfEccgZHwxBWGEybjPEmKY85Iw7P1d2bN2WJb3rOhN
2UhHbjUOkiSSBjYhOBpVWWeyJcfajhO6rVzYgyKanPhSz4k0Bt6ffMUH2GGA4s8tz+GRyKFcRF+W
TKMpp7AbBh0CZvZEfvbisc0LWHsPOJvgG2ZNTkh6RnEMT3y3n0dZUC6jGo2PWUNFX02xU9IFogJu
CpVAzomCmJATuDEAGKBruHQ1dxwaHJsYYXzGwB3KzGR6PPYmK9xa7txU84TFBoVsHiBn6eVLj90F
lRHUMC0fUUBfXqsxDtW92NCG1qGARiWL1DYhBubopK660EFG9EQI+cC2OUO4C+NgyiBYIVDXl/ep
Z1obBckmXm+lV2WuleYuRCD7y6beYtufDhmqdzghbZCi+YPcZkmyBW94RnUbuRyCozwmZ+XiU24n
TEyAOkmz/+oNseLmV8gw/p5uWyPlSo13g3jBWsIoNzL3vI2A8evEw/48uAqRwtQps24Ze+nfk7UW
jbD+2R7s+596bm9dR8STzzidik9nlkDvOHF6Grc22RT/7E9S8AcQ1Djm9JQph6XrksIoN3Ru4h3r
7uoWsLcnNSsP7zo6Ra7tE2HtziIGSa1pfidDM0quQJjSyGnv7aXOeWvQXyHL3WeoR+JPqm49FOfB
C6QSMlwt8Hhm1RKScfY7kQLpHxI4G/tJZe2a71Y3+m/ZFQHJVHre4EIKjcDpmJsP/+pMjrgOcvxu
ojSTXq2HeW+8loMd4Qswuow9Mtu9iIhgQdjo+XrS/hxb0NHDdDZhlf2A3lJ53GFf5rQw6ZA4ZExc
sMx7RN23HXmRYnSE3bxDOkuA/8V5f83lRFTD6dGMnAFgrpz2lVCOX57tPWsq2bx6m3i8IZiGLxoE
cTZTzFc3zNONocGibQ1b0noN/q/kTAyqXUUUv+PaMiBk4rtB5mPJENC39HL3saOZLMRmYqAOEc46
kdZgYVpoM2UzUdvIqTDcb/9bpCpG4w/ymOyKVYhgF30ct6ZKcmdxIWPPiOMvkZIoy6Gax5wHdL0z
e3KFGwh3CoabjKWOb1I++Vlgrxbm7b7EbAxVMi0Suexqf86SSLtsZXU9SCej4FvX754RJCJ+EfZm
mLA6FSEZhLWc+O0VS50EmefQMtFsdQgMAUAy5UDtMs1qU+Cl4Sp2VHF+yc4JR1NyxekM86YXyGcC
Mf58xjid+hjou84d17Z6oG9zmL9FQMAHMqXgrTE6gdKfde5jhikUHHKdekHsUzem4ILVJhO6Y1hL
0qPIC8lurrf/+5aoswsb3fgcnkezkM6sIPipRG2oMh6bXdigJHHisvc6sOUWBFzuMpZSs5iz5xkL
xk2GqU5zV5B7WUfOhtp0S9slgo06thYkNDz0pOIMeTqn2DTCL6L0KdN4d2hmg3FqagRv4nJ9W8Hq
T2mFHP29KUfHK5Yyxtzo+jSuaeETtU+H7OjitcYKh1/PHv3yzM5HCUCKhF05AK1cYqDiYqzGMvKv
2PhfFDOKbMDm52SeraMCI4WT1KuA5D+EKaXPYxCKAtBmbF2dfoulAufojmSyK3pbdQn1XBbtQE03
vKKniarf3QLjiz+BD7wn2c7JLwsySehv2qrtozG1IjCmByZp8zkhrRojir1g8YyPcggHIxUj0VvP
WeQTqcEn4FTeJ/HxzDpMX3Ir4pJqqvqpkC1vPgmb3+fkZT/Co+NfCjd+udSrsdvxL7nf8rpsZg/+
f3GEEwIfFWPGlRBQTOWMow/6pmCzmrZatZe7Q+oS9+XILJbCGJp/fznhgHq/+GdBV7YmyFPuHqt1
MtBVdPpAcu0o8SzCtjoqtgor+WyyC/12OzT0h4ZvZ+iu6zWLfK1+FZiNkOeK6wJLBECDrAc80HYu
Ne4qaMM7AQQ6/CKThuqkgf5AKPm2p7E+Cd+9+BY/uj4Dgf7eHwtHsDTS/T88N9eL1rMR6VK6KLwH
1TVW729LI3O/0UL9+MgeFyHTrm0o2pVpROG3U9969QKhuUYB4vUYp/4PV/ulTxhkIbpbeG50X/z4
dY+GB5pTSN7+ONI7TO4YHKHXWdXy9AmXpUyRhmvMTGC9pwvSdfk0SoR/8iKql8NxS035eMlgxIEh
KPg5+/F7Qai9OwE6JTYoOHE0L0NdRb8926Fwlhrgn15vUm8ZScFtOy/TyezPz0WlEyNQbU0ZQHiM
ZCOpa+NmqxrJ8bhQ3vEyDN7LdaGwUuulhVI+ez/xzGEKOaSPPQpTloaPTNhpwca+db9zaKOs/eMT
zYMw/aHk/HzvJqHcJuet7jEDcv9Gk8aaQ1unzSpJP4T/xmh/0IzYSKKqOpmZUDdCPSvDEHCoVJ5X
Xbh+VVZXco1Udvi3hOWvENalwHZUc39Lmh9BruU7i7T4GZv8SLfuzaWuuf2i9BHT35ywCnkGJijT
zZz8An+2iBIPryOcSgYm5MBBnGece5SVlxEfzq3e0Q6CltVh3QGGd026NRInuCDlwgLFMnk/hn90
B8kXL6F/UFc/LIFTSL7ETLLeXD7Rk+/5/5N2QpnpVGGKEPaRwRpfu2LFcmJh9bMQQN13ACqvN92Y
UxysCrB7XnoPbIwygj1vsBBJQpsO5vUAN1y1v6z+3QjhfATqtpClYGh63rPe8KbVtrmoO2s9Lw1w
Ee+ItrZTRzV2w6jzpHvfwNM+5PFu2iCPEegFC1dgNRL+WpORE5HUq+SGlrvKxZGuA3q0BcnDrwFB
8LYOu6AObHtFqaSyQ1xANh8V9v4dDgvd802xRqAw/P1/QjQZ5vxZjX4WQkYNLKtn9LR2V+xjjKSl
+Zf7WdRX/8+DTlyXdfU/b9wIXlonmb8tTaSQgo4QwOLoqnW8BdMhZbSKPoxj9inMadgsNRAeQ5aC
fA+3RrGSQvLzlbRCpi1j+HIYRjDoluuveqt3PkvqL6j2RunHyTRF5DOWplGBiyXhlBNKQaMd96dh
tumsKTghrI6WGXmMcsdFVCMaFPxbfMjNQ64aX9OfR+3GbmQ06NWteGkCbOG0CJPtj/jwOt/FyjgI
sDrZn/I6o88wFOIVpMTb2ji1ryI0hogTqjAK21ccTcgEuZUsfnaaTN5xV6ApNNvSk5DBu9evxjtI
P1gDghZFUHFuCKcTDWqtXFVcXwmBuiNAmDQmtBBaRrBhof1e7Y31CCr7z8zoi/obCxY0/gjs7GEh
cdgSGBaL/Qkj1vp1iaU3c1zMipwgr+Wpg2h4XYsB3kmgYNpyD593WnTaOm+d7LAeJahZmvxwA29K
xJOhUb1+jaKNeh59+v9+vjarl2RnlNNo3FBbDJcfq+0ZbnxRHzzk3db5kXAS6pkoR+0087THo2z/
NO9P47ETEm7Co75QzJNaGi/mPFhHj1KceG7U4t7uFFNl54yI2lROYNrhFqoJE5y0QmLds+JztXcA
8j0H3tQGmSesWJ7Qk01iynBz72ekvXR1spk1iZ1OPGcKL6IVfK1W1Dy9fYCxjbuGe/pyvzMnPUAh
58V3x/zbDvnBo/DKl5kXaHiPiw7w4Fx1W+/qMwWIdB1EC+zqumplL/tTL/Pq6/2gcjkokslsGsro
ZSW7d3fWSBxqGhcHX913ZAtF3eTm/Kx9F89ifmmWZPY2BzObzRikl4YynpPh981SYFWC/z60yikM
36Q7oGB9Y1KbOke1xJh3dZ/4c29cm5WVNFco7KbqJN3hEF6thZKgxX2mfUm7dKnsaiheMwG4jywC
oDuszG5hXb0MJAerkRkKXzoOf5US5uAIEqrxib7J9CwM7jLmNYuc4RXtwgIx2BAsc9GXH+1PzTuw
Vbtg4OXBF+iUVKtF5trgO0YkXdCuKgi0NI2DgmdYfq6Gj0riGfs6Xzl/76eoX9ozeTljVThYYJYe
6GlZncMyNcmbyJy6bbV+swVzAnKY29AjNK4ROCtpQPrCCRIFtfjITnVO02rW7ctZdPGAJRSkn+BJ
AvQzoqqbxRoD8Kc9R+njWgIx9a12hQgyhCU0eJ2n23sr1R1NLweNZxKUh96cQeDooTAnap42GGPO
lpd9I8WLzhZHri/gaE/a71/gr/GmeKfO3C58dfrRDsbB3zLKKgLqfHYUT4xn09sm9O+oH3CN/JmF
ZfuhG8lKHMBtJp1PVxIgpw2s2gfwbkb+fqvKfgJokXXQxh/IZ70/g4hjIuYw6kIvx+HbQpMEfwAm
CI8sd8aDKiO9OniyCJD4E1Up3iExYCSxmpPzJ2e3ZXhj2e+WNMscRbWCnt+5AXNJVHhgsUDajQL5
WgphbzIHyMIDyNwLbMdaiRMjlhSahUZKurK/VnDitny5iRNxhP/7L3OYRlTIdLeiKiP78poJI37x
I/kp0RV67904Zp72l95enGjT1uX/4aV5YdZwadg+RIK4ZOhVJlIvcT3DYo4Tw6OCeL2cogg5TjXQ
Ktk3kce3vyo1WJyvqqqg88toX9jBSEr/SSMcIh9k4JGpV5kHYnH9YRIySeuiop0LyFFUBh+0USvU
w5ngCtLFZIrud2aCXwUIv4k1j9GhJhUvBqyxJOCdwN4MClnId7OqPv4RWQsIImPGxeIbVY4w9d/e
DnSmt6bRHTinCWZPaLgQvAWRBm/uGWQIG+2LARfJJla+90rqpZYzwatpCkHh6AHkLEclLzfTR30H
KZR9/1pQjYRshDvSBMqk5rg5A0+2sWSwF0P6Qio7XEi5hKJWA+16Cf10qmEJcQ9U6J8vd0NScqvM
+3XcsnUhPIGyuVkYnmbd+Z8aShwMk9V/UXB8nUNOkWIRqCiKC2Zww8iOzQsChi6nqOAz+P4Xl3CS
gcfq3UZ0cHgbpOE4dsbJKG4FZ/uWeEJtRHUKQ6EjtrSoQ+7aXeVsqBvJZrI3yBV1oSuWA/6xT1+Q
H0tvxOlVd/unjqqdMt2fDx7W+uBkzGcTPjp0bCpU1TJ4O6LLhG1TDlBbH6inFu5oOTtDf08UqVp1
Co2d7cQFOgZUQaDraniWwdrAgXJuDp5cqY4Yakcyb/77l1r+yiSK0tsRBjEKj99WOwxxMb5VWAJT
qaufWp/qUymQog5T3q6wFQeuhfUBOnd6czM6gtWR5hN+FRZjWhN5lX3XPMCxo+FtluHHrlv0Nm01
foXH0OClcFelRCS90inaetRzbm8DqcVyVSNBTNc0iOiFhe8qD0EPfc9MI/4LWXN65XY7Qnyngz8o
P2QoGZsNqT8+DPXlKzSVQun8yLDV6+/0pfcy/NORhic0if4IBvhOp7SK82Nkl5S/ET79G35J6tDN
z938YmTYY83nbR+AO05Ly/3BGjn4sgcf+HOo39F7tLgZ0151jnV3SJQvml2jgqdouiVG7SdwQRY7
EuaP/ADWMGgW1AFPDWuAPUuD5DT0iIhjqMUN/WIGzShMiEoIBjHzCY4m4f2rjMZ42tCo0aWymKw9
NqUsAfrAxWankfd1po4ZCEqPORZ7OKRWlxHcGD42iSEfWFBdwMwIuzb3geZZU9M5ijfCESjm/m72
+Mq/Rjmg2u4YF7763SPzkTDGGi8rrhUCy/IDt1yqzQkUUCdZlBOJsIy31pWpazYaGdZSgnpXgWLu
OvapLrisvfjqbmewLEHg2u1ZnfpEvr7ciMqqJ+Ss3OGEGaXOOiE3W896VKSpoLBvpuXhhjlRF63Z
5fU3e4evstgaDLkxgozlZDWls5GnlVO7r7P6P2xKegwxnYOBMngpyvVnrK82I/DzSxqKkc1r50iq
OQQ/TkNUCqiushCQe8alqQbf8M878MwnC9snKFVQ7UEzw8z/vzJl4sMuT3IaePhA+RSqZ015P9wl
E3XEatoCOxB6Jt4ns7FSAtmXVomvebsHD3tnYe9/fsW7DpI9ElPr0WbttJ6dxyD52LBXHxeMABMB
twIipvrQmWI0g5gaZD9wap5DWVG0qrnRHMiLOT03+s7nlH+iDmfP/ZKtHg38it2BipKmpCS9lT/E
lYL+M+6slDi0RTX2AoY6newttTNhvPBlCKmR140gZku9rDwVgw0UjznaqJZ27lM8Fe7LsGsTCYcy
2dcMlc3n8D1bVwP/96FBmTdRQr35oDaUlz76DQVQWrrZ+sXi1knWJBigX86rjm4lhTVVJNnRDH+q
o53CU/jp6GZ4NgudRgVpU5tkzWBpmiLTT9VV4iDaWCjX+Q2U1g9/atww6xDI9ezVdi2YuzWra46F
cVwtXhmk7vWWbh25V3Xpba09FIT0ryP9i62cGS/o26zMEVnPWGdmSCl3xcIIWZa2KojfwCG9b+/j
+R9MQepFGYHw+w1e7u+YZBf9KAoPjIuQND7ViqIFxTlDI+Vl2vcpavi5cqVUsqArz8Xdw69T8B+d
dJHKFF5b0DGi/rRSONYsbUswl0MQE9sBeQJ5imB/b3yIHj3qlEpvADKw0jdra4b8ln71Hm9QASgv
yL5WTjiTQ/0pVQ23/dZwdT8QiyXRUwrkMq2F16ylUxLwbdFSrdWI8iSXbj4mtsCfCkQl3tR99FS7
t3KGYLPTN0NSwjED6d4LuMaN8qjWyGS4qqpK54Ew35cKQZ9Mw0BuIFm/muNsquR76NwdXnJlDjE+
ZfXQMjV1src++YdlhRo9HoMLBz5nYljopNRlHVDIwqol0VKeYhY/gywXCLWWKvjnstvW1j2dLo6H
PljVZqg7rcWUWM3Dlyzb/6tiLMu6tp+kyJ1skMssPwFg3MTKPmDQ+inr500rZC3AiTP9TrWdnlef
NTmTlC8v2GyP2l++pB1iiYKsxT+5QjdFgKePLBOEO2Obj0YILSx9woB8vPVhjQrEM7B2PPkWOoFe
awUhLaraYDZoDW9QX4wGYNGHxR9qCcmPBmPXYbwFkOXghgoI8I4LbyVyWk5JP0c7qvQYcfSc1mir
2J9ZACWl/jfa55d2NK68GLeCtg39CJdh5/xrBW8ZHRsnMecyzc7i+jsP2lk6e56UMsZfnuvGfNHD
Ve5jF3T/SeaUI2lOqKGXik/T3wk/mcBTJ1yu7MbSkZH6nIVC21Mu89JCmnqlOnJScUnPCUnp0mpO
YO7j+Fr/Dq+zmI553/53IJ1fJH5xChGlyJGimDCnIfaxTZFTFlNPXg0iiAD4zsNUFgX3sqkd9Gn3
WwRmfM7Vqt/7n+Idn42tckoShn/WyhIzj7smyn/JcpJVLZcfgbb4Ob8otHZmkZ01ZQTCRhdlSixs
MzfiIU/T1poPmIZCqLWGmqLbuQjCs079wTFTdbX4eTRk6ZfUP94EukdaLuSk8Lou7xd5J+7gNS8g
sqM+ejW6tQ1talGN+foQifoHXHuIONRCfAViVoZKTXR2ZWa5v9jigdqUtUm7k4LwyLQ2Em8890wx
5m7YO5xDbW1iLNeKqwWEDZ2lOEu7VoV54vXCIHTf407qJmjDVsa8dQZBecHUjMXDP7ollmkev1/5
6DSsJIPT+ReWgaZxMaQnJwvkotvJ9p9yV2lgRC32+goUZieY8xwcb1vcmtban0zA5w0vwb07L+DO
1SM3+zB3SBGKt1RPZfNsjpaCwBYOQ7KzGwezb4Gqc3OvIxrTEC5UHJj3i/N9N1PCpBGHr8nT0HQS
9KsW2fv5z8iakuiEWSjsUSa5ac5uUvv+ir7hAfagXVzv2Ff1f1AHpnqcqKnMw8dfwCCuiW7c0lET
yhKhMIh2nB1S/MxQx0nH13O1TVGUtNXcKPqrPf/VpXrVMUCI+R4O+qx0TRAqFbYgnSbjSMWYc0ZS
Uh0/v8JqEvotXQqLOZdJwfEYk7Ad99b20plXbs9uFCq8Zscel2P0cCfhKpYh6/dQKxDfQLbDHIbh
krtpU9OiK07Ci7th520Tr7X9R7hm1JlFtkEttMP25C5ovOTkNxmBF0xO9yJctNMJdOUMmjh6jcer
RiqH3p5l/htB1IwHLYQUTz4hmZiBgiPHkH/4wmS8tUscQl+5HA+9FhvBCFfgOd1ROcEzZQolJooI
ftWDD8w2WAsHzEs4sL7WI/55tmLAsRvedDROfQeuEjUnLzd+1D6topqj84Vg7PKOw946XNaEYFKJ
MSvJpbZI7A7Eij7MliiaCqJErxZHFtPsO+4V5XS0iq4sJ9AvPbg8Iqn/SWKvJ1wInRWDUfyFikJ4
6CbAC12H2Ke9kRt+6sU7jYMPiXLDHqa2KYzYtB052hgdec8ij0Ovnn0ihlnxR+ZCXlgdPgEoXKLC
YJGzWQlhc1cva3mOspjr9s1Cn0tu/Cbi+nbIGUl9qiLo2X+qTN5IUAsuCV8HqXCqIeJ3M34dlDhN
jQZTUQ0ApVd6sqF6wd1mY4/xDssuzUYkWQuS+4R+RahevxSSjmVazFZRMxeiG2Ii5qsJvwHWe0xz
QUzPohH+Q5fY5L/BbHTXphBlTMiWf1TChaZGiauRk3THhBGCiatKYf5OyL3BQIxoI1MR7lSypOfr
OLvStmk/HsI/ns2hBteiwm4R4g4M4tRWBFdSc815zAAqbaVqE1RD+WRzRTpcBcMFD0Ivn2ZYTWGs
6mF0sl5NW95CuDGjMmFHte2oECl7SJ6QzHOX5pe72LWtIPj2tCys+Pw54ts7ebtt9MSxX/HS37sw
qtVC9Fc7GeBPvJ+v6DL7mzjFNZRg145CtQN5kUi/6XFFl3oPNw2l8FFoMM92tjXZEepQPA23dIjm
i73Foh6kGEbz0GDUdd2RKEyGC5Zhjr5NG5ARBl0N/qu2AC3LQ+BXP5vA27NXyOWDh8cfAxcr84F6
j5bODbm/dvrnx0UafKXSeN06bETi9NGNbftD1xjnZQBCuij3A90iFSGKroMW4gMbgpPKvtHhhyb6
tIH9seHHNVIc/9u843dcx4lVBtyZvLSJzBoM6J2t1CRaBuTeyn1XleyUcvUe+xBjO3Y9+EZyTTV1
M/YNf4ZLEQKsZQOCsJepZD/ke7GcbKkuU1vT60lfBs8a53Pv3DT4IqYBHgPTP0zXt+19tGk7zhek
FTCxS+mQsgE6q0iRhTxrUOAcBQqN3wjE6RElkBMKN1YeRmq+p9WmzMuLEldwteqCBoA5amsYkKEu
0TAdnDKHBKzVcbNQ0Y8O0VWbtql6tM20KJmC7sjTw6oOX1n9pr4mL+4QyKTYbchIJqQDMh4boRBN
COZVC9POAXy3koyZ+74so1YVNIXZH16BPwU+HeVX1bxbBqBGiMwZZbLx2nrPdHRTrslAG6lPuEP7
9MLeJX0/fo9dGD66aXG9uWcnBhXfDt3u2pQx3c/rD9HyQaN84uaoDNeFRjSYWA9ic2z1+PamwNsb
ykhRedoZj+09JTij0ljhipGlwY2N/UtmMYKIsxv7icbD4NrN4s4Lj068BSZihcGeFkyfQP26EBpN
YKT4KIN3el9d3PygSFHqaMC0kPvg2nMjRSl4+hESLWBnA2EzL/JMRgcpNLr2LwIkshnfg+qglBDd
gyukz0dFeWxsanVCG11+pkdEiWbdj8RCMyyjReKojLRCu82UyhSuuqdmWnFo1KTpZASJEGYcQ0pK
VajTu3Gka96owihpIfpoz6S7gUwwjnpAidUpomcgfTEDI8VjsEEO24nOj+FGB8Iy3K0cJ75Ryao9
GuQKG+btro/SYNkL2MGlxY3AL8wMmY5EKzPOEqq5rxqtcUmVjAewpSnd/uP+hWpbf+gMwvL9xIdp
N2q6j4pCUeby5BNnY9zWrM97KXOZ6gU1iKGKdH6+DVvGrZGP9MBa5rM9y2lmJe3nV3f8BWDWrlaT
C0+SsiMGIoUrMX3KFQHIZf76QwegeTnbUqUghrfRfH4Emn9Jy5AqvduPsOP4k/V7vOFULrBPu9LB
JYd8FnE+gnOrvUaWLh5SOAiudRqu+aM7TUe7iu+qoLoTtxQgMDt0J3ssoYf7xtZodR/cwKEDOyqO
fgR64u4iP0o07KQ9Ufh/6biigEPLwrZo20bS5Aa7CSpd5JKYIgmncCm1IxAopCFIgyPCmROTXtwO
+RWLRlfDTfgl/1aGxGAJiakpsMrSPxrwa2TspGQV15Ah9XsinK8qh5uH71Nyfrmovk03RPJTNj6+
nq/sJfJBAvGDPlH8fQYyR+lLVaA5TPDYLfjYOQweUljDbtq9OcPyEu8LKt8463P3KuFPtsrSBWKC
lShzuWqgLHoUXJbIE2jjD09tIvXeM9tOgWL+cjjYmdnvK3XmnAoQOrX8a531Ij1xUQBzc08XkdVC
viKwExaWBJTPABLX0vOkNBIbzShprLoFRja/PiKNDUt3K8bWYFOEdRWLlpgRGXSmHyA2O7tLFy73
RMULGdEtWDNXupRjSDm29D6XDWUP9vk6oslPObNEEV/Wi8TMt5bqE5CunrR4WkkUmAHa28bLpnfn
Lfh3z5pLx/WtIHut0ZOQpXC7iwsPzoCBmqerMsMW4ygLDCjRPiRPFDYemGlSihYqjwfOw2eP6RJ7
4AYntbxmzLMykfxurRanJaFO80U6+E0XuWhKdDW8cAqqfXARIaCtPom+hJGeEr08xdd6/1TK+tLC
uCXAge/rl8moCrqjuIMBKiamy3OufyhoEjXf+1fWSjjJo2CU14B8ftGDddy4dJZ01NceoIeHuuV4
76XaAli8t1Ea0m7OqfLuWEiNWiW2/WHcCTa9KeKZlTIs5MQg565z/9jB3QXuQRZ8DTLqUuPYLJVa
JMytqtNCQfWRC1skvCmbQ5G0V94h47xPfF1M0qMGQP19ErQd0nwezMB8VmHEDi1alBHTI/Pt+23B
OpAb51tsyK+Ontldc+B3WBD2BTGiS+QC5B5LpPgEUlAgUZRlxyt25TM2kt5rx33yi8BpUqc8/RZS
ICRuG9U3mQAnGqFe/EBsBkdL/PVtydyv1Ule9RhSO5GCIVZeD84jEw0aazB0AxjTog+wtwKjNJWV
1n9l+LBrRNd45uufRVGqIY5donMbEPNlBgredTm4M2HTopC9uCT2SxR98b3FP2o5oisS6uaGTIim
7QS7cbxOX8g6r1GJBI9n1tiIZ/S3P0+yq+aFSdPTHVUb/4ayscpIgf6RVD+D+6VDBGYURttqo4ez
ef8GrG7kmgcVYERY8Ci8qfY/jSkFHMN+JBtwX7v828kMvPblgoZE6eUBfyraluNfSVDECLHdGPN9
DTNA87tudfwNgPC9yssNMjPGxsPj5KpoIfIWyjKxxjMdwOSVGpXZumBlI6m/CWizRLO6Sg951Qgd
BY1E729LqHoB2y6lTW3CK+KUtYGjJviy93ovJWEzi36C4EEJUXT1GcwHc5ArgRFG2Mwr7BCqwx82
soJklSClPqaRyAOcPIpVPV44idqrlnZzg5jIic+vcyesF7QjGz374sfAGCsZZNVcvl/vl0tyk4Im
jhInzusFpt9MY7TVNU6ajcqQu9CvePY8qwUQ9jidVgkYA/drAryWOSu/lLXn3nRUaHPd0uMfhBXJ
0Uewmrs4HuB2CDYNOds28GJD411dokobABkEC1PNBVOTeVzSd8ljZFzb9sS7zHrcJNxVBZYVHzLc
8Tsi9eMUdYLyQln0LNCMAQF0nHSMO4haQGeTBveZEohzx0Y93P7xr8PlCzMVJdI1Tep2lC8b2Nz6
vHvlcpZq2VIET3CelrVzgGTXips1N2sbQg/oj1H/cC6bxnUPbAY1h17Q5lrIy2PgErFke2JzmCxx
aHg9GSTwnFJ+0MF/jvoCqZtSmKmIigBZ/XtD/xW5X6P7UAK5Em4AVeOn9Vs666MOZb2A/ojr9crH
AJsnfGTW0a3uIcN5JWGWULzDEHtsrcArJYCobARZI0xF71L946KMeRCWkaWmoQhU2hvLbfFjzW86
8/qE+j3RuXPqwAyktykeL6CdyOSs46NtczscMDEEpC/OeROui0nhQQUcThmQ4tCRiHjllAzCdqHm
KSFuSCOmXgTvyevuO2TOG+0F5nt+nFJlqrwptPWz8IZxCrg9O8oW7rNnv68CZd76c+n1wF4Iweeo
URWk/Wrh+WdNBPF1f8TzdSqvhK9praDKFqZztGN+JFqsa6xzb8iXmCr0uLvfPNqIascuxcs0t4H3
+ukwTe/Pm4S0JvX5WCNa/5Dj8XGfsKyZgSUXr3NO1GwvVWcI1HRqwNXMijLiXy+6Kcd3BaRz+RXU
xGfUELn32C6QP4/rUpZFlypeyKPX5flxx2z4L2EkV8QXyw3P+ZdWElFQJblP/fCpzRgEaGu/t6FM
v3QGltkZaQMkYNb7Cxcg8zbJSGag3TfVLp4OLRNTTZTdCcO+UTIyilitmnbqz5cnNG6ilGkU5ifK
axY6Jcr7YKxDwiSfrVVvSqkPDfBkenomzCzevWMF1rDFBgpK0GyfaDAPuLHRZcW0aV0W/o7UZhZi
BVSSn7kZVgakNQxYspTKXesohk8fSdgtAkB9i0pdRdzl29mwQvpWAYff5IshvcDXZJgc61tMH6+1
xKMEICGpP+qD+IB9aekr6BBnAK/aXbZ27PCsUDqlwL0pVYS2z6y9KP35pAsw0J7BYa0ynDK605/u
flD6SV6nMsbP+1v2H4bG5MG7FdqzYyy3CzP82hq5C1/kbCiXhTA+qxHiFmHUFpvnQJ41fmJKac8/
MjFP33Yt3LLDznDfzQBNF+vWm9I6KzfjXEjK/iMxJtxdB+G6EASuxe3JFX75FFUWKl2jZx0ZWpwO
mk8TV4F1oRi6Gl/0nJBQ3IVaBdjB187XZEZMkSZ5SWwUbpcXot4XkgZMjlaeD75s0J2yeFOND1mE
DhVNFTr9XeY/V23qOx7p/m6jYsx/bfCzI8IJLL8U9KXfODAuismXBJFPgyfhX7ptJhSZntDGHuqS
/lfPxmMzfqQ74HF7mhblji4F1khfUR3JfEdAF9V7U6sBLI+Z3Zj0cmMX7H2c5gEQNmmOx6CWuiso
xlwyiY0fH0CMp5I0GNNP0TLbzvJjX4zsiWa3MeSgw7pWrodlZW+6OykSIF86tOvu3l1wPz+1Uvj5
hIt6S9GnVHpXtPwhxmcxv7Jd0S8jInvGrwAvNZ8VRbSo+eEHHtVMLWYHSvOiK/2/6EduMRV0gB/F
bCKS4YPV97hqQBWA59yKAePznU4VSKBDi3fCY0tXGNKUGMmUm2i3sORfc74umjZiB3mB2vImn/JC
ostVi172u7UI6AI9bzg+84FyCvftPXNiwgfD+KHsX5Mb3wWwkn4f/wGt00DhLbdgREf+xeLCMQ0U
VViFZyhp8vE6A0IbjWtsUkYqzK8o8UVae02YxQBgW8xhzSDnRC/yTgMXCK87K9rYGYoJZUyQwHgY
qkxdpm5gzYG6q11fNKCKUUW1a6u9Wdjo1iCrpY1uF/OxJBrSncAYhgmXGgiACtDJwCF74FtjLDJQ
UJSAWkFkghfOPy5OEC26dCkbwqlUZ58bS6Zui0x4vHLDqAwqZtBbR/7u9EchQ6slFR2IkvEQTTll
gUDFH1z4M7ko//RNUJEBiYHn6gBkfScb6nqkWh8a22Kc/2ngtCUuXYG9WtdWjUAe8vWZsCuo45Jv
WQVy6UDW1INpzRuZvON/e11crDgwc3r5pM2gD8OMyWY+WtJDTNnrObWh9bKIhbIMnfndG+k+wPJY
5OEw5g8pjQKC9wDBjO1CZGQaFHG6y2s0xrmP30AfqmggkGH5dMg+JhJRXCMhQZ2rVInbSwfxyRZN
AQk+NISp7iArkG8/Rh3GVAjlv7FTt4KOoqogrBGEWc5073qFag9/FhJlLvmVgcSbYj1DfiGeZCCe
VDG8Y82VpU/7lClg7CKg3O17EdbsA240Adfk1JUQV1I1I9gwRsSKFsBLH1wlo84W1ax9kjta1NkR
GQZltgauwwHeYrT/MA6YN55WmOeAQ5BK0M0a+wGdznkyBVEj1mItB2tGSauaO8etVyU2VHn69+26
NAGKq/+mFM9ll5NfbHIX0u0A5oPfncikDhfSTVH6HQccBs91s1PqOSk0ewbC9GoApn4UlK7Pihqx
zlD3TLdagTb1Eo4dzWmeO6smoQX+uFVSDznpq/6KXL+S0C1XIeYQGjQHfDWKDgtgUB5Jbovpn+a5
Ovx/APCQJM7zGF5bXhj7JxBIQCzkOAtq8xY6i5jjfMBTm0dwv/rfbWZlS7mB9av7LYq0pwatn9Oh
2rQKGU2MdSfXCpfvpC/DpNzgdQNGEmkJfQ+sxKQpqCXZo3lcxERXDInqFrk4Fzr+QV9WKMoODPN3
wAGBGxg49cU1O0Vz6zK1G6rHkXez+Ctty75fX3x3YtbFYnAlP/cPej6amelc2MZ2YlH/A7l6rsAY
abHXaFFc6oKGGHwuLuYIoJKlEJ77TI73EO6uILVwI+U7sPTgwHXYw8/tQR93J1CG/PZ8O1TctanQ
4cihykIg7PYW9+JTu6P8eMECFMxyKwCkAzjLSQkCJb8bQDTCpNXYG/nVNob1ZQLqjzZV6QSiyu3z
MU8fkP+2Hh5ZMUJdjQW9a8WSMH0y+DSv/MxwRAxdXUBlnnY4k2S5Hpypuv2i4QtCDuMsAjpofOT2
aFQ9uM2OLeVj1DVJeXuSabAgW8TRLJ3k+TjslLNoZ9Gih0kw0JStJQ69gsfZLjlJZcJ2Ymhmquis
q+EQZog+WxuFzd6OvAF66PSWkazx2WtcbpM/Ou7d17NL8i3STScfaad6Rkph0fMO3vJFVFVo/aB6
N2nbmKbfA/cZnBH9HEk2gnkbNaGLgjouKPjID/vlKpaur1FGOKbP8FLwGOJqrb6gO/lqpa2zYXsg
eGxWd8OhNwzwZ7Gbx/eljPetjb2o9WeYXEP/hlyyP/NR3GSASALmxJLCR+s7L+aOybXpEcxwhZwD
OlAtfU/Wc5WY1wJWte3gMuD95aFxXIQEE7MFLTn8qulsLapnM12iTzDJs3r2yVtopUVXzdOIWo+o
rZxBFErEj/eij8ow9P8IOrxtmDi7TIY+akjgDVs/aYJEiCOaEi+vSO7XVRS55euXuwUK8ypPCTGu
cp0DDWVcJYnCwUMg8V1hL/VOoGo9j9AUk67XG6g5oyIVQCvt7E4pew3IOn/JJPwEzKhCot59twBS
NH3MjNI6Er7H7UZXKiXfeB6gbRfp3wEADU3teh1IY4M7CIye7CpU1nwSPeWM0SK+rwhd4xOE1SxX
qc0hSB1B3UcFNSnCNQVg7W2nTItLv+deaw8ps5EF6l94c7hLgKZanCDnSeM8WdjUUyUeAIPMaE9/
/gyNtht+FpeBWt2G0IiESnskRTDmWXqnx8ftZJb0izhVX4NzJjwuOzlqmuno9OflHL+NOWIsrkzH
o1eE2UYkhFXLzhr7IuiCWo3Re+W0lvcGVkgXa2uPEb9/k35BK7Z1WpXW+cjwzC6ivvfzpWst3Wib
kieuzSuHG5CZSnE1poWsCeU2jRwQmUvbC1tIy5+h3Pg3zvArZI2FkKJcn336DQd5ahwEQ2FLepNv
iwg78S7WA8GmzMkHZFzFjTQnPMSK4jApvT/RAbe1IID1bTRmV2iEULeDAdYwnRUEbeTBPoYCkhdR
WMaBevcPkQM9CDucCglZ2nRbBJ3CeDtmbHFF1DoVAX+BkSYxQTy4EJGrQ1OM5ZLR2fM2/25aoLbG
6CFxJ40puecT3JsEAZ0Kxx7JdHTXLq14SVeqb55VS5zW/QTFlII0qmfNc5XhowVhEovYwy5Y4XdA
puahmXvnkhQpGPB69s32P6k/ySWSK8QqA3nRTzcM3y51PoUY5ygDDfuP3VvQZGrkwJRpznEYjoSJ
5zRdts0he58hg0aNfxM2Fkb3A9xzxeZ4MkjsNlT2wthjif/E5iCp261yzFFd/LgXJbAnuXMzXM7q
JmAhdNMHeKxOpJBvYszwFu5kKi1R2HaNM8GR0Gbc+RWJfjWSHqJDRpyO4Qp2/pMunvKRK6pWTdP6
ONR8HnvfxiMRwIH8qGdNex5ydFT1FfBxWwAML8hPdqyb4FsM84nNA5ltAoJDZXY9JQbzLeS2ulnq
aBgZW6Cej+EB09E+FmxR1JAhmEcKLopzmw33dCW2BgePOeeFlH2B1jVK9JtXecBgWqyLIW/sKkR4
iFpZhfR+EA9LVY0VVZbFtxod5PwmPoCCOPNV/QB0uzpdg8ABvOHKeAmJu3vyoi2IDNGavWHOK+Fk
eXW7ygbGodSpXkpabcckpdDj9i5r0RA1WoELdzgDA3mrpwXgPUcys96mjQ/buBGCLTOBotHSNgfl
1l4hS1Ko2808Hzgjjdxp580Msu/Z5smP8kBSEte+MsLqtquv8YXk97WuQHfY2jkVkgHaPPAH8WsP
r4/BVXHK9wyAHec6uoG9g2KiQmZ1t7bUGYTpwvhuSp10MlcImgoFrrqf8KFqcxNZBIZfomo0mBnD
oN4DwhXlKNTnrbpw8pjqA9SB10xofxrxls9X8A77rxdoniGXXbfqYounbRwQ+Kqh55fNqXWqAnnf
hWTXVCOiZJgVR749CdrccJeGDvQjwM6tnmYKeIX/Vwlzi73bXlZpGMVLAVzP3V5t4ye7It0S3FrJ
PMTfpsVPzEIdI3P+7XaRYmGXWzQpzPKGJLPnsYzBLF6hrdW0EolVREuhEJvkBaNnWHfgXiGjicMQ
w6b4cbxU6v3kXpPE2apceOW7MZi0Jiwb/v6Ew2JCk/VtjkWEUVJh3ZfAZ/un4m8pEa7U+jUEjG50
AwWmlKbGL2fpghInMVCFE/ZNNa/uKFMvM5SUa5TvnvCmsM1dFSyNoTwv/7lUhlvkWt7//KDAPNZ6
hDYicsvNVGxjSQ3qZgaGWoVM7Ds7xqqZ7fc9oha2CsBnbRssRXtxDQPfXW0avZ+GZavs6wwzp9xe
5icd9MBWBqS05FZ9HF3cTaJ4JQJR1KskCVoHeu7HXgU91HeiUsFb6hyktwThtzwfkXGPOXOgHoVQ
sdyA84ZEBJMhIjChzauchwEeqUbwDHLHQJOhWxZwaOmM+73tEJ4KKHlw97WUtDLO+iVkquNyngzh
8+fFQuSTn+Yn07Xt1qMlErqndpzSjCXBUArsu4U9FrsI10gKn+Lju1KvZmtlR9cjpfkyOlupoXXU
qXB2Dhmokt6ogh+60WDs/ooR6xh7+h7dn8gjoOCR9JR0mHeMwJV3fSKKt+WHemgk8fTINdKWKX2e
snDeh2UV+4+D3tvaHlCaLlGgtpWtEjcZ/YitZY/O+o/hJRpdpfzyd0lIuPh0Fv1g0ns33BujvxJe
vuncwaptYwir5OEZJoF3aHCRXuYMF9le6+hLlIqJlLeYzjrVque+hLY+7W0e7WI8gYpaRXVKlm9I
54YhDAS0QwoPxaLBeYFfFldMUa42mKVjLaX8HPjisX+jJd1YNGx4AhmniUTfq+zbcPRHFsfBOU1h
nDWBfqvms83aouuHweuAbO1XosLddTfLJTcXomlN+Y+pGlhOVKzEXD9H3kSUsuxulWAMCiVzHOE4
lHZP8BJZI6nik79/x1Ek6qPATFYtpqzhI68Qa5ZM9mySN5otgb3ApISgWQG8BIPHcR9IUqb4ZmcN
51A41lrq+cODVEGOu1Wy5iyPWAVuWzQC+muBu52WkQaBSVoVkoRQFLwJzILHwmA6XyajM5M76+bv
hNad9tjm4PW6C+6Ojmmnw469446lkcuIE0eGfkobk6Uy3LH8uQ5Z7Dcan7FKhDJACOakPsjttlWg
oEwlxarciS7NP/Gr8mw3U2LgI1LCKJv4VpbY4d/4dx3ab8jicpPkMHJQQXL/6ki4SGjWxQuK/ICz
kNZfNG2JfG4r9awTYH0uEmx7ZNDbX7ECcJC9BHuMJmf1GExD7i4aKXZ5387vPL63EoptEQdchF81
SWqdC7q6W8efMCzMGu4ITOZRKXIhp78rDyt6MrliWVyLrjbOFu90HXPh4jFPYBTOugQBToXvkeyc
L870FuseSDARf0JaGjHX4hyrHO96FgkQgn1eRX9iNZ5sz/e7fhMyRQsF/aRk8GtADX0t8U5ZhQ20
VbSgzZK711a+LXz7n77Jcbi6Kt3qaf7Els6yovsoe7ZCrwI+VG6IBGSW+9H0qsyiD34OP/FJNB91
6ppJ6dUQbqtAb+hI7dZ/XUNQPcT3hNafD1gHjCEszP+z6eXeY3HPSLw7nqjfhOpc1nceKRiy77aC
wPrmxiWdsM3pvEFYELrHr/9N0RUnJZ58TfV8zq9MYoX6DlvqtwcbuoWRpYfWEVxUk7mDHPwQIZ0f
x9FVrTCfqv2gnEM9YrqhzUtn1iEdrrZJodchlJDdiiKYMOtLJzAfwD9514CuLkM69NH7IiWbq34A
OyzdMLrBDK7+uWjsx3N055JQMXQVQYTeZ47xbFcKJq0ebvpfPxpg73V4skCG+vC9QJqUoS6w0kbM
6afYuvmWH2YPWz1ah3A2zIVeA2DPCEgFVSvAhM4IOoVJmteWU1CPOe1gfLcvjB7eqseboJWabmU9
Lzba8B9kVcFGJehj6F+0xnPDPOytdN6STBsBWzn3yrAUH8C0S0PDPPUBuC1J5YGunW2l0tnDsgs4
HLvIOuBRGOToLWqHAQUdbNzLhggejU06jcdj12c0QKe/ts/LfdKau9ShoD8np+dk8akx+Z0CdPLp
lD8sRqLe62Xm/sjfaaIzL9isIez2YVL4SrvUwTr2qGJ9tJRpkhZtKVnq9sitr5OUA6pJYNyr6V+k
piwclkzR9BNnBrFzNcm645BpkK34NgAlSvwozNpvvT73ktJIMDYkIw97jYvwC01OPl3Okn9kWWrw
RRRvneGgRVG/u1KKseEDxQkTB2Xzi23bfze6JZvXjVGeWczbvQ0iDJhrB7alB1Db0Rcs+sOOMXun
oOYrfH8TMcak4ytV7M7LMof+EzUApeRbCBHOJUcQi/6j22VeqT3/+p8/lYYEuhTMnIYnBN294Lzr
3I5laEHsTqdDO4Z6M7Mr++f8ffwADcadOQ/AvlzO2F0yKtKbnM8Yi0M1WGq/zn3gXnUzXaPv+Oax
bZHA3i00e/VMemLN6mgblcTn1e/CHpEP+zJbJ1aaaVXWjCTmMJSaqK5iQSvRvhsbYTfdz4rS2bWF
SbCcDHvNVTIW0Q78ZVKvOkGp7VQ6mEBFPBZUFx30kVj/Vglkpq1XoSP2IP3ISUnEyT5XH0WgaXzD
VMDztdg7k1JPkqum7OxuCJL7i/nAB8VzyOPkFGCoewjNW5bo5COubaD+fq9pcQW+WDS/RVAlLfis
v/UaFL6rmcysuTfn77prSL4PddFPNgsfYSC8ErkHpXKjBhEbkrmvroIuPDnF8U83HdleeBNF76jN
wXb3uDmQ1yGoobOgQYgXoD0j5bTsCqFIdJQzZQbiCWXBhU7RE+MLB3pZqr+bqWbAs0fFfhsRbuhS
dELpz5EuJ0uPqIKcobrP/O6lsBdU3FcJg6RRfoMjbXCEdjJYtuI2jDklxwtc0/Qmz5vSvxhdRkVS
6sWpdEFQhzDlVMNJIwehBORshfYzAccq+Bt3CvkeAbSBr/wC8yargXXF1BStT+TfTgPeu78hNedo
8dpmCdb6qZG5XCWM8UW+6J3abj/++Di5qB+17wzt83qAA+wxzcPW7LiMXBYh7egWVcJSCyLSAlC/
jLRsP2JhME/5Hh6EgeFppTMYypgc0lM3/ms1FXFLKQ+ub0cHcTxHUELGIzdA5GKK+vw8DbPYr1oZ
pB3XPGVz64RK2nPRNymVDlyCb4sZW08Q7ZdKTKW68aXcvO3eMH6BVE0H0+7Oj6IJsbwl/7fHfh2f
DCJdFgMEFGWc/F4RJa88yTmE1DERj66B+uozzMTo3jVJKS5X7FTgbfjr27QrdD5LQIEQ1mXLbOty
IrM4wGDvpXG/bH0aOFYWqhPWNsE7k+5U/rSfzqQWIVrXI9rTv6wrZywNlAeWzerXAuRunsNxg1mt
PgZjowysPPV2ttdXg4nv5nfOTb+ob9SUhhQKvHLCpgNdTpLckq8I+aSbJHqIR9U8bCzuL6ithKVH
l29G2JPKBIULW/tYy8DyHKiR58feC9uNeFpfhEJ+4sT6SntqOd4+B0eTHt10aKTr/uVjwPHuZHKV
nDSNz5llVacim4ofq6+rD21p0zHf+EvgyS/2w1m7XQVnzJzclF7EpAVPTei9qceydUM9r8EcfvG7
xHs+RSscTPWk/jgyTbG9nYt3x+x8FnlgGDZsikyqJ7ltStL5xQmzQFnYehQqmoWjovNriVdFGKw2
vF3WyUQpBVbV9yfQs7Shi6qZZggyowk0MuvLLy6BlRVH7C0ceVmahU3X7VA6qjnyUtd9thh9ipVY
RCxngeF0MwwRgQ+OyD4tuUVe6Vk1CGdMaJoiQU0myyFBByyfl6M5P7muQdq3UcMnWdP9Wx8gyGNo
cc0FOjt+TOEup9vJqFjOqxyNTsfUj6w2Ot5TcQPWonz48MOfogtwn+Ux4dPhNeb0hcTuBfdbvdd1
g0zfAFuGQy4KREOARLt/V2rUvhyKQNhk/WhS4vo4BXKQH5EKtyI7rWRl18m0Wv+nsi+j9LcORyq4
n6s9ln8Cw78tNbOk994I0o4OhPObW0blB38wV2oHcNnrT5E/n0fMaSRlWQKVTITLsvuIwfNNN9En
Qm1kxNSL/XRB/DII1J1zlqON8fvTTtz2MNRaC7TdB/pkkTsPTWBH0AsD2YfkQYybGa8OAb3nU+/6
jycGQpYO1KlbgXkU8HTa89OZt1r9VVfC+XNV9bHsVDmBwGSR86etKoJP7b1Lh52kzpA1mE11uwll
y/nAPFrrHVMyd8FOYC5UlYDhGzn094WDo5flIgpZ9Qbwwr31JQggROl0YeQZubx84f2ZG+FcYyIQ
CG7tbbcQNMATfXtvCUxnjRkKALNX4C86QqUH0k6P6w+jI9ZX7LD6UlUit1a6wePyGorj9Mi37phL
Mjaj/hvycg/gnUfDkaydBzUJ+aZS39Zt45NXr5b29gp0X/J6mFmdVwAKYrlB8IbOHdcn3m64oLG6
3dS3IJgpudktYpGhxR7mwnRW9ddiDO4T9lglWjI2v10MNhvAeEfXsUSKls9PUqyUU3qJHBFQYjrk
QTX3YLP5DMmMEvQndvNDhwGMlXEyVOO8vkiMtaGSmT4l8vb30Sw829Bgq5qA2FvQgP5+LinfgSt7
eAq3cN3oqDNRRI0tSiZeRKpCrcsCzbeANJ10vT26mvYobi8DQebnILEaIqwbKriSpx8/sfKbhpMg
4DqVVtJEJLx4PbJQYbD7EqAiNsfldFNGZKmSedT447gk6wglo4UaqvGLNaAYCHbwH6wT7lW2wAnm
1KXwvFX91D94RZtxtPklZduv82lLc5r39y8BMLtScj1Js/TjuzruMPSMnPN8ofkFwDStVAcqFm4u
A+YohWI2nq6RnjLKDovLsi08aj4Eg2meVboqjIIttHJacKME3lY5DGG6TwhxFTu/ofY4gmGZqToT
Icmaia2aKMBO3TplHoy+r18Dv7TRVj2C05ZFZ1HSf0xRZw9L+tGDAFYSObQq6RjGswZv3zUFgscB
45BX9e8P/fo5+6IC1/btRQbi8rUl/2YpwWoaxfFQU8EgtpKlhIWpbFGyvqrc6pnoL8spIghPQbH2
ZURoBJXx6GEPb+Ytr3rwLu0D+jE0oMrn9gUzXvewsiyFUKVuzfRUcj1GzqDjBWtBn0XQEgSv6/R/
wLehLHa6jG2tqDdSnPJW+HwtfSG8KOKTtCo7Ny94V4aMf0Xnrjcs5BPkKbe1E3t8O29OQSJGaUHF
9Vhhwktj7KsTEI76ku0YS6o8u7V7HdE/XV/TbH0/Or87X8qySiv46RN1whhW0ZfcJCb88UVggzlk
38VAVEepjyvier8uc6shPM5h2BZlcYy6O5+2yBJnswuh/jem7oc67/c8Ao/E3wr2QgdgxBoIO/k0
WZDxZFwfixpEDhHwr5+j420g9i2UptKj8OLUh0V7f2Qjeik7aJMPAWijDz5mm6PPAa+xk6Z+6fzf
uvB0ow37JDnG6kAA+hecQ9IW5kif6tqKPAYNeCMe/Lnm/haqSoP7Gd+4vj/xU/B6SI8SzdypdgEu
glIJgIq0xkw9AEluHwSFu8w4G6i5f31pJa34w9eC1shlLAf+9HCjrz0oGq8l3mPgZ9zM1rzH5M4L
EBtLoXlBL7QXdKDoc6kzdg4EUlTHuh31xVFpH+x+rec2hsajMPOwloZm5tc4pcPmQw1pcdRAVP2N
e5XjlsAriz+oXmYN0iDwAR4O2pB8h036648wo2HGIEYog9v1f0Bz5b6gwhOIsRPLL34aDKV+Hy/H
X1+BZRZvGhZ90c62Xq2wlIzefivFycLH8xZqjac3mVDxAlKm/VL/AzUwoiZAD/1b2rEuCVQHyyvP
kWKvxQ7i2CCL2JbahJnWfW7bExjnIwej4JK+gpexsaodWEYewaKkfFFz/HZKKZ/XUIIFdkzlmkN+
9OpNhAxVJfIOegHlpMbYsPxA43rYD9t8xbOJjA1S4/shkdQz9sgVmnT3yizMc1lNHH0Tp7UETIfJ
koZ0b2WFUMVonrYompSIhJtYMASGfMuQ2JVLLmMbkLhwM/WesR0Q0f1ayQfc0vjMOjA9kyDu+fPG
oAQIa6vZuAC8MnX9CxQVXztx0EbVguia73rWvEvnnP9eF5eCC3oqB8S8N0w/PII8V92umOzPWl5B
EighEbU1k28KRI/U/PWJ/jjIW4NhurkzMbqWzpq+I+1l0pY+nxMkdOPkXoTAgjl2ehE7u67rdp4e
nf2OOzIch1czoOmnr3SW6AwRzW1llA7xDK36pzDpF7XBtCQZrpOoNU6bU5Xr3eI90o1ZWkWy2b1k
VLXA7LQyZufth/UF5Embp+f6FyVo8tpwSjHksLwQaExdGl6bvz4BrFPOtqfdgxzD4FY3QhW54elW
bUyDNIBwju+IUNHb+kAo/7ihPPypgjSkJ28tPiH8R2elwRAosZ/PKOMvG0SEnQvHuQIO780VhHVj
FTRvyWNRXuE9s6ZwkNd/hNVxHrhLbluDPseGlWFMMqMK6/2+X5C33cFw5Ywd8oaREHL7G9YjjzvC
dC4S17su7ieNmcYB/+HvaokOKvHCnalNvC2p1BUgAh89Fym9TmucD4zUTf89W/+KaNpqS27dtQL2
Y4EcUR/3hcD6S5TliXqONBO/saG+e71y/j9Z7MwzaMU/inOomGeyYdFlLzvRB6GSAZl1lMT/VCIp
GQMXBizRp4lO5TQkD0o69/62gCdKFoAYSdxp+lZ3NY9uKjwyFCpiqJca4Yvjp/QMxhfp7GiJEQEf
elbVg3O0URNIVFQJtnbJxxjFvQUd/cYfjl6uEdK2bU3c1N9SMulo/M0uy9cDm3Q7z6TIDK071VuF
nB/PSzPxmW6U0xGmRJVU3FVNJbk+UjNFNNBjUT/kZWLIo96NMbSI4zSi7zgSxd/ohvG3R53kxYXV
FivvgZ5bFGa9ab2prw+plMGTxzlXK8hhaMToAP5iXKPYkGdGdsaxDgVwq2qL1T5uaMd56vdO67MT
bN29LtgCOIPn3BqAGeCUgIkK6cu2ioOTdkEJIWl90p4/R6mby34aRP5lzing1LtEZMLoronBD91v
BfAwvgm0WT4JKUwGeXPvSCrsJ/4EB9UFMEUKlnJwqMbQiRIgfypELsbOEhrgkyl8gs9ECZI00wgO
cnjf3N5Yn1jqGoAZdJLkQOZ1MVBbFwkrLUuXpg29IxiWUqTL/oilKcarND4tmOzPjxndaOcTeSRz
UtHk4iKCuq0uVkkG4Tn0TNn5bk35/JuhllhcwDXeUjxHXNlT+oyOqbykRTvW9Z97DJUV+PGeg9qu
8bJeKVe7IeImiguoKQFqqUuNpSPVLVVQzHPVgBo4XYeJ5VmOUAXeY4YbFsvAV++U1myzZJO2EWxw
9nyLmFJy175WshgzSbfT2QuhGO+OUlYTZgbQPCRQCDlyqaFDYJ/XZdy2Ad8SsW7jwfFbSvGKZ2O+
ih53ca9cx/UwUdJ1c+y02quAfiVahu4n1EeyHcneK3cX/ecskbEB88SVtr9QNylJCw81wVE0T9a6
7suyQQdjsk60SgJOkoZh4sr4w0WlGYGaGH04bBMet/QRnKJBZZP1My9ttB8COmv8IQDM094dKKA1
JpPbL3DLd1JM7sAoeI9cGFIMzHPFzAji1TifI7/lSkAYt49RSlL5xSJNOPb8cDZxfUGwGfrvnCEO
a1mzrtjlyOqMFDLqQXWgWxVa7loZrfGRnDa3vGyXQqKrAXnssBdF/YIysBXMJe4DxZJpk0tLaBv8
TWv3JHkMDRWWY+GLMeqTJMZFZo0Ur/MXLfuIIQ8YJj0ZcDUJI1Nac5hQCBlZ4fON8aPjohtlVVuR
k/B1c+co096H0M8t5w2YjxU3UlCr2VDboFCeaMT74LSSl7fW+a4CZWUcyzY6kYEE2gPZWcryoe+T
kXfee8fak4R5nP9cyAUxqqciBupqJQAmGxBMM9z/S1Mz7quRXYKdAQKWoYt4WNoLv9oOqFROVYnp
lTZbPwUmmakvcweBfRwU/+M4X6Bx8ZVZgkqtignTbJBJqhHom9onTqwmFSvrHEm4svGO4wYAYzOy
26PtPYDEnNUs8wKzOmlCnNuOBGUoLiGdLpI3vx02c+lOzOKiceHxUwgKVdOB7xp7zbcmmH6TkjFj
MBEi+5Uyfv2dssBycNznRfF3sF56Czx5vDhSMTwzVdWvZw9p8A7YzOsgUp4oHBibR2YoHxCM2HD8
ZYBkqf0JsnlWPkzngiLmVXYyrgw3ISA/soNxr/ov1bIln/cI3Z8RJWucvEweHFstDf2O9E0nMYDY
3C54enKHrfDFF39FvFLJYRcLl8Mpl/egu34HblOf0ISnI9V4gAtn1MqYb2VIaQ1iTbbUY/4oMyrh
XssCMFSXLJL4QFrn5LF5e+jKKj1fWYTZ2IBYp54otxPibf75DCkGvJzGhxPChRFc/TsGxymF0kfa
Ybd7PADRBcw+dREOSO346MZWoVLUnhpm1oZMtSioYVRImDILBxdjANvNXy5RySH++r08KOvCvrhy
rPXwNZF9p2oMm66rNKHa8sPJli3LNxDQGyg9/iaqV0NzUM+iyo0DzM0scpCs8IpID2U9eAF9GpVz
HLLl/7rkFHYxhHaolxJUq5Bl9gPiLu9X4GMcAakljlHGy3KHrWZqbVImlQLSJmYLv3ifrnhVU9KK
N5CP6LoYf6HrXz9+Wshptyo9kbBavBVWX04ZUdRrfIocUpFcksfPaYiVRuwIxGpSGFLisHWSM9OA
DvWdTEgIRSof1wjcJNkdFdSKuQKsM3hr3qZJQ1dMcShiNvV8dTYg3yyXlj9AdEOZslzcG7BHHubw
S23EDXQej4XO9CW2uAHes8nKuLc9ZmgYMEbWmgpABCCjE+vh2Y7lE6fkDbIP70u5K7Pz5FUcNsVx
RdGIFKjQHyi98pVOK33tfgl/i8oZOBqFJSnP0xhCaMSs05P2CpsSTecxYBRq0NpfUKZAbwEvrYB5
7Ur6eUL0bTgkTjCnHCPhfNPHBBvujvlhVn9BaOVhhPtDIUmi8oPDXNKh3gJPKDZPxtlbYQ/zwHtF
igj8QI9h+YrkRLKE9zXGQ6UV0xboXadJqnGxoAWbbgQ1/V23IgiDVgVYGTT0C4pw7q4/3P+H6W2E
vZWg88GAA5XYzgTlDzDt+XY7/nMlkGMFpdaJvocwJ5i79eNtQtg0Us5WmMh1vNhPNO+7oEAoz4Gv
ddJ8wIGWm+j0trx+JN9ESbnk261uq89nhsX7mgniXoE3DVdHhOXHAED+zryCJGcSlI2PmqyMN9Db
a55/nWqU0lTvjGAlNfGk/eGd8Z/f22MQdwWnw09nYMDgBgLFS3kJKCJAiHiHPOK/OBbpCBipQ7xq
3RKNgwAjGZ9PfGzfobcFTkGz27FVrcWKSlOCO6fwj86gM7V8N2Xea2ZINRqjJBR4wAegB/iFZlsY
FZTUlCBpI3y7eyBehgAn5syIz0i3SAiLNVYVK5adZCMVon1akWYARe7Ae2WPLEoDEUu42RtnsIq9
XrnYdISdTuwRHvg7j8/6s+iF4IxhBT3Y/aQAUIQe1UgfJoFV5QBuUXDqyKa2k/MOc/rz00JMHaYT
ZBTS23DD1mlX+K+L5C9sYwDrjqliB3Bl3w5u/myMqFCYcMxjtKtX1NZCv3LCJS/kE8sD8+PFfRdH
bkMpDI+AKTBA6awEjfCN/atk7K+82Erw2crSN3/zbvxS3IkWG6EYaYwK5dT6dePeZxMmDAyVyAHl
wVXtIPfrVvaB0LqA04LlQwL+W09zNKe1M2/Zt8mJDDDMTzplfcyDaZjPfv4mbyx/wril7832uZda
VOcYSqbWG88ekvwcqI/B9eqQASrmzfFtOoTAdLoyyASq3gwWqfHrQ9/mPey6IY32YE9cDgXnarJ0
K8O2EhgzW7JCHwvKe7ruiD5nXA6h8lqkOHYXWVWMH3yj7FDnkArDV3ODtGhPfvic4ifYPpk8eAT6
KU9djSpfiPNCtXpr3HuosNtuZoM24NdFC5YRgbAM8J3CpVjb5bw51rlIkb6asJXByiT8HYs06WyN
K5u9FnbCSPhh7TtQBH7QyhxcFbTbk9AWRp52QJroEQTdPnqzZlaLAqGuafEH0RrstLerdG3XF/XZ
aubFCvLbLTRU3dJth6eLKs0sdgPsoEub9jkQy5GIO8L56dOxoaK2B0PuWhBrMvMafqHB29hKMafG
Pyc+EWXHHbVEPhHAo1nRIe0C9v91qp2QaMqKRsWKRM4GnJLnv5gNvk3yG8/EfY9feNUF1bIQoFEH
qcthvre3zAZiSD7Y6qpFBmVyaefHBvRWTpyk8tA1AB79ZSl+vdJ3OVuhCoNYSbbVJX2Rw4QvWKdy
HsCC7t2KLBzEHsG0rW2wcLmiKASYjqRlu6lQ/qBCkiU3Hu3n2gxsQnNA01ekRRQCAXWqS2YwdUGP
3Z84U4nxVRjZV9bqIAbWi/Vo2JREdtdruLu39SVkc49SSwv9wEgJ6gOAa4wl2XogQl2nGPh7/NsK
JemkPXY6gCNhwQbiCNJ6GyIgDhwvQM4az0UJ0tleQgLXkNhOcCZ3DI7KRZZscrIRGNwzXsnBGPOm
J5B4LK5HhfDTqAWpSk8ja8oe9nARd5NY19EOGIRGXsX7WSIPlrNM9TUVnmYhEWXcavzlJPRJAlv4
EHxPya6OkQucDDinOOfkdFfymUzL81Y9joFlcFQvkg/CrH9BZKIMmqpcU6/NN/95l3n6+94WGjSJ
0tvrKbIKLAgZdzjmVmNGr1Jvi0SZzKfNnA15E/JqfITAXbCOgjUBur3ax2Vwak4oe+8Ahpb1U5LQ
jIKvFMtQkJ+rM5XpIpAG2XQ6QM1t6GpqMtZOzqj2vDLAYU6TCmHk1y7tH2jK/t3tTVgVYJjYalUz
Znnun8F2OS0Ky2WtK9PjDK/6yxeKOLGRg5TOEaWPEjRatfzXftfmaXnmw6jeyG90ljaai5K4nF7N
mX7CdJgHuj4i5bjZy+ZYPRuRBjBQc0+tmAOOIh8Roh4e1bvKqke83RpkztEBjw/E5GS/iu7Oy+R2
VvMi+1mOvCybLqhRr5IFZYXA5vpQoPbB4ldCFp6RR5wmMIYF1Ae2OiZ75Ujx0MxHowDLbBRQW6n0
GM41mNThbcy+0DvieQDXobj7puHJ6SrdLL65UkWWdI3kmWG3xDO6zYPnc47aoVtVUGawhz6Q65iP
+nQdVI7UPyTlJcTtZINeMEYH2VQiGn5XBMg5GlIKRCwXwIskVkdderLlnvhwf9Y4Y0siqcV+Erru
2dlo7nspQtsXvn5X6wWgd79bu1JZxGHW+vztieapmp+tHXO91b4/1mnSOBQZGGDdhNFhw3RDZlB7
LaJKbGu3G73iPmbzXEViURy+lP7b7AwLZz/sKcouUHw+A4SnnF68xHrU4hdsKrRsBZWK2e3zQGPW
ru8sjYgwXE+GcfbFhwRr89+pOgNZCPoSafn7gaIk2Uc5XtEwJWGFCaggaA5XDWHR107fAUXmNRLb
fR2qk1PuDZphCdn/yWUq+gw0FUPDS24cYzrvgPfflJzR5Et87aVY2MUntV4uJReVfRkOf5Pcdgb4
ZjvWFLZ8zkWNaKjkWuo4BuKObdiOCg+sjX9iPX2wcZQaF5Lr0m8qnVLRVkxIHbdmarxU2eywNCqq
R69SjIi5apVii24x4Wl8CP6rpzE0yhKzw5ESIUbwOeS6uNC2x7g2dRKagNyssxmVk7XoFnZsvwaA
t6gyIs3hlr8SUblKVMWo70vw+07yqCYySGqA4o8srxXy1a915yVFhE0D3E4Yi5Om0wfRAUHbfdFG
dr/SV8kIRFdm5xpE12yJ3g2x4m/OA9YSwmeWGiKKiNXksJnoJtRdMYDPCE0fYb18ecHBOltkpU2k
43NYkGVXrboKEQL+Nl6hk28hjn9se5DSUjfPsY+qZ11CWCDRIvTsUfGOmKP3fzvHOk9B8Bz2X/dr
01MBpqdajxA3oVyNKExXP2010fC9b+GJYJHrVVtF9iUq/+5LQGGu8FMSkK1Pv9xr/kRYfSco8LRa
gvhHashWdidujA91srQJ1aqymc8LX0DjFVm3I8plqxim5i3z04ZYNd06XgAeuFEfFkEjGIO3QWVR
XGtjXkbroCKi25DIMRLz6g6wIxrgvaHchRWPi+t4FpOmPjtc+AZbeN8bIgBrxotlWEHXs6WhnFul
/l1Mez39wkdQZu/iEsD3+b+cp9g+LgScg9FYC0FQX5f9BypCD1I3TFo0p8pWfwTIO2I7D3dAIgL+
7FZuXpVJbs29alkEnAg3tLampQu3jn/E6Q2SPtNoEuC9Z1eKsk3FhjWMnWnUGHenMWxotPQ7Weil
N5tXEHfiYRGY1U/h+WE66XbXAY6b0sLPh2NZgZlnm6QbZa92s7OaJKeXyfrCI3AMNRHCWhluNB0y
zI9DL3vbLX9/QaMzwDEqkBAAqIKkLA/2qF6B0UODExL2ULUJyoy+sEckf39vhXxpf4old/lrpSFl
oonDTIyDujqeOIlTq5jzkoF0ogQuj9AlIp06kKXbeBq3sFdepwSBxEvCaC08T41wLTaHpx9RTcaf
zBen9UYU60hAKpkh6PdwIsNJHemwlh4TJ7h90jWZumQEQ5Y3lVMUE80QOJNCEVwsysPL3rBn8Rwq
31Ruh0S+KLmWjhRssLcCE4DyQLnK88kfENCpnjii6iwdCdFdjfkALn/m+oVSnJsp5AlDNLtcrzsc
rBJy6EJM8sMhXvdYeJ/Hv5qF0KcvCWt+HMB+Km7x4addVYH28jv8q3BHi0QTz5ZwXChfTDSrjxzk
la2B9j1Nq+8NgsZBNYrPpCaoWsGljjTQiSrRsfhGDdCEArwzHXIXiYIob5adfDo/5KNBOcXTOkCv
8ZpbLhUWMO5PSIp5yABwqLuMyt+pRZRLEL7dyqPChhIa6Di8T3Om2OLrxeWLlRyDDIF0Q1to3zNP
WezU1jDXQKJKVw+jR8L7leklj/MkoxqQlRj1f9zThSk+Q4fUaGv9QoPHf04MB+VJIjscH3t9YpMT
SlPoblSrroZYN5YM4uwedUj3J7zS9ki6T+Z7QLnFSjtDunveWS8Qe4as9Q+HUx7ua5cv6crHYoQN
kYi1k2EfCHAT1Ian2Mqa/iKuU3haUSn6Lltm1esJF1wpWXAYuRN1o6ogIwh+Lmm7Gs3/iCaLSuOW
HvmusOijyop4uZOuU54BOTNCeF2EwbjWLH0AQI9YKgJxmAFFp0OZsqJJQSQjtn+Lgds+bAKVDZ6Q
2uDbDZjOH0Gt5Fxm7RkcbLTXzPJZWSYY2h+aHPpO8brXLFy9YZAtQSv2wCW4YyT2kbAWtN9ZNt0F
oZCne4AOvwNhB4UhQ3BFv1hiH59nz0hCb/wU6StzqzMeNUAYUh3WIfS/QZ0fIVUr0z0bdKnj6HEw
q56oE3P/kVtDEWF01XQ5c3A5eDisWp5GncAePlFriATWgF+XtLD3HcXRFdqBNRbqRuyvNuHXa8is
OuYoN4mpy4lcA1BIZLQaRM46mmFCSnMT1REZEFRSmM8b19NY046sZSn7DB16+UcqcLArUcGj/tDe
IqF6PKmpQVpYjkCb1f6z7w0XOFy2y7CrwOf92a2aunouGkM5YwnGQZvWi1lDETF7h30AFtl7gNx9
kWNP/kWGf3k8xcAqkOekbrLnUnlCFoqkVPIgrN38ILlI4491+lw9RNY+LsDLAgQEj4NFMA7aPxFk
JUym5suUGFr5ARLPchnuTdBxkC1RDaSDQM/p+gQghr9mOqnLVZLaHMOgXZFevs6IAmj6db4uUGgE
HBtv0dQsqq4sNfsjVZuZ68AfSEYp2bEqzkLbVpDkS3WeyJH5Apv7Q8TNOSGzDkUiW4Uqxc6svYVH
/F9U5i2fMzMEhxHOZiSbD5khRKUkWK5yp2amLuu5PePGYREHlHZWCgTGdtFIlPJF3X1E8mydGGDV
b6dmEV7Xh8B3qVyML6Os5lQzpP/8ZD3OePIAdAlpYNej1lFon+SBJ7b6eb8cWJgFbRrX3qRraQ8G
eAkBKX3LSmzZdyT4KrQbk9HyOs2ExwkPnnmLPWKG2OzmtCYlMDmUaCZmmNHvJs30kPmhth+oSd/c
ULAi3+EAoJarVTVYhkN+I/VSDcl8UA6s1TjPPfN+CRk4WHm4cSuoYY7QDYRQQiAWYF1kueYlKz20
suEw5jtdDQ4eSrXClkTSqzOsTKVbzecvbrt8AAie+KnS3NlK23lpi3PBDcg29wsly/dEG+LqqBMj
p3Gezy9B0ugvWe1KjjD3I4EH6neHKap1oONRzjfX9o5kIsmj9Q44xbRKT0rFkyEVV2rshd3jLM0V
Y3zwjsq0Ks0nLIsOfGZW74l/7h9DHFkmYzYx/NQHexYGPySaG0hkYnI7FkoIvHiyRaOFSkc/NWIJ
kVnEEgme6/fO0bgH1Xf5w5kSkcAMrF/8eRSWkq4mPCyhBgneuxfUDlEacMEHvIl9RLlT0RXhhc63
7zlAeehwQtGfvKneITKGvbJe5Vp1TZP55OO/E2LzlmELiUIpniL2yOyZHRXxrq4buSS1/SKtqQ6z
n5fS9ZzZTX24gIbkqwZ332mvFJs80ZHPQEBIb1p/9Kr7oV7HBwsEBGWZt+DM41F6O1Uxzb06oqYC
FAvZFU1BpMweWNhHjGIfkrFYLzV1MveoRIcRa44976f71f2z+tXSL6Ydj7ePNC97fAyo016Co5aP
X0UJcKrNhevUZDY08CAK8x5gDFpB553jIPafXZEl6t7d5AaM+RGZQbj4z3pQdsyuGEUa/WewL3m/
IO2fgvXzDxtKtWKPt49tXhHzN0FQKp2KX2y5nMnB/EU2hs5/k1eDDsI8/J9Vn95b92bYoHdp2hUs
91/TuemwEINmPux0tfnm96AOneQoa1cQeN3kh2gPMlNGPRX2sr/5Xebn5ZqWQWIq8C78yQrSIJfd
KnulgRe52ZwJc57ESZaVX4UHNkbt7rsSYY9vyHjZr9D9NfAlLWsRsZ6v8RKcItpEQMQsxV5Vj+th
s+xcZN5HT+uRUdX9R5sIrguLkN1zbjyui9DRDU/r3ViqFe82sPBX3Bk1J6ZjxHSeDtjWfUojl2HR
7Cd7MvTvau3PLtdXZimCGjRq0SqyeX88dFM46UbwptACpmKnckY6a4McclOMan3ss1NaPD/e7/yl
2R+EPYD27znPlO8P4mLzPmf3aHT6jMHcF3itMWp0TTpW0RXqvJJcTwwzfaRbTUBdkPDQP6HlhVOI
JbMMRdG9rHjSsaxTZX3Bt7/b8iwHgVxI7vwmpPMw/eTuZzMQTatBq3WxLk4rfYHBAhKMuEhBlFfj
r1vj3nwJBC1aoA8Xzvq5xI+uv8d+XNPucTrgkoA3jX8f43qPjTgoggg/5aucdAKnabDXQyvjqEBY
eXCxptfRneFXZg88kiLxjELOVhtl8Uz3tLsz0B2C6ce6fZnzp+7Tul16TQ238587ukYJxiFCh+aK
8k3oWThpNe+018BI8+tiagogEa9Bm72qvNVvrzySvWLO3CVtuZl1w+Jaim9jWUWdPI7RGiYw8xY2
KjY2fBte/8GexEHFyS73QsCCfg3zpnGi4UuWmKhoe4C6HW1nKoMuD4J4jtIQFV8wdBb0zX4MZ6as
cOWqtjdE0AtRwqNq7bcVbF+CiyreI1A1M+nGh5idE1YMRcPEOCIyr9eVmqzWwjQ3Rj15PPsaD0rz
51w1oxSsoqrVmuH8+6yudXBGhROsO6hjkHVU0pyjPbXm3tXzw5Io2sNakGlsfuPmQ8N5C3vbTXA4
C4JPnsYiv1j+4zMqX3vX5RH/7Z+kTmZeSOCdD76IxjyfymAn+sBKP1UVFdhRJ0UU3eb4n9NEPwaQ
N2czqpDZzC2S8g9JzgqDeRFEEVHWzYfHAY48wKZt37/fxW89DX1DzmiIyVnQxbEnHDlMUXY1QMc/
ETLivbZ8cFQjYefuYBFmHqj+iSrvETCV8X8TnrCOaB6U8nmZFryt+Q2rWgW5efgTs3fSfd7MYRkf
qCVlQxM1itKeBVfgFtiwAC2eb1SoOO3l0KGMSGXYNxRUXtoAb3B4vFmheoIbdcuqmJJi4CnYtVAp
ym9+CIS/JP2jGEDKYq7ztUWQsNPO4+OjtkKIOoCXIeoblX5mGz5/muiar5uemTnA5GyBH+HEgJ65
cLD7SHRPVm8KtX1jg07K35YNLL4NXFvjy5B4fwDF6HjmACUo4xLMov5UR0vg4u41VVRobsMWaoa+
8WRU1nXJmezHgaxd/LrXdbPIqhfOhANTQPvN1HqtQuivRai96ZLYibNPMgG3tXNPdl79XJWU1cvl
2PpgTNWpsBJFfWm3t/nH1a12TQqTnoVHRbeJv44kSUjpYzRQRTxM36l9O01Q27hKkaIos6928aRi
YNivqiLn6wSUG6h4GrnwL8aRmC32bxjyxLR5FM6oDmH4cIWG8uwT5VoXCcleqMD0txq6m7Nv1MaO
OQvdqoWEsPA0gNcbv7VLjkSRhSTpjPvuV5mjqWkEaK4c34OLE6PhG/LTyJbFCEct1NCCmeuxwVO1
q8rVFmYI+8HqQApnTKGL+jv7YUwrqIk8rzlZykNjl6XM66df8vQE+mHHXdtqJ6dsNMUL0TDhDT3U
jSi/1uKXyXKbU3lLpUgICm0Vj+i+YrUR33dEV2rTaH46pyqIo0pDzurtAJ/cCj9dJxdxV4feZRGl
mG/lHYn+QHA4P8Iy9Y2ZJVMaxiZ36F7UCJpJcI6i5VRGr+cTanU62vT1jWHTbixYm1jHHS5hA9os
EC/so0eQrrNMgekhJq/A89vdCKaMu2snpHcA1MG9gstVeEvsQRZFkT2Uh/uD9MUdNROnldzwvQj/
Gqc2EyEikgo8TwanBHxnShTGS+7bal2+rJhJKKJ4VVcvqEOgf9UVcPSB634jdIO0ejw/mBLkkYP4
1QQrt/0MxFByj8aqQdsZ1Xgvrm/o46wujHWUAXRsF6wLKsHmSyGa++Hs8JgDVwu6xQac3CS68Bm4
eiwqzpr2+a95ss+wd201EbyINU6e2kxYNqr4zVfeR63TvV7ECY1baB6JzsM99MEHlR69HE4XSNEZ
fXadOW0zfcZkPbqKpXP7GnvJuAywHYk+cQ+8JSNvYgIxPZl7kTl+17M80lKkVWUZ8OgKzvO8mjAY
Ruc9uD8nntVzTN1SWJoSUE89nUAEllXIZN98XOs4EwDv/JJFW6vVJ8zDAcrkqNc+1Wq3YM0a/I9U
3g9PB2IQLkYbzjeT/72JFwpaCZ73QT+ebjksigM6pFFbxHPJnRb1NlN1phQEWhbjvsh2Er25EJLR
qAsMXLUnK3cCd/NNDG3nFqQf67A5fqeZhbSIeIGL2rP/ikK1cdMumuE5l3DhXOsk71nErsEygONW
O2dIf5/Wo84RGnFz9Lu6R5WaJ5ZzczbEn3rJApOWVwd8Ryz/MOAVQqyXRG/ItZUU8VtcUQL0W4ra
9P38ewmvX1V6QnBpoVafTs4KTUdxepA2ZPqUUKrFwoR3gli7Ik1vbOhdxYkg9ZT2XKiW7EMCGzTF
yP+BSI50lv7ZDgxuASboghZbSfmO3Onmrczmy//u0Wna1ZFkC1uivpnzkfMPjEe7i2lHYQA7T2Yc
QDTHPHSewEHZT9T+1VUKxhz7UTI7By9hPACdIZIDkzk2qpBtYZ5u9YhEl0fazCdApSwoomaInhsW
925WzFEM/Vo8XU4BhyV8JRtgbKkp/xTzZ60tKJA7pck17F3gvQiSj5AE29rjC/P+MZD7fr5QFBsc
xLyhV77xk6sREtxd/WwaWGdpfmRsCnqJTfOB2CznI8di4QMvliEGWO7jnZR44DMEN9QE/BdDBU3O
9KZx3S+lxLEVikwiY6atx0HkHEHfL6pnyLxHEl/dZb3oKr2k9e9IPVxR+8vS4UN+UY+pR9E+AV3/
pdX6K/ZjYFmfJKtagr59M/GT5lUNWBL9hUZzDzKDh9Vinmub5yj6zYLR7oxyDRKvneFZIQPm8eb6
EqqYC+QAM6BsMoBbOkG8j7a/Cq/l9/n06bQOfYmlmQIVCoq3ZXKLiCnwTV//oxYobErVG5UjaFc0
1ltjGorgeTMCQbhe9+ASRN6VCF42IAXB+40pukVtw57iFFcARh4mUj1S18lwobYiqpyFHvpX98Sn
E3pOW0eY/U6a8y0tcFUvZPw5yXsGo3l4gStlkBuSsrxXKqTLEEv4CcJi3PlUmB7HOoPcLh1y1MqI
9d0Wlfv3g7QXgdOQlWUAhIRwEesI/8V06hUjZBEzHakRBMfVkG/uxkOJlzKAuLAJWBgd4/jKszVQ
KS1ELXXOBNl56ZmK8chZuBzWza+5iAo5MD1xRMZKjnOyPeuRoAqQ6680nFx6ImYXcNX2DVB4K5zO
O/v45IXxkJDsBV2qaDG4Q0VfMDK1d/uX0rn/xXbYYtjip4tHHyKxslfRHN7Ov77EEHEJlJHqEhmK
7Rc/J9q66t3YUSoFUH4SQywdW8ClEFyJDZA13mhbDd6/8/Is3vFIN9vWfpiAbmkLs396PdzcBTMY
Tmf0K2D/BNkgGIN6eYgadDuDzSIGRibLfHjpsqBPo8/707GQo5D6o+j4FredFBEZOR193KALaxxm
IVU+LToq4nJ4Mc8dwzQZXNtj73FZjoppxMy+VWxqUoKXyt7J3b6ZXssle8/NMTosiYW8GGu3o8G0
oM30iVtLxmgIbfpK7XEl4aRs+Xuo3VVuuMZzracKRAyWjr0Du56fy1cAI1RUyxpiKP1Ohmyv+Fit
0PaYWW0xO7oR5kpmjv1Tr1pkGjTW2p59+B7LPbOB0bhVg6lgGYnzjdzusOM1tX8dYS3o2Ta6qlrl
g/LKSx7f5rEqgKwCTQIRhuLp04gMH9tsqTTp+9EvRInSkJWGC05P8F3KrtKhrA84IGAZA1awYjWO
U/+RtAKO7n45XtlUs3Ipe2+MehJJhAJEQHYRiCFdvD9KEVjzFnwhqany55pFjQp5mTflnIxSXlJ2
zukBjmfe3XdA+ab3ieJYfWRzn7a26G28gOWHRX/1YdN/n0qDJ4tuXFiygtkmp1MWUuJJx1cDMwPa
NyePTDifQQCn16zxiFrRszPUfkEThM4NmPCUu/WgHj7QlawhCac6HZOn3kFQpL2n0BWVah0wTMoT
Sy6qJ+eHFvUVmKmH+QrepkxADBdjc+WEd9C7i4a5pblm93F5wYCy8UXmJcqIzJbBsuVJ4EZTYe0e
EbfimX2y6TacG4bYYvrZs6wROfQsACRMtvFXCBLk/1DNAlMtgpnJAr1EKHB9s3d2ZMP0QEl2FuNF
NpJlZhAugqwNF3qh0uu7tCFoCa9kVEL5kCCh2cTp/2P5GZhzgSG1LRVF1SxWbzRGxzE8bJqDexQ0
bQH8uQxje4kPFME45aSuzSxExcs2A8fMVGGMyEsYVvS6MFIfITguQm5r0pJkHZPyqCu4/OC+NADq
hVYe6ZvBZo4m9JepQSNkS+RaCz/uhSIIVZiYP4RlzJE4slsY5T9cdnSLh4BGweqjuUA/wUV6QPVd
ri6hpiYS06LvdB1n9TWit5aqUGqFsWmY2SDfrNDqkj2JxhMZdS5KA3MPmUyuV7A1gS+/Wv7WrVcn
AG61kO+f91XKMiBXQ3Q+gnU4pPE1hPoGUN3Nf5xOiQ55FGIyDuQITD4NphEEtLLe3oZ6GHJdB1G8
xD73jcVNrBPtoLzuC2agl1RtLMwOU6PsJByusIg1aa/WEBaE3MPJEk1Zc8OM5vkQ6RA5zlWnR5KZ
4h4U3g7OKX6/lipktRCmFW2efxMyI2Qg+nppxelFMGhWri9o5CqQBAtbZ6M9DUlrI+D26l8VNs86
Jg76oCS1hAJ9N0udzN8/HUyWAVWXxLmbO/wiMGuRT6J8w10O9Eg2jq7MkRAZRshH6dg45GgsbkEO
SaAjxSESu8gzYuzrSRUoVSQBa6ui2z4+HkfrJRlzoZxZ8ZuK9MRtcV0uA6LE5GGFJGpDcEee0GAW
kaOaTO4wrXEFWGKGtykQg/+t6zPYppIHsfq/kGG66iMQYwNV5BosazxLt13JxIvymPrQq9OhJcTv
KXy5pz5ZGZW8yLa5hTyS7r65/wPJtuTQ7+yKAxb5w7/fQIYI8xLfKuD9QJ9J4MLDxNTUALreq36m
015gncTwC4SNM9yogfSWhLyEzmMGmRBXy4/jYgCI3d/g6GoZnTICJ8yylIIw9FEv6VdDPOJTTjoO
rqcziTnfzuwicmAD9bj2rEAvyXhAd243q2qJH9X1yYp8JW0xHvtTSBsIEEqc4bABvR2Ew8i0cso3
WKgiWNJGm1vBwT/3fwGTExj07uxGbC0KxUT6Chtj/3fdm6uuhsKDrPJGyS7coBoUmyN0rKMj8MtM
v22xSb+Dw6p7Tkpz8QQfn2eyUDIroYiG2v7lv2YuB4CWegDJ/OPxPfJ8LyZM6ibjSRlZxKEJCTDi
kfVtFeOVvdbiYlq4Foq3qZZnUjrCgNm22g2rA2X8pn57H9MwU/8DWtNfmvd2vRnK3ofomfpTfwqZ
mbpVhwl+nwm3eGAPVus2bxRo1X6mmxaUvpABvUP0wYkBMqPb549miFLq6Ka4hGWPNVuRpPWii4kE
vJMTZxwAVAYJHktL+UMMkuz5Kj/MGrL0uVHd3Df4pw6ivB1je4ymet72373BZt0Tw2o6A6QRu62T
Grq6GPqaCve1t3yOjSohhUy4XXMNLxZv1GcidI96YtTTcdptLz+qS9z7dFi58ajdeGjm9t0wkGt1
wJXay9hNGw4HLVYm0QfGcOMGQy9JOxV7CBcw5rIPQCyjxn0LeZYjAsTyG6SttvJAfAozsh5VmeHS
DHQZPn7o676fOGxrXlB8WB7ojRJvRjKtcDmMHmL7rwmCD8Y0rt7w7gbJlXL0/Tf5EUApukZXWdcz
dbgW4o7rUwoZChsqquo9M1f3Ir3rz1nj6BVvxggxndKifgsLtw9OZOezydsZG0e9/okMsQP2QEGW
9spvMKkrY607seftNkR5OKSvZGAqAsd3Ec5dRaG8aurNLijnErjrWScA6GE7o4e4G8RNY1Wv3/lj
8aq5GBWXPqvhoS11oNlfnJbGu2+tPez4leGc6a9nYE3lXT3rCVzEnfuHEOdYu1v3DruIUFbCMdCU
CqIPGdAvwbnEhvesSrBvGa7QCLIjZHEC1YPJBYZ0XZMp+2nLjwK2ZlblQxxC14VsKn+/MIQ679Vu
4bRiVL72Rv0uvsakYyd7HM10s2LemEXVU/0KYn84ow7a8/r1P4iJMbMI3IcM9WiUUi3onRbh+w+k
6rxedkRNtp09jp101cjE/mZznIX1WSYcRvL0LQERFEXxWae+sC5ywu43sLQt1hfx4p+gmhU+JN8g
tmG+uA3v0uR1rYqA2chAyYzkkDw5oAiKRVybQ+HIb+5n/WORpuBQXJuJQI1IfD0nRp30U6fItmUo
+m0wOxZV95u0bkcE+fZb/vy2DXVJgA4NkXJgXKppwa/9GHI+kVMiYdgV4o7yKrlEqXwb1+LD4I9v
N43RBfR6V1CHzgRLsj5SUOuPQDRgZ+6LZci2d7PPDrUt8pqqwtzWNW1MdmFNTeVmBJov9OPPeQhc
4tzWbXPtRyoPkRKqBy3tC8itHj7JBEXpkzNP/zmF+jbA8QyPPjWPua3tI9RjLaBSB5q1/Dh2uNGR
+kfcTpR/3BDGWQ6aVb79Ox1fCJQ4dK8tkAmLw2Z+jt+99pVhre/43HZD8i16EOYNBcK1/aXkyUyE
eWztEIiQK2IWyFuGicA2Ch1ckbhl3L0pT1lZ4Z/wh7f6owUlJKSuN5ASjhfvk+jBENa+FHVPzAhr
/SlHdwoWG4hN94VAT2VRHX49X5Wua05RF3pbn1p2tQSwvwrEe/+RTME0aIHIXrWpPkEAkJ/flU2B
6TlcjNTzsQSpO6cynvQy13I2+a5MQuJOX0KNYgqtDqxUjhjGHjHnqzg4L+0idhDtLTEkW8rDvxkM
3d3eEfuFmk5s8b6f/zA7a58urqINYO5NUZSzCkT+RxVTVvw0TjAkUt72hMheMvLuCC+OMOZogeJC
ZYjW4xucVmi5a5Itr4cogKGIysta62gooJro7cor0AFX0aWOSARXXHuA7apoPJM/YJaXS+DZB40M
UYq9IHSrxlz8QAqvRS0+XDzQSvWZPSUTmzTDHx5dICHQatLpk0CXDoPSE2erJIqKCNN53WPWTU+3
Hr+eHFJynBq96qx08ODurLTMfwETJ8OAWJBTpfs3MpmuJjWrdDqKmSMB6qSeknj3b/tkXG3Su50v
wE8Tsj0fNDh7ktkMUvEYPqBZdCfuxwX0S9uPNxggcPsoBfhOKmT7fpdd81IRjMpvr97TkD4iXZA5
Al1NPbCAMFuw3Ne5vph5gUOVe/tnIUVPlG34bFwnj0aKpvL7wj00Jyv2vdz26Mxw8odFGP53ZK2l
jskT5IiFb8TQfkqD1Zoh6d5AQzMKE5zoRCQSTH4Gbrbbaj5bk2yjI8rK65oVRqEhwBKeDTOlISLS
4qJUG9KJ9HJeuM0b0NDcmXGQ/VvuV2pFJzYXYapYOfu++zu7qZckMEJZd4ahxKBXwwlndVhLVn8L
nHyN3v08IiGJi4uN+yRtpCCuXzaJkjdmK8LEm6Z1PDGLZorc7o4xi4mLbWKObHvSF2UhpE9M3jSo
Lx3tz/wcnQpIPGICk8sZTsMTv9WNdXU1raJpPJSOIWprkzVktg2Alf+J9JWED1iV/5HzYvvUGjPr
/8ozMzbIQRkcyTcxTkZ+3/T+2XnOHp+v4Z/x8XcEYvYv8jOYXGL0lwNgo+Naw0jN+4yJj6xjOnGI
XniSnwA2PRdU1WD4/A0g+zQg0vnSFf47sWcA4DyGOh/nZq1InCt6vjAmsVkzH5S1Dhg9wkzf+yVw
sn/w60WoL/E7W6lpfL5Hj/CGvw4nfqR0COypV/VcmTDv+T3xfw6TLBWGbNAYRAYBDcIyOzIk+eR+
SG+uC5O2X64wtwPeF4a7IoLcAIctlfQGTNHhuuau/eaeYJsiW5B2cXAiJVJpxQv0WyWVutW4RbNT
61HYplsBIHgTU3IHM2/X5Uw6UWxUFJJf5/MlVNt4QaygXxNYRgAvedZ92OxHBu/1DJ8P8S2cDuc8
vRjxzwpfPrS3TCyg0Kpim8p50lYAta/l39/2o+zDdTfkaJY7Aj6Xi7W5GwJAet72tFcGGf3a37DP
UA4EQ6FpUnUH4FJt2hqzx/JUt+6w9oCMeZvDb19Zv7pFLVSDRxnMZI51NiKqcdtRyFonwtLj0eNo
Azc8zg/d/52fpOWlAHImFMH6WYV6J/U//yRgpMeQL1/975/jrH2Ho8D/Ob01i6sqWesQiAfmUY23
+1bGyUstOR9zCmsiBNfiUL0uy4tFuC4EaLoBKYa59MjyxyKJpFzkxGddMf92pPnU1TuPwX7AG/MT
Ng89fw9HmvvaOsoXGq4Kk30Hp28gv/USnuu2pVbwqmklW4RvQOy2Gd8+ZhuMWZklvYsYs6359++Q
Bb0Jv7wk4HVrXE6nAW9m9XEa/rvTKvahZu+CF3ESDzqhU2hcCsTzdr73IVBE4xV5XhRqOCX9gXeW
FBMnsyxaRpYM1GKSnZKNlCowdVcNjXTyRKzyr1dqnEu5KdapV4gGYKdYCaNkmOw5PV2+5i1nhARF
rJPY6XQAz8FX8RCxV9b2e7Ox7UHw4eSutADSbVNFX9372qZoP31Pz7oVz0s+ceTUQhonJ640Iu7O
MfbnAWhBgC0joFSYa61aM/Tx3sBO9w60SU1MjK+/4Qt4QaJ77ydsb88gMIunOQH1QIc5sgp9Uuf7
v7gUSJ+BR1/lq0dy8sDOuvbXL/dJxhwwGDuc5jVS7O9hMa5b2AHjah5ES8bQOWd8c2w2LnzY+X+j
FDTcZchMhE7klGfmPe0xVURpWBhhtOAOmRglUCTpgs1WTK2dlizsYlUsmW8nk/mk5eJCL2ekkPUx
KzephRwiF5a1ywRkKuBc+4/84Gr6imPcpDMGAxbXsapyK/XLvdprBmizHXqBXaRIHu04MNspApHj
ygIwCG+AYWVFqteK0yDGyxnkGN9Cd9oxbBwQ31AyIZLmcEzZtE4Y+IK+ND5vilps8erm1mL4tjJN
VqcFgHVpShcb/hxM9V3UC6F9UHFtqvm6pFvrKylks3eF7wh54JKUoTu9OhJo0DxxMG5/W9K0tBIb
3Fme0GkVLI84wWO3G7K+zINhAbsvCN/60xHnwTbB06R7uokBceQGgBv6OvVJgwZLpJsyAnzuniO0
BtJmfjwIgyG+pTxtFzJr7GUF1ziuEV2Cd1lqTKaD8zkCiP4Ly/ErIDQugDMCux+uGhdvXTmXCaW2
em8UxpKjsv9r7Kx6ykyyj+hZwLhr6jxcJhoRfdREADV4kHsP0E7RmS3kNeZ6irZ2RYpFyMfhKA4L
XHZNDA7cNhERzGY12wtdVYreev/JIPG6oYZHchk8WAqt6tP5WxV0PGuH8/+aLjNBodboYJwWI54P
hh5bP8wzWEHbQct1XAPRF/MZky0dZd3LUPBDwTMYcjUTGyBURU9490DPT9hOVn7i8gHOctTj+6PF
adBo3haeUwTmRhGaGzvF4T3m15ISckmsvJRfIrlcWzbH9NH4BM54zHWufGe4pwIzQrmUdVsWo4CL
JJB6Cj1+jC0fjzLJ34shYXegmRb4+2aQjSMWZVyS53Spbg2AiSL38z1B+/TvE+6dNbTL2CymHA8p
/3fcr0wiZ9cZJaD899PLy3O/URBY0/1npxwXZVBUUwAgvOUUk78TPaAQ5gEMq1j7SFX19N6SarO0
0y9L8IgypOttV7WnJDqoZ/nQchGlUxkq+oYqvLS4fipd409F+YWZ2OsCVJ2gjfSpYGgUCN4sml/N
mqyx5lw/retOf5lEHHVEyChSs1/E2KwBReEZxbFuYM0uEuUAYEPCn7GCyNGVZVdq8uLxZ+tA1efY
qN6dAFl551TyhpFHbhLkFKBtsgLC8U2ucaFpTnPhT01y4o0XxVSDBAuQgto584e/RnhuzNrPUBHe
+PHc9INdLtlvYneo8mS4VCxhOJ+MJjW6K14un65gV+HHX3KcTZgdOozh0pIaMqvQ3Ts0IoSoB+uo
WfS4u97LZD+fle4mAllCiAMs5REsNquOEjbWcOcTCme9kWOqNeRUA+aaq5W3m9PtwhxoaF6xSjEx
G+kjXNi4UxrRQqRRkE+RAFWfaOFaW0MZ+56dyrE39oa9bahiyKmemRtMcYTXEHfuN7EyEGnNPYu7
xAifLa7d462yVt3BbgJhannTDoPapDc0SUvdYuoP2V0RQ85zxk+frdowQQNX4EkjWvoDltgyQytx
nlabW+df+GfQ2Gcj/HkdvlpJ1BeIj1S+f8XwxDz/i6w94pdw18pdvTy66PCNVA9ISSA70XWALSG5
IKjFfUiHz5ywnJ2FpwTONbHrJv6ZiUpG/QbkoGFBIrZ1ae5FOQhssJkkELwy0aYojUUUkVyDgEho
JH0tr14PaMSP1//FmT2T8l/DM54zGG5gWwYb4Vf0pH2zeHLRSVOAidW2Fzbjx+V8UkIOTAbI6ndh
wweOMnze49PjSWr6EsKNnNqRQ6jyyjp06FNPSyRwvHjheEWGpjwYSMJVcm4cfJsLpPQqrsPhqAyP
fJtDk9mf3bEdUfrT7C6Sp7EVxLd2AkXmWODQthT3r4fAl37XcCd4cpm0j49U2lAJXJGk3IWz36kU
4EAdlbuiA5KpYcMvjqhHqJfpPzSyeRyPBBxdrxybfJ4x0G8JjQhOA3GQJNIpDkwDQBBqGcO0z4IZ
2NV8cpY4zKCjANlBxd9/eo2Z4nIwy3lV9ZALxFs0qurRBBLw7zGxDS+BV3byoLAl5JpXI2q4bqxM
4xViDzb1Rvk1kErw32oAGmgPkQ+UyDXsbQ7J8W4y5vqTIHrYQICveXSOzCjl7uDSPWJb/blY7qic
z9Qgj+XyGyPO+7W0O0EwK5Ycf+NSnaZ1DprlCIlvhZC+8KmeIEC5eYxTTsNTv3iaG+Z0MGtplqyX
WmQ77cfW9dz632WaxAwmhtF8hAHms9z0nFsV2VVzChH9yEknv7dXFVg2jOz0exsmMwaePKOGNpaD
HTXBR6r8tpcAXu/2SeJDOGHHmCu6WCiCNpBtwIIDKUyj50zNA7Jyk8KX4hlooleYIyK19DAYmFP9
z2ZZXJe+I6Tw2/knO8H3KQnlcECFh6iIbEsqaM99d3LaMH38mqiNhtv/+D9cX4CiIu+H9edJQQeR
SIgH6KvYB482E/+LMnHHUHfvjiKE/OMTHiAKrMFKLe3RZr+z6lduFnaqrsPHL6MhDzJjV5B1yi4L
b3N4pmidqnrRGw1U9hCa7k/2tDindgtRREdpAyqj6Gus6huk0/gnV0fZtImuyXGP3sVJ0TeXG8Mk
Oc9ENYc21AEr7sTUd8fuEV/djUv8032mtv2CJ0+rpqXykIseXKjPhD0+wnbXrMml+8ciggPCzpBA
Cu1vw/4bFEMD6Zb4P/ZOOTlZBrO2XJS3DYHSwgRbSgwW8wBTb+4t5i1kKlPgX7/XkSnMTxY60F8i
mHmXsbF9TzgVAQxVg0tX1Su6MCgHZeVwxHFmujS7ZfL/AXQy4/rprUO7xxtQhIQ8C+kAgIPey5So
PoYaRS0+7UQj+Ux/ZwDk8oyUj60oefEQ5/gA5p87eQluNGXy702fZlZiCVP5S31eCyWSIlqPFEX9
qUHwx/auHMyg/LEyav/A+0ZCCjv+VAP3cwzGTupcfltQmLm3sXF2vEN9U/KRhn+9J+I6czqXrPxP
dxYNeOm9zxXlc7+3IRCPYdN213AF8fU7MvjtoajF56FPDbvHTgS6C8VNXBvciVE0TaASWxp4dhL8
y6vRhcFCidEW1Bx+N3E7SknbfdiST4DwUSvQsbbdnfASI8yrDIuJbFrWmZmsnkLSWVglGCMqj7Hc
gXzmvCK/9507FdLqVh52ey7haguWX+i6Iv+N3ke4zg5veO4QHtNaLvlezTINz9iePeHJs9K7L1Yh
IPhhih0v//qx0jcDCKY0PXaVuWHouumlr7xKezg7V2LYjQgfmV+dG6NLjIrCyk2yfqtp33boILrz
ZZAl0yo+ejcQjQUw7NU//cuJjxOx2OSfCtuXW9KCnAJHSASAypNj4udyvMRCCKgZyQ027oHtNyHy
Fp2ETGpHa66z7aZu4/Gc8lRyyCWvAl/xAu54yETyiqYPz0q/9wIw0BNa6qs5YvnxeEYnrC0UcN2x
/X7cmPeqk4C1YGsg2M5VNYNNoGaqKPtQhz2sPVc4PLVtCGS58WRPUfcO/XILHXcurxzN1jMgRFw1
7T+26iuqxQAon3+h83MUPwiSy1lHX9sstrcLmf0zZ0mI1VJ/rKps62aWEy32eUKGCKF/L7W6U8XD
Fzx31YvgBdacvijGZbekLUPG96tGkqnlaRJGsFEvKUwgk5K8D3a4CAy1LKFkcMb9EuQt7bls4OII
6jY6MPQuLF3WO7vUHkiZiSnbHiBHlhg2/RTxwFxBhxF772VT+9SyEiMo2d4NQ6TKUMil1FFfMZjZ
PUA7BYiIU4pw07iEm5oqw8sCjqhS4tQ8L1SXciSty7JoVS9Ov1NImZX0yF7oJ7nF51lfyKeTIW+f
S6jNrSgdBTbtjp+kiJEWEwhL7JH6IJm0cj9h+CBbzdwna1f0Yr+UaC6J/Om5VG646Be/dpmNklL5
nKab91D/K2tCoKLqyY/hNTADSvKtCn2P5NdQKHHTOTAZGYHspDGc5LhAXse8qMkLw1by5FULI1no
SQkvskLE37ifuW0Cd0iHRXnn0Nlu7c9okkLdRbVh2acb+tPJtVNiuafe5X4ztQPZ57027E2OLiT5
bFQtv9gYdXYfBBpFHk19ydnxsiKsPFStflYuc9teTWoxDvJSDjiIiedcc7VxPrEFU1AG6lkyLave
0oXUsv94PzU34YEBzsT2gmqLieRIKf0nM6GKzFVJdHJ1eCb9Ky18G8eZNW/b+QzT+V+z/CUErdKR
i2haHrMXT2Red7BlkiEv6vFXZGrYHtnBHxbEmTef5oq5vkuhnQdxAYYjhEI0KB6dfDmPcB1N8ehk
djwsiORkaQcTiVTpyb7nHRyxL4DDH2Gz26MAdac3F8/+iEAHVU9S/ZeOgGxbi6wedrbsqp7Q4R+w
WYdXXywYZRaZOQxIYtCFjfyJ1Ny0O4/IlPl+e4HsL9T3Nj0h5lxxZK411Fxv0UQp0pZlCI/4cLR5
JiCBj+nX5n8pbD+hGqMjwgYPonX/H5w1qpGnqTv8oMMnViYTpVNKw15gdGscz3iVvsB2m6ltwqMj
7chzjQM/8yslDZ2GGdva0IufPNY5BtxsPEzADDNGsLb2qF+OwMMqzpSejbLIqY2WM8cRNCWynQ3G
LXiq6laDAZ4VVz5+oB5MQduaZGgm0tKyjNcH3URTWny9QbKISE25yJl8b4xherYOn6EKBBX40gtn
WNSxjy1eP+Vhof5rHCwW4Okoda8X5iO6syCWOUTiEhFH5DfBYjVi9L0ZcfhP7flEIwfGT+GUpBOa
6cOv712rv2grorF0IUePbl7FCHOLhrBkKy82Ygw/Q8E6JfBSmpLQ6nI8FuBGOw1uctHfX5uMGuz9
T63VcH9vgsl4w51sYzF2jcl98F3bD6DS6fKWG5tiak6gp1n18C6wqPL/COpQ+29VMLTy/WUYgGjb
sfnyinxjZNbFst9Ch+SLV+mWs9sRCq2D2LN7aALGMW7ZRkAFun2fXMDMdNX9l6FPWrhI2KPkhvde
TKrKCexm+AKObUHuFbXHMQqopWm5lSxcH2FCft4DVnHIF/+bni4SuMp9G2TuQEZuPwvjSf78tat3
d6DK/KfB/vaVWgcsqkYPf6VrSTD4HIVxK7CBLYVMdiOqkegYVOJkUjv2IopJW95U2UNkmyYkToPM
UcvIEs8uf2WVlLABpPQuGIRkZvhMb0lEpjms9ad74/nQ+L2CHIhNmwzV6w8MnIT85/8x2Utie2yd
HAzj/iBFbzIvNWYpyM1iSr8sM9GDc6dlmMk8nhq6iBoRnLUV1uQCT17zkDd34lHrmD6UqboJ5qGR
rWu8KH5WnbfkahV3lO3q3fiFdgunspU+Xas/sheBDkArveDDti/HpwLqhNTYxOY4cxXehiKKeWRG
KIwx+9u/R82RUR86Xh4y0uDExshwVrpjRXg3dARVJWgZZgE03GkG/afD5FlPiiZVQxrv5eKhFNdq
2L7bVp2PZps9ttZd4fJte324BUt2iRn6+KW6r18yWYCnFy6nkDomqHg/zMbIvONDPe6rUw09GAUY
tUz63hWZJtXvLW6f6Scri9Aw96p5mD3EnQujpD2iZU+n4iDVpT9nlGvV+BkwryQ/Bi046kO5zUKr
Jfl+fHIXxBjGydt9nYRpgkWhCER47r49legAfU4cq1Nu2/RB79IwKEofKT6SbT5rc1vcC9p1KSi9
lz2XMx5iRd2s9B7V7guFPa3Wvz6TdeTasXOiwrNNPEpN25Tk5deZIFBgwgaRcw+/R0DLYwmWOgaM
1WgyYZTPecn4jDWUq9rZBRqhXY5K/3Q/Sq5DpZtHGqkLIMG9N57bAd3V3D0v69PeyE/M3BFxcoGJ
QIgjua2VA5GfU8D5VrYN7lC47Z/EsCI8U0AmrfOuEEtAmNxgw9TlpgJDQgJoshnIscuh/yJn7HlE
CyB0nFs/oiJTbD0AjHdQDYwoZK2DX9G/U/hDSk2sZE+/xMuQt+tyeZybqZqYZ65rbnmTRA/Rflb8
4Gi66Qz3abJCJkQv6dAYEC7b6mQ2tLVbLpDk4SJCopB1JGATjesRPckE8NXokbTnqcCUZt/rLNCn
jd6AQilUO0h+I2BlFVTwoNGr+WeJj+jmAes8AR+KyXCmVwEJYARf3A/EM3mVtR4Ib5lhUr8jwykf
ZKUrb84LMmY/ycEibIF/lSW3rOYsqyBAkbIm7j4QpkNuGSo/td1AFCj7NlbDGErAAZwRl0RMq3Lg
FLIrRfi4dG4Y/5xxgxoqCfmhB2AMYnQy8/H6Yff0SXawdtaKYjBOcKKTYIdopG9hqCGJXVzEO4R/
7zyMdDQKUlwwhtE8+tRNpFvnZwvPHsdPq5lpYCrhJakZ2FFY1pQPaVcIdaP+jyV86dLLEG9CWIcl
SBBON5eGGAtD9mN6GNhyfhRpfhKHEClPGA09ZO+F45nqbBgq5oDR59aZ2ZWmJqDkjM9aAhDl7TRz
4PpwUElxn6HIbcNSI7nI/m1/+eHSIKq8wVVTz9pzJiygkuAsKhXxv4KS6JnnuRKBO9hE1gjg6ve4
X9o+nua+3R1/zolpWNqNniQ3/jW7IRdQpqX5xV4dQKm7EDapGC1e73FUfEf6uyFUU/nOl0MrjyYG
2GQ8JNbNvs0BKOxbAERGahFlaf2InF5zLE8mdBl/y+RKojWwwLX1bFcmXQjBb53cbHywOaM7/2B7
xBW2Hog3KkwuX2tXCw2ZRYYfJOfdpbew2GMnWwDJLMmjmcXUqZRTYRlsdxqmduCj30rXqEYoiuJe
r7jjTKGMaBypYbTsmW4YjPXvTQDMw57dZ2YQJkPn85qza/zOaqRKNt2TDTGGkVhPLp97ZRrqDK4x
xoBOdbAmRZIkROf8tWE4NjvqUokE2Hwq3HsncHM/UkTyeS0eSFoDyP0dFIwT+sc1dRvQCRlADVE2
G9A5DfrEY0GSMysZBC9qR1Qn+dWnZjAbbRfWnL6NhXdZ44lErAdiW21o5zc+qLRIEgI/pbMItVSz
1r8bERgZVEjbRubHm3+P4/Ql6pnuSyUrpG0eaLseVNveUNaQXJldJPu8TancsfTQqr4rufK0Fx4m
HZyJjRjgSdnTxXO5B0PYDqaq3W4F5Vc67u6FZe5HyXGJbb0SWYE6+ChAbeJhoG6tgv6o0uclER++
1G3zf0MqcBU++SFKaf7TnYP66wAq0gq28bpqEuCekKDp8z8qTBBk93i/mMLh6pbyj3m5gUoiggCe
sTTxwrLvYFdzAIs6I5XmZ2FO1WzNhYGTTbBbXbE/LlNwlcN4IXY76CT1dHSnht+J0567gTS/0fIU
p1sWWKl7dBd4W2JRs5jy7JdJU9pEnG1XfdKG7YaobMrlbZPZ2/s5FiFX2/txXIf3yLEaTAHTSysD
jVg0uM26OJBzwsVz10dBvI9n6gyvBck3EKNVKp6xchKgvWYnxk3dtfOpwO0gD5kshmuTuMYZ7YBo
ijurSWJ9Nwsglpxaex7jdeH3xa1BkcfcmMRwC4xNRvT/i50DlV4+Dd/W6hl/QzEcmCSrkTTo+mor
lPXyC1PcNJuvqVBX6u5Cm9ROUBF8oORm20QrDh5Yt62mM2JAhLXccaylDm0EKRtIZEeuY9rL+Hgs
wlIToxmcKpphLhIUs0C0OacSsFQUa6dxaWVgt8B9y3wCPNmVMfeluaBsGUr7r+Gpu9ZIhv0AXyDu
APISs7gBMWeNdwMkT8P9rgwGsnnKf5LW/79YZyrcEWE0njKePzwSKHeSxndebEG3qV2y53KgGZKC
cKg5/dXa3Ly+iCxZLCsR3Jn2S82UWPH43VlbtRZz/WPOgoeOS11fDwSRJpvt6sfcW8flB7KkXTJH
vMf8Wpi/D/lUf9iOOmSK2UFNO2Xlh9EXJ+mOo53Xlm/VA+skRUKQTTbCeEEvByiV7xSaHZ+Py7iu
hAklWH/0sA9re834vIlC2na/YN7a84ZGfq4hoFAUeY9kUcMdf6S5Xs1/6/Kza1NjK1d4dRPp09Ls
L2vToCAsgodENwOEt8L+cqcpzpXRRm+tUNGPrTkT79QnebNnzUDGtcv8HQO70ekA7nDuu9T2lJu+
zdOx2jBAXIt1d4ypem3ZMMQ2tCpr6Qe5Lg/cRi4nYr/1dCwNQLn9/t6LLccP+f5zEsraa0y6ZEuL
Ydo6NXAs8WeD1vPJ/OLw5VfGeBt0zLKNMZIP4avTBl5GjRVtAlp1lJUpk7zX8ufypQo+l8pgfwVw
NFI2SL2o5wOcL4GnpVhhKRmDQdnS+gTpNP9lyb55G67YrPz2FWTpMzzgKVoZPFw6FNHn59XBphr2
V88lgNZxkWbeRWIpQZlJbPOj6v8Lbb6THkqxwsf5Ra+UDCnlf2urN+V+HM5uGxie7YJw8zBakTLA
/G+fRFdE7/Gaj0Q2SrehkIH42RQBSfLiGOEvEc/fss9qYC5BmK+ET4YPKwg+y6HlL/7Cm9FYYSwx
f+c3IMQCgzpyPa5HfgwXrkgzQ2Oply4fCWloL5xON+Qj6KM7gsgFuyX3PwvHTefy9hdaGs6JxMx5
tS7eFOyLcW6SZVQieY/Gpn1cT6J+bKjbH1F9ufGc69V2olWBbiDMq4LZu45IMrOZ4zqJwbWR7gP/
mY3srBvo8JG2lhZzmPqsJgBNlSNwOHbZiR+hAQUQ0LkLxVdlLd4P/g886JbTJ+Q7cnqJxHecfG6+
THH7FFjgtv8QUlfSu7NSdBQFMGU90Y5ibMIlWNuvwLJWvGSOukLkycjMtsHL+fB4ek+1I1rRmm5H
CDcV9iPMDn+KvMTDbxG7ezlVSXXgbWTcHfMPyQ3NL4ZUOxBuiwnGbo1xoxkBuWOLMwMqhWZBrMgU
Gi/31f1hbWScQkLvAXbHpRW+/7AESIl1VO4TeMPupsUxfTN78hvW5+JSYeSWj6BKUF8j8LdH3MRy
VJiMafsK+5WZJBRw4hCaxq0iYLos0su5fNcUEE9McjlqPXgk0IR3aoSIG7sWh2Ca3DS0zSY9KWgx
uaK3zYZhFSZT6YJEwC/pVQLFHjB39mo7+RxUsxSBhf2WT9huZ12jhWAnSuaXw+gslas4x4k5WOR5
UeS0zkeesG49hxtpPAzbuYEUlCFcMWkO0l1u4urp/hkIrbjIMDe58LLXbF8u3PzFkOczcl+44bQC
n+oKn1TD1qIJKOxH6AjT75sU4WszX7S8LuKInGav70LYcH05HTFpVf2Nb3pTPmMNe3+E86E/Jetx
MlRnRIqtW2NerymVuAxTcWF2A2eL2Vs86fHL78Okn06BipYTncrn9FJgVBnr6KILmtlKer3dW6Fc
vElu2h6shRigjg6Rz6PoNremtwy93LTRxT7eMgDYSGVLwAQ0pqzYbNs0KC59Uuof+XeJNn+ccC+E
Yze6XB/+yWbTKzL3mwcO7ZZAFGDHHsP8D3rHcBC0/welmlEEf2N6uhDhKk7wj6ABOt1SdpUy11zK
gjBQzfk155oFFvOnZU0+MF+vRIQXIosiNz5Obn7uxqPorh03s90YBlIItzKD+M/bI38tSxhA7sOY
P7W7T3G4DAmNeQu7xILXGDmKSlEz4Mmbo1Z227saNnNJn6HlF/xl2rihjoXf5f5PbiF86onIfKqT
ca1lyU5O8IRW860mXLjVPIklHJZztLi0fwD2ghUvUh2ooaklvgqrR3ZB+l+ffYzepYUTXhbZ2n8k
9oBlradKCGdmo6zbqERZcuLqhTYegf+PH300ZdTG3O7Xh77MxSJtA6v5Q8vew8JUp4gu9MpCgUZq
RhWGPEx4KDOaDnApZz9gz7rDkt4S3/LODn2ai33P2SQvR4QOBt4s+VKOcgXBBFGXjeX4Qo+uu5H8
SqKO1iZussiVwhXcyPauDPUq76BrpXyh7xjtx9NE7cU1BLOyXHZisYLgW1bhdGIKKdpCGL+th0ie
x4L1JlC6WE6aqHS/bIRwhR2XAWWGiOmij+VrL7Jqgc52Hq0l+Zr3p7+wCAcXOyoL7vI/KUMOUubm
FlFXG1QOMTfdXkBOMyeRIAvfo4DwpmxtvxGgz81ankbGmVQpDrjxz6FnWfvaDFvh1/1QBXjaKKKh
9MCgHHMQBEyIYp8sPbjFnY2FqcVGCamHCCTFwggj49ngfvVpdDPthmVKJ8QReGmY1qlCYIyIFcu3
9Yc45z4rPa9ej+uiHDpmjKxyJj7dy8AUlfjkBxhQfU4+s0+AZRZE1R/RcYhmgr7dlHg1ECoyqoeU
U5qH4LbxhjYOIMsx7/MKeQQsf4xtGa0rQFurSUbp68/RcIKynj15TzJujteMC/J1lwLAUckwM8xn
gcmoyRc1349Kz2Li1tdfH+loQI/A/PwhYKtdVxJLkeWDoHrXqHPlrW/ja1lW3zS07zre5tloiWLk
SMY7oK5qgKZoYAHrFJLkhsTSuKmjx4WV9w+AF5RDXirxBHHfvkhBxquEfqxZCREbsEUd87GVNFd9
pu87NFdYtbb9RzKVpvClEmbXk1idU7/RxdsutAjMBgxdC/SBPNYX+LshpKCSAfAJuWHTv4l9kHpL
GuAX+Z8zTkam3n7psvZCAOTKJDqcOHEPm4+HElDeblnnPluPQ26azAobD0M5XfOtDBr777ygbx/q
P1VpGEz6lhScP9x3E7zWNydVe5FHs/mKR+ENPXk0lSeGT4rS6PG0RBFGtqB7qv1KUuh0HZEKEz2V
7jXsaj472WChZymuEG5DBmpQQ/tCBAJbtMkxnvWPjZY3TtG/DN/i0xwImhRAwUV4ROghcl0p/AI0
LWaiXOhbEJ0Pq3GPAYzbQVJwgTmUf2EfCAajizJgFhvBdDIWrd24Z70Iw3BCaPj5YXXKe6853Sbp
ntPwphHp1IRDwog/WErSHj8asi0qv81HAM6OmcR0k5XZEAwgtBXeMslmVTMouRK4H7NLLkuPp55T
rfIaVKh2Ljl1KQEGr/nEsvqCYHDq0bj4U5Js70SVVQ1aErx8v9aHQKEqw9jSPRF5023303/EzPRp
Yl+aCiENzeMddr8XypCOzH0nO7BQUCjuvWj57srKcdjaR2JS8K4pF9NYV4I1+5anAX2rW2CH3vQN
F1PT/X1eF5IF7lCxO3vqUK87mYOAs1tlvELOnWWLVtVpDvgLUqvrc2C4tCaZcptq4m0ptHDSkgkI
lBQtaH/t9Y+9WBn7vRm7W/JEOmsSzU33dzn4dh+phBh1wAItxaFOJ5HM9GGyxYOTpBQ/D1TYfrWs
xb5GljYpSyDpTeezNGZjN2KvHYNZbBHw99L0SKPMtrJYmA6F1DuITLWR0GgUKhPJcUoatg+hXJTi
A1GTaCNw1ooT69KvgaQWAZ99vtq1Ngzgh0gw2Qv+Th4lmO6d/lFOTV21v2a+65bVDVqggiuHHwds
/Bu1XMoQjzss5WbZ7yl9bVnDUWPmXW9VnruP2v4sjd43cHadcEnf5L3DwbYpzfK0V2DWVlIqPY1w
e15YJY4JeeGzVVqjXZgKxR1NYw9OljArNDEbRma/Kf+uEbq6XMOZq8s+kPtHK23jjHxgGuv1WZ2Q
BwOLE5JHiNMiKrih3lHvx/JrojnUrZOfEDa2zZ/ZvUp6DyelyUN0fa2hR6Q2gZAQPnBU3tyjPP77
W/WIYV4o1sTXnAqXpVZOOdklC2fVXiSsNe32hcRf76xJpG7qLAMDK/tXxXXqhOTGAnTI8Mqsd11C
ZspMvLiqhui8zZEinZMuy9vPteombd2tJ5/JLLjfaedu1twBSpsDu6KIEx9ge+CMDmjKoQED0JIL
U73+HIPGxjcZoKxiNirWlZyjXevBB7tn5mQur6kD1pyTRMnwX74J1V3QE2pbBerW9BDeCoJQaZsE
z0py2cYcjnAjHEMQeGmJ6zurWD3q/X/2GNmYUwB01bCG+GWKEZ9qR26bXSRhOH4/5C5BAHq68zDJ
20d4bCTWP1ww7zaNd1rqc0QVgVU/AQToAc/XRCGcGOuTzVqQGMD73DwhASLeKHWE+u/QZF71hZpV
u+hwuMOK11eKpIiEjUuAN27+AQHVgSf0sAHFeSkpTATDy2cUExMqr/UMKEG+8hRHiy8FxbKnMXEn
6QZtyIz7CDb4ELKo8VGZamgpIe6y/qwuatpZQ7qwANzHB4U4G2SgcZHTH5lGBT055qyZ6Y9ORbby
YGyv7tvUOfPUCg/AkwuqeJshjtLYtvFj/2baV6Ab2KZnh78tXPbeHTLotRlnMPNLPwD3Tlc5/dgb
H1O4On2Clt6k7V60zG/VCDmM/ZAkcdCEad/Ktz/LEgayixJwONro1J7MlfNHOt6X7ydxSGu0p4jV
EIDzkG6yycf3dZdWbReS6TG00ujmQkLAv7MhHaXIb6C2K7QTzZtu0klAgAKemxiKkDulEbe0WbJJ
WrkR4tN89F8gjDVvSwE80RAMoJewsIbF4RY/ODYgr0Uf8lrjV2ozp8o1khfYxx9fezLCT+IEh/P0
DC4ZataA8s/DVUkcvDpxLpIadIrz8mmnBt6IqxckmNcH7g8ouOued3NMzGOsHRzH6Gaq1rQfqXlK
AnCYkzQw41e/ytyaXx+4oojqMtQrAua61JGqGt/sWidBx1TgD5cBQMRRZmm1TdTSZYzXmejImFco
IZyt4XwkTqez0dpQFH10g+c/wrxTWKHdMEnbMCbrfntwZ2RGVMXg6sZ/oudtG3AjsR8gZWw3FxzN
vvx+JuAawzIIT1GWqMiGYwcoCce6aKGfRQFLvKFhSDg4H1MzUtIEeut3Sgvx+CLexCPLBc+OYzyU
SHaw1kLq0gvo4PSFZzwbzKEF5aCIXoNfOYbKBgOC/DQN1jRdPe38XwBfl1biW6Xt3OJMQSeJ5n7n
AJUdtdwNoV83xASS9Nk7ohtzuEg5BcWcDRQhx87o5+I0IYdXpDBYGIDXFeXMvWf/MTyDqrhkLZHt
pS12glavLbZkk7qUrTo/S87b2wlIBfmbhkYv0TYB9LwU13ul4J0M9c8mMmr9PommbfTj2KMGnaWB
qC719crPWS8DVXyYltu1oj0dVU+N+s61HXJq/Se0rC/prG6jlh8VfHvsGE9t4Om8a7O2M3Iqlv42
yUjeAdbSSdsKsuX6fom82bzRgxyHLjdBpjQBFZKIFr4mq54BL/3okC+gt0kPlWrbXrBVpWcR+0m5
UxJpeQRjNJZh8+l86RpqqSizTJde/mMh+qO7LWbtzNgAzjtSrXwpUMYLariB1lGTiNRd77QPCRrm
9wqYZ9el+W7xiObWYt0IMzKYz6u3+4SKgjiAIVpo3MSm9OMo67tpviYJGJhzA8QIB1kyMd4AtbLs
ojkM+1ENtWKtVwFOv5cQHiRO2Mr1u3W489vtOYXdnm3/DK9TG7eP3ZC3aUwc+irhDspxr9oETak8
gGzrVZnYKUBBvY2fVBcrCQO3T/qJdTGGfVZrznqTi714Qz4ng2JYhiAyuzsPPKiibOMkJqrSGsxM
ELy35f0cLa3BrqmqsuSX+J7tqaKlrh5DXRROSsMV4xHw7PxqUiM2SYB6qJ2XzrBGRGDVQFORRC3P
DExyZWlV78x8EAIoD3c8C7rodMu4Yg75EYEuvsgHcSkaY3PszR5bn+co62ig4tlrRIlBvsffz8Wo
NvbTA3tAKv+r5WSjYZoAU1W1LKVjsrrtrxMuGCy2JP3ygVhbxvf07cZd/aghFR6xlqrK0D3EnQa5
eizbLaogdvcnCmcVmI8kmlwdUk/mYfhMtslrzQj3nR/85Eas5r7h8nGyGtYD0wx5KmiArldHFtZh
XLBF/u488+AT6SZm0BOK/tTt6amosp76OB/tMNf8ueA2xP3c9QjYaevClyK2HsKjcnbCB1Lg+xMy
Qq4ij4zqiks/K6PfLIYgoZeeRFjMGwPl2M7CPY5OUx6KJVcUIuWOcqnSROJwSwS1vWJLQdbt9JIr
BiotGYw0/hD80+5kCtf9tlvVRzvFtnBz+osxQMPB+WCbxVlpnt1BwxKpjSJ7REvY2tC6silx/0x5
Apt65mtL8B0F7TXW0dOGEK0+Ud3Ge84UljUz5JcFDqaE9Z5+fDp0Y8cGXi+hJjr0C44aL3pOxrXV
Iv/Z3D/4cx01ytvrS3PXIQXDRepgQHLXEnHeVtq1jHVprFywmRkhBjdzw5yyI8s8XMgcgRmtOQ1P
p/3YAJOyrmW3VpekUPj0hzpLflVPFRkvtdxsqytFxVS8mJ+oH9oThCDXdMcWp4wyzhFvcOmEhwCM
elISwi3e26CJ6B+TiqRZG7P6K5XKv7esaGdqnFcunF2GqtMFI3N4hi+u4J/FqEhcmONoXNiPrHGQ
cXOIQIn2VQwxPDl7UzZf9pVXx9sZEByhGwKWSlJc9AfyAI7ZlUUlKhDoMJKkoySk8FSp806mqFoQ
7VtGrD14aLMrHFU/xx3WORJAZp/1Vixe12qItClvpN3S01k0ErknTtTWamsPDTP/hSUb7okK6+Li
woMTKpwbEhy929dNIV693QIWilX+oL20J7TPoNDfB15UZBvitUIsHneoMjCGyexqfmyWPX5jrdpr
HQ8Cw01W1/wYkng30slZ/r0lpStKOVpEHcAj2x9bx4/QundO9HhpytMChzzDnkRXehu53inteWib
kX7sb16WN27KKigX8nyvdo1Srmp81h2BWHqgMG+t1AkC7JL6fvD5C2pSJif1OF7UktCWZAN360ji
aEr9AvIxG4BB01dmJgm1RIbaF0RGJUsFgKll7uTlnYqcMwWYHpQtp3F6uPammHYmZN/bVK40T97v
yRycden1EFXR63CW+kDwvjZ3cg2P2ThBgXGBh4njvN9hU1yCSUHmbBRj6UXm+5iJuYuyQHzDqksG
DSMVMeQUfi7wH9El7aE8ZdcZYZgHxyG1xCI1viaV+o8QJPV3vBFNrjHOD1SW1F/L1TnFT+aI7pZJ
AcdnEZLROzjLIYsxXIEp6gu320gIgnJYl9qYDjjqDvvi74ERLcimsmGsImfgp8vKb3k2ZZQW+9/O
WxDJAsYsE5MRXKWmKyGyEpj+m2dlfTg8sMC9b6pGvkOnT5nfzKsgEYQBw0KUL/fSY75jIw+CgGWk
PNNInxDrsZObaM7MJhuh2lV76vJ5J7hVA++JbiA22gP/kKp1tjXoKCTKHt1KFW40zF7fFtif9ufW
oMuTSQyZOB93+NN5PTsFQ8yG7pZhfgLVNmzNmpd0DArAZaI1yofPDbLtAhx7LqXPZwrjipU4Ayb5
im1heUu7mSlyfCNDAkB3yiD24Rywxxp+r5/S47jBcYpuZY2cmRRoWPSpBC1Qp/bN/eArK1uBbUwr
kbJhv4iKBxsHW+7upm28m9FhnJ4OzM99KK8sSJVJMrgi2i0b1mSVb0byJzog3dlLliruNA0aEFd9
OQ5ZoH0nm+fyazf38sxf099jeOKav5HU6xuY/JtkwKgV120/XccCCHLhrcVT/4cIxJaKLTXcKQty
xIjNeA020I8RNGXMpjmCUzlplfhrOJXXe2yXTcvHBBQqc9Rmuj6eaLcnwcK3eQmp3Us20j7ndP5K
+agGIM02Gi0Z6GAWwsB0a5aFDt9dfuQa2XnuafZnIU8orKdbtDZFypWcV5tFJ12G72KgTaRGh/Mg
V8b2yEMbTKBDU4q9s6cwZL9e1KF83tXq0BypV2gF100KBmZ0BP/qLCGrNhSiLBTXY0yMyZ8s2DCb
3FYPM6o4n/JH47J5OOeND9dSeMHD4R6z0iI66oGVb/vXtJHZU+qX8QpeXSrZnnwDqBFHYrBRh+on
ATrvo+L3fspby2+hW/E8Bv4Nfq7j/aaciNfupM4fRlwY9pPsKSOb1i2Ru88bIvJJxX2I5ijdO9kK
z21lgbOpnvuFtmBt3keBRw1ppjwtK6BkSUeOzZwebdOlkJB9Xx8fEytvwIlHyKkuhRpYxC8xFWL+
mo883g7IbAt/3Ls8UUUahkAaJldKRgWnOsboockaNgWN1olxPrbIVWkYiDDE1jTkvkMS3GrhM/LL
j9ATlYNHgDujt9j2PptKysauQVZ2ki2KppMNWOPOhXMfD8AnoF3SSCq/+9srfgewtmHV0Srrxg1l
zgMCNxcFnMXfknZGpAaWA9rWax45QIpo990zTZOJ3g6jIoMMWKlwYYunNQgbs7WNGr1znrCRqm/a
MxAcsjBjbaWA+Ma/moYJXVTGPPiQ+o3G5/e5Ff0gUVbvj3Ohv1bFmdu1gA7BkCFNd0oGee+dhWhv
rUTo/y/b6w4tuT+5SnSwcokNv5OgUF76QjMbszGkMdPKBBwiNAmwnCwXx22U7gx9e/VA0htMnZlH
35plkHCdHCTMSlJ6WhmrN3XoJtOwLjlk9zkS1cYNvBOxtaPRQRCu/5fx5OMMdfqjHHgUAUf88NE9
Q1lp50oSo0hQU15NTULP9lDe4dX5CL49uQnpwBx14PJyb6f7e0wYKWjf3TmNLPjXbRUzAwVtGuAz
CyUT5YvqN4eugIzHC5puU2TxV0MZ7pUySlcTro/0YzrFYOtGWjheCLGtkSJ/A3QSjV9b+U3D2FbP
TnzTvAzgFXmvIGPWV5JETXMnAJLhYbrOESoqiJUcn9klLshPLkhkOMuCBsU0OKM9r7YbjW1WbFTt
3JkI5TfKZwtI2o1ZtBNxWWmff7ba/Wn0NRWY42K0kWxG5xLJemMGRQiaCpGUb8Bvf0o6LvgK6MIZ
xZQ/rIyQYEnipCZ+fh4sQGFdan7KozLNEtfxvOtkJ+DLyCbuAQwQOZlZpZpsnHb40teudtwwdHS0
TEhvJpDtZayxVUuHynFvklAJuo/2XbSpUSOm3NyMT89xYzOk5fkfYgFVk1H26j8Kc3lnakhNoec5
3+v5Yw33NcAu/w0MxwfTZH8dGmM4HI7GXkHh7NvUffNOkzCKDssMSmgLpcUgix/vXP6pXMNCRLll
kK9Ljfz359yCTbm1XS78HIJYy7xFAaQxPfh/ktVd3JGjubeAkL5GFO+fnS6K3KITmcund3ZQuY6Q
24xV4vKUocFEQgdXiErmZf2lkbttPs/4pkYX/TM5AN+kDbaFyKFCXVY4CPhafYtGsvNwaWhA4jfx
hGSl2zyu/q6TX5yhFFQQ3AITKXz90jPuXcg53OBLpRr6mb5ZEB9MU6QkLlj1hQotfe3JX94cKkm1
Le7il1FyF2wXUFSIB2Ua7hwlyWjQSt5NpqxKRA0ct8mpfFPH+Ar6cZa2LgAVDz4Tatxk2L+iuzl5
zkE9GSovuSKAoGSCkwtGfFxcCwenF0t1rKfyw72MjLvRVWrw7WB2CL6YUGCyIy6plhdzmRJG8pz1
DkzQ4ze/HjI40pKaPr2X6eiiV0m1YRJqOTkrpfGPis9FguM4z86YO3emoaPJ82F6qeVplDUX56w4
nFJkSAdfHtKT3vUXO7b9nuiN86Z6CUf+oaWp/UDVkgLMKa5fx6QIO0ot5GVp8F7f66qM/tN0xYbB
SqU0CVrZ1YhiSILJX/dtUaLB7hZ7BbPJfIJeIzkclNV5kDKzmiKwG+aoQfpMeHjCqLFQwRBAMeQp
+P5dabkw6Gk6wLIVFEfJWa22a9iJ33KYKv/OtR6i2TRKndqQdm6+iE+Hc4Sxt2KvstAQXD21LJ6I
tnD6PVp+DCltFrm5xcvqdV+MUtuqMz5kGpTgej9lNOKLqgYTjvG0LLVCSiR4b25C3Twi2F2bp3DM
rinLCgJ1cm0eswmwXQSGSs5Z1/71jornvjmz/D9T/fP/ABpIJr+CRizyCUPgTMv7l+zcq3bRiAHQ
PypSoBkLPANb0gQ7dnCHRVwfxi/9ibM2/WWkD0AZJ1lJkoqPWiAqUEozT1brukd07Ox3VBVjR0qt
7txgnCwlSccgqwA3PXt0FpwoXbxBvOKVHet94pRyKS/xmkrT+zgEAG3mAvN/ltWc/RnPOnwviI1z
iq7T6maRzfX2S6Ph7e6l36S2+7emOl+0B4e9bkKZy4LRlm2Qe6vqSnlCDkV2ZWgFeOPYWJGNCBs/
RYVpki9Ii7NxSxBKmMJNPuaIXHUe2hf8PSqzIf+iIUUFXzcqsCkCXtnWOycIwrdKKvAB5SRLssrV
c00bEtelD8H1xd0VUV47d57MO0ILndUuRfoAPpKpuVXr9Y0QXxwLa3qeU29ie82Dt41JxKKkObNH
Cu4eU14mmH4GnDGfAlouFnFYiBeDFj7AailtV8vLDALC4YahTHHqPTzWG5i+BugzOWgD/oVcfVmg
nl1seMd+CmtWQzy9HwuXHIfwBIKjsSuYItSecUY5edPUlaITKrikIHCzFXRwytnNm/NsbEIBxcvT
ijyRxVFSaLREwtExRn9CKx6aVAf/5dqU6Q4UIgaGGdYPc/PsVeveKGWcw7Ebw8I5/OZRlyJt6JEN
O2wmlkuWcpyUfO8y0BsZeSzMY8fujAc5bajBlmZd1r3moCL/JbbJHLME/QBlvAZFFkmWBtOrqcZ5
Z/ZQyirrT054Fjs/umHW7q1s0E/ZaxBsuUs7BavJbuPvniYaD9Aj/1jxn/ZrEPk2xYg9Cez+/oOS
jPhx0LX3djUvEOdPNNld69Oww9zE8KjpEWVjG2IRIJrbG5knSeqHLd3nsXPshvGenjEIAnErXT53
LDoBczQtSlFpVEB1O5JqUG41oXnhHcqyy6//uaFT/zqPyozL84XRhOB7xkuebUdvsJiF4jigPg9J
wNsxE80JzZMfbISCCjSvQkANRhdcNPJ3cTrzKr+YFMZ5GAJN698EZ99ZJETc2LMTd873Lv03LHCW
eheH9P43AGpZzk1pMpWkwmXZ3SzmThKyM8s0Y++2D++oHmj0mKijUcOGRQE7dkVRKzlH+PfEMmv3
Gj/l+Nr/3k+YubCbvESDV8ip1q1babV97c4Xw7aMlQ8t2QcjtUwtdyFBo7y6ZzmTzWd0xgAEL4nR
4nhVPROfHs/F9m7I0aIeJdV1X/3XktBRAeEcRBw4f7EdjA6Xu53tVHr9EvRhHjVYP9rjJ8uJWRhy
793YBe+qNpp4OOkEE8hTi3CacLuTIBjtC37kUafQPR6extgpHyp0kfSeF9tiL94Aqq4AnWUzl2PZ
K+zNArG2l6zfNYrrCFWBxBUEsjCxM0HGybnL1/M5xSTNN6r6jAeS2MdQi3Ah2tbED1deTHR/8X19
0XE/SnChKIkGSSxTY/sfbRSU4RRmkAyD6iL4K4hNLo/7+m7GJdQxhNjvQ78+PzJ97E4Kj678sOon
dr+giyEmcJmv72FEkinvgyju2fn+3RotioKeff6wjfkRInS+9UKOhfb+89ZG/stW4i2Lagw/BCJY
QUj7KxrbvJ5bQ9UjVrbVuJubLkqrN/QBmnc+v1yYhhaXknJem12PewBqc8krHaofxUVOfk21dG5S
AsEK0YjwkGOIdN2O9gp9qUKX11l9VsOcsj6QY5gf8pTLdpYr47iOHK4TEnGlSQVzX4l2Us0po5kr
OSDZk+vmCIDYrbzMnfrA9r3psraQpYErfBHO8RWC2cFgn5ml4EbW13Bex28HPIc04SrRe5joHuCV
6bVH3NKxYBaAn+XbLFQMMauiZTi6v9o2XnbLmGWGLZRoNenQ2/OO+HdK+/debp9U0EjunaPz5yHF
BQYd3BB09lFkn/3RBgGnaCMSZTNzsG7WI4jMt1tY4Uoa8EwUEIEijSOjJfKcTkIUMzSJ9bvtQDW2
hMXNTXYO7Q4TahaUMusIcocBf713Sa56EN2QfKVG/zkRSXEU2vA1SdyfumeDasEfeRhBZpQdVoag
8ukC8Yc0gpvhxcmnJWNaIHCRc8sYsbEKdg0D7HZ9y5xMjA2DbS/2r9YczFaTCpXZgVGPJMEIgVM7
NdHXy5tr8cHVhtfKJX6gcUA/ZHWHsfHoIYi4R2uJiVMlFaaOWFgH03uOUooxlS0fPJstlLEKTedk
PVHDFCNHY7+2kAEpoqJ3GNNSgRCl6KsRdz8fVtZrUwsaKM5h5Xtr6co15k/Z+ZsczhVB8mQjzUAv
KD06LhArMgnXiuUM4Sy/KhgrMmaIJpASA+BfDeBtvEeFAnIenkLzCOVeWtvZu+IeAVHI+ShBCxpx
5+VKWahpL7aKyHkWQJm/ygbkkqy3zY35N/5qlZDKYKQi9XJr3ChtbHIAGWU6LvXC1M1sGGYCedET
9NFMqers1wkyBlnGgspGmptlztK2THVIXg+gVxcTUgG+fWTZ/zGxiJUBE9SdrgVrlbrrQyqot+HV
BRJc3HiQD0KXNMMiD0tjMJxICCeUhnIDpOOfn2g5GIA/hGZZkHRclBStzBty1LP25+0uI4j2khuZ
PDI7FiPBZ/REqo/oqWfa0UHYV9vMsuRvlO1P+KTtm3l6arglJs54TOygsunE/fp4yQotZm6ZGgNl
pEzOoESmZfED3x90N2dhVDNgqKlIb7z9GcYKY+rYuN82kLLoLgH3754nV3FmzhwN9jhvPZ2z1Ati
c7+eNxQ4oBfvGMVdAwOkywXa9Y0Jkbyl9Y3kS9kCWhGhNVAwREGcIzx+d52QNoOYRcebNLi4Eo2I
itmEvmq+jLk3aIEJEV9Kynew5V9OXyPvlaf50RQFGQzuMx1Vk1YnP/YLisn7lvZLcurhPsmGAE4L
GjaiZe9N1hvwua06qkTi1MNg6Zl89ekKsTjFhhHKKIZ7/olf3udhkOjcV1yhIHu3pRW7bTW1+EV0
wnVkeOx7dgy4RwsEkSxrDXNVBiaGaZaoryLAvWK1Rra2EgcYloJyk8MYjrt9Bz7MMQ4yY4aDOqHW
a4GR4waqBo9J5v6pV1ixV+U=
%%% protect end_protected
