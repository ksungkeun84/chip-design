%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
As+6sq0UwmScPswU1JrQWLLW8hNOhQh2cnKyiPBwCQKU4EAfc8kkMZBJ0IRa7+n3xWMKqUB45iw/
aYrZjju6m1wtY8y9CRLYhlM4x2GzmK4e5QpV4u/hL1CWlsgmox7pS58k4tHtrSDkcwYEXKqq/kcb
EplYmCdzMC/+yNWkPANf+Xo6A25DPt2jxeWHNOOHrIS63l8qV6OfahwyMN19zwZ2aIXFRS6ojWQk
d4wvh1QThO+5gbJ31jHGBujhn5oJ4iyrQM7ji1k4Pqk/947WQleTuTE4x9GyLaRjHdfjU1Xly9hH
0t9R9BdcYr4UAxG+G5EMGULIMxumGy7R3v+7TQ==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
Mu/djnJQuq2SG/qalcYbIgjNpN7t3jxupCGgY66EqbbNvczHIKe8ikWREMoN9JJiGczGwpJXEG64
AAatVFHcJM17c00FT73yziqsnSPdjnYrP8n2vc9LcUdEAMPDDCawUkZ5B5HI63wTJPRGezbXCvuM
6hGgX6vPjB2vJIZ27jxnF8tacKcXLcpnPZj/yR6NKF3zuLBjPXk4vwjnbIArCD4esRL4t+wz2f6v
UyMJ4H5GNVlELcVrEs/JJTMYgyrhyweCD7U6qIRuB6NB46EMTJCb0IuPW810tIsuG8sGehf7IJHe
iPoEbeFoow31QrkclpH8g2Lf7YkeOH3VR7eZ5HtRm9HMdu4xJqcLxI5AeKb3CNfmYmN93JLzlkg4
aVEezN5dj3X3I377wJZs05LmERinjERhXzv7+rJnSIt0TniPFsfjggeyO/melN57ASLTtcZHtHrl
ytEgpk5dGQvoMCaOOM7YUc80QoB2M5Af/7wCDLwIQuHVJW66DUVKBC/X+xD58W83bbIBeNaNV8j/
YbCEogTczf0HvRKCPhQJPySN1YWH7aUnQ6McOq2THCLEP0neBboYiunCB7kBZifWj1EoBupbO5aH
ZKKvQJ3FuiTExMa4ab0k1VqbUTMvoRCws1xwcau5kSLj6D52CEgFd+B3v4frFePrhB4VZLArd8ON
u53pSQ3XiWdgVL6Mjrtq7mPF6PyrZ1oLp7vQXVd/y67QoSc0NZUbLJzkarfpRzPr84hOHYOownE7
+SLem/KhWwD6a1CTZNfsV7uLbOUAAFkUaH+K/v59MDChskUeolOoPRHODZvrrWQYZ5r7TI/xOfw6
UWDkBlmWfiT6MkQXYlDWrG4dIAwqcAX8ZxaZkBsL7sTn126QtD1Ri4hf+lm8PbtZ8dYuu68q760E
7D1xe2gn9p4nYCJtUNHSu3YQ2d4Corl4hhwy6Jtxl255HU5WinfT9Le7SbGxQXrOSPev/OnViE12
4OvkPtpljK6aK9hvbLDdhIH/dkyfI9hzFx4ansJaT6XmcyNUcw96lSpKq6qUywerEWiQnGmx2yYb
3rjJohBChLKr9Gak+M9ExLfoJSnksA0aLbAwE5dSpaibgSUvEjlEdiJhy8Brj6/J25EZHmGcj7QE
vxqTqB5mSc9q8/Vg7G3F09ja46xhbkrD63+JGQe3MeSLUdI4ZOQhDxDUEBL+NJSLtDoekqnOH6w2
7A7/JkIo/Fau+GuOBQhA9v9XzyVlfYRvcV3A5ZzGtSWPZ53COPaR7Prhq8i+QcEbr3SZW6UTrE+l
6W8j2unNe3iVjCHVR3edz10URK751EC3oGuNES5V/atspaG7TOCHmhuOFBGwBncPhj1IjYFNXsEe
gJR4YFj/JZtDVPKUKu4fwU2U44nzsEcpmlPqXEImxcG7VWNTZ8hM77jFNEHrSi0+gkNcecYwKZnO
87ix7ACCpplzv3k6bR2onUvEzKkUSezX2wsfajnkv4rc4Zp0o5mgG0ZL2Xz150bxdteVrQAHEw9J
0D6q1nn1Z7AdzJAaASSsG3/0EiEGc9adShS/+Yhxdz6WJUOOwgluNjvBxuql0rDySyDsnkKrRagT
DK1T3vDP7hNLPbE+9xRGSme+gCVHW3CeWdP5S9rqfRKVAfyADfigfRkpTEHFZEGonFsAdqX2/9z5
HQo9thpKhqVNLKqD5X5I1IHHfIFRrfDy6FyQGvRnKqi3RWrGzvz7YITuTkXMgKEYP9ILWjvBmjd1
TDYkaTeNf2v9YClcrj6+JyA+GQhU564jVbZ6igBgyJk2nzu8Ib7DJOQ6ySsdzij3fbfIM744VOf0
cjeT2e5JHQ29PX8B7/JS7l9SrA7IDrQ7au8pW1mbDlHLOVA3BA0tlbIPIwTx7yH1eJ5JBZ4hfST5
gskdpQUuLZaFjkQghTwY2PUVofEwymfYHO/m/kITDUVcgcr6fwVpY7+vJPHqS4bGMpei6SqVGRX5
ZgrQcLU478rHmU3oFAcno1nuTyk/pOfNXAtg9XK3j1ter4A9LGAKEbNTuOwkoYbIGfJmeMRBtlJi
6aEuRoVkBemn81sodp/isdqQKlg4qXJgXYmC3tQQvCc2AMWtzoSPDyII4fO7yyx5NZplAPSs0kQZ
+pYurCoIMz4aydGqsMs5++wcuglc/ko76PzCJ4YuMJOarJkaeVMsyayZgDEDe4B6+YJbIQa/D9SI
t82LkNzWd1+KC4t6zdWueQpDQHCMnrkLAPiRxUXBzbm36lhyIf/uJrm0yhltJ9R05h45KvtYV5yV
bsZbP+QnMURDCcjf/QQPbkhLpvGAfBvhOfsOWBtmoPL9qcTHwr9R74e6JKOM8kF4N+Scfj20e2U4
Bxhz3mpIzxcWt7Wf2sxLvrpmIZhcqhBsk6S0lWurAf98eHwrG/9P2xL6j4kVsx6KKs1vbPCROOv9
J1DXWNpY6mb4ODsuFkxp5I+advo8CBaGGYHutt2IxAwe8irEOyoQ2/GR8GXNQ5GbFMuOIo9WNNsk
c5WKpjpMDPHVZAVArpPaXcjHPEYJ8GKXPSiZctxpVVVOsgEv8NIlFthA3c0rrAneEKFFuCCN29Vw
5pYn0Pj/KC3BI9WrtJFSQs4Gcvkw3LijQNBvNEOK3EZEbrVKMIyxdOEupOmNVY0l91UjQPh3OCfP
c7igu07rSiUP5fGofDpZbp5kW5Osic9dAuTqkXEissDLwqohVixLVlGTbtKX0O/yGqBu6Kc23xHT
lhAAzNjxa7IcxvUbyrSeEa6Iai6pelyCao/4tRdVcj4Y4rH3IuxulnKYyrHJue+S63AzlWSFFQYZ
trj2Os+zzyVMIMAxt0cvO4/u+UcNSvirAxC2mnp6AU7oNC31Z6CvFoJT9ZLRd6YpOzHmuUeZuWYz
JtS4Wl/WU+euPDwP8JOwmC3igYSQq3kD3kBxF2rnUXINRETdXx5XKp5KLoAJVPCmybwHrhrJigRJ
so3AwcQvlEAqYfsIHBRyooFWkK9xIfEYOWBpMs5MBzBUUlV57ObLJH5Ruo2XwvIkK0rCQvn6Bwjf
toJUSyd9cT67WriOKVyAGYmit4BTDU8gQaXTEWYaEz/hNS+LT1K9b4ZtqivrLiQYAHdNa0liOZnu
3p5npxXza8soLnG98YrFCd7s9/c/tsXUVIJVW0cKhIuA2forVUqoYH9mitkKJeLtrZLv/Rq7yOGR
Pe0bTuDk0MikUHiSKPHgrx2qFpK9pbfON4GaxsVZeOX8fQ72fTxCn4zH8PXStb7pNQA8FxH3x/wb
P7TKg9nz/Lk7bw6o5xkC+Zfax7uj0sAGcBe8sXINMcQUxHOLICRUhFFj6kWJphtH71KK3ly7e+Xz
8OJcO9Mc7qOLQsipt7ab+wqp07IBG8b2yAFkUQMYBJ34oqTM8wMP691mTlgVCSNzYil95u6EgFao
Ik6UWNkM+HlFUoOufQgRWkhDiy5abM9E0gjaxVMdEXyuC5chRS5tN3yuMfwUjQ3764BAe48ekHeC
GGPEcaU6yMr+C+Iu4mUgaFOEO0Z+KkPEppz8TZVaPJo5TwB0AtN9PQTaRjDw+dG3u/987hNZ3db7
ihsGLxE2iQIIdr98ptd7J8ooj1HlqOfPR6N9glakTA0I7qZ4bm05BJ1Au0pDcQ5jbFJM3VpUx+a7
EsAlyvhfjv2lXH+4WvxEVlQ7+qYO5E+86uLMnupfYwZlD1ShCWj5mNxAp2M57gHwlqzA6L0pNk8F
Xgil/bwb70WV1C/aMjp+m5OPp3LAlYwd+6WklVXoU/lPhFxmDQLc0CdoNKuBY6ee3DNjn2ByCBQ8
BlCMVs3q0diGdFGl1Fk/6VRtAa/D3h7eM7fW19scnP5XdK/bV+G+v/FUU2oAIB43hONlVRq8GM0p
plYvfk3F2vRlWJnmFPHz50OPOsTGOn8Lmb7GnNvnJmkTy6EmpsGOW8JyAi/RuQO7QNwE9r+C2gGy
/XDKFsypdxrMKm3do6NXdypqNOLm7kKy+VDEQ056HTa1SuTppuXdm2xjCWOHCHiJYjPBQ3AUd8Px
hm80vGIuM5rG2rZGTgAhPdiefrA5HcIxxFxxRZr85nl0aCrj1/V+HQ+JSB0+nxlqaS4phlbPwJAu
nz1gB2L3aT7r3lqaq0yYaeB984XwiNRQHW+j82MAuMvTex+2f9pJ5SZVE9DD0b5H2z71MzQSxQ5w
mUwHDscOSsJ1fKiU3FcavjclHDIMNpnlHXtxeE0Un9i7tNBKnMU/eqC0gsnKiA5+jWSTVLmNVVAA
+A9mNYRZ0QL/Yn7wacTujhPyc2f8+2ziWeF6XeAzEErjKn2BDHBRX4RLOsRhPDAThD/DangJ3CRp
dTiRyok77RZCOpC7K5SZifUKDfS4CGkuRzHIiZzTo85ZB3oQ0wNQox8agjd1EPWuC+tjozeTuNhP
bcS6m+FAucXM8QeAxUG2doct9mTg1nroXrmF97lfq0LvR5hp18TXrC4CvuCJjwUsbODJ3X3HzAI3
8f+f6B4kAFKajGJYCzIBtbs5wyVlZrd5iXNALRUJxMC2WSDcLHcZDpm1Is9pezx9ZjBonxZD4Ayk
ecy5yCZJQ1r6WwFsRSdOLBivjbs5hfFQBHKHCALsZM7XThJpWlD4SiHnYIK5+Vz0YRINvuauE8kJ
vIItL2DIR5ZoSAAMdt6NY1oWYRIKJxy/il7Pwi9k9a/CKTTgNV/njRloCFmxqQJrVKIrjNSQ5OF3
Lpgsq97cfNPwMdiGD6gh3QZBCN4s+5vY8zBHBSBT2jxyged58O6tuOexD2P6PaoRhZY09fRZPtLJ
n7Pj3aBVynlE0UOqyFr3MRQcgovC59o46pScAu7Fql3dphMZiNcdHqwdIprj+iQJs0XZSdGBnxLR
BaE6m51tjOURD3UmoovKiDLOMlrMXc9RY+LSuQOt/kysWjc03zQqk1CHl6t8KAdNlG/yFbLxdHdF
RNu+lk7f8OiiyTjmFRsXyVqSOOC1WVHw3owTqJnz3kEZlHx8sf9n18VWSSkO8U01jfMcPHckIyIt
QKXu38m8GU4pgcICBh6JEsA2kXjvMLfYO/f6mPluogzIMbbnXmaQJumHm6SEF3PSJ4qGF8xJ+HKI
hGij80rnmj8lAQqpGo+L5pgMfyrjquwAVxdG8IEwUdXxlD5gZZb7UgDANNzcobSZ6R8NFbyxcWtG
aB2ZXGvQSji9nBgHF5/OtIl4KbuBjfry/3I9HUlCBoZvDkDY6LfqCvYeu4t+TL0f/utmbreEM1PB
HvRGI7sJ6EkNATApD9BKHgpcwE+aDFQY3Ot2F1zxwDP1EbW3ZPygOnsNpevGijwtgO0wsZBaOJxD
jA2RBg13MqQ/1EQ++y9m3gWK/jRH0rhU4wpwnkksdt09ZVd6D/e2s8THqpLrr7o0nv3WbGJ9e80Q
SgzIJaR3DW6bmMxVkEft7PRhAk/ZekwfrFCw0FHr8yHKeDIVSdO4/H0rI9fHEtMXXhV/nl3PLddB
Q7zXa7uaXVdEs7XcdzgIqUgnfRualq5yw/lLnEhhgW6UH9kN42yctMXOLc6Mfjy9Klw6g5g+rEqa
1VWk+iI29dH52Y33H2zEsNUE9arkQrljaqVUQdnCFxG4MEJyn2ilPgSpuqQLmrHsHU4l14naG3tQ
uPgfZcgvHjFJEUQY2erkfGWjy9t+S+z3BIZburJVO8uvidCyh38RPwDo5sP0HG7LEXncm3Aa1YvH
r7te0T18G5Fq+LqX6zkFS+UgKQClc1CD5P/CsWCHIgKQkLWQtqc3xo5CoPHhPokRK0dbDFtGSf8P
V/VEx3BDeUDPfVjTV2Z/fCq+DwfUp8u8tS1y98ssI/TmAWOWPybgDwIcXFRAotLqZZgIYxOKFHRv
XKN9FLTp+wA1Z+fdZ9t0LD7ps2vldfdzurRfpKlL6EtfkkGai87HMXVFjwkyAVECzBF19/MuJYYd
5uRqMBnzH4CQRHXctb1i2koO3pdRj/QpxRCTkh0C11UT5sUMXddfExy9RUQDMNUtvJ3jV/HFRXqo
BtCkMXmfKE2i1m/CxgV2VyXrnb2B9+rOqkgkwIST8z7dFPz8XDegHyYnzX04jqNBK/oJQkgVcbed
Q+b/HmAKfTU991R9ZHmUFPRFUG73sAsfe1diirLD6oZtUKdzLLBMslee4YLNalfQDsmmaRH5GWHT
d+CfSsa3n2txvt9zmoREgLYoBmQJaHhb6juz44KMrCcYvIYh+C6IH8Qb0YER/JxSU6G+CpBx7o0J
RcCvFcU5KtHG6PTZ19TBaG+23ieocBqWxrteV0JAMOWvKD8TwMESGtAFxYFCu6VUJAI/kuDrzzx5
T0CtznACEGrZJN/KDQQe0yRzCLWJF/StVmHTN0mToqocq8t3uNUWINglJ8N/EkhkBewsPFXNl5Do
02S3ldmk5C53xdV4fOoZ5dJTfVqd2A1HRvggsjJxFnElxPCY0ezeFU+4RYn0uf/u971K/4te3eVu
7d4o2gnodFlfJJySGyu6298hL+BS+DRSp54u+qw6WM8DzPDugJE2KpXf3pLXZAjhQlNlflUi4yCe
KXr7876tUOE6s6BaIn8wypegf2shmdlI5kQbDN7ymuEM1IjuP0mDjUa6BEocvmf8i9lPfF+6+0+w
cPNFwyBwei8x6Akr2Ci0rNnawJV2a5tcZLOo1airKdIQImivsaEd8WXRwgtpSxXqbthft5FL431H
OOfD3UqHyV12+sUMszajrllnZNB/r92F42KHKh+cL7onbuS8CZJNJYJvZMEtR2JZR7yfYUszIuNJ
qZ9UDQhy5xghRzGvSMwl6NVyFSGrOPMo55tiLzHX7Ci/TzaK/EmlGGl+0pFKi0CvXyFMF9GkjTcw
ddVT15VlCjw1YXopYA/4THye+Q/HnhNjsKquJ9qCbSxGX8GHekNGCKY7SX7iSl9sfAor53BG5Wuk
tG3E0K5z1/1SbewaiRzvHVb7deVhp/rOXdZ8x2B0qpnGu80AO9KupXQN1sbid6UnmsL+6IiutVnL
2IJsMpH7nixtEwz8e+SpJEKxCc89M/CkyXngHMvfowqewBx1lM61v/dWDR+Fly9K42LeuW0eQ/2I
1eHNuU5+9X090SHYIk5hqxJCoPJg7r7R/ZuPLR0ziew5wKIgj1AAZwArmUYCfX8+JjuPqbe95POX
amH3FG6kcnseBucYW4uNK60JUdpqb4D+eLUDgMi3KgIBomH3yxWkQO+NQeAt5ZcsHQU3gzGRVNQY
nqZs0yzIfjWVuCnZcNZBkNtV6jdl6fRrnKTL6VS1WXyrzT4WGbvi9i+AnbUvGmKI+d1mClYn1VXg
EugWLEbb2MQ6k7ww6kHdRO90YY8PyshY8R2bzbP9rPR6EWDGwv6kso7UJ+vLkn1UESPUYNkzZt67
P5KBLOx3uGQmDrcJHegvMtmOCkE+p/S3L2v+4LHJg46SgX0tzkoTQyN7/cNA7L63qqOkPEW1SoUU
/8hPFE6pD2qT5UIC35ODT3eRvAqb6KrTySrRtXeTcGfl8m7PLDYELKeht30E1VPPjSA73IWRo+EV
yK/Exx7hZxZiw7tMA5FFlgrsbLMLiy59UkpaS1N6dvuwKY7a1GTjrHtYX5esfyF2gVXGYxQZxlb1
TkzybwLI/wtVwW0AXp+gTu//KDoEWvK8JufQ/EcXw+tJjI4kJE4ZQmSo1DE+fOqPdtMsDmWJMAJW
mnDQdMj0uLXeDFD4l5YUoVKX3SFJokkDhWVYx91HaOuA28UgPbJOthX1GEKgPH4QeptoRQJXT2Ao
PDyuSOf4wqjAlecRAH3Cgn59Uj1LJn2mHEns72YtaWQfoWwHovLeKOY0uFoaNL6pcA1/0nfAVL8D
FzSNs1F5xt0zU3WZ3EujMPGqyRe0FPS9Y9To7Uu0aayGYN7YIz0/v+6So2WovimAHhsaHQzDiIM8
XkOgPJYkQXazTBXaclCRfM540CVf3eaIDBojSJqZlVafXJVwDCVhGx2WeL94fuK7bIsrtf2B0OXf
9vLPCpqxEnPdAj+RUISbRu9vbUlQbi1vdzgMBp/4aaD0/9dp8amj8RjJXpj2GybmIjuQD3UiWaB8
cA6mrN9d1HZhygznNfXIrqVLcGmvqNpv9e5gn4zeLQYjxb95dCyFPwedLGJ5ObRdg2JPD+LGPCr8
m/FTS8Xqudg7bcJhY+Odo2f0GCutY7wx7dYzBA847cTAWPns/1WfYBfn4gfNwu27VilwxzUTFXgI
fdmVKIqcCDxCj86TgG068pLFXiYY8FNTf5GfYla6SiYZe/ahGyQU5Eh8EtBrSUg2Qme6JdHt9OdB
BIc3X4XfDC/oRSxFgF5dFwr6SGAXIZicPF8I33DNs95MEwnUHJNm7TXh9FG3DGX7vKo8rsI3v7aI
C0JOwQBhB8thyXyESL3dO8ymaV2N43JyXsHqTKgWR4ylqxlZ8rb3+lPbKCFvjIHFu5feUHlZHHKU
WNp2IB6Oz7fsup8+oMklZc/RbNc8ZYvQhLpcyiKIxEUGm6sejc7LfjrDIvbiGuAH8XVYO8RfUHwL
goXVEbDffYWR1H9L7tmBU1vUJqK/ygIyUo9wZ4dGKUA5cTx8QizySOEPWHaWRqtEvrNNf1Tf1wNz
UPip9bFXBPnPith2xYaCRLdEWQBcfO6HDvi8TfEMbHtRfGJzk2sYSwhv5cQDHnHhGbtT8owaHZi7
TUiEKzSOoXA7UkOaSXDyB7LuiZsdSCWSG3oB6Spxs/m80Qic0nh3tNlgYRLtojPSJGUORfc+JHY9
ErbIArDYUK/gvSaW6rUROTw7aG6gr+hnBMWM2sHC3uSwK1W+oYmO1wslCptM2oFX6rlBqjtbkTgP
tzrx4rM7bIWt7fGohk1qAUfw4qGosrtQeMlhvd+vXHdzfhwFWiuZ2L12uJXd6S3osGR05MQiN1ju
NepZlOrzLqi2kM4y0xjTUtFboOtSf5tz2yxW917MUp+YnrF1Dd6IlufuyvukdM5UEX5g9YR+psZD
72iNEiGRgbGP1WnPxs95GNoVUFTrm9RHd4NSq6tTmR1OYa1iCXWPtb3WUZ9Ujn9wpZ7PPLxu7FWN
43+gHCuoJQ8jD394lUF+rMUGMg8pcF+bTR88D6ijnAckxH07siGOEvCGxUIGqFp+TAbRLqcLQban
DmqA8S8/aFm9WcjraE91hYWsbq41VOyehxyMGluHCX1ohClEaM814oGAn4NGXQSk5MTOhm3+8tDl
jZ05EMLBhemXeGOqbG76IjZYq+D1HqbU6KzY2LGt3wKkfl2s5aFM000ni5NIBmGHQoi8VGH0MuI9
GFEmvNmTsHkcomhKsEcezYcGpPddwKz8HWizPgNfqnoKxFY7/9JZQgFKY63SZI/agERd5hIgAE5+
3rCAe2yZdj6kE2PYdSYwJfYS1tBan+3IhHUkDnuZj8RxGI4JCncSkN4fHc23kYOEo41iI8eNLsFG
73P0Tz6Pfnx0m3Ao/PpF/CjwiqVE5oveEouk/yg1vXE+KeD0/LpdIiiJ2q8IuSKnWoLTgd91rJ3/
Kl8mSNbZpcsLj8Uh6iIMchJA5g2Gh548Co02NI6FQBvJDhNgbd3vnjCCtoAUoVV5BbtlI4pBBsN8
5ktIrQ4ouJz6D60PXdW49Uhck3OBGmzrb6eINt+s/d4Wy62wNXVRfdlgT/aMD3v908qaJ4StaRc2
ZQrKujSLQr6891TBNIeQyQmRUqt80aiB4LixQh8m65oNubuH2guZT2DeNGPwqroHgr8TbL+zRSYW
IBbDGqjn2bfZ1C0tHmiKbLrbE7lEtV6Gpz5AL1ltcZVnzRMaU9XAhm1gSkGUVohTYFr5OI0XBB2G
aaNG76tQLipzbzd/h5KzkgucvvuTYSc/Rpgod72qYWBDBrNd7qugwIZx+j1J6oeaFcwECpXwm3+q
3lgS2U7ycbqo1/pM59A8whqOcRSjBD69OXvXPi/xr9QgFAWsFEvmrCyzXzrW7SKx5Psi1jY6KALS
r69GmsIFjnxFa/C+C4B38HzbjbboCDV7haM5L4mieLY3v6dFUUMzN1jafUKSL87TcEEnZXjEedWY
m9J48u7M6oDbn+qI0+FrRRAh+y8Gwc5hbf4P0eAu34aJMwEyg6T9kh4a1t/gqpiJ9iWiM1M9LRfo
ztu3NTDOZrUP+4IEeGyYNCIt2jjGRf17ccCjfyJUhQebDjqfs58fIGlloRVwjzzKHFvSarRH6sfS
T+9lf5GoEzPJyRFJI4Pzy14a2dWdrjjzItWIGRdfzNIaJHsQAHbDG+ttxGCpNtgU1fS7SaxSbyHQ
1winJr0X/6NQ9d5OH9kQ1eaY1ep4oSmq67/dj5T4Xqt4fK7QwLbb5RYnCvDubrNouaCBr2gtSwP5
rCKGZe0920kdA0y46h2P3+qgaqhnKpkiYqutKG9pYJp7A8u0vKpv5X56QChSfjRwU6sjn7P/iGLk
28z8Uy3s4Wum2EOxlTQCbcG88fjO0k6Ow83Rkmy1LcN9ZM2wFI0SnBpoqJDWt5Ah5/zH5HQH/B3E
T9N2BuzTcAIGDR+YORwkmNvD+NouI0C3DODB/WuC46U+V1qPwbOsi15gohX+oMO8TnC2I//31GcZ
MYO+c8jebqcLb6PNjzpyYtWbE7t+4EgoMGV8AXN8TnvURRkLCCgrV5ar3cNWh7xoOHySkStmZrmP
z+38wDr6LRVJWw/qls4pwGB+zWmKEwO/1FIGfgs+WHjC7GriM/89DpPT/1PXIkmjNpwZCS3HINtw
7/uY6LLsPkAy0A8qAbEjWr7H9vwgMelP5qum8y+P2czIc9mvC5kdVAzHNDD/MpCLzxMmNgQqVYtq
3Ite2/39irrXPkAO65P0KRQJAeY9NBIiomJEiJ/JlRHpTzbxZ5ifl+X2VUkTtQwfLysF5BU3PhXz
dWh9cEMqDqhTPmxAP+O1ZwVqMEKce+T2AojjPeywvB5ejiDzwdmOQiE57Gyv6iSUQP/V2SNWjY31
tuwfeOVzWCavy30Mj901+f6um9E4CZ17pg47JR1A20e4fsm5PgggfVvI9fMtSrbmc4NZYAnhDCQz
VCeMK6Qg/xIpVI6Iokj6YI+POwHqNIO4ym424eQzq//rlaRJLgYzkZCBOWU8+FMitkF/B6ar66Ve
YQe3GWO/xWZZldhiifj7FJrB4mXU2XzR6J30KTGmcYuBEOVq2VFaYTA9mRoO6xNw1bEN9/fAEvAI
+TJHUdSlV9rfsf5zCt56FpXf6ZKMDmmhbxoju737gkcfaTN80g++mxwyqmaVWJ1I1mk7diw5+hO7
7zLQYJWHEMc249OuLFzVxUKLzVUgA9ZS1EaqnMTHnbgdg+YSxSnaNCcho3098ht15aSw1wyoctdp
E1R161T0+Qa4eXmCIAWVSfLpN9SLxi26Y3gHBqlRijEGWwZPMYSqVsu8+T6SXsUiyRFJ1LoZiCA2
/x90BEn6BTes826xn29qmqAiZzOhY9iDcSnl2TYnicg4fyee/mJaJcfmgqmUSgPci8IXpGAzaWQ7
B3W1Y99vmwJU0HaUrr3tONr6643n83ef2lU0q93h5b/6ghEAkDaKY6vOfVyDQEeLHW/l/GmcCUKP
IP6Bk0KoCPeLEwLvNlNUENpImo/YfRLJqZJybHiOj/0Rg+pNpUKdTIpFPk1intXjjn0YnrpNKPzj
fbnu1QcgZN67D0dpZjrFNID8D+r+4yw/gNsNesFjlcYvjz4DJfZWtNa9M26FYIPTbCw5yuxaVXCD
s9AzhovV1s5LlOTZQPXKP2H4NmqPsQoKSGhlhxRmkGEMTD7a4YQdnqsgXPLGeaJZAz7mKWVdgqJ9
DhEwSEqV6Yz7f1wdc99etMFaFQWW5P28DXa1gpJ2mAqI4cdWKz/nGzlCe0T8Lk7BZD6cpFV43uQ1
rHwx5y+BSa2/r8hk/xWm1bWD7BsGX10QFJkJ7jEcjQLci1fsb+Fl6pSDMio7gPT7CSn3tl7Egmyy
zOjp+t2lmo86cBcRpuivinvaJNanx8toW49ptXslJgedr6HYYmscHuFlaowfPrm/4oX9vy3sYw7L
2w4RpolzBTxlIyFE7cNc6AovBkypbP5tpIYLNku2vXmRDpkoCDovjffCEEqSX26/XRB4e9lMI+TT
P2kku3l5AC2jWDDGY1Mt3MfyBbZuCf9Z5HL3pIPhSaRkzOIc1pLcaA6CSK3HqEnzMymEdgaA3XYw
Y+mmFBQoWiUL0+v14zAKalJlOuzc3xRKfEIrp91cVVbgY6355dWOjc79SxkM8LobkTBrdKl2bNDE
ygc2CVGdrxYDRin0bs8kgkguEfJDhijE9g/NzaG5AX23rr8/Djlx4wczNAXvxBAGhUdB3zWOEABE
ttR3hTVEVWpVEtpwvKu5O7IIUtBHURyy1X4NCIfOYaeuWAyqJXW+0o8Ao1heWwXT+KjPydH+VDAy
HvsozSl6lJOoRqPAId3rbCYdT7RfxQIoX3sQB4vVu/dyXi2FR4YEifp3H1oMlGbE3AzxG+HNQFYU
kSqFE02rH2AG0fzNezBbv1so7gsIQyxT7m1yj75iDGcdLEa1jZ26MFCTc5+VAZJrNwkBmmDve8Fi
YkYY4vS24Qa1txbQ9W92QNI8U9tWxM0qERewrzVmHFm+TtTP5uLprHoOmAw0Ngzad55MoXUBs/ub
yumUF1j+j2LDFb89pjicG7R1ipCD7CsY6COgUxnCuRkXpecx32cGvMJ9Zmos2aOCnAMoR0XkBfJH
c6eT3UKvbAktAi9YIFQM8C+8gXj4aZLF7thtHJjcQcPVaqU0Bsc/+yEiH1idesE5Ta3tqQNEuad/
2krhoSdjidtx87ESob00EDRRnMwU2kaKNv8FEZ4holQwGPmFO1NO5Isyy2jpX7YwZzz30f6EBkwr
FKyLOrkJrFwqCHCZp2o+vmDjm0am7DgKhgGyENWlLHK7s2a6MrrtUHUPUO5v4FXRe2NKCwcgiwRZ
NGW/NyGwOAk+xjAN58vkqZXYjUdcENci1feZSnjj/k0ZYncdOqynGnMn+G38gbWK395AyymaXm3Q
AGHz/T4p3LX66l12+L0fDMHSi8B5mXXOcl25FTB9feZUnlS0sN7BkKYkD3w3o0RSKH0plvt/ujUe
UGuqgr3Ed+balKE5B03gQDhWlQasDSWV7MfVKyaV4ot5b1MEpgzq4WawLGzOpRZRYIvoO+tfyWMl
FnDjPwq/3n/o7Tk7lN/yfIIIJ8OHnsZbxmM6PhOm9KoHqFGQOkPwbvGYLYIlHmjLXC8kjYIucXYZ
FBd32KI93COkq5yNf/Lh+M7F7y+zdgCS6w9/wnIFFFdv7E2o6gezkza8LCrhoaSCIgl5XGjtx3NP
UhmW1awiuJyCjKt3FTD1WMziSgGDQv9j8svRrX80L/bNu2Ji+w6VV4Rqi7A3UbronlFwU1kV/0KP
6CczOaDkgMow056wcH407j0OsWnqv5ACD5G40sA6bAbGNtq2SPOSq9KqOlEvv+a6rK7G2mT+G1r9
H+O3ooedgL8AoVP2RvNfncCV3b4JwXKr6pA7/uc0CvUf6WhJ1Bo6CentmI78V8yeV8gDYcrN2o/Y
Fb/Ao0QBqVt0lDjpPMvsavS0GXsNHX91LlllouiadpZJo0ytEoRS9NI7v0diqVOgKOsZap4vN1IK
s1+ESdSqUX5HuVPaRhWxsT57MSpIQTMRdza2FBqYXTMbi7UWmgzBDiNBhfffXayjfHf49fsNg5Hq
gFY5BUWeZ/1ZFEv9oDm/mzHIfNsWdFbmXHXkvL4RoXhL2vLGTCMi53T+zcKOtf/8gD1IBVCDRl+P
kUpOExkM88ZZmjxRAm1FYsfqevggoJpAwL7z1JrcYxxBWgU5SWRK6BAZQBFJkt3ms3fWJJTiC4RE
sxyUdR87FTQJaUn4YHUpOZlSm51XoPR0JPuDJYuGt+BNwcfQKDPMYzw5jZ4ePjLsG+yDa1oyCioO
gL8vPEEZdziLf5RmmyCRNA08eZPW0GNdhAAKSoFYf/4vSUq/07ktg6KPDQVQa7Gz5vqq/yCna6mw
SwVCpuJ7PL+nYJZAwm7tuPDK4WSneTArwIDRZs2qksmpP7dowo8PaQnq3yBbKGJgrLEGq5c0ver+
gyhPHrDPVauq+uVru8PbF4WiJ/WqsUskLvbT0aZ3C2+PwxaFBtvSVIWe2/3i2QsmlWm6tJ4igud/
2omrKPG99ZTDXZ0cYfYaMO9uHmwr4qMFYzdcInsJmjVcD/5+Mj2WhcWGFhRy4UK02eEBjrtTe/FJ
Bve383fMd8x4DktfqJQdKI9TTU8ntYUJSm2Js6WjEru00DxTSonD/HiqNwWLuKlWk9ESw7p/hTcy
HEIm/V11mpvLjlYdXk7WISX7FvFDIKySI9GYjCTtJl+42LSN4TLrDDe4YcwKC9rfHdIj02nUQvfP
oF19033SGhTM0mpqnm0yExbsL0gOCig81F9dZE7yYQIJjjtVaidWcdhLrurbzdd9RcCl/unQVuCK
O8g5WdTge5lHTMyVqzBbLND8khN0LE1Ta8Qq9o79yo3811LJSs2zKp78DrJ+U9Crx6kfFHtr2ddL
d0c0BYHAwlliP8D4pLTpaa/XM3/qxlBqmrywwkyA57F3xxNDfmjJE0qb9r96JSklJC5wa+PEZ64G
3/p+1VhXJno/ra4zLGqpfkDTVkckDfuBIJkgcqfxp+0/d768wKVZ51Hd1M+CXbvny7gywmf4nuP6
XDVS76+12cC2+DfG5P1aaCtCnbz0A8B4Ct+BIhmfCd5BqEMqNlV0J8okfuJDtkxYpil0UbSuS1og
QvwAucMRr7iEawamWZKFjYcGJqSKjl96gqyCXSui8/RxY9IgxmJ7y+lgj1wMfeCQ3BV1FKyob8xU
m7qaQiWMsflUDaQfFf7FJCyy7HbQT49+RlhsI/qlVgZEtaZT4PEAF1zh5AUEOsqqnfOKnWCQq1u7
+ABuu2b3Dd0eU2zksUCbPkxXeqHDs/3keFQ1XbHBhUVbz0SEmJgGw77dSt6kmEXORGZNPgFnk79V
HpSsIpcsFuCiApR+TffLLSoZ2l0F+Hps/r0AjDIXb+HqfzFMsWYFfiFnVGoozEPiYD06PdymXmIO
qV3iH87eMPT6M37vNqbqq1Nrs2lQ1rarXT2ekyRxWIEfRIct3IUHR2o4EReafAFEgIEFBCZrWNTn
33sN5YkMytnRmLMYzwCMLOPDGoL8MOt8StrtIq/MTcaNPCMJTaeUPqgLZqxMHzpWkMj5p4ABrGzN
xPw2NZaFy7cH0NLYfiuvzadZxzuJHzBXe0iw7hHwe6LyqfFf5X5pPRb/3VOmHbn7BeKcmPKpm4+F
4TSLNMBd2lDxfiMhE20agDIASzZR6juylblUIbA4lBYo0vWNE60Wnz3AwF6Gd1XTeRE/W9Zlx5pa
GwbOn89IZFBmlV0ONnLQPe/VoNpT+1VbfOi76iG8LtEktmMSyHMIX/9HxdgIYYfuk5THYxxRTJ9B
2JbtAvt05Yu7CqbR7CLaeLEPoksm3+HiOxlOReyiWqsY/0XsLmvXSTq+n8VOkrLFWj1vg7PA2H52
GeSjLMceatg7P4/PqRkY6/GD4I7s2827CFtzeiE56KTszzjvW1y580QOT9Ggiqms3GclIq2UaxJ3
CY6pauASVIxNMisSJ5h6RLFWO7UQ/6SNZOi4YC6+ArVzYq8AgPh0x0YaABfysap9d+feL+EY35Q5
VysaWPXb3nbt34Wym0dR1nlNxDDzKVJGdM3i8C6i7ex/vSACyJuqZRvlevF9xNMKdKwGX0Gfolda
joBM8zuRZorXQ+1xm8rhWnhhrWokdj1nBaf0zFR5SPnijBZrxilNLwUEmQY9CJD6/vZPaR/3zgYR
lFWhTv0ppfBmwj9qw8J32YSfDWhFe4BlcqnxburVdXgHdFULZngqfRHYuQjWAObkY4/2xTOnsA+2
VqzL+HUkmiDAz9cTtK6GYASI0WqfeRkxzYwd3njCUH95NAQf+EN0GDVs4FWqZRygxeSmhroLq6oY
aplS1psT+uw2NPLS5FKO+DuHG698IAg4AI65cpzdcTJ+oFJMSoj3RUDsQAHdq4IGXXa11/jFeNlU
nr733nu/pLCe1NoDREXuOn3nAGFd3Vc8cTFUvk2lfgzkqApTB0Pn37lffKH7vyLqPgTAIbPA679/
OXEv0alpSPRPvtXCA0Bf+xrojzHXJtVtLSWdz7PiLHRMXwwN692y86swH0Booe9YBlatajiPPHXr
91+Zcnfil6aI4No5a2SzjK5C/zJiZlpI50JD1JRP4W7b8UgEhzZSGAl2cmZ/hUCLwazisacT8mk0
Um7ewRJRSqKP6hwOyekzLXFB04nIm26Wtc63eyoODlCYg+VQR9gzTFo5U6pNewn/6wHV/05PWspn
3BstvDFFtUJ8C3f8C3F/U3O+HIxcBIxzQEwJWKndFCr2JU25ff7nvVX84sH48aX1iCH0IHYH9O73
GmVkEdvR6onmcAN463PDYCDWiXoVoLZyIPXUS3nSWZOL6cbT5UVs4HYfY3Pm5qWnyQ73/oHhuQJe
C5gZ3XVy4Fcb/N0IDvVLj9g+udNT+Jjm58OYkGjlO4xUMgzcSt+42E8M3XQsTysOgBjFybZOar5w
b5flaj8q0Fyva0iqXLE1aZyyI5GvDU4VZxR6bCi05z4/UjJ1LVd2ju70TM0DOYLotrqWSszQTDcA
/0o3WfvEfJKEScwMp+JrIW+/93LTOBR0j3nuVoIuhfRYp9OPJqxLUVMiLVgg5670wyQVz5ZZMqOV
Otwk6yrccciZqlhJd/FVAa4oXTlok+w5W9ArDKhslZX5BkIOQXChBz8XyRnnbs7Fuy1cneHEw2Li
/QSApp/yCtXJqNSfZlc8CIrwcQArYH8GrdXyepMY8v5RNadl2jm/6nwLFBlIT/Dwc/4HK4AaVQin
iASaGYjvfpHCUd+8qJz1WZrWAj57Reb/0eYhaLFDu1NMvKdux5aGLcYhdnI0UoLaJUfKGOfRZGNN
SU8bN54m1K4OQOkCHdgNVSjNxLPA4kYj1rbDqO9a5phB+Cd4jIdPN86aqu16kQQ6+I5RNBNLmgJf
IBN1hZdyQrittboELmCMPWeI1j2kc+zRVUfukRR0e0pwhKHgIOgZel9iJB52aW4Zlw/1vkvJGCps
XvSAbihXZ73jzygiKUPDj355SkyfJgRLEyLkAiZYw35SxkF3E8wWsWPDzNzf3w6B+C2MvAmxm/Il
tYXKXeF41eIJt9RV+BmkisjwtL9aKod5lShQRBqxxT4IrZtopXyPQ3jsJdavTBZs2ifb4C3fQAGP
ByxTY8Jb8CYaz5iVaNQ2aWPmG2SMvS7wowe4RGzlfi8Z2ZirEAX9QEzEeDXIDac9B5SjVDkLOgM8
YOJ0yteWtgY7OZ+hhe95yorRX4UGpdbnVaXeV2uUY6SXhd4AhWBdc6LoRA+52mG/lr7dOyNuTJfT
edRnHpjS0IBRhLyeRCadHtx4sq0VrtmrBw1m/YSEyUkn5bdh//CH6cgB8HJQ5uh6eKF0PYJcEbEg
9T+M3TnuQAb+9a9z0ut2rP6fsaYDrhg0tfttiP7y2VjQA2WcH66SzWILBeiUKBqX9Uya94tPJK1H
znQniM/1D8W6I24n7ktHiu4ENSml6btuW6gw7wyidw9Wc3oTAE2+3I5/av61WejrypcFcRoTlgc5
g02DsCSdXxhsuhO/PtsyYkDB0LjJ2tTQjqNiWhL4l7DAq36ZK9AWr5W5v66sf439jPjgaOEb4wcL
2i1PPOwHc463O+prtbeJxw/C2eEk/ye+sESDNpeSrzxGG7vEW6o2vl+JeSrCFVLvP9qzzDICq4Vd
7RoAU5HOWhieS+Iqk2bhurohRKRieqh+369navGIAGDf2ZpN2yjHAmhPzO3tyIyGokhvd6TP1fnL
ipsSV8Q48Onr4fgBfReNTDkVzPkDvjmBS70k8OU8rw9w7bQTHC1GygMVb+zhbRE9glcia6SnYm7u
oYQ1/ucw33oxmcy8yWzUbWFTcrE1QuR2N4HBm6QWaR84HisTOe/m4Wsw+6+3gV6dPX2GoPhHLM33
PS362gAIt2R1fsflRfvLxI9X0XQ6OvbE7mAHQDvlpbtxp7ZSjr1ZyR7jz/tI69DyWvwVnHgcajPT
6anbu3fq6bSHS4aN/dknLvAyaRKJZQcdd+hzj2v//AbWWyuglJQgrw2ZNaiguw2EHaIJP8SND9I8
ps/Q34WKkcu/esgj5azOhv1ZvCv5lKQBWNGZfVrsmx2hAyMKJJA3z/YRVzWDHLh4co9Mlk5irgGm
SN9EQ99EBcdfq+5uMhmul/DfAnirRYzd9aTqkoVNYEc6/l6gZN9p47BPziyvNo3wRGEK+8qfWmqV
m9f3dAQ23DGUme0lts2TWHzXGT1hOMbcDc1lFivNgR0yLUGj3/FyXbSMwz8GxsLmkuZ3HLxZp5MK
Y8M8CSeFcYE7bmlcC9GIb0r7YoKihYlMQc5mwacwGTub6wlSg03J+oAWUeakptpcoC/eR5LdEe8G
Or+FvJU1r9GYyzlawKV1atLiOtgixRDtSCezeaTBEMkMh40ym6eicogPeDd6cnL/iOuOFk1q/ykB
2C0Iy8CoQii6gtUqCWDpq5bDFaMjancJLULJlF2TX2bSuZerde4qQQrsLwz9bi+vQLE0gbTkeK3E
s0psMVmuG6VWDKSxohMApkRmunY1L1OK/Yw5b4dG1S+k735VdRGh1zAZA3YZbvFyNylxa/53JcIs
265aKRXy5ujIXdxGYC6oOBTgvYkj/u/LHhFgpo/XaDdh4i4aL/YzOv9TJWdIyvoo4WkSWUInGQqM
RO67IdPWULRyOt64bYt4qIXtBPW9gIlnDxplPFh+EDUInWu2ceHxSxlyXCyiYcFJRSmAIf6BA2On
blQf3zoMNxNU3apR4yfdy4jYkdnuKrE+VHBQOl51elIp7EM5zE6o7vw+PYmRJpKVpiDSNx+H7P8R
Da/rnGmc5XSyNm37HmlN0enZQIKp5kcqWw7kCE/TVnWWDnlnXUhcXHUoJ/do72yHEmicEw7CB+XH
/3GrBiYoce8BODRjJpuXT3u/k04/pUebnPw1MylVQBmF2EuWKGvBXoBgfTP9EJ/q06kVq2CGFExp
n6nFbfxbUEdDAW90a6qJjZcPKBN8Q/RgPtU15gRw3xQOw43o16ruPF7b3otCADEgq9IACq1IqFPR
VSEuVQxsZptl8PfgouVK8W+nj06g/zYY0ZQTTVvHNu+OU+WDJsvAzkduPhFAbR9+ujNHsNfqSqsf
bvy1BQnuK0ur/9u6wTNNM/gHuaUHH5ninPp23+dqxzx16hWecFASb/2AsnyNdXudlpiI8SrN8xWH
1awsrW7zFfIBpkR+eI4WP6dOIj+c3aaxn1+ndLCtHRNEywJxrq8miRwO48tGujglCyTbCWVr31Ru
Yp3lcDSw3VC/hDhOSQV0BmB413/wxbVpz4HASfGVVkd5Yta99WJSnvsjtoQ4aMwpnImgPUH/cEPW
ntrkir4G18np9vr+ou+DVC9u4vfpyJqng51Wo1EfrDzoAq+afnfFaR5I885nPDRY3NbVnIQHmoz0
c3PFqs83ivA6U/UjO7uDpw+vEox/BF6sEjeR4ZIcWKtkCxblwEJwACYrcKyLSneINHuSk45XrghP
0zbgAvI99IMkcoGIVluyhxuwJfoQDH7aLftg8IYvjZmTpumsf/g1m70Ta3iAixqNy5KqDqgxD8G1
12HILRZ8v8AkSRUi9LL6tgKJDOFAISACwajellwPCf+nAX7pCwBiAAeHh/KQC5EyEZaqY603NqVg
seAAUDC7caD5YdXm7gWuwu4uNFfAkfv2n/OSRE5A/2PiWNV0e4ncfnAtdBKXtCcHzFvKkFcr/RHo
+XySKuvpQDVT3jqiLbo758XRmESSdAyhVeX12BnnrhzEP9/KHBDwS4ncL4SzeT3X887wMZYUZaol
UHJF07oBot2hTQ82myxBAYk8R5xI71dWVZYpRmGrbgDa7gYiyTEeL2toEoqf0XRnKyQTQx0JtxJC
rvzId0vh5cv1nYicOleYpfC3y2vLRxvMHRayh4GbV3vGM6biNTGqvYuWSOqrPU6VByCXaAxXTPON
a+KxP7Y2V/e59Vr1ARZq9f8xC0iUYwOgVDymVn3tBI5wbqS9e372Vo4c2Whdn8Y85mkgVmLjWQnl
na4/mi41ZmNnqP0d46OSRO1TkYudTsoVvpbHodN9tP7TWE9yV9QCeKExZMHqNWbvQO1d5OOZ0HlZ
WST1qMxbPu3afyue7wgbx4q8S0LV3Yk8gm/sMbZpOKw+FQGG0AHG6GlwymnoBP1nXG1WZ28cUz10
eljyCyHiQ95R5UIwsFZQohZ+x2VovX+5MVUDuo70OEcrdsI4DuYVTT/VFNM4VzAZ4FtlOYnfFCj/
2BN1xBv6VYTvcG/YPU1n/S94hpZM+UdpvBox156UDUOz9oS8ojBiCWT5xBjjfFMnvs+vPHIoqdBZ
Cq2mVEUaz2sZW/KqpaCHuK1dasISyT13EMa+ZBfWdxJY0lw6r8sInyVqiXttJriMaUomrGuE4fDL
4CMZitqTUUD/CUYGmM0ILUnrllphhbv0YH8OW5gYccyp7iHoc5jAX5dFC+1uyjy0oyDaFcKJngST
ALUJCIRgXXeyOpkAPgRItSFz/Ls2X6cxQQq28ovAT0D/yrpHX98vEJZ5gPKj6SgX1fOv3Onw0wSJ
mDo8dlTWpaA2+fQG7HCsqwFGPuNCKxsvym1r0+OroQSkDtGsbInehcScQGfz6IRFT/tCN+rz7WxC
738i3sdUrjM/EZpYNFfTS2DZZNKQ88LJ4v7ffnDs0n6zqutZpAkAX8UoY1+co0mB0svEqhUITmYa
uORtuICcVvqj1yT8Jq27Guj5nX8y6coj5ViH8kEh6EREzjbFR4babvD5+zS+rToFqflmM9QdHMxx
TLeT77YCr4anYA4w32HfHhasws415uqQsAa/nGG6Yv6bPyub+fjJt24dae8M7PyPGo27zTUyov60
3A6Jne97NMfNTB/l+Y5xCZhXsf0k0tgfh/1HGt11Cs+TqMA5kDgPGxfMs0HIlpVpsKuB8ih5Zoqj
rcunwGLqCFYOqEEbHs2nvldYrGgsQfn7KY+kzcsgouGijC9xdIrSNyfSbZeIHuWkBCEsuHy9mbkq
fyurQU5MquK4+Xf49C6g3h6kKTJTT3yvMOLcM0A5V1etyz3osLaCMVe0sUer8oh2p1/Pi/sW4lVo
T0nxJc61iGjfEBIYUlnjWwfhS9XZgXnGNSb7pcPPZF5h81YWUjKrOiyDysQ2+sTJnOa2K7sjGURZ
cWSZ5jIn9vU9XDp03NMauGQ976J0KZe30E04SGDULKUBEeNRvVUoxrqwArHJsLmNPGFuykUKba+B
ddRhLaOKxkkyXVkRoMQ1hScFksF16oiyNpWEv1bxILx++jLkBYxSM1ZEAToCp8O4QfP1iTtZk0zf
dM4Vzu4aay49ApL2zOOmfp7FE49xF6LibMt/BXzGSULnrs0POnVbccTsCfoYubNN6dfCE/KohT/9
Ipo27HLT0jpYGUhi1rC/eATf6c8AX86eXkivJTgPrdVX+ylDOrd0eVayuDYV3CMfMpHiAgrfZDAb
m9zLQcgDE/tzWlv3oBz83FdgqcxMLjdHsPL6EPyGpIFL5AW9G6LujtfvOnYEDkv+o9/5ZVPrHQ7g
tj2SsaBeIJl5S1Zy5sXKXutry/x305Ljw6Lqm08EkTrUzgOc3MiRez6Iv2De1VaPZCb3iDqMdRBc
64qEIkwRWMUX1bd3A9tPDIcENzCudVA+D8iu5fNBKmHF7ABhtnOhkUBEwcez6/HHDuxaUJ/lMQr0
tJmjQm9Sff2p1Irasjx4LgGwXbyPs+M/1mIeKGaaF5F6Y0Um0urJHphW4Yrr8wgSJk5L8y7IoB84
kTF/nvpY2X1NjEvS7fEOcnVIP40ouBhmZBNwHdO4Djv467qjdThvGp3YfsdSEZlaIYu4uJPKsbS8
ZvxlEKrfArOf3qo2l+/I2iei2JJ2QupJqzGnm2rzp6snsqSyYQJHTsWZzJp+rBG5KA6IJcMCJF6m
KDN5CQKiAKEIO7FOQ/fEo1wfhJeKIneVj17VCGQJIBC72BjE44BaWexNtYDbbghDTBtEOS2VqGZE
n+vxaSwZPnS5Y4xbtjlefY6BIMCEyRekRRooxAbX+z2gH7Q1karTCCP0eyY4R/Y2oyV9dIoTk6q5
UQ+gfjztjnoZ6WHjjpyg01Zwen2fgZK7+OwCwVAbuliVoEBi9MmJG8cfB+miV3rAclm071Wpao3C
pwacH/nQ408dp6dlUMuprnHq/AnM/FzHkrA1GZcQjuRcMMDHvJHT/TCfGz1k8NHX8HPVdM9L83j8
Lls2BjWyFqDFlXnHEKUHY5gA5uv82kguwtgfKp22JUCDoqcV71kZEhyYCZNxU+Cu515ViXI4BaEJ
ytqCJw7bIL+NE52DwK8pPNAIUQcyz22FZA/7dXOqMRT62cN6qrEeYRIC0KvNDcyWmDpLEYiRBY4X
Gh1HMKErrnBM90RQev+6jgF2pRq0DieyRamcpA4VqQ6U7324x5iNrNaugwc2ujiDmRAeUI1Xmna7
h8yo19XoVsqnQ7RV6WTZo7gcqnQpPPFljAv28k/LTI4nhvdQo6Er85PgbZJZUBKlgI5SvC3B3KVn
l2l40LqO1nuWqtfRyNVimdIGIuHimBdM1jOLiEZEteEjEwhmw2v2m+XVZ8AmyerkmA1XeEkZolQ9
OYA6m7RSSZ+aZVY9wgsSBfjEGf3PGL8oEoblALXEd2z1kkp72xWSJqdaadsBe5nou5HFFWEr+nUi
SER6RZbNOvj9Qc8ffmW/lX9KOPSqse2WYA+OrAGQ89cmOwixusAqfYXU5tGzCgRsEjipHCkgYxEX
xNe39aXKXHzREHuCtCh8uhrViL+eULs0PQpgcvoFMvBZLCdZY1ZLCNUuxHSAPIvqwlZtqeJJ6uYi
E3YOlRinVJFHogP3drUAHf4aIAnulEUMdmUREVfK9D1BjrQHuAZhsffmURHwZwNM/8HZEDmMKcZ6
GAr45IQ+RRoqegsT+myvzU1VLaoorhI6RDWyCTly4kteNXL2+3GiY1+nW5IO7A3kbX3PnJ02AnBo
57Nueamr7d51DCEqB3CNyWkgtQnEG1gtKhvVzyHRG/OdyXCaV/DdcvKnn9DUbj2aRp7aA1NZo3R+
V0JzsqNQF7ImFDauce9T839CCw8IHJradJerLRlj2cFoua2sTXkdgtskPtAFMWm6AICgcrss3HRl
KipNfiNTm5Luo6LWEOBiVG9pvHl1eouyTKpTafOYzUm+4xMfXi2yjxpFteiUnOxijaCmJLO83FgB
nGRR05uBsv5rHKqNlDjJGiWYRsK30iQP29YT5zet9RkBdDYLrpnHKx3fShXo21OxBgSD9E7ZDzMn
Gj8I7wepUYRTiNhBjjkd09QsBZ5w3yFqG9vQ6GUkNE0X2Sa8LCsyfs8GPOmA6PiMatyXhSkJQ1m4
6M4OlNSustfa74BDqF1TQsBhKWulMAKWaVlebjLTGmNFUae9iNTqepY9qTltB2nugp8sbwmemV/j
lMrTVWQvHcz4uRzlug/NUQd2I8iYQStNnr0XCY37Fb9TcxB/B3ZLNSRcI9efP6bSuT2hijExuL5y
uwDkNXQCDtYF2+8ERvrqm3ljO8pDF7Nn3uzqioxO+HRTzUVkadHUtUNEFxgL63N3IeFT70ob0OC7
BCZUR5z1trhkfxnNhY49BvD1MBFEczxqKrxU6IL6TPEixn5wW1ZSIIwDekVoBU6HmRh3eEeQXkYe
69v8Rw2mDuFsFjBm84HVYNW4vfKs6HmfyFD2H/i5ZZFN08icwP1nO8FZpCSsAtGFGen6lrKBiYpZ
xCVK+kvZ8i8EsvBUh8U9k38ktTDvZXdHfN7Z+k9o5yL21/kJYshjvpjxCWT6B6li6KUNUoOD3SUj
5kuP72TimUBRI02u5rKsUVVMpm6F+NRoHnunNdfpBXVzC0vmeXmCV1d5zoXI6nHMzN/Wki2gvN9e
aKb5C7+EJx1iQvyHFHNgglY8HbYFkmT05Uv7SwAWcSQTiLhD+/rzG9dkvGp/iQt/mfkBsxw758LG
X+ovf0x58tiqf5rt5I5X8HVhl/KkTQLS7QUJCsMQX3xftGs3lIxKoIIAw7sQyqnaAwsRThSfik4j
Odrzp4N+GimDAgJA3tFOJi/+vAPlWrCXcq2vNtZ3ylL2n6ViqowWm0puze4Z1TOtSAYEN0mv89VQ
nbLXJvod+jef9kkitN2yqddFPgnCSVVXEs+gO6UAccqM9RSipj+eSlnmJ4j2AiBeKhpsrmDiIAJG
6HjXBuN7tQjbIeqEW9jibAOBEJZykFAyHJDEDP62y1Zf/ivk8mtGfIsuWVvLmRY69j/v9Vp2HMi0
Oz4CygFKkcf0Cu2j+Pv5GGATle3M47dLzQI7rwkng81SMLuwCb6zvqQ1y68O1ErJM5zKvuYphrnk
qj3ep7/0ArvFQsBirSyXf7MuLMExl9lKW5ACD8bxdiSb7eNZDsisb8Q8n7OAYIAZpRwKL8XzsQSv
2YW9OGSIDFwwUVIsKOwZ3snxyzkFVOzDji1pM2BafXcVXl9lik+koMuhzCrZ17S4glLcHYsWIzW0
pkBnaG5O1zD6FDC5ZlsJ2CCf1uSQGR4C6u1gFrau7oBfGmhHoh4Kd3KAFUExLqrG+tAmg8IzulXh
dUdxn2BmcAO3LAN8F2XX+YWmLWxZFcn/1AqPG3B60lo+tKwqqgmZMSuJkXY+6/aGjRBLkPPYzHco
E1Gvzi7DWQfHRIxXE7fE5i/Y3QLVYUI1zsuhpXiheB3xStPyG9U7NcRGkpXdyOebDxp6SvjQOltt
2vhOW7vc9/z1SOgGA2N/9aydVVyG+//+0NLQrcFklDoInrJCcKfNOAzze1HGIqQhE37jHNC7Yoid
7KOvDeOVKpBiloCuFxj8ttM7bWqPBjsLgIj8dp7R9ebpa78nH79fdGFbdTedQekjuMb4JkrDFlgI
fGJIo41ZAqBshne4/msoSnhrsq2gDKG0WAqwMvWaItBKkx/dM9QsJuJHD8YMoD/tdsqR/6zkWbqm
nl3cckXOr9elUJ0FsaPuLfSBmL4uh453bBXJ7nwoE0sgzpv82c6He856fFraKGiUMhtkwJtZU0es
pbauAO7m/A4y+iA9RmZAGNPiid0SizJIUT/tZz32JTIoHt6PArUwJRLHGaebKc0AhQFH9Rd7qa2u
XegaQlcELR88rVGPu5szQHL9aiF+48KyRu92mwe/M2IcO7mJCMgIjwgWhI0XNa0uqQOJH6ndgOEk
g3IKJIJ6+THFwS9bWDIdehADi9gZC2FOCnQBlP0iEJHMjOMjoydfzPFnDMiqkq39ZU4YV5cRm0Tm
4+6y3VJir2fb2vg4LmO89GDIBxtIgfeTtEZ86rKtkZL2uhCbx5ZMSryOfdrIXE+7kLkCnFjO1TpR
2rWW5X0E8GS40x87SQY2/HcU78rxnYkv40eOm21YHRWIzHnXHLDC5BNpavsvY0LMQVBXot0ZyFA6
bQKEjg2M0JLqo/FWAWin8uJjR68wt6WjrA+eJSwBZOyInHhvWnAQ1ddAbRg95PQh8NxlXr3zWyVw
dT/34QZm5j5Q78LcjJixIAdcSQf6M9lE3yvpdEIi++ghSJkA2a70iFGT9Y/PxGIwFZHobaObcpYL
esK12D035qVJ/3sI0NVNvBQo522qcDSqx1GwFbG61RZ3E6Kno86uuAUmubNkl4NLM8HtZuxZXqGN
EC3Rw3Zb9LIkwHeDhNZOzJAXojSpk9VMzGBObwbz+Y2vbncEftkjd9xBBA0MpLpmYhZrzfk9kwz+
p2mmBA2DQT+mxiY/9xHhamaNOaP2hyynVHAC736Pn+sAErmDaUVslnW3yyHo8VyucM5hBSoh2JoS
7r5vzApfyCEBtc8xq9vuFcH7MvHoI3P6+rGYBtZlFpkmcO2SY3U/rQEPs0yRS+S4g55bamEAhStK
8goe1o06BvHqSCd2b+2v7JJgiDJxNDgHsORG/PPGOFGw6FMyjOBFj99BDM8YCPOEGkyKa7YzHHw7
b66Ei2IyKovKSGAytefNWWTFm8PNILetx+S50LrIxM3z8M0GgB5BgcvbuA5MOU/Av4bgVVIanVtO
DbOFhxNNBwMnIqR4wJSVOM5lV33tXEhYirvn3/lYrI6Vt5UYYeL/o4Wrl5xtWKRf6Fj5nmYZPaTo
BNQsHDDXJUSIw1r41klyFDbySHIyxfuc6l/HLPUp0YlyO7CMkEREQLmbwnKwsv5mCbOilOZxiBGo
ht5o8cHZ4aMi9SLowl0Ivj5urrq3bBN9yi1yyGOJYDt9HOr4cihO5TwfMwPS5CxIKA438bm4MmVk
o8cckl91SmZHFiHF9W0spwZ5I0y9pNH48Ms/ZGtus/KBa9qpKTzVAIbJWu5gtPqOqXpNXEc3XtS1
xSZLzcoRHcE7QFh8iUIJMuMO14/MyG9M3q32ORSaPHK6cyCXmeF4K3RzTdfXcnhMnxI872UnZ48p
4OyGUEi/zuImYspvyR4kZfXXG9OT5A0D3gpD1VaOuA3LZ5chndaju62RjepAfQdVcOB7wjRP5ng6
9kiij0TjCKeTVhV498fki853UVgtAXX15/a9JDSCXvrkgq3DO8i5HNjJP5iMEK0Ny22v4tOcZYxB
zuMczbdEUTT4AZW98xGy695MPznyOKBjDPL8m28EB61+kbzg/FDjeIfZ43NCNccfZBv+MvST9ii9
L9WM05dpH4n0rohLojmUF5DSJECOljd4TbEDIETgSxSsKUG6lkMRQeEdcPgC7sObIakoEzhquCyy
CR8yBAPcPYra6cKqzqY8M5XyUm8rMDVpx9HLCBPEFt38oEy3PMyTp/mImpId20vVsimBD8HkaAGx
j2Z01raV6Kw+VJj8sBja7I5uQJFPRfywyfKFHTSfroyTAAmjVRmxP4wImE3M2I3YDN1euXk5APK2
FrtcOU9ZzCpJ1ntAmAUdzUrh/b6mOi2VoUNPP9F48BJJ+C2sfRA8+Ul0gRNK+JAoDyQXnqZ1fyMo
jidjepWRrWhyagUU96Q+/6S17ysWPjcZreVwTQob2QX2FLM13LHPLyIptnqB1d4cdRT34n9xxs5r
PNySXdVEXnwRPkV35ohXa/nLozStnXQ8zRkDLeEkymU+n8siZPHsIFtZ/HFIveuaDcnPQRwlCcCC
VEekgbsifu6gEKrCaZo12BJMvcqcCwX3n0enVCoi5Jb06Mq1PmxfwBEiTTFqLYlpZNdQ0v+uxSY/
eVafkUYHTGh2WTHS/5aXYjH3WuyeVQRwV2uhDJpeyyl1EwCaGODSgOEX1PSp6hw1qWVJ+H2x8unU
HluhTzlFU10WNj1Hp2KW5L+twfjZczKmWyPp+cAjE6IXdmzU9G+Kcn+2r18LMITUxfn9S3Kx2bvD
sVP4MZybPl0xMR2owKxW+KaPg6pUiIK7smSq1fEJ8JpK1yRF4iioNrnPJ56co1AUwZwaEu4jg71Y
dPyOLKL4PAG9JlDc+jG8TaBcVIbqQu10YDMzr6c06X9I6RfPGd669GrKiCJk0GvFoIeBRdIh0UO3
vkJzLq4zejIJ24nFLRuoIOhvYXY+UhrNQd84POMetI6h2FU+C3miyUe8/BbcLFZUYC4wFQ5xwRey
72e6yD7QWlh//lda+T3N4A0DGZ7KHSeLd80S5U2NzYNJnygxpX7Zf0n/yyi/tX4KqHF/yU77oTY3
48fl33ESITMFA0WagZ2cwn4dqavpzlMuYGZo7KVYk9rQ0VVuJ3k8pmUsvNABiS1kMdEuiKseb6rB
2SX7npFtk6wPbVO3Qrm0leU0Ty8YiKxH1CZG36DpApCbsRPJsUj7jOCP8jElyuu7kEn2AL86vU50
gKcDBrfHs+5DR89+ZETTb9nvcylZmLpYcsiid5GZE1y/2lEIVABXHio1ecXnR3S1bjdjp1Z/+n/t
MfWC9awWcQJeDPQJkbeo7MapzBW8CwBT7rblMgD47MSZGYrbPOrFrI9WerVOay8OjNlnANvG77vy
bf2OKV9b4J0EdYYSKczd0DRREfht1AiRZmJeFnSLntzSfYyWSdRm+WwqQUoW6kXDFfFQgAPQawno
kLLqtn0DpFMlUQMBCRgQZUNhzgtSqJ4k41hGIXfLVObsPHdZaXQf6LwVf0B/qoLT65aax+1yXHuI
Z3cErkdRULGCsDrZb/WwdFz1v9DkkqMbS1N1iQnx/0b49cP/8rcysDv6De3B9UGGiXwKEaXb/D64
1RHJFouQvkGsuSHNhR28/jVkHsj0h4XJWJbagbNFURy+XYYclbLD7KEYAhp4Q0rhibv4LCiD7+s+
ZgFZ8B/pe5JSCjuDHSDhRyaExbh/hUv+VoG8lQEzI1p6VX1hINfcHtmvRguHIqd9HFK8nBOWHjl7
ZApKI/KQypySbT8QHCLY2zQXU0gT4mdz7YAlzCkQL+dE/ruoWuM2w6SAj4Hugk1MzFGRL9u7e4z1
M7rqKf6gNK+cwu9FQ8D1douXBI7jXQpUHd5Tl7SiBH8z3OzkIFgqIBm7mdHb0uQJpfkBnjo76pmH
+c1ppPxtcF++6I5wu5Nc4COdnuugNOjXJYrwG7VMiR+gA4VfvM7+PUhKvDzsG2CKwmLFAJyhGoCI
dQAQ4J7dvg78wo5QfJQyIpdIrC3XI/UEa4Ys7m54clE/aplawCBv+rU6DFG7qe5PmVk194vRfuzS
eg49Rffmc6VUDvSB1abT3F+93CVA273bbBGrJU5hrhUGxVdLL3bKNBNBVBxgjZ/Vd5u5cFhUNrVN
Ml9tmBrKE45T6r5M96esVRPvQosEdaC6PFk3oFoyZWMQ/uMCigqBKyeW/7vvJdcKIwPymIrn1dE9
f56wYreY+/gHmmWJgF6I1560Nusdhozulw+ylplH1x0niOu8eGD3QaLTOHnyPX2olWEKEi1qw0zL
9gu64XBsGozhSwYl51WvtqZG2RAePPa1on0nLAS0RztVjMV0TqR0TQhPqzdGvDi/Z2J3LWDPzwMy
3BZuV1IjTUgnZ22MzHLrnsi3s+jzpxEe5RYMlyz4TFQdUxlW2Ufb342ifwz8k4s7quLcnBgp5dki
1yTUBEXmmD1NBJUIro/SiIZ7Qr58smj8F3BDHrj1F2DgibvSI0QvqXm1pm1hzQDQLS2r0CVP+bZq
/xi6ZJH+qlaI22RQok+oqPFPS/f2b+vl5ViiGD1PXkRJRvXLEGK2j+2NpGxMacKtJfwlfGN1erDy
I6BG11PWa7TDOQ/Fes9FY2hfqvJMuMXI+jY2mbQd2Pu6Vh6aie6Lf1R/qpdkzCWmWDa65KvrDcwP
7IbFRxNu/xTJZHABL8B1MEsV4rlFbwiGsTTeo2jIz4v2WCaUxG3WwYuON970AJ2FiPv2hulKxhrD
uMzp9FJamaa8t2PS1iXTf6nJLmwEKdeSYMdqPezGeBzvOSHeTf8MZ38deCHqkkpqbGe9Bi8UCyba
6W2CROKpLhVFlIxyyrN6Iwq66+3MRmzu/Z3K/7y7M4D4fv3D6CyN0gw5mRC42M9x5r0gRa8hxtjJ
60IbNz3y2Lz11x4wYF6wGT+zks+5jSNWKN23nEFY1obvkGhcX2vrTK5vaL+ZLLBLqtmrMd2Q0tKU
PrIduCRSdd5Udky2iIOaINzFVbGTjjDjpTHc6Smgwvoyj2xfokpWpTMLlAgCR4jJwkAF98JKw+WC
tC03anvHz3AxdjYK0wZoQSkoW0033/jF1wblqVGqt8DPxfoNc1H8wLB6fySQXfBOhCouZfyP8ZLR
AcVkwSP0Q1C3P8YWv+d3Nnuen9+WTHxUHOIciO9Dev99gAg8DHzkHW3GNESvxf/4O6bkG8QBmzKt
/I/td88eV3QFTbo/gG+L1Ee9edKH69wLkcTReGKeKg0bh298VnzNkXwSeD38c38SpxdvlDc7phX7
5lKj/Fo2CRXDBxiEIo3+ad+s5isIgoyz68xY37x+ro7Enuwohf90ib8pTR6GFOXGzutE8ioqVLLl
OlDE9RYw1D2JPz6OkxMNUgB1X1YCE9OBJpJuF2Bqcr+P7boVpos75vgMHdI+V0YKkQqx9sVqQLIt
dBNQ2sopoS6lftOrknfTmm09QC/2dokyzqqMrTAr1nU2a7ndN24Q5EyKGXZR1XpCbDR1LtWoHBDf
lQZZIaPj8/8OAELDa2ZWJRx6ftJYgfTuDPWzX/5Tfw9eEGX0OPY8Vo7HGk9mPAlvsYNdw/3TQreB
n7gJXRYzqCmIH8gXRKaStYu9mQcsrnUThBZVYfLb1fOBhSN/2jaUstzsh1aVoiqoNqcjloBopcnt
1jpgM8eTnRUA6arIgYIYEAzaTVnr/qpxSJrZqV8z/mAeKZr/0Z/oQmE6ps6S+C0vngaMG7XG/d1q
BbWjNEY5V7U+HlCbYXSWi8bj/g3yJRMIgChplUDWJhyH8ZTeHf/XBY//quyUQ3sjKcYB4yMQCYRB
EBf/m8UUwDiSRMc2HfUfYSqk7pfWiqxxdR1ewHuTXvCI8HtqXR2oXsY8GhV2JtPL3EF8HqIAeeXO
JagAkAG7S6RO/EFD55Kqn//ev/D91iVDDYbk77xcyuvg+R0vWJrGnpc+8LD+QptVD9n9wbofTlrc
JiMTjksaTxD/1woPxBO2Dw1fFCKqHRiXxwlJUsZ1bM0C9UpEVWam3Wsu57Mu7WWa4nhUiQT2LdTC
x+BG/7ANRul34l7NTZM2jmQ6yt1PfXr+tYv+Vx92/oHkv4Sijc+AMDmGjtRDYb8mnXa0pDQFSvjR
lMrFNnt1VlrEdpuZIUlQjKNGloPtx3/g2jBeuC9TK5qbCQARIiWX4VU+C5tXzfsCjOBmJ2nmV6Hn
/CsEa3JHT8NCCqRKlfdZocBnw2Du2GX4FawJKneIncrMPe75nsVjv5Bbuo8u0W9pU7rWDiytKgy8
R1UrpaO1u3Gub2WHvwXrAr33C6royPQ6yqCiG6xtcn1EF5bp4iDti9hnt6vbtONYsVwhcYR//5GQ
5bdybDMdhy5MV2YD+aLwpoCHbNvja7TL+qPQPtNidnArYqGKXbQ6MXI+j7y4KnREZv1+euqMKdSM
ekCaxfQ8yQ7FlpdSyXmwet3Ss6zGt4O+zQCdiY7p5cLEI3Rg+GqQoot2xm4AyBkPSvz/UXv0v1Fk
EY7N9FFrve5QSwUclrrBFyaC3MIPmo0mIW0X+vhlfEE4iXOZB294OFgd8o5y4Amt9vxRZc3NykB+
dAYfkQ/YtLQUGXgGuioY4q+YvnZJXQ+0E/mL786cWO+vtygG9Z0hq/1wPzXpf60QbGh2IpC1IL2k
sW17c5hkKQmMIU0/UvJWUcGQVEqr5AmEh4CSgPgqz+ySgN+/1aSxplG40D/nJX2XJ6paLQJyZ8/i
f1Blpj2rtlgXqo7bHReSu//VS0VdZ7Ef0/lW+xp+7Hi5l7hAsgFOTpC8vRT8LqgdqS6boseQde2Y
wwTcLA2lkUfoTjo6YumDQtKYS+1J7w+iXvwMEpo9xtlV+MTmGr2y55LDWSRXYEYP82teMU6MbmYX
c1s+Pyw1fcM8nXD7Id7ZPiezRpUxShD/+XsrpkoVk0UmZepXhz53kn/0iHKpzt+DqCAm3CfjKWBi
3og6I1GydePhKqniQLVmOqRrsv8+eKqmYQPwpPk+FeXDxIREU9PPoydYyc88cunAe00yL9TKA0Bv
p/xRkSq2wafXqL26ccZSt2Q7bwy2ToNvCobBZLlQD9MxTOQukhME2j8otM38fHxvTcgSOw5HjKq1
0Za9PrB3vWV3mBwtfp40QR0vidm2/c+kxiosW19syB/wT+32DIxvOYKZxqH9awr7FH+6xgQisB6M
8NYsI3gZHQY/fpSGnWD2bHblBaqaTpEqeyFirH720HFRRPfeGWSxeEzzou7yg5LK7xVo339IYY2+
jKiHv7x+ny8fTympovpDR1c7DTANkocLA6KGacodAxExRQmazMCYkMtnF94SnuM5SjngfXRpDv5+
VsXyx/R+bK0hQgatP0yZWCohLr3tdCJnPFZhzrlbelhnotFnHavUzP8m7vFw11AysJqW9v1HQJLb
SjXvO6T+IJmNeP9bbeNPPbec1NP2t26QKqqYqbrKaUjp0kwGHMxY7fabviWWATz+ZRvEzFOpOHrk
ojlo1s+KtqrFmR/QGSE42X0RWKlgdJnZqu/05IRk6kL6TGqsFTycp6G/yBQE/rNdP/kniI6vCdc+
GfcbPn47BPUWaROXeVy0gFmDcirB64nb3OrkGu9CKa5EITTjOfjU0NrbYdnUU12Y36GqMUqPmtHC
vIoTpp/lmoJU9VEaH4pKoO02xx5cl6JzZG+MmhmCUJ0WYgJYSAvshunYFxB5OSKT4wpZGoXxUJtU
1FpfCn91bboRhrb36UPTPaKrLwzx8cwC6qmMcWMQcEkfpxtCyTxDJ/bIEe4OVKHR8VMehLUri0u3
LrOETh4XJlAfQkBFEmcp042R+YII0BvMmrlORkIJHagCtEQmUs5mNVCzMxrwnF3SPxAbQlThIIiq
Xu4y0AYZKYTkBPtw8zKCN6xiy5b58mlcKMVHCnuKFJpDfB0WIix+XNcmMggtz1GhMB+AZ+uwwgQt
rG0VSE8eGFa0561OIQSmlJ9az+FHPGYSRiDIZNNb8sDnjfxsS8GkgxnwODMEjDkgTg5GfqayJHdR
q9Fn5OVXa/VbEpmXGxC17sVViT57PI4HS8pREaXNBSfFuKDaHDx1avwjpRTYtvxX+cUBC2KEVSPs
iiJq9GDPG4VW96x7C+Oq9ousa9sumETfLYbZsyZZGHxJbQ4HnSLDrEtwXWw+3VSdLCxShVdZP+p5
rZjxaeXdLquzDMst7oPzJESUd4IKzrJskmCIpxYrYLM4c/Zt9oWJ5FeauQb1foGxegxVHRMKr59+
iSIGBtGJWP25TPmjJUBK33TX4H0DNvVA8TlgPVhgaUK8aPYUM/orGBvimxpdGNuUtiJiPNsNbBcx
lenDif5LBTw6WoxlpakfdMkNvk8YvC6pc9bsHkQL5RdHGiGjzSU4Or9pf4aGPS9dSMAzGFxAXdyk
uQne7/q6jdRkLb203Z6Ob/h14IZ3MXqk5JhMujUKQ+VMwOnqnH+ocgjO8pGcVNQPiQh1YGLtN5Wo
oURT16ihBB5j9MPjrngiUES9o3fbNSSZ1hbzcxybKj+cHB8uDCqXC+19dYx7CyLd/z13g6nspT1q
xbaozbgHdgk4ldqp7OXxP/UXUK0x6eCuE20uNasp9IHumhrZjxzI2bBtcCA80Jv+l2MXDmo+XNcU
suv7JX3qSg1M1W7DHuRxdlkoJfkOWp75wm4fWDuq+lvv45/zR6kgkYie8HauElUEUctXNUP9GzUp
bvhm70AXmbCQxYnZwdxE/NRDUBJkz3gi8Aiuvk6y5yvgwRXeIXX9Cl6OaT3zBgFRX9JD2KzcHLL1
TBO7LpjlX/NjWviMrn13leUnyGYPDMRSiRfdyrgNGszFWfAqEpFzt/7AXyPnnEJiNoOdmyLXY75u
GxuZ+XV9S5W7WGCP2SlreO4lMXxJB/w71C2b3Fge9EoEDk/DXXFdyBazuAzgZ+6KVXsjZZjvYfi7
XzPNIk5QdzTilL8IEFGGNVsLSVcqV3FKSqJgoW5VbB0up0TT2IFSP4kcnmeFlZwpKWIsG0mUTP99
GgZ974cYpkTlnc3PQt9WPW6ogJsyLsWtYt5XdZcXDvZ6ODq2QqvhZDD9JHiBprx7AKtuOA/zeox+
PQiKxOw4KMwSZJmuCPUHIvhwJ6eA48kb9b+X/W1bShsVS9e4dWzN2WnRFd5raRVXhm3/ytcbuEVd
CyJxojv9FozLbn2pVuW1JGt4INT/bcN70TDfoiThFClNC9XHVhQgwM7dr4OL9f0ZtBSVDQg+yUsU
TVm82RcxgbXWAa6l0kqLEqmRotf+ihrrrqht1eZiYGE89Skwy8mzCph1ip8I2rBenWQLQqSPMII4
yN48f0EEJYL1p1PYZe3Jk3MtYGhOPCMKPUmSe6Vb3hhyLOeqrcxogoXht8rU5rE+/948T7fYgkHW
Lxw9hUc0g0qFxGaqXDw0Dzxke8SX2i55qW8Rmmi51ug8UMwtvgfAn6DQmASK2/2QZjJ6rSGqa23l
PVVRbAJgh9FjNQOrcgdxsN/roNaHFxftil+kCns7zXFXqd1Q3lyf8C94hjoqJk+pGB2TZeWapbZG
dHVsPwomID2NufyApeiHJWsw+crd943fc6sSEQ2xP9nDSATuELh2WfTf5rGQqQU3Z2CLek1rmGkN
uJI8Tz2bLrctJHEdxS+2QCKxJwjjsQQ0j/AEi9IYUqTE0/5B8sU43JIrDoQ+xcZ8YQZGS/akSg7+
u9g4GKOCOgzrVkanri3QTJCwnujJ7+kJxFKj/z9jY1S3cK6kTdMFb2Idns9k3vAqKvMVdz8od19A
WUmG705N2YWwdDF0D7r9FD8+08WhUiUD3fSG5B7fSE9xiIbVzgmWdNv5SMC7sqNliYB2A+FcYthd
oubzIMGkUSvfbmX12NtY89m8hWlIKv+aBfb4T2lqxQsoItGh1e3l7SaDQ1lxLpenkGZeBKgDUQr6
rSY5jvDhZ7rzLzQ3hLpJotQ0g5q4bSP3ApzWhqYLSJvCVLV4AFgrGrjcgk6fblfFw3YMRzGLuHfz
Orov0P9dpeKspUyiZJohGdyclaZb1cRPsGusiLpbkPDk5hIiIfMsR7wjLBjVaVVsYLrjM0UycoLk
2Yn4ctx8gvNznQR8eVTGnbqqSvILrIZe2+viE1FiKbG4vu42pfiX5lMjzR7i7wr1K9yz7FKKNvGA
RsP9/gtHqy5CQguLlytHXE3jKzlzuz/u0Bb5q14SKTxRXdbiyzqpGAYHTQT+4tgVbI29nzh3fXWI
QuDOgBi3Ie+yH+1Fkm7jWheCV3Rmtd0+IQ8mT1XaMbuZ8jQIxW1iO4cLi00qxQyzr/3dQczA6acN
H2yxm+kZn6PWdTuTmuDfAxzJED9nUtmF4vwPI8FboCnBkmOFJBgyHCaAKGfJsmPQ+i3isyFQKaar
YjH0dgDbzFSqqsstr+dhCU+iLA==
%%% protect end_protected
