%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
qJ4Ep7SYsEk5sMQHv0EL7qn3iDzNexhGkI6YkJ3ah1y/OJeMKAZxmAhN5vecgDDG5tmmip/yiNBA
5GPhO8Ny5KetVjlLX6EiFvpxcJtauo9Nw4/4AtkKtQKJ8Y4pA6R0TIAvtHDfcKrYoAkWTSUz6rwC
ivPO49m6amJMmISg4mcPMJkeWlwU6aQPMIRvAUEtaLlnpDcFccCXnChZm+FSNl2nyZtWNhttUQaj
h5Eoicp3dsohNACSqW8rUNUijro9z2SN6S5U0PpZQ1lNNeSLb4zIAiH3xen4boF17wZ2ggj7TFGM
GwljSYaou5ZLmxL4O8rPUiiJPckCrkTd3LB0+A==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
7xfQKKcRHsyvH+5Fe2ASUqsVnXoi4NtCOvEsDf68frjhxEfxKtgWDNN2E3/TCVe2DnGLrSzC412k
sGwF+869MSBpBa9sXPZ1Jv99EfAY2BcSWTBjg5tI8PQy83YLi598dolcd7acNs6wWFSt80YrGdwM
pRaVjxnz0eG6E5Dwl1V8xGEwx9LukkymLfoaDaCGPDnkzqTVHMVRV0byfDbjgS1jm3vLtH6vz4Wm
uOWPb7+VRlqnG84HskCk3tsDt1xU/NMFX2AmqczO30tJ/gx8DGiEX4ycia9boff6ZECWuIjhkket
NY8vrzeS7jVFOfGv6JlovQcLq5Q6w4sBxUTkP0FZB1Ur1uy+Hmhu1oZ14dCGVNywwsATen/CPhaE
jClVKZP7tb6olEBmRkQKNVn5Bp2V7b890pghE1I5EHe8fp/IzecFNt6SjDx5hHcXRoqVo/IhTLO2
JsJPcscHS5WFb/EfLE+DcaHIxWORb8QPe/nxKOQY/O6pnZ2I2vNoku5gSIARyXDDisQehkqaJl/l
G6nusxf8cqFEmrrnQBFdmjA7w0HUt0pBvFsqNJFCQl6zq6jBfFfydiu//IE1CWkrUUo8JTPK3Lxw
K3EWuQW0LTKqOPQ4Tl6Xyxse5iS5Buf9KUcNqD2JjmvDguEbpxzcYz5ytnB8Yd1fpYfQQ5IehQH/
okt1zVRZYmhI5nhDdoA+vQOUEdI67tO+E50orJnAz9dgpvwCDep0iH7PZU70eVaLK4QVr48TXpFI
8gbWcIOEyuFcykeXlMGrNXzawqhX57sYyqyCaKiDSb7FOhLfVBdZfx5kL71YCerEzQVBZFL7uxnV
SbzhWlrKdUMUwKq9d7vJGVleXCqEADqggEfhhGKwjf4/CRrMeItdvtK3VQU94ft81taN54jUUeqV
sByWhS6m/y6/fVsIjY9MuKd/yAdnM+iysYjYWq05QU+pKuc6NhC0iVATdyE/gVQMyUG2L66I6mir
myWwCTVIAe3uU7rkIHUPuByyprKj8djT+eUBWSxeGM85GYhSBnOPj5VNALV68qoHR9/MB/jc5l7H
OXsiL7IL2dIW90EkdYK1TBIet0xc6j0TuZ2fKvkyDmBmId5H1HOvqzHVcKFFhffGtqsqzjAi2n7c
+fx9ZXi+fchhBzb362jmHP28shitnjJyL/GemBFVhQstELW8qU1gjmTBVMx5uS2UZPH24vmlECrH
q5WAqJEBtdivspDdwiJzd/mWiM+pYvy4xIdFOvWfCXSpE5t4vjn0lJw1gtqfr+Q1CsfJBJPOPS2h
+9HvkRI536MNDcoY3O9uAr5bLiCy88oLjc4ZaJJF/eP3pfSbEl+SBTcDq8ReR3SIaXk1bona1b6W
qE1R81sgosnY/+mZkSfn9rvL9vGeBm+7iLUDRBIUxydINEH2bR+xxN0Wrn/vY34P0F5xOMpGWoDK
sFvbLVR/HeIT2TU7gcHuuttBxBALfVFHafHnMa2Ay4vjI/jrbzkdGOlyPaWLC5J/pXbBllzJ29IM
AsZspWKKx0QiO7GN+butIZ6Z+5F0DL6f+CAkRhg1k1nFTEv+I0iHwnlBRH4vasX+SOC+V3tPgPI9
p/kKmby3tbVthzKrTE1ilzEewMymXZjVmXgrHtQDM9hXPFzCUl0CTtkVHjxhK/SXy80JWq6hha3X
mJCD07S4b3p8e/Zcsg3OP4j8AFIphC6FHZVA7rK0hR2zjbr7Hr5Y69FVVTDengIbsQ3wLwLoNBc3
g+IdVt0rCd/WIViNIbB2AvlFVKzDjvkTpYpnWin80FNFM2d2Ze839/yEkd+fJB9SiAbCPkOLCXnk
sY5fi+Yj4Web7XLvp/rNBnprRPkDGKHBFgyLwv6Uk5NnZB+k+8pJ4bsXCDTfgDYzGxV5ngfHqjrn
wC7FOrVm2PEqJDNfEND7zX2vihAaOeME/wxA24RxU/3ugtDI0WCCzDAD8yedkW4+M/dS9uXqD8VN
urc4hUHN44pFF4K26d1MfaZGRbz78wsHLfR/eFOb9vXHelahTIl9puQnKqZmVJMy22IWRRRPs+01
z57qdCHIHzVu9pKhJ8CAqmmzz9Vt38xqHpnFY/ovyZVGl6Q72J40OO5Xk6fTY/8rNNPM5wvcJWww
Z5YhxlUGK0ziURvVIUGqm/J7ONFostK1LyfE5ztP2/NG9O0BtUl0mgZwH7AqDy3uuEDDJVWPv4+6
bG5tC3xlNxtgCetZypZSO07RLlJJa6wCRmYXI9Y8AsfdzRxuTAY9Nwp5btUnv+q27yQdfq37YWE8
hVmZTuTiOWPzpZ92HCBlWLDJKX0KFSeN4/zUNwfluqnyMQNcrHzTFth66IJbsBk9vRTuaTMO/7Hg
PvgqhYQPx1jtv7jxTsCmTPbPjgNAIG8y2Z/ZLKGQRvVimY4pJ9hCe0HyaF4a92EyN84NX8nn6rqx
X6VgMTymYKdP+ufxTuiaiKmEO1k4FhIGbLTSPWy9IXYDl/0D+E5jtrlYzjVRyMVPQHGLt5VQB530
O37TBV9YyIdG1Csea3MjJiZGX6THJ7+cPiIyEaaejS7AvWM79/1wFQ6c78w5ZGEm40eaJHfZ03mt
kNX0cUVwceYBFV++T6TlmrOz3CahPP8t18wMcPnx8ZFjK8/JpQLiWzqNQbnX7/QP/G1MC3NVpHT2
amP6AfxWXX/kY+wKyJYxdlzavwZbt64ADg0Hxh4IxHvzNIqmunq8Gyr9wWTP7RuvTBJ/SRVTebg7
+1UtcfHG4MGQcvNPI9ZSUOf101n24bADQstPOVfEOtaM7dgZXM47PVclUdoBqalspOz95vMJ4jMd
od/mUiuTcpU30SJKTxSdeVwraYZc+r/FCpSjg7w1xwVlZrUvkPqZy1oBrE6D0/uJsaLPSsTt7RSG
/R4YUuNrKpWCut0DfB62vhCAtJ2Vq8RTPnZQD+Gyq7D7CWoCTBC2o52dt08VMT0evfmpp021JTo/
94TF5Yg4soixMasHShb5AU4QYYMKe1qpDpWPrlDcW15+5hdduX0JEv4ePGKAaKc71akdkVDDoVDK
eUC1vylUwPL/UJ/3FRCXfHM5iJIh+PmuMjq0NiFkB+AXJG5I/8y1C380WScoH/cNaN7yWHjHQu7D
Yjbnhrr1t28200RfeOB3s3Yx4t7C6mmny84do4X+pf0uR4/BSXMCr2dib7tuVU+n1CFKYKZwmB5G
q6Xef1T27wFzLBPNfi6MbSDgKsh5XrG7eftMA2FXrs46bN13KVIuY6QbaB1e+PYL5/av/APZXi5I
huBS6PJ5bqReCvqUSPKuscvI/yz7Y9u4DBuMeyQw3I6f/3RuKzB+5PUAx+Aq/8lUZLV0KYr7nuEu
ZxbQZ/w9579/C0AMHVrZyyeV3ELvUcpg6bCcAss7jw8j4sSusSEWYqF9k6XxHtTUSuhYr3zTpDJM
IBcyRfzeaZhgRUNIUdt4gmCU/tmXaV7IfJk3DfDQQm5oG2S2as2SP4kPmZ/6iTzehxbFRLJNQUoF
20vng+URcFd6W4vrHYfNkVomPRd0LIQP7jSMC7gJ0WEAzGXdEm9Aw5JZiey7sp3cOMXzmRmcV13B
IWWVLr8x/PhmURSim1GVjRaYfwFBnDxXEYMfpAf+HTWojvaBJ3X47zbi8ROqdkPE7TONXH79FFXM
2fGZPLWRaHpE9SwZywFDOpb2q/j1WpFWKQm4+zJD2BXNXjj7IXQj4Nwm4Ttu1NGxVxIb7BZ6Pgob
OXc6pJGFXM8FYj+gQlwKvrX09sCEB2bsULvPdRT1hcbImeaQqJuxd05y8iy6fzPLdrS2YDa6qMcz
KH88LX0C6Ngc1gxvKJ5tAmULB+OGwHXut5I7syZdny6GrZJDF/QyKtzC43fx/fxqWedpbkfU15sj
QW/XomZlrI/5wce4AV5aB+OOm/ONKaJlrrd1/VZ6FcNqD9vhgCjggKiuwqRCVoO8EOJ4sGJcAsgD
KV7evquH44LpZhHnhE2EXL7BCTE9uc4k8LP4D+fBTX3NB5NimXu14sFIuokJy5hJT4qKv2XyZ0g2
teFuCfDc7delSvU9EzbTYsJjf9qH1RcKR17kpaOvDN/lyJOu7BUfMBHzLIcAUE8bWT4o0yEKO55H
LOLNUuqHVl4sMnLkl3iKHRZs2bZb0gEK9Op8yvHfDC3CelfncFv+QKBMTCsFQ0QN9pIYHo2aXN+n
H1PLB1sed7efmKOZPUNgq2Ds2xNQG/4kDo5FHrXZCGrlnVsfp4QWShKmvep6htM+CYS0OndBooai
7+L5Mvisz0Vq7ehL0sAI5YYPCg7SF/6Z77/gxSNk0euSAbPGwwaBXIysZzuiA6a02YQPYFqGYtlP
gXyFjcQ4GFLUaVWq/wyJOdBUAQRvO+XSvP7T136ONp4GUqZSss5dZHXBRd6JdrQoqhEGsWUQZFQ7
jmbCruLGeKecW4S+7nGgLVVLh1Wdre3mn/r11bOVDtJUUSBSTkynU/s0B9SI41PlFfWxm1NRr+Jw
9wdOW0ku2oRJhaX6u+a5u8XvZzTVxp+RZtAvRHoPiKJLgUwHvJnKeJ0D7IMi1Oz8H2IiFbJLmEOx
Oa3dWzdyD1w/WDmbkr499wsQESau8iMlI7/dgtrLn0u93yNA1xLSRCYk+8JWxd9se5rPkX5lBEFu
mM5omTDbOrWgRqXq3BKook4nKukaIH9byb3qUUNis3rkcayktqQejjGY0UqBkvMiDMgUBCo2fxcn
EtawHzXVtbrdZYcfNGwd95xejOyAUqjRWHRuPq51PdGiSw/fetdMlZhQibu+8SsRICTGynUVMtrN
nAbtHFvqcFRIkJcRiNFKxBjE8uSbUd76CNe4geL1jhLiXVr0fsT3ZSwdXgD6jS6UXI+f1mfSMfV4
YNtXyNIn5q0Kq6rOfR/Fr84C7Mbr0+h1OBhC6RKRYn9TilaWgwCYLr6b/eZxdoUJbAzOhtB4MAKj
xJjo0HkSqvJfoCRscAfiNWqR4Gm92T0xOFQXHm/LyHz6Pqmc5XJmbfSY+NglkhrVLOR9Qw/9iFcB
ux8smOCkp10g9PiPxJaKLoPh/THdPrVo28dVpG1F+icUXUmP5hKVOOdiPfxdcjGNvULaT8a583C6
cIAF2c2Qi4vpXzeybgL45b0wJg2dq5B86MEf/qCLWQ/WWXPa2KqT1Uruql7XhAPgl8ABCNI8W8fI
0YfutDTR/DrKsOerOv39cCVWdEwWiAGfb3hetpBbyjXkK8p2x40Q/6HS18dEC+r6oBRfezvEV0gX
NdBlMWXD7HrM8uVQBXBYo0M1UQLR3GTCoQqL5CvG30G20KwuqfzcXMUePjrvPI+Mx07DRHTc2rm7
u6kef7wIZ8iyTk8AtzXPmVwQBfqYZy5tPHseMrCHBKSj8e7NRYogUziAz5Njt9xBpX32fCyFLiqH
WJK6YP4YtMWv/qn0lZbL/Rm6pFopdLiioUFy36ET5g8dtCKVEK4HubKWxf2k5kfQbJAtTDiu6Ndd
TU9fqo1MghQxzINZHVbbctna2OcLhI4vr5WIXsnDwdxNustucaTbtTP2NIwgideZIQ1tsa5xYS5g
iCt4r1x3aoPPZer5wXEZTwQCBQmTStPRTXYg6+q4rbutmsvMRbSsExr/Fso73CjXtd9a2aOTk6KI
Md5gXJPa6AN4vfu/j9UQAPf5wiA9z71E/CzcjHVdQJc894XHKwiZc/RUChaF95OFXJzGwCIx3hHv
I50lTd5HXhH8Tnn6R95fWrQRjJPY+kVgrPxcTmeP/zNvK0+rJDez9STGlTIhVui2vHcm2w3qVS1Y
ZgOjy3JXb/UaZdm6dNPx2Fd4ZHjRai6RhgK66VomaBhZb9OZlqUup1SZvaU1Fw0bG0gO0VRX/h++
01Nib/6astUsb8byvWV7690EZ0abON/TkmTPdZZxUg1EcqwSD1ir4wQ9BvcTfLGnQPg1Fp8hi2UF
KaWohcIKiEJV0LnYBUy84tS9OG51kKqIq2d7dL0i0Tisi8ZMTNhVdtNCedD88jGOSaUs21jjHizO
DsJgpVcvPkxyLxJTWYGtmJR1VbwEYKGjDuIPl/BbC1so16FoIdOOgq9ZhrmBkfV7W8oQlh3KiruQ
obyJhzI39stPeKLjg6BzqYKMvGw2eDXlCehtfoS82wtpsWDOi4smLSMtC8sn3nXZXnuUJ/LSsok8
3LHnTv0R/rP9YDT8t5puH34DqLREoP5IM2nfI9ymAXGYRO7y16mPfCY2sjPekkdguS42H73yY1LR
wzBPK5YZDIqUx0vLkWF81Byp3HBleQjgMjoaGHtOw15dwGht2pO1KREq3VnARVPO41NwYMv2FAfx
3++puk2mchOa1WsXD4GhbtoPtjP+XK1TLxpX3snndxDHhGX1kM8oVmOLtGPq4+SY9JJJWUrWw/Fo
nAghboFJfLc6/ihQGKmSmMJSnrPEG8rgPEUSiJLKUUK4tgRVPPtDPE4fyA01Ow0kKC9KPU0+Ywp2
0mLf/MbfwO+lL0D3iuq8gJ6Ghe16c0RIPknUaTd83uDAJEfwVpLM1PvTrzhjw0+ekdbS4KO9IOaM
3U8HUPRUy6HGyBVxemtlZksbC9BINKbaFIupPYfbNPvKYxLLL+yr1azeEnnNu2FN5gyVhsV/BKE8
V8S99PcgOAr5DrTKbVGymRvWZnse0LF6hh5NU8n/5GHIUcSNOG+Y3myWj4Ae8+ZcCq6nWiWjmaFb
tWl+NjjaLFSnUa7FQRnTVlfhpsihkIkBclNKlneO752v8p6jPs3CrKswan1a7VCa5S/lKXKXCkGC
G/kptVz0GhEY5ZyiLW5r3f19k2U6H/xnRwJvXkQ3ZnU3N55Qb6Y2tDy+XjVZWfqmomjL5binKLpd
smjFIQjGNTFFyjM3FmQ4JZn0nuB/Ka6f9LPU/c1+C7I0FRhI4tU9U/OW7V8EQeLZip94/YcLrp7j
/y5otfwO1vmiLrhTc4LoYOjY4vrzejpWz6ftVQLKQ5saqbr36uOKK+Zg3pIETUxYRIz1iZxeavTx
cL1ULc4rDbFPfIR+sgTxV4lc39xPcbMUwrJ1lhrk3QoFtcRwKvRR+j629n/GxWbidETtiYtqPm9C
J15N45Qe/MHqeI1xI30dXRZH19pKlNVUVzeHabQPP5CX8GpfCAjU70W+7rdOZaEr3UpvgDkHAGUB
Dc1m29I2uPupEDoOGMRdOWEqsZNg+3H9uKt+R4x3EuKdyDK9ubEX53T1HRxm+B3B90WL252a5a4K
bgVZMFLTbedj62bFJgoZ2DQpz1OxE4pxyLRUBkzN9Khky5AfPZhvDPpU52vpt1oFgdx49ArPYrxu
Znsx6Do4gB2ZO6s1ibCKXcSSOp2hDEn+arOsriLvjG3DJfv+ieYW/Q0RD+eYbCvUFRuhXmqONzdb
Eq3Q4bMr/BQPdEJiVRE8EtFqMhvsqFulu7P1ty+32R3cN1qupGraQAuDdAkTbr+Uex7R5x8N/gP4
Rf2UNQAdS5/SllDdTcBlSKYKzWGPEQdVUA8Pbh3DZmIqAUgR5AqJWwo2MROK8T1+K9lgOKg4170k
1PxTlooNH/ZoZLfedI7+bnJ9o03jahHa1nNqCouc5Ie8UYi53iZhd2tjGLavV7px59+uK1nB/uQK
xHUINlEtae30fbtZVhx+tNioQGnP545Z/MvpyyJyL6JhDeZQ5a3q9kCFu1VdMqHVrztxgXZ87RCD
3Bzcs32uozEAQYOYMYulLMncqwiJoMAak1c5RBnGrYVyjDHLd3Yb4w1k4FChtSpZChBICT2I+FHx
ngGVGinnGHGHH+y7Z3J2GvpZpWyko6yQaqhD0vSpO7MQO7CD+fGJOHi7YM2MLUgQtXL2iuPZr725
wZ6GvhorUt+1iYwzkcpPDhfeypBNZl+GaJgMXpPJodv9uqhpqdgA5R3jQFX++ZHNRgsTqLnwA6OU
9MwOjVjkADvqsw0Sz1YxDxR/FlBhsB1PT6OZqigPBls5Ujjmg5IoN6pu5QxXGP0BqzTwO5HAOtUX
793f4YwrM2xwAn2dcRGbXtudiHQuzwWLD1OYnFVR5xhqbNNeo9k4THvzmemkDhXN9tpRR+cbopf4
Jc3IGDmTL3DQWaVyyOd34kudtGz45neFerSXimpCQyL8ENezKiNjycaHj0YMWeBPEIVF7m5+mrH7
dhis0F30nGTc6Rk8vqGGy/+0vNLpjS+s1nAaxnDpo3ydEEmzeRBxU26qIgltlBlzue9UMvsNdL9Y
6p4dmVBt24Y/iYNcbOjRhIK0IhlXMVXMGmlt3mu6+ksCl3oo6Jxb2ZzWfGTb4EAa6dWUaPxq7FJ/
gpON34A82sXhqHYoenLgXME+BXYOXXpmNYdDffRIn+a12KDj4ENRn3AedrDVRM+ULUy9MNfyyd5O
XPH+MBo8V+fGXFhwSE+yfy5NMi6sIlKEVoIbzTcqYSDeur7V+3S88/LkfQx6eHf+in2YHYLGr5Bt
5QQRXb2D4JsTrHqu/2Z/Gl05UjYveqq6ddENnKJlYzSzLTNV5FL3Frqd9ltU2txRKdgsyF1w+Fmp
adIk1mi7/4NBsJx5v5xfMZxoodL3ek347xT8RMZaQ5Uq/6VXOr2UEhjo9PK2Hr5pn7Z5Frxkz1XB
psuGNPvtDok/wMhj9Vll1nv3mjpGwBokclB6QN/oktZWoJmOcx/hgSliK+6eY4GZXLdQNPTqwk9b
ALZkf/NH+BFPzhKQnwd3XN3z/jEU5STq4drvHWNdSJkStMjrwn4Rw5BKZh4ztqFx+NhmF+Q1Aeh9
wEoE2Ni3zDk9zzILh9seeAuA458+BVPv6RxVwgAaGMJEIWIRoP4UZb0LuYoi3dmrn7TDctItqxMM
smOUc8PJT3OY/uNO03kV4yXI7FovPBlxYMBf3VmCZFYS6ci7RCAjDrMOhVAaab5d4V6NewFWIJhh
VjVvXXtahoEJ0w60jydCvXeSZWa4Z8XTNhr1WvyFSr8O8z/TJzfqs68i6oh8ersQuSyQRPTa0WRJ
gqcLsbPTMExcs4mzOowQwMNI+mmaS9AjLUZh9ewMlGXuT/DbS99VtHsOBA51jt9t4RrLRrv77/E5
VwQAPBXDxv18yHANVXoFHSlFZ60yca32eG4APOHNTCcrcC3x1Dky6cOVYxsHJ2VKmbcCQLkLn5CF
PaxGeocZReksXPxJW7xl/6Vvz0PV3Br31fm6E1AqzNU+gvJyCLKELu/FXLY02vr44Qr25y5xvKW4
cdclzHTHfhgnQTIoBYaktSs0KEVQFUXqrRUDXFkuUbGLfxnLGKYx88gmvVhK/kbfaJGpJ9jrTlms
FPfZQ+QgPXXelT6aEgPtrrZTJ0z96lQlwBw03zkLxCBdLi5xZ/jVA1+RwVI/a0FJa5Meekes02L0
6bOmEpcwvyRqnJF5s/OEi45Obu0+kmerIxZlkMXlB8SuZJwc1R4O3tt4BQ5V0IMzgku/hj/byonR
PJllRxiROMaHB0+QtxCDSHntWpCiN+r9HqZgpXLAGMwBMYp80ZW/SmvAN7NvfWgIUrGIxRbXATFL
JvpG2OCatdqioIutgTEaGo1c1k1PypnaCGBDy4gkiqEL2tZJ3GkDheCU+yGTGO79/cFUaBsTFZZN
+WSNC7uWq/WTl+0dJMBDSIdgAXa/AaWIz0INkEZS9N06Jb/YZ3m4OZHvAgXlkirtKb8vXvFwSu9j
uV2/5RsFQUycCYLt6s2/8nSdVjS/ZLvYzPAIwtePPG0vx8e1YNit9/2a+3PsL1vz8h9/zaHNDaRQ
FSKmc6asQ/Psq7ZDYHqoJkHccMR3jvGAdKclKL+DxueOu0odZyklcX0t+ni0+S7PCHzHR6/Le3R+
WC9viBPUeT+iPt8m400TPjU/UTr6pbBf7MO4pOV7ac+G8F+LKOtlizyhBSv8W2r8BqZgf51VhMVx
1FUk56n5Vj5JYRtRG0waEydraNcmvLfdTgejjBo8MWJ00Vjqw1MRonaBuyosjrGc6z1dItKccXby
d2kCwv3h0uNTYDmXVdRuNUHzYP9oMOhVgrots/CrX3iCCMRLr3/73UWSYF7xmb3qq+YBYhqbx9+K
oRdmlq6dzBauKemoDdVlh64C2jIw9kueva4gGuJvnqf41wTZENsMoremu4Z+eA2ZOos1JIMK4bfH
CXiZ7tlSS7fOxXSH+vMWJe5Qia5yojEQrnN3kTY11H3ZQ0vzw5F9OdppRLXfDfCj0ut1ilU0IJZK
5jOE5k0bXUw/y2WRcMB7ptZSECBCbFaGUfMO9v8/8s48UH76AK/TjxnC41GqSkYrbobM232QIhxk
+fH50NHuxCyBx56quD/iJoLXDcM9Bv/4ldDpEDNEvN/RUAFqExfCZgsA21tUkvyPaPx/o20zyw1M
MFGlX+zdKVzRKe7Ur0vX/0JEIjLH08jv1KlpHTPEFV9klbg21Obgdpgdsg6OHekT4ZPAqJL8YZXV
F2v2jkiTaXU05rxI/d8jjX6HLEnWvv1EruBNdK974tZIwb3Ex6iwbbwu7ezjO/o2aeXhq3iCQOJL
ByVOTh6Agpv4Xjqh20Rv9Wr+Bn/Uzxvqf83y5UDNef8PZuvigQYmaSZ51kmO1EWVyo0ktMAcFBWt
BtQjNaunQkHOl5rzFu/O0l4ez66jbGqVt5OJY30mQK4i/+K0q5l+LT64Dh35RvIn188erSYbsNuf
o5XZBI7Z8HlmrR1fC8HxYqEiCD/pOlkfYCsxUzFvp88V35jEntmwGi3lz4oojzC6UX2pPRlM/Rwy
QlCKbSfpwpS5JPy0OChek7FVzVew3Mj8+0Y1KXeabb15STqcsozPGNXDHYfsnkEET4tZZrzpYHzF
noYjxoLfvK+QIoT3bzZJJHrtiGa7oDFSz+HgWiLW7xgVbbkjeg8fHWu8vo19IHyiqfMP+yYj76I0
mQz0MoYcH4zuYxzTL6jX/qUTcQ7sqf4W1sWFgf07+SMNOIWU0mXG5RBFPAh92ydkJLdSMdfUC5+P
FXZVJIRQBO6b8j9sPVnfBZ1+taCKtanX4+gjhnimMxPoh5KDG9apRJzFpx4Oz7yURE2N7DxP8VIR
cvvJ9DQARJXKBwqUnETJmRnS+xggGY9NIFbDvNYu11kxD7g9K9sQL5kR5545ATPocYJGUrRVOSoi
bnkWAD7V+25BtoY50E+DtkVhnwnpL2EKLweYX4OUUYVD2tNYJJoQFoBnnZAZveenUwtUzO3cIRH4
ben9GOjKuaZ/SB1OQVyH1rG4+qW8tctWa565Z9DQMCnmzR5TJ7hj0H67hziTTL/3gdRjgmLp3Ph2
h9NIflENOTpps5+6cnRNz0ibEkN6OxwAs+GFIlrq1K0ZFbBF2Ga9QGd9e96R1h0L3x4wXzf/1Hyc
/tJB9uQQTajk2yiSey7Uoqp25N27Ex+JVKANTMj48tvdh9jXrmjAgr2OCJzB0ApTTj0cgxl31RVV
++1j+1ONaL6FUe9/TxTtuH22PMWBL5FKe65P/bgfySm26J4fM4Yy6ypyydJeoStqs+mneKAiH6o+
QZUFd1rVXgsTlqkWDjcyEyREt5cM1TDkuR9aTXtrWY42aG93t3tUeDqJ4Se+3BpKcZ0FXr1KpdXa
unhggGumQ9BEFoKNs8YlofYsSXMdaK8r2LmbRfphNCy4hrJyPTnMXyOGnY9/KGgUk3pRQ5SQi00O
DQgINNZATdUjjso4fXOxC5nu0yjS/BZuKl4ZerV8re3lsfQxpdbTMiJ0S/gt5/H34TBIMwOph2CN
PE3R3RUypDn2AjpcmG/vn+034ZkOLHHICbeZ8XrjZbA26h6t475uue+Lllzx0YrwLdBT/FpKVEDm
0dwP25Xx2Pkm4qlv+VXOnDfSKOKT3LtFOHplvLv3LETVCzzj2D0TMCKNF8HHrGBTsvK8xGy5L1f2
bRK10QzmFw4M4nWBtmtO/wYNUXQGKEHgWa/G2n0xnF0CXLvUcU0Si69YS3xYmnkkVc+bz4/lejgP
FYRS4MorNbYOYWYsVoZkVMyImkKFtDU892bxlizL72IM6gPk+lMM8LkNBYLT7hxRAhzepmkW/bG1
9tfVQbrAHMGDmD0zQ5XU5kmE79yLZper/8F+l4yHHQbQt41TJK99BzSPQrNQtAJTzKsyNoeg9dSy
WeGZdNSLXYFBl8njl0Qi2UeveXrT6/MdDFS+VZ1BUR/Z5/69EZVGzVB8Gyuf57qjgnMf9bi6kUQW
65/6C71OPnWYOm6tYksKdNxgWAXFq6X09E61M2g2W8+0NXSXlNRmVvmj0GHV2YXg2Z3RLNs3Ybys
zUZAKel1WfOs6zqAksxX6YYBst9nJYE5XjazVbnBQ9UvqBhqSZu7WFLER31nuZlQSomuuJCvxxq+
+q8pLTILKPQKol8esWs5393wYdflJ60XqenHyP9UHynaCQz3KSNPZVRIVVybM7up/FoMTYNpxTOD
kaz1d/HRWrhUBca5P0zgSo7zjmODLH/6VF/v5bsQIhWJndL/WBsKwwvcu088YAmch5QQ5OVEea94
Zpz4lNdhyNPAgURefbWGvX6rCVCp1XOvT2vCoW2k+PAcyOnivPbqwRo4/8z1lhHknp8Xacqi0G9k
6frIR0yElV5DG8D9e1mJkKMQUN2MQufSjekj2KSLaULUEfsIWrq93tLs1Vm7oih7cHrFeWTrg0Lh
Ams4VF0eaJW7ACLAmr4i0bv5OP7Li1VgH0JXqCbfGbZ6kSneRbzkBcjYnuHuthi+gZAL8rCMdv91
1TMh5rENH9i2EGPpFci3qr4B+6HWf7YPTWNKJd1Fhpl5a+hKZoPBtu5AAn5pOr45lwBcynlrQsJH
h/yasO8H2cT9P1t/x7CGSjfdm+m2nchlRAe0KiB9BfeZVrzs4IGJMe39KxZfjps9Jx2YL0WrptNI
pm/TiHavdjXTjEOP8Msnf0QqWivZAT77hNFtHVjHyG2AP/S4f+P0Ju+1li5ndKApyej3iR67QwOR
NOq8acanNC62NqpvswBTHj+Arp2+ZooLB2nUH518up+DCJrLlf8M0apF0mXmI6YFDuvU7k6N3exr
9twPtZUVyQJPNFIHuiWrgqLR24T9XNTCkfj2AWKydQOmd28N5wUuF/iSUFc3ODWO/mFI/6hO6nzQ
kQ5K1tZ2Pi1rnhGFUHr+VAmOo5tA8kAyxBNWhxywJQj4MOtyKE8R95HrIWX3OQuZriHbHB2gNVMJ
zSW5UKF6csyQZgjZOfiM1i5UvS7VKtXjSZJKzpbrX4d7YjoxwEq/SkUBH+Gh2BzNRdQXsc841Txv
c4ldSvoJNHGmY++allZFDOb1JQM60d3mU5+6TLGENn3iIlDKX+86RKCdNds63adcUhZWBn9SONSM
r7tR8tUR4BTow3eU7RlicX6Q4LQjO1iJfF9riOPNc5jWMq9ZYvHU6+0BkxwhGFySMQhw+z7UBbpK
QOEh/1nisJ/7Jzrsfc2KmrkI/Mft0dKmEzaWXNIQsvnBUnrKemZKSUKGn8UeP54CUKnsFdbOth4C
VEiTrfUqaak1mJy/7GPNzKeP1KD7SxZWzN7yczqsMrCH4qlLgaBFCwK0ciRYxQsqSGmYcr4mzfcE
5lTdkTRC8IOdG+CoirllH3R12qnu9uEgYmPNe97AK2Y5q01irMJBTwBMWdQZmI4jdLE9kCFwpeSm
m1i9aieu/l8i56unPGR0CttHB7TmyqpafJDqTmUNkkEhjDSaxNsQB63r54rCN9ES0RU3H7lxfyyp
EV+zZZQhJcury/HJR6Y5ZbzUPTkvkTAsq9Mhtb4J9tFtZ/mmHQo0NZ+CE46k7aADDNmGqKOPFFia
xJ6BWz+jcI+K/xtRx5B3iCHrCmHCVcWyQP3a7UwpmrBEBImDl9k6iFwx9k+GtnCYnEDQfxPzKnSf
Aph5AzLiQQi64DGwJLFtl+1FQHQNhMVTk0d3fKXbZUZumxwoTbyJoncqvVPPpm71UzAf4GuDFhoq
AIUFyJ0dvb3LAaQmP1WlcK7CvGx55WzhAH7i3gMeGdHK6uoHxAVzaDK6GXzpyHrOwBf85j6D2uCh
OV3e7hMebG6iv8L+WT/jQxE24hTn0ChVbWJmfp/cOH3WW9G8jHZq6VWsw0o/6XlDQ6H9muJ1+7xQ
ModUHMwTvznZHox3aCvP32ZrGnDuKRV7iY/EO1W3N9arEWnJU4nLCai8TfeNbWt7gi4lyALamPjA
mtw3EOdgGE2jnVj8MHTkDKI7KxNTZVQDWpD6IS5NyPXKujnd1k1f0Uyc3yMpfZYbJ3E8Rv/1bfld
v3OVnetPJK2O56ZU8u/4fBnOI22uwy4Dozcd0OVUhwXCzEOckDJK/XS9F4i23arHkAmtsQReVtZM
6bwypFNravm/zua03qIl1ZEQ0XSsgK6VkJIR512N0RZirnKJ+iAk9MXhVk4QNSCnIklTD0Aj/E9f
l3OYNJmptP/WeI53z25R+qwVJPLBS8xfuhgpMyqTzqLwcu/ezLtDfr2QlCt4hqf+rQye1esxydxN
TglJ7y8zK1Ln3Uj5adawYbeoN/qU5YsjONrA7CgB39uyxOYLiHb1qipmyvPaM8k1rOKUyzD+xPgf
P2qgSpnOs+KM8OGD8KHHWmN4CIrLWaKTPvr8b3aPMNL1cM4VdfcJ+jgXU7SyUYTsZOifPhiadx0+
A2TC/L8BfIh8yHKw9jEl63mHSefrK8wIxiDO2s2Pe3jsUKA0cjnd4amVgIU7yxMC2KufG1ymcMUS
QcBd6NdZdmaqWg7ZsFyJCXlfuIvmeRsrruvwa+UQ1KrzE4ZH/IHIOXgHT5oZu403VPTAr/as1Wl1
wWJqWWrW94YNUs7D2sqSCq6Q+GLWzsniZq7RDNhDe6Okk8q+p6rS5iGXOq3CHMLDy2BorG/oXz62
anJMVq+GvHZPGvQr0IWpG2RQeH5MDONvwvsqX0e7Sq2WYdz9wHROx7oYvmTf5BkUlpaO0gNlPEV3
8jjs5JXas07F3g7HgfcyVXWOK9Xal9zZfsmOzejg+kw4cSA7TTBElCT2blmgVagQ6EIq/cmprKdq
81npAET3YlpiOdxaeFJTh80AWx5mu6XJr7AbjJf9jljP6PihTPxT+sws6psIaxXKK3TWyE7bpT42
AdHoeI/h4bvSt7bwIe4mLECz6Z7Skfn0c86lbe1mfqaYo9qM8WbvUXh2aVXtugvaCIo1I7A9BDHM
2u9wN8/LlQSMJXSuPPo8liPA2yyOnuziEpq+ZYXVkBIbRvAF+otu2YHAEUbMV084iAkkQ9fEpnhW
A/1FYtysQQHAPqC9wnScrDYlylC506YhuX20Gie6nvMmAX7oU7qeX3u6whN2czlMKvTyxRvwGlaL
UqwSHQ1rHQuddZmT3eHmylvYvlebdxbDeRr8G4ceP3ljMV4OqXLRG5Ht8GldGD8vQW6vNAklpVsl
DKyz7sV2SVOY4fT0h13wl+GxYbE9ADrXpJL3ercNuc/WoNjwEd5CsXLImzKbMQHNLMWgtUl0H5f/
m3K/hNLPhIvHy6+u+gE5wASMmfwtayw6xd0RLmcJagyDN4D5oTcu7lAzWJQzEcCRj2wqwmZHGd/d
SSZs8vGGu4huTow+F/80ofl02gUZFeUjscs89hWrBqRrkv9uPj0vmCppRb5i7P2hqGD74zWW9J4M
pm46Ytc1C1JGZMrSYIH6ljP21G4AwjhdbHMMaTIHfW2iLSLka9i/8Qcm+cile9YtwB0hktRJYjsM
cOWaud5i/AKWwIvzSg0XYHvsYNdI8IbW8abHcY2Avsjc1cEgRHtqxW2w3N7vOzv+3SFouPIHhAO/
WKV/H44g1AkeqTqzOEF/HHqC9Avkb7wWLBw1naSTEkqA3iOo5rBtLv7JG3+oRlWFtEuCDWzv54oB
MRSsSJwMUvb5krJJ8y50Nn5O5QmJxkbMXvYwxOHEJRHthXSzBjc6KnEny2D2k5N5IBeGMBMJx8f7
uJPcRV5AZPCesnyIjq8uFJlrt0REiaC8+XuMOWtWuVHU7U4Aml/GlphYZRV6FQEH4i4JIXf+CZym
HA8PlGcbwqZcBQjXwpoiDGEmdVhhB/GXMOjgwIVLyunkRsWFfI1nb4Gso9Ta2u9GgKVkMr5ty1VU
fgEMU2k4ex0gfT1Wlb5Ikc+sUMINZtqVsQi2o6lXcbQ+YIk5NBNb32AtZse5wFEOlZYYZWVikeUU
5E8VR0zkhi6GsC79X6CI6BCL/x6X/w4noblmFRTosdqeIh5sMJZgSjjEFsmI8K9fhcEWVMgQoAAu
s8KpWGsg9MiTzkj8THjNchERf2f3iGDdCQr5iSOocvMHYVLktxdn6uDD1/VYJDt1SKaOucK6TqJ4
3VW/KaDGBbl+zNd9nlzvdqrjySIECRm8vdvHj6TTBjSMA1dM8Nx9QRSLbwRM61n1d3JniP7dBEtI
piYbC2CknOemZrNXGNPEeNjijQjMhaOFfsNvz1MtITqLBQghEzogmBjSoyzTq9ilfCx82+wOvi+p
lvbaV5p7MLderdpnkwusDtMYFwgtFM+PvtV0TFGfiTY6T0iHA6XC5jDkH5V6fy1hNLr+nF6K6uI0
YvLnusFROKPmVWx+keFdGIVgcK9cVTpxFVRum0R6naAqVXrlJO6gqxSbAma3AP0hQBoQyRmJP9rP
q3iPRUmB4ZfRmqL+5eNBPlrrNUJcUhdmxMSPjCJ7kXpCoQVY3rQJaNXij97jkQUESTfgNd4j5dhu
mHrNp0XAHe5onn1UKhB9x704PgThfjBXbirCH6guYhCvp724Kdw9/ZkXErnOTg/L5APxrBPD5lWk
/Ry72MFknzTAuEUnG7MkCImtgNiTS6HSgoDfVt0ImzKdysPYOq/QOVa0Y2KUwGR35HFs+iGEkWWk
ADhKZdfK7apZm6lTKW0mq6DpNhdaQCeRWOBFsM2sUvTDmyGgmlHAymbKDicVWYWUYhf4uGJisbuP
GLcDj3MoTnwWShwfQ3WC4xp4RgaPWikkv/CkiSuftPLnsmI9DLAmsfzG05odImsdB+qTwu+/V6+K
3/wbEEnwGQLfaC3dvo0vod97SOvMvuNi19OzVijkC+U1BussbzMKz2m/aN32yRz5SxSgNwM5um4d
t4iAk4yWcP3dtc0HtQasVvlNY6cGssvn5vsvagBF5hSz4kjTNwSvf/vaQqPW9C5Fj7WEaVzgxbZ2
/Sk8WnMS3HW9bCJFuoFv8FD+lE11ei1GOUvWYXyT85f4VJBl8ZIjie2CtH794uiJGAbKNM1R2UL8
Gi/4qmsp/lkboDME4e5ckMDQq9YVFCn+xB9QhEpTWXnSSF51v+vMv6GuD5KzlYDO+shUczKkkBLE
OxR9TfCVtwvWN+7SSs8xkKM2lKia11UPLR+bpSRCclieXBFd2Ypy9fyc5g109e0wM6Y6RhAZucaK
CBSxg7J0inzWziPKTJtQt0DcFMWAQqrw6FPJ25elI3KSa7hITj/IWG0jU9MYt29CI98AAoAlzbxN
uNO0wUeZI3o8bsTc4Pdzdiid+0ML0E//AM6NBDQ0aAAf+atNTCRuAu5ofQ/njNm669n5kvg2mLa1
wubed3WSdSiglQsOOoIJauaAHEKC2iVNS2rrqr3BDe6EkbdvFYRb82zACdoRt0OVPqN1azVGreJb
HA8FYRIZ95W0UlhLZBYg5BYD6x6Vtmy6VA8BHClRuOt4DqxgetKsJw6q/Kuv4QfdrQyzofd86uBi
g/V1HYPuvwFDeEpzwycWozAaQqDrqtsRLK37d2pVGVldEiuX7/4JlhFa/jW4B+FERKgHC6KlXa1e
/sFCXYp2gXXbjfue+2VOT9n3F5uL5K15OTUYyZuBXsHZydp4oWWi3YF0nBt2YBuuzGXMocqZlya6
CLle76TZ9I5Q6YUNmMWSVo+/BPVGVDKLL3f/pVclgvbWjP7xCVWIQFTU7M6YTFZWHnbJE1kpfPsn
K9bb5/luxy1fDUOlmjwyDIscX4TmdzLBRWcok2ie1lv/4vmfr4nvc/Q0T6PNN/j1kW+Hfn1W2gAJ
0KQQYgYWUNIq6CDEFFu7U9r4mlSI8oRCgImvA4qnpf6ukObMe7LzSVeNUKLGEBigoEBU/jWg1b98
5JxfM83beH9KRHyA9SXFrXGbfn/JyzwASFwQgZNA572p4muycPOSyZ+9KN3Y0Uj4IPF21vQiU+lp
jJu9lsIfYGdXRDciAbetBaTjEubV8zNZP+7sTamdafX0GJj4fv1MrDZZ9Q+hsulJ2h1n7cfOJrQQ
g0zgegu9DXRjCvuNBQU6GcRf5Vqx5s2/zRfi0FRXAX+3TdNlkzq9m+EKllkeJ1jidU/QcMesNG1W
XE+vECqqKPliNQvjfvk8aNt7tlAIfx5D9aN2Wie07anuJtbaP/aNqB3Sb+0E9idT/ByUz9Frz0Ml
zdPJy0DkQ/wX7lImH9ayx1373U5dPDL/zFRplN3VAUUNEaAUxkbABqk0k306dErt5hxFX7ZALxSV
e7GYxDqIgyn5/o8uf/vPgT3Izr7a0zummRwYBEcX4QbuZi44+YlezUbk7wpqsEBw2sAqeyHXjy5V
+8B0gSyL4IOxAVp/wi1xt6qc4tHkSqJbkDv7hDGv1pRUBwDzRiocH0FyUw/vLuJk9na0flT7aTnq
IhsDRBrubAD8P+JAX9vXW7Ap8PpgohkvVUz5V+PPUtIorSEyFKld4H0g14yEY779jh5Y7/UQ5FSC
UCEAe5/yot8Cq2697qGB70ZpqcjHa2VfJwMQq7aKUnABJAPepGBALcInz17bqrgwK0uIuTYIOMge
R3fu+EvCXa1rJqc3JbkFxG10nlXcOkKvu9HiwUkZ5sTFls2SHbEvyZcGYV1Oam7uoa8AXwukRXa9
nMLIX7njdw1NzBsE3LTqZPcQuNSbgw9WRgz7MDaYA46QVDEW5Yl0nhDLkvN5+Ji5Mqpj5UhHEZ9E
g8WIev9Rq9R5qNkMMF+oPZa3y36RCYH/Ulq9eXbZCW0hUbU/mhcufLUcZJo+uljoOWmKKesvU3Vz
hdotnE25Mb0JUl7VOfpVsaE0IUW6GuLMK8ZlFnun+lOGPQtOKovMxf8FiqA+4ez1ZrFJu8lrxx52
DSFqG2Xb6ZiXBMxHrrmIMNcSPb+reLA30UUEF1zgj0H2bolvcyLDyxuFKrQinz98tB1BDUJFbZ4C
sboyKAYuu5BouvvIX78ZF0o7DlFJlz22CDWs8rDDFVdkMCZV5rSKRGg21Bcel0cOhS5UOTH5C9cF
LVKzoot6ajR9ct7mNi73oxpIpV2ZbfbsNFjtEcLMN6exzYie4d0Vghd7HqZsA2WaY4zEFXuZoBrI
qnobck/cB3dilOd3FiJ4QPJqarg4khecBibKgZrvFiIg2dTZh13qPzgTREORXxPp0trl959Dtn7O
eNt+O55+S/0n5xN4YX+Kxb2+vWNvXqxMR8uxAzxNUI2de/6ADg1k9djJlP1JYzFNjrUE45f1EWtV
wQ2FtpdWQtkcas4fZYzJ3ppaSW2fJWMDeV6HbCTOzOP0SDYHejG/i/nZH7xyztGPLlegZaSSglVP
KkP55L36inBnCyPIyx43LAVi7OIaKPrxlTBqrHIzVN/IEG+eQ4EQ+qNKAZbFayXVfTINY63G0y89
QPHVfEpMs6Ogll63oo97Z13Nq1hFlDpbAq9vEyW3SNz74QiDZl22iWO6MUF9j/ipPu2+buCcPVmX
bLCZGKSA3FLTyqRjZis3THwEg2ni0FSAAPIB11rCY0B8FDAL+LTmEdzfYC2Wnx0uzHdPAsXM3+sY
NMFr0MEXdP8nJ9qaxDHw++PNVzgI/3TWJjK4WeFozENHwep7UqX1Lg98Q2bLEh1t+ohTsmcCRm8t
M5jyjkmY+xuc9bQfZMROD0uCgYxrH1YHZEGwP93TOBa03Q3v+Xz1abq5vJVN5FvPq6iIOaCcto1K
0Xs5pC/oqgTvW0ux/W/iZNKW9OdnhLwYWe14keqFLAdy7OFTcMtnEmtbDr5gd8LabXPK9HpBnNkr
SSF7xU2VdQuWVhzP2uLYy3OkeWYjYJ3q69CiraVqTgDJfIvRvbb9OQaojW5K2q+qZdo4bgcNs8F/
CmJtaDFlUXqNX4/7Im082pdwJERi6Ol/YirTB7FOm2yCW+cxRMtAzynLeX8lvu0tjuxD4lPymu/V
wkkgKG0X1vJ5QDr8ev1BO3RdNjmQeeCDgJWsHG02a5MtLPln+kX+EPTWVfPFzx96rel0v9/+Bae0
4+gTdR7PY0sWrZQZFPDR8pt4sGfyhefNps1h3WMpBu4eGPuroxeNnsea+3ArguccCGUwUaaDNRDQ
CLFrKdSl9w2JFtOOe82+Y1ZDZTXn20TrUZcnqi3+BY3vP33ePO2GHrHpLTwHUbf4PNpz3bc+CqgB
ABiNd/BZajPwj6h8lUUZ1sMr3npkbBqV0Ez2Z6RNjIBbslKLSu3GGi+8/MtT6PkMx5aMxMq6j3Zp
H07pxrbfmEwk5ThBWbuLtd0OW2p7X9mG6fRk2FRAwZ4+8+8oJjtX4s7QVkln9SAcQI3RSmV5wNLw
37b1b9G2hgI8r/qQ7y5llPKuL9DsgFX8zmFJ9QAxT7TnT5BGVS+i+5Gq1ioZvC6onK5QqqWjVSY8
qd6aFhID4D6LF7moiWtZffdUXWp1Hqe66B3Y44WD3RAWMetMgayAZOueDOD5ONyCOr+QX8f5d53u
SZLsEscstKS7LjnidnRgozimtSGrHQq9Dztr63QDGksSdj8L96emEiWd9zrRMrTnY8mlY/dOPkg8
OmGQZ6vh4s5S8AXpOMhDNXolMJGlhxzlwFeCQAI6/Zju6uHwbcZuLRTLd5FtNgnsFzehZHnlunt2
xTTqLJ2DgFnsQ1+qyes29r3J019ohq9yHIKM2cjGa5h/sBkppPnqRl/WgdIADQm39f6UnkYhG+HY
GWZ3PGC6vFdgBTdaAGP+afG5WgkJrGCGXTu9KR3axMNz4ddClQ4IHkh5wJu1sD9J5UEcS7NZ7r6D
1PVmInNsradYgDP7754DvNUeVOedI0dTVR4FvjMbm6Dldi3wO8FaxbcHBtZgzpitOBhvwxMI+OVy
+2sGz2v9h0q/ERT3vXw38304It3nAhv/OkrRwgnbSv08dQazJVGzE4lXHhiRaVhXzSGvgvVBV4jQ
vG6g5uaWfXo9A+8MpsOkDG19jmxMDpUEOhp0gg9Z9TsrwmmcmsD8Fe5cZhWm0GzmaimpPVB7PfZs
nCQDzHJKkTMdIWFBIqQVn5fGTjqXgT3b88pBa4A3AFBnP6fHaMGGlGl71rht/Fm+tp/zSXkG4sV9
TVvW2SA4N65cN999Fb+eIpOmE/LnOTMcfA5WV/QyGzoBBL76DzpDfG4RJsLXNjfSpyFttLo+LGZf
5sbXaSbb/VNC8U+bQZtRFk+72UEh0+3lBajnJKDYT7+J+NZ5YQ/rCRNAkxkytoF+CxtWpl7Z+Z7B
q2dWG0a2e/Opv9Mpz4MLE0fdi9zTJ7dQxjIFVquSkHVxHMWStd2LpFWb1NhmzxpWT3YbCFFBvQdF
yXml1Kvf7/Kx/vnwLpIqyoCjuYBd2Xeu31yyk8AyOnszTz8aLG97BFHdUS8X+Dv0B9HlHHkGpf/l
bgQ+SLCUKcIZfLQp0TFy2xJ57no9tUyC8Fovo5YOnnCnNaQ35+0Q/tfRjp2eN7FpwTQUBjihVmVQ
QDiMmTpojCIoEmGDoIfgQmAcC6zxTbSeERlintJQsRvQWqMmdl48lWkn2cM45h2FpE0+zeGDL7xc
ZZO8UigbPO9AUI13p7suek8ScteP9ixMpmajnw/duaYnyLxLRhYslqZNrli9aL1WymnqIYjtnxNe
1BjRZdhDTiiPemCvD5+klIPudLhy7wNLEhDWsUlouTLar3/NxeXxfLoXlg0Mhq+OC3BkOEdy8BD6
HlXZrQtKLkarOpDUC5Z1rMM5Km5Psz3mtil/72mGDaxw+FliaVoNvVb0HRSGgKO+aNb9jRLfUhVH
s2cpeANilhy+oqB+qfVhP++ozY5hlEzAbGSYj/dRuDjqWduhv3AcMqAI+RquOWQrwf8Tw66PuIPa
atpjup+Q7AqrMwfsQr2VJB6SCW5KjUWXmOWqygT7OhpA+GpYK1KspN79vUL3Kxy6V/BnhsJ12kty
9ostO0xF64q3izKEdq8tC5EUzX6RFuairNBZKuvz8Qr2knVjdTLrnSK/znqgoqKGo8PSVeVR3j2x
j/AIdFdSdcx4WGEBs4IW94eXj2MEK+8GOsMCu4dtGeopT9osdV6pXhK5K33kYVmIJqElqBghebNI
sXq77eWehv6BnDCU+gJY0Tnn1BQYza8YBUh18z5lRxw4We8jNh9FmVV5C9OzI6PfgSYjBP61N1Ok
Y0r3TKnDIsxmfzZCdyQufXAU8UEYSaniI9BbpW3nUkNN088gXT5rGkvWuQ6C+hEtCje/u5qJIxM+
8rexrfvbbaFbQiUUtZzvEmrriXtnfyyjuhAXVZoxoO2Mlpbd5wH2MC8N7l10lYC8kP2myQvs2Bi4
OjyEDYoHaHu6aMBpdtwzIcG3s3m/qJSVVd/HFEgCy1aUY2fjkUqRFSxxBqrTHalT+cnRrpYjsJEs
rH59moE4uAagCMXafMVYISCiTQO5CvYnk9AEfXFfFw0605b8Rjv/smEyCGSO2b4ktEjopJ7vZFfR
RrpvHxRiawAjETYts2RCuGecilCNsxT7stMLx2nCgYOSbmwcq/ShLw9jbq0mX90wSWxYq5WkmUO6
Pro2iMmT2gW1nH+rFrdVXT83toSs8gy+3Vzt1H1tbNFutOZhEtkoNniAWr3ihKB7H8lQ76Ywievv
ZVnirTI/ytOvs1etnrroxiDIVzaTR+iFxZo7GhYQW8Yz10WtG4fbE0FIREB3mglihMA6tHUtmsZa
nxvnzzuLMYHc4svXtSnEmNzxKv83cGZYrm3WVzo7RRas5/ML3DqIvy8HwlKDZl+FqBRkAhvVf9uo
kbP8xKVnR7ZUYQqk6XGxUY5q0rr/Ue89G1Mc+21SY5UNq4PDwjSa4CtYndBMP1hbrJ7p4GDAI2pE
Frmrzk1TEPp3g8MpxPz8luXpUwbhxfXN5vBbK3ZHjcGdXc8zb9N8SO8cl2L/q6L9dE/kTx1Bm+ZY
mH+SdLf0or7wM2Eyd/I7VAIgpyQ9FTH+suG0W9C9BrMeCqhDOeTFKxkBm6Giwy/YMqx0ut0ceHKH
kJO8O6umcSF/EFB0KlXq27DCz+hWm+Fuld0tQWxbbfSZrC8y6BS/m4fAFUuYg8wLve+WKzzZ4Ub5
y9tGjcXN7B1Pf3FEo/90wxV6MuG7KtxCLV/KjxHddQJa+fsqWx945j5vPxdskCah4gS+xeyZ+Rsf
uW0Vi45gsoJabhBrvWsD6GISb4BfkZaBRI1WVU0wL1bRDLUIOFwi1M6A4sfdjCpStS8Z4jUBnBW/
/c7cwJu69UzD4uSUyXWPTL8C0lep7BFieJTSc+p3mm6yymB9VdJIcRaLdw0gNI3EeqeBW3W+eIYN
ujQ1A4AtYAtQVP7Ui8XmhKXvZ5dqcOG/UPpZ0jQ199Pnh0rl0sttVpZ8aid/Fst8gF3/8IEATd9X
TdQjKx+L4mJt9ir7vMG9piIGv74l4GmW4lauA31YrIuybvIaJgb+bvTDYHfNaqAmT2Esn/jmMziG
Rv4hrUTk0mRHcVSCeRk7qusAy+paY7eUwojouFCt77znGrGktRXYquH7Mel+/3vWULg8PlCEgrvG
WhOlv2aqfCvbZsGRS8MTnDJkLaLkECe65aB9ooCgGVufFU/oJT9sVzDfLLN1xTc2NZVbTK9vXq6G
Krmc3KNGl3h1jCDUAGTCW5KAQzdmYs+Ya/lZPia0UtCQ9uIHSUh8s58CLM+x7NXlFLTL21SmZdTH
LKM5WBL9Yt0Qyw9at1PdgB9pclnID2H9FpVtiDr9iUza+EUAJC+vd+knQrmLWeCLmwKYa9zOdEqK
SCX3flj7U3ZQwJuKK6FWsUUf2BfAkhEK2J4L1QqD9Np82+PAApOyV1lgsRKF4wmItbUM82ILKBKO
1Vn7aplXdwFy6DjizR0l0xg4iGjpMC/yRoE5SfWeNDCTvehoun6umKhdjfujb++cXSPXi67GyTzF
VBNpoKS+oJ0UmKKJCn9xwhpJ99VztAS/W2M+60xMc9o+IMItgB3REYx8hq6DOQrEhGvatYmza2yI
r8Bz3tb1qjczg8usg1Q2bhiripudsomhMKMXX8E8iCdXsaZczlJS1pSxSjAovHVWM+PqiLRSR/FV
bWBJlcO7gFZLFFF/MgrFxYe9l386gAxgoHCUQz3z76xUpoerjhLT/v2TwDNfs6G1vzC2gUUoanEo
ehXfhygaZ1rrUURCtCDkW+Av3euDfWblnUDHPhMRY9UXFtYEQf++t2HnIoA6CmkFrswsqy1XWghB
mbo+OLdNP8IY/qTG/tj4LS1ttXTJ9DNe3OFYWBiFQkKQWxoPfXv5d8D4xktanyg6zvjx0D4oQwKP
od5x84xHVCjVW4E92q1ThLtvVUUZ8ilbKl4Cw4M1DxU3wV3GqrcfLwjQnEjgGTtRstMZ4NPxSf1Z
1VKzQ0wYzBOGWXxVC5P2oEQDz2Xk/uGM3h+KdhRYIURrmyCbwjNbG+MATO9fUjrFbOA1TcesJRV8
Oyu9IkHGH5L//glyOWnzbYdli4GOmZMc4nADcj/tvKoIR6xvsRJH/wk4sBhw2q43Xaf2g3SE0e0e
vV+ing1CdcJuiukHOR8Ifc7BgB5Eogg+dOuKnmTXUwuShG0ABuprMBJS37HLiUda6xvmw983QUo0
RBLjCq3hOyf/S0H0sZwlZEmgfsL8YaYqV0WTPZSdqvX7yA4lkaNOQJViY0BPsA/4lbVg5Ua0+E60
bxG95ZZl8OZfdssAV44tqyzKhekFZUg7iGzhHV9PFKuQagaMh9F7uWIOMJzawSEVQOZs4L6fLyRz
ki9x/itus3V119VDN+lfj7iGVyYIU2nac1kJ9zFRd+LG4OAtiZymllD2B/a+ESNBi57zhIMmpwq/
Ga81qqijapY+X7mlpyFkD5hmdAiI3teJvbQEqodYqYtRvFIoynBMH7QJ8eHytcXhqYWOvIQ9PhEc
C42zSGaqCHqW0p7ogVC4j8SYFdMbgEzHcUpkRJtAjGOC/1123xDh1ijX4Ay/lnDa4ePUxyCV+e97
6OaIZy00D41wGrdy2TFsSflGkI83ta6qjTNwvsHU6MKhNAjlmS53Hob1N/OopPyZUpa4DUElf7DN
0if7PnPmeAgI+49YCVfWIpQ/1pPDcLbDHIj33NZKNcO/xhGGmuOEbK4jklP6HXf8JwrJ96a82//3
EZhrZMe3ZDHHIwZXreaED5Pl/csnZC/6z2ePrU4k5M7tmRP9f1bXGSOv6Kzgy8I+xX/HWPB+H/Lu
lNJ5HwLfE0jfmTf4kppjMOSAYk91F3bK4WMJZcQn2XfCwdBlyYK9xc6NgpGnzlhRk1iN0am9pSDz
ZRrlv34hJYObAObQjUElxHvFyRFHhKxVHcXohgBlRbA00kOSkAYqgy3GK0+R07l9FXTP5fpgE/fN
UZHnFvIAuDoVf471dyFynWsFLjXFZUkvmIio/p6J1DKdufRbEWr4U/8zteeWXLkcc/n1J6491tvj
EgC5Yf95PPd9PN/O7E4sfMFmiMleWWye60qBS3Z8UKv8rcOlCBCpbDeg1Cr+gX3ebGeyTjNBHmYU
jSOWQGML9QOlQjIKKSYnzune6BRwmkiHHXcLDM1J4Uk14uOO9dje+AIvAHV/Y3SzA8GjpD6gInt0
ek/46tnWqzPNiJ/Iinb4gX3BUxr8w3RkI2F12k87F1WC5aWpc7JVNgiF4R6m547VAaFgDpNvK2tN
ViDExOsEyu/Kz4qUNyTLL0/p4RDa6q3xhqrR0gDZNSQ5R5Vz+WlPD/6sBKswzHuI519znHOID9vB
Qrw8mTYuysm/yxQExaLQmurYNuKMaEoRVepcr1g7uuSJuzoKEfo9sAkTpji+mA6bG8kZ9Ko2pkC7
31hjs3YxVv73N8BMqrQB5W61LXI07e2ZaQxq+8fMc5FWteMMvArzHI894vxTKsGQa0KgDjTHbYmx
p7CBCjHMsiiwkgOKteJBEAOVfX8BXiTbIcXcE7d4wGeG6PhlM5PKv1Se8WuWE79/BrA7FiJUkOUl
ldQXbHIWdx9YwA1YCLUXC3HvKlE4O/OomN7TYzsf8TyQnk78FTqdAWWr2vHgwDTHeRsKK7FAaYGB
bcJ3SoyXrooLp8gCCRzIglMBgF/XM9YLtFabA+TE7EtR0R3eaYEjfQVdo6Cddy+uNICyl2VxGE+C
VQ7Ls5Mi4h9HobAoYoxME7l1U6aSpgZXaNOo/64niieDz7DYq0Yl60Qew5FE6ysWRIdcTkK+nIO9
yujKqdGT1eeQ+HVxM4EnhaGKzczh5K9L/z+7LkYUqtft/mhMl6Ut0S95l9mMA4glGUxtdbtUGQ3N
9wuSlqS2VKmaHSw4JNzAIp9e086SQGnl57a+DkgK+iMuMQDnnR/zfwl6PjIgUX+Nu/R3zIEfzDYh
WaEz6R0nII+mUDiIsLy8uMYc8ciRajm4CjufRb6iQXoRSgGRN70ZRThK1pCfIsYCmzHrxcvUuYy9
sge4rXsNMrHZ1UqE5+bh+P66FRqNUIQvoztl1z41DrV5Ef+hxpxgh8stnrZYpjRmObI2Oaagcrtd
DUyhKrDur6C3zAbrKVST4851JzS3NTPC0qk7f9y2L19ITlcpu8qM6IfD/90T8BoOQ8BRek25J2pn
TxRqIPQ/QN9q89Jcxg0LLK86ZT04mulfRCa8xXnVhj/ZS/BGpn9x5LuzquGcJCxmukizumJ3zGp1
a+fZMHIPT7kmnvHohQaaoNSvv4T10klZoWrQec2zuWThGygcqCTqrXRIWRq4ZCWgBbbzOQVjmy+/
nxdKGoCSs9+jqilmmOjddIZZrJBuJu8/ouDT58xwjnT/Tx6N1Tx6+E15zRoZ5roG7VoLMnl0g1wF
ZtLvGEW9aWcryjSkPalzKlm14Ggz801R/hxHIXSGKLCISO88BZArstBTD0KUQoBqCckQfSMVo92Q
gJd3eRw4VtHlYEGgc5056L/0Eo426Yozxaih7veJ1n4emtElC35BZSOm9oSgH/YJZIqmEK9SauxX
qGVnD8RPKFME1H2crR5IfwDof/WiBHfZX3kqcyuPmYjPgmCL00ZuQVeVUIxw9dndsG5qO30DQVxE
OjDhDU9y+xBD7VloKwA72H7uqeSZHRCmTcjP/VMssdk8gn0IVb0SzafsA/K3K8Ki+yUFs0u9cJnr
w/gbFG95g22kkHJiRHsg5T3J0R488dlSJfDfXEFnhMOhPxpzdNMbzawhHR/N5biIMj3mKvOa/U+V
ekfkXALZeO2W/DFn0+JEgN2LYYofmKZ62GMWdiZk8Gxt8F35qUt6Jxl8LMC1p9SKln5GRfVsY6mL
fJwMQB9UhVVaPmz3SXns6Hsam88kKGp1r687ZnWhe8+xZ08s2zx6xKEiVzp8aYVvez6wySr56qEr
waxrymGIEh6eUE7EwIR1A2ONEEVRJ/fCA/RVZ0H+7Kle3YaaIFmUudeZ4pSShWUfaHdakenA5Itj
wFFpjd9I1OJXlUpu+pxslSoGbfDjkZq9ebC16ri19XJtcI5rQCbIQf6xx4qv0X10pDFECyfcot4x
UEkEsb4g4BEAxlrz9oRr2fB40q+WbVu4Z5aavM4CsdyhWkMyZn4OHLtzsBO3utZ+t+12kXxa5scR
pnF2BMXCuOxXW6WKRYcLQk9SU7I5YyspgiNWFv9LoJZJ9sydhUAov/dQAtva0VwfIZ9dAw86KlVv
wpbxvfYsVGJEVqBCw2B/KQOIn/iu5rZarPC4xqCdPYsE5Kb1vl7l4aImGrmMnq501NCSwCUPoxIn
puibJIPEH91tElU/Vkma6aH7UduPHppKatdebTnKaCzZ3Ge0sbKGL5DBFc+Q3mcdSCddO7DBsXtw
8xs2v7Lei9CGegaIcmgQHuAIl9n/1ltHNcbW3nQ3jPBmiocTCWmGdzT0Kfd/48s0qhMbU8tlvie4
m8uWedCkpsyTxf1fDJfDDr5D2TI6bI8PD13rm1Hbxo9I2JTVycM+eGVLsbgN3efQYPaQzUudQ2n9
j56GfgwPtr43kca90PRXuHX98vOMS4zLqVezcPelunj7DlPwsQ6RLgvRRw4ZV2MAfFbXNAfibxKX
RUst4ZeFTkPVNb+U0UilpqK97MVd5pIiRpHiLLkW+rmRzTYwbul+xvOq+dcyzK+f9lCQFA+gaORw
hMsw+xR6nlfalMKhzBOCL+ZBpCjY8951tH0dJbXf0XvTjo0xrEXtyWgumpXegCWkltzvb6LCUHrr
q82eSsLWP2dPzkQw2OKb7evQagDQ4DbALkJqz67ZeeOBaWIKzrrU/46AOnnf0t+mM+arzjgXeHCH
Od0V01k6uDWax+dE9ep0xMfoya07fL+RGW1WYw0Mg+25Z44u2xazDeCD/pXdpaqNzV/JELggvZit
J3Dn5i1ztWRnjqOOyn8WKnbUVGKPdJggsJ3reh9ukosSPgKhZmIpelJSXCLDmdOGACcCfbB/Awtj
nSTbEQMdClHJdT4ptMPdNd23eObgeDAcZO4puQTrvFe7kOGwK0813E/G8idtGVhXXO4RGQSAfvhP
YoBMqNG0h2usg+1qZI51nYmhqtiGhxz09PtKaEtRVMZTsgOW+QyDUXQXG8q/DTmGd8N+BbYXTCa2
BWERoPAxcAghVFDMLBwH/dzCR+BffvVSCQAymfSPyRs5+YQnNVRG+Ps+coSSPRUC8lqcL3gfxU/7
40weCBf8vluX1Mlpjmv8x/ceDIX8zGeS6hCwEz6NOjGm1xHm57pp+yxYwZWAhz6EG//PzvPmWsQ9
lL17kQSWvFFtafmyziv2gKlSFcuAS4Ga0DgDmjR6ipz4I8WacDGL5TAGEMRoXicQUcO5BDyvesBR
XFStsGxlbQdyg0C5aCJSAgunzAzOeAheE3RKYmXfhMK+RVTIFx5J/aPbjscgKwZMHU9+RhM9f1Bo
8pELH9s/VSgI64ODqcKZaRC7nolBkDSRmOv4lohha+vMYKPxjT6Bfn5bMIdWrr98qk/m5kC5Wzro
bLeZHEcUq6+fMjxIGqEKpyiNaXWI36eE/dXbnPyOj9jkBiFsrToG+ytiD9u3AhoC3pmMIBb8vTrN
GqP2aQDf3sReTNwbjFAM/PVOrUsqvlxSNeK7TmMsuHYI7G9kAotW3b90q5jl832THHMnQZhjSLYw
L2UzCKPwn+B4MZNbZNicISVthq0WqDjfxyyckl5r5QQxe/WzVOZfZxsaDVBAAiubG/axmpp7cwYq
P4JJEbfvOtlBgkELDW7aOAuJjSl5SaK8DIFqanVFIjGIBNDCR7id76q+wX3L40nqGvYrZhg8Yed+
4h99rNkhg81rQTC1Ku5egNbLHZTFHyRvHGTvZgbc6k9nwPUfT1OzVHVdSC/Nc7VdTacLzMBNbGdf
aIrutyDksq2FMDuy911LPXwOAhx4jyzXfLLPFcdB2fIfYeCQYaXqgTO9WbNRlua3rNmzRfbVk2/K
stWnOWNfB0pT69CPmG97hkjadSnBXT7h0+L7hGUumcvj23WGy5wi0DZTXvXKl4bqR9AuyF7RcYB6
HCWIAapmscp+JEVy+IispbpPkSA2CYrGBYJIJUFht+rZtgZGM5GXAL0HVgvg0MtYjzOPeHkRN4/0
hp5LWe9SmzgHvzVYZvRzPwz6w4aHDGFIwB0Q5kYz6pT9yTYNPZflrN/om6hDhhr+VQXBoTdQB3nx
YLBQ4xkpd+z/03C457kUceNrl7KiHugrkBFxrWio/esHqmQ7DVYFznfirm92UTLG50e0R//JwDiG
7q9zCeTtjjyxkOiwA3QOWMdfSxn9sMubxjRRXjcx7l49BuZSTeG/D40ijaJwGtxQjff7TdVGei14
GyTPXkr0PiBrS5KtV7AbCat5R2GXxnayYFB5vW0l3BW0LvYJlZEK5z3wvYXoTQxy/QmUs5O+u1/+
w4La3gZyKb2No+3VLoMgpFVAceBnjxHsC16K8GlHg/g0KsrYt3YfuaHsfDETufd/dmaopLUwpUNb
p+OG9jOYgkzbrLc7jo1QOX6SlEKqEa+iuiQ+QXcbFnieioRspUJwJA2DzAcB+aOzxzq73Q+KOMg8
5A0bzS3DFOUr2uyT6P/8wsHeUspMI5uSbGIrP/UV19fijX+tRA/RGykNacZL2lm551/du1BDmuhF
4+X0ujVTpPeU2pAkM9Yo1Dcm+SnSiafqo1AZIBZdRbXizojC7WMdUR05xx/K+mizCd4KqWKHDy4/
bsCrNA23tPtzTcZxAuW0ACBsOBv5zZ/qefvVI8CW7v00ffOa3cYvuMBvXG7ye7XCW8lFFYl2yQ72
nB8VKi3/lxMxIdsNHI0WFj6o0O+Kbq9wVL+9AXa/+szG8d1LHcEerfRJOWSO6Ky5v+I5lHVtYH8+
t2m3KK5zvg0nfqvr048fKKIZXmaVk5Xa6BSqRlOIJR6DKP27L3oSly4f5iFKYoa9v4boLVRze3tt
Y/obPx/tFIBElcfER7O+yQh6WQB1d9ZxC3nQj23xZSskEYDasv7LJBTBJ7YSiRUWFi0OvVZWH5gN
FvxSi4X8mTXIzLNGoH+W0cM845K2LU4kqTButMrbqwAoF01afd4HPyoaWP+3SgEgOosMBJFJNIZS
Yqq3VLgsanLX1zQD5oQN831OkD5X4U92ulWGsSKFnf2MDKi1CZ39qqUq40byQK9GSH/LnpsotsvU
Sx71t8wmVUhv+rBtyMBrsuwt2oUZ48Oam5PsjVsDShucO7mig7CREDEZgqre/t2Dd7chaHT+HH/s
JUu25RpqpSFXu69QEfsymul3wopmzJy9MdbLIA0ZmQFPGOsX99g5br1uA9qWKSKZbHXLOFdW+mT1
NzdP69QPpbnwpirA75eLj1xi2ImFoRWCjrTAHbOXoQEX5o0b66aRn+6P51GxUyQIVy0jPI4YyHkN
DMG8QjgyR7p6aubtkV3cLTyI+tyuif8BvCHi+sjoIB3Yw0T8LccIqXmlvV4115uyaFT31Vy3wuQ1
0VJQ7UgnueWPgApLL4yPmXJqrMSquSdVcZLJb5hfCu3twy7IEfndwbLVCprCzd1SP1lopRpI+LT6
WxBoNKD7Jcsjc8gjvzyrP0nFsOq+DGDfVKFYKWNh9hfYmhPNz4jLYlD6gpK39kFcbVf/8quxTz1l
HcS443AG9zLZosDQtWVd6Vj9J9JXVi+MSoFEniP5Vf8ZR1wTUxwXn30cz6Ig/NtFwBTWdX3crhLD
LIAvI6vMBa83fq5gQzSJCGNWJTBHuaTr1iZVw4i1aPnxvbL6QhNJA6j8wP3uNuc7exo01cVIr8P+
MEYF7lIHVKhZJOeSTx2Xi1bx9GsoOUmCmanDEKJMakghwy3b40tyC95UExRylORWIvgTNDxHXQ2D
R7FrUqzgjzC3tgRKwy27xJkcaZ/ZOfSicarOywFoET90SajPZYLYk00YIHPBVOK5SdBFgzdlm5X7
DG9X05aoUmuiJqEfcvNxncbjO/+lIY6AO1tR/1oMBNExVJFWCJ8Cqp6ov1oZeT4jpy2whcmB7uKH
zL3HLOp1CsBIzDvSeuppVPbqd9SMkwo7K6y4UCwmLrPUUqFVMfuaZVYK8qvR9tBPzoJE+eID+9c9
prlDhI+c4qC3xTsifSsqKCL4WyOIrzXk8Wsbelh9uZb2GoD+PWQwK871ImKkIV+SkrlFO9m32o+y
XbFLEhyljEKIH9PJrm1/kU7F9u0ijMaLjLTz9J3p+Gq5KptnWjz7omHGVmByZ270e5SLci1zzyxy
GeyjLZeQ+P58hK6XdbK5+ZiKXqRyi3AafiATSVk3qZr/2+q/XIX8ACK6P/Xdffpr/f4sFr8pJmyb
KVwcl4WPvelScPTf30HmdNk8top1V7CoArb3TcjnA8F5u99XeVgvkz7X9Dc5VBnjNP2BPcdeZiT+
6hDdoZ2A8BYAulcd+/efFcrjCGcpunm6Z0WLlvZE70ulhMq1MpPGDqGdK1xZP4fsLFNdHoLOqGa+
XneliZfkd4jeqB9yH3Lnsq7I3JCxOkmd3c6poOpAECXS/BA=
%%% protect end_protected
