%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
EB2ZJJEBsjWE50HKoU29ak7C95cPcYfnAFAsu2vJElUtcQM24Dyz2YgoTFQ7IFrO3DYWnJm8Guz9
O0a3yLagNxcEZLah50+TEUfw2Awd9oup4pDXDnLbp4RMTHsuMm9eltDX4prjnF+bs5N6G1w18Dwu
xQTgNXZUkZBI7Fr5/lKJdr+8BQIybANPQm1WkgLbBKFQrPOuAb78qPKa9XKskHytxnksJL/9t9oE
5DgEXYAstMz7KxA+8SOys9ZwKCYzPgL7utciPewyf5AAnt1+wuOnQDispxSNP/+OV90cHAui957O
5exj24NP1v2ybf7EBbslwoct+W0sQI8DN5l6QQ==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
uztTqls32+j0EquYCpkD/ch1Qhut74rDT3zyKRp+PlqZR7k38IAdyzS388I6x0oyoZ/G1iamuniA
RwS2p5fS1ZZ5PAl52eaoEF0dlgRvBkWollttkrmv5IO4dO7U4P5mluwQCYK1hktbczjxlhoLgyHD
0BzwZyISxd/n4T5n9WQel2wG5X1SoShPkRQ4DpDVlR8pAkktSfDA+349X2G3p5O3rYYFi3I+bain
Bm9nm14O9vz83R67C9d2wF1UXxjNAsWxzXUQ+JoqIaYTi13QWPtc9JeZ4tLpw7aM1GcVxy3Usvn7
vg/JonqcPSTp25NfyMcPPvKiH/wKv7Y7NA3TyycyI8V6q1l0vNfmp8MeLAKnQp0ZanaiS1QlhDUS
88ICcOVAwBxY9+VX7TBfY6l8jI9P20kehimPgF5AVe+0sy7Mo/UL+cDF+JtnmPxEeKlrIT/OqbSI
Djq0F2SvLFI3/kKLie8QeuKsXJZVLl0m0ANx2rGMnZlb5G++8+EfWHsYtTRtuYtAZpHS4nWjajmQ
A1DT7mdb/0OfoguZJuiPCVyvqg0fH2Vb9xwt482rgFbKj8j1XLR3EuXQQse0F/nDgYojb1DqNP78
jNZO/8E7g8c8VJi0rjVM1Wy5n68MoLM1HEFlGrxwk+VB6TNZ178udp8iij351t10Ds63AelRCekR
upcW+5/MBNwkcCFfdb7W9ZCCE4hbn6dWSwxJzX5TnLuaMeIm70sbeS4uz7QlWM+IEYQQl7TuA3cS
9DRyLgVD3jbwnonRfez+NFGM+6mFfXefb4M4zgX2QSmOrr9ioG4HVZ/zkUs2u8F++ibsFM5JX8ie
8xN9Yxrru5OCvk0WiCqF97qsXyvcdZ3DuYaff2XEAbaURkQ0Hjs5I0p0aQr5aHSllwHpnGdZ4K6e
LKtxnxIINXL/vaZgk1ti+kAdLZp49bxGN+lKhFO87K2MhZDnw05UzJshIukHoejoNWDARBlrvlMn
OAj9K8sWvHvs9GDj/MXs34q7HPUKBsFeqj2MY7FWSZPkvcRNuubmx6uEQnXjQ4M93n8Dgg/u259E
3/+il8zRfTLJO3KuPQ6P2Lbxgzjf0u4zawtJgsoBPEoNCK/W8XxIueOf4oZb04D+cRgDfZQeWmSi
EO12o7kVEuQRUpIeaO+qWzp0MUUlemSvvtCWxfdBg8gEJfDqrWaP02mFVMWQfB+by/VZBIaAmxXk
RMQOpyq5WkDj8xDsl6H5fXpngoMep//AQXatxmWwTIpQRBHFAEntr0nqALsDq9/2BIb3XUFlqIIB
6uKbB7EXMEGToGw7nxodFfJR9PwJc0BQ+f5D4Oe2JT3pxyN0O1nus4vnKX9tt6AqeSAz8tkOo8hk
aPP+hAk+F3IrCdqYitTtAulgnBrP7XYLfOUOPKvms/e5vlV2lGU/LKvZlwyCr3Gfv4n17W5RpeNw
5elq13DSlH9Hy/HeMGjSeuFJ35w+MvyIkR6tfBIPSlEC8nGgvxYWwsleaAW+t62FFWkt9Mt3I5Wc
YLOkBReoRFmQUSDhJNPugTqEtMGRwZ9U/MQfxMbRUsrF5u/UUZ+3vHn4cYP+hBpAZ5Va0PaZ4onP
w2FySB/sFG5r5wY94B2z5InPHXwqc1Y0JV77oqSQtpEgs+MQwTD40CdWWgkzrEBvymuluYOOHqug
drx1VgbHH3iKL0LYRb116nhmbqtQ00E3bgYuE8gkC7vhtAuLefKGWpQP+IiuBnufvkDZbDJr+Yr3
TpYx0v35JWHrH3hy7FkjZGl7mwJBq1/aSrNmFMhKddtpWbzRL5r4ogMUwMBJoVCkkG8Fq8vo4rNn
3YYNVQq26GJR07nwhyfgI3lvVN3EbVY8FRymC70iTAzN27zzH4JlQu2wSoigmm+8J8cu12cdU1UQ
iN4h5GRXxx1FZPh0cFEFbOOZlEZf9odZ7MndIJfOZW5Rctf/D+xc91xi5EuYBVA2xu6rIWIB6gtE
FRNZBDcxumCwG6qvh7e+64fNtMKd9y8qzlhkGSwsdiEGAqt6dAaq++cMxSUewlvVqXiljtE8fGLG
DV5IgYJcQrLCfjzwKn3f/DPK6Gdxx/fgN5C2OtA27LArMQKIhazSRNq7TiAndB9KGdMd0uNvv8JC
TE0sOnMB5xVeHhRc+7g9cSg6aDRgLtRMWIRtJFKz5IsS3ySmHgbc1RvRiPSx71ge/uwiZx18XyIO
rTnGe4d1iCEOIEHb9V3DwAEqz8svrHY/vCOUXL5M7RQfKffXsX0o3ZNuP+WY/3YB2UWB/SZ4+5qm
pgknL7DpF4yTEdfMDOyoMZQrtXkXpM8nthvYB+Xruofg0qnfNSSBcQMOJob73Sl3C+yhtaae8uJo
xhXx0hAE8Txp5koq/8oQNNaD9JiPKg/ID+C9UFJXfsrX4zB0JXPxg+ohboF78IKyfveEKwGIAe2I
AQY4Qzx7DPIXz6ac1J+mwjrJbpOi7LWb/ZCN6PWt5/nA9nYwlWVzGinmLaS009r4yNl4LBAwGEvm
BScUwHvMKrjE/RlGQ155PkGvfIvXMCdHiH6ZOOKUA4gTXNqdzh+P7uw3lkObRBZNvB08GoyVe29A
9Sqja3I6ustZDOTxCKR9+OouPk0rJ3Imi0NC2lj8dTxRnV1oF3c8B//rOzxF/7Y98A6dvio/9Ecv
weZ6XjnvIeReGoa3wGud7p96h4uHRnJfpj7Eds4f9tSt5XUqAv4Ks0umufWYTQtitjPBNIORDdpj
tgZe4zyX1R6/sRZCjBKBiHDDsHRN8YlMzX7NbSQ7GGOUuyN1z5hBmHsLoJleFe+HbTOs7zCXofom
ybdCEdidmAMfzDQiMUkAMCi1q34S6wRcGeLHLEw1YGWgggNa3Qb0pZ7E1iiMJHl+CHH6WlLwD+lk
lfehzwkj9yhFOqoDTJcomB8GJBSKUygmxnGtFjzSNrKAMD3jX9If9rXDYba20RUQGmiZMldteOaZ
ajAzLkrSSk7xzPhjaTFDkKGILwYWwVwoFKJ7e9rFZDdKjU2xfxkyuZBb+YEhXXuV60cYHxgIcyEA
e8C8JHOjAJ5/ke0MoJIO2pF3lEjBr/V9FmModIuJIScUjWJ0OGHFZygDXTigLP/LX4yXR7jdNt1O
zgTO2gqZCwPxdoVb0LfiTamXoeugTnpD/hoIvgEgIfPtPH26lYkYxeeRwlaHYfemh0RZsrICkEyy
HxGAuUk5Rjy/RjFqXfyY6IAqyKxlj5YdUDkqNmylXTtVigxMtnExIFJLGXFS6dSYBO2VhhVu/LNX
qGyZBwQE8ht7RBC7EK04bCNiKl47/VXp6ALhiHVmDHdxyJFeKyHfmotzstzjI7hfXN4zkcaaK5Uv
4xdAEGaj/SbecZQKXwRF6PXlBIRMyC7ZlxXfwvrx1cho15hMmrN8TyaGd31Q1FxA0x5KVkKHUUQu
yH6lne8QwxjaYaR139LwW1cCYBg4Ow8J0Inhg73hcqbFzCBKcOo/m1T4Uk5TzsFeVlUk9S7FhMhE
aWljY6Eul72ooCzRxMKCjtjYV352ES9iaHutLkKPYdLuiqhJqndibrsgaqkw3QjhuVVdw105gewE
YBhr64ko6AFvLahG4XTrMtr66yPf5vOCWQOoL9xquxwRhwXkyEPKspUsHpgtUX9jh50zt6mGYtN3
jSuVhfWZiQsX2oL8SoMlYKFHbEtRjTgF/JKlPPF/GIToixhJmmLs0d76mAf9CcjVokUU0dbD5XR3
Lvw3XEBPYrpkFPGGWvs/QCJBpKxlxwaOrcy7GJYDw3XJHxGuTvjJu9nJq00IpY7WCJmB4/+OHqrU
ZHBdqbCKlaNaS/1KAfYfctj2gz/6YooJNmOZ8lnrNOKs0SI5yyDqN5bi5JUUlGaexHAYh540GCYv
vWXecwgK6tvoNc8n8yhzdlsvzIqnCb8s4OmofG+N13ZVhLxbdBn+922FcJAIHBCANw9buCVP5DO9
mZscchZmGBkcX6jaTOv4BIYxTKcVBltp3DZCUrxhetBD7m0wPe6hdA+EY1f0ELGGoKZ9a1zGjPLp
RQGLvvsdNIBq4cXX2qL6PRsXxjcTf1WCiYngOoP4Qv5uMIZdLhNHWm8D5WRiz+JEuNA+qklmCYcV
mdQzTgILEBh/xcowEG2lTB29u4FCYNfXpuftC2yEuSckrZ/61pUQbfNyU9JRCzpdB++/SYE4rhMH
vr5G8OZKpgikDFzTEf5niqx05hQeBSrnpfwkHbVxS9bCVZwEoJ8hNVC8Hld7X5K9tzsSaY8G5GD6
42+Eo0CwxPrgSeXv/Oa1CO/eiXUjxcZ5DDQf7u3vA+hCRxJt6N0PcvgEo+cntNeab4rtgHkROP2E
zFHUx4cc3ezmVq+/8z/gmyKP23oVivjcRI/tCQ7j/uT69w+4Yz+TUk15JCgCwfnZtQ5LFqC85Qd9
LifKqAP64KuTwNPhvvGz5rUuZwUPL5jkJlndyjmZ8r+lxuVZf30DvokcwDcEe6xMpZnbo1LB8z9F
/NEEoWIrbCUMQgc70cYLV/gN3l8JwmIbdU5Z0MbLnD1KEZ+r5woRqYE8oWYRj2pjzLEqZ/8I4ddC
8LqmbCckxlaQu0vkImrP9IwFcK6kcLPZkmw0L9l2+98nbbUd4pEXfF72LfGtKUqM3eW9uG8bVl8d
1fTuWupQNg2UsUiEp+0EEpjYEDQHYnvotRnhbXd21gzKqiYnxHUgNZx1BAWa28KApAQil2NF9q/7
x85VffwZSRLxrGd1nOI/QZ1tVRNF8UOwuvZ720lYS48n4aOJt9InRytUUqJY/RWR0O0tXVhB4wRl
II15YenDGxWNxKhEMj5Hv0HpiNZYEvL4hFKspxQ2LxJ7wp0RxAslYS1CCB5cj/5CQ2G6aQo0UvU8
OsIIM6617MGGGCLL20CdtGDF5baZ5hIucr/9I8klaR/xmeaXbfpULRIyN0Pgl3w1jgwiJmBvllQs
/YNVGEzL+Ns1XFi3JtqQDRsfML7jCnBrUCZf+X5H1AAIo/hV0Ry8G5cmJO5AMYVqZuA92xVsZWat
iRYkTZiYG2m7au2nYRAg2ViDC1LdQknrJZu5TkLjC+ccRN4mXwv/lw5fCbOBfW9dIuHxy5Z+xZkj
uDm05ttX0nH7wLV3Sdt3jo7W8TD5eIfJDncFkm8LN2HDX73NjmI16+F+G31k0mgrlllid4mNiww7
U/dm28Y/shxo0wcmxCwG/pnJUcq+4Av0oVjGVCBR9Ky8PadwkTJp5x3GeWd6LvV+m76NAg9p56S2
FKbSY1TsXlj4b6MD5Lql/dGE6lhlRU13IgjWFzgBKUsMNtwBS8m0IAIp0jRQvnbQpnP02C1Z8nHh
/o4UghGGOC/RPrCnikO6YQmGuVuITuc1BTHMo6v8WioxNKQLuKZ5EyUrn63aPenb8f7JW5G8ueTB
A/J8ZL0MHM8a318U1Dks5azS5JBsLottHVf4oR9uBkrFSwLV8D9W+j3ZIWYgNpOewzEXPHaiwJec
zRjqVtMSWxgS9bZbmbBbsomKDPuFJmh8rZWk1rgkfs5eaJf5ITXRabsCZSYhwmAKmKZqi4egOdgN
WzZpq+D7sshdf+fTlNeVH/BcF4IjzF6NBRQ+heJ4r16+UzKX0oLHnh6OlOu6Ltuyu4NGTFxl62XD
3VjWCeSBPL00OiKDRkjyvWoSMD/CZ5Uw75CJdX3Kqd6CXnZ+Dg488RFTll9Dgr5q8IDE9V1+1ekQ
YDLdnNX9WXo3dPn7Lt20OJbLFOHT7+1OqarGMAZuiMyYDPi6J/CeubzrB/x35YTCKOa7N4QQn2Al
rNFLx5Q3Hdaie0JsHnIym/eEf8pbQGSDjXYR7VjBSy7w5vgT+nh43/+P6nsBZDGxDOmB7sCw9R81
o1DovHp3oDCGDIWlDNAO2YEi2az3h799mcIArx7nA1NsmTx76zn9veZABcINpNtKf0f8ZPLViO6T
tT2t5G5ZgFEhRwlMnMqEdXDQpkKV93JssaR01J+slzldvnVA+3YrWb3eH4ljUtsv0CYnrPTwkDt+
/HzbMaZj+oxG1bySDpLCRWrW3wKSSWksKOhZ8fhPGyp+AxJ+2GNskodk0YVHpaVyBi8bNCx/MbpO
A0NShKS1K5O4h9Ow7+juB6YdFdGYZynnuaY1iVJrc5/wD30OgNVzE+m63Jejgza3nK40hLAX4oqT
GGjnCHmHxmmUNr+1QEBHSt6QZpYo8SC3CMG9N4JswBcUHiCxfDLrHUUl02zpJFobW43Qhej8bawx
Dv1yCBjJhaharpo7g96oRnBOE3s+C1YwzA1cCaSb58B5mm7Nd8CB0Zhzawv42ytyL/CTRuKzoVNH
dz/T60GI1HJeT6PsrzPkMYqlVEUyXo4xNlvfRLUQv/tLP1tGebeBHULLhybJSFggB8pEhkb6dw3R
952F3MgFYs3pmVvOZ1tQjZnZXNnbSyhPRZ9CpzQnXjaD5MKEDXwvSuqJ368FLemCCm9GHZt8DAvX
oxKSFSs8fAmWqAEKlOes2w5fhDCEMnLYrtFjJdtTIYYaM5K9iL0WH4cDFuS+ZxDa2rLIR773z+po
ZtKJ4AroGKNtLjBbGHP+2tTSdCJvZQ3MjGfVE8/RWJVfr7qhuuMkBRcjjrVBtahChmTPYUUHOaix
eIMHjtyZ2cd4498o+uwyivNQPcOdC4cbXd1Ig0m3K0pW4oLQKL+785Az5lzCmnDl4xtSvmL8e+Ea
GaLbwdgagmY7Gsmwbdz9ey11RHRB201f47wW9/AFPIqA40JAPhBRbYRnjZrf/7NqgHNQAgUzqjpx
NQVn54nC1HqkXtQwYxvUe7fSJFx3WeEiIu+RaYP/VQ1ydWftXNAT9xMb1Xi7IQliNlNVa/vgyjZm
ajWKaopY547yU41bxjSkcmdhcwLhL6ENpeaa00jj+jNOPNq3uKg3QKI7q216kb7sp47l9BI0byg+
XoXSxkFSIf6D0HvHmuRj1xwmU3BkY1+nl2vGSL7GKyCjLRw76nlis9j00wj2zMXlBSjhi+I3VoT5
Ew4tAD0Zwc4Lwx7ey2BzMM92HSHefh0dEtdrLCjnLzzDmVf2KCBfdQG2CIvex6ldUSuSvXxpAETN
Wppx/FD8fHWtvypuvxJMRT4w0YEmTLSYDncHwHhYhniGKSzIZQBVMuV4SB30VXJzf6EmQPffy+9d
lFnV2IXa0MZntIPTI4V5NmjeBMMVfwrU2/c5H1MaAPlckdy+BHXOy7JQc8wKmSFpV4H3gb43V2A6
kOSeYqNeBnsFt5TnjKUqt+pk+jBfwuFb8fjO9ZFLrz2IoKK2Gu8LeIhNHxJKNsUIrl2Ih2UgWEO3
ODbmx+KCFg5yDypnS4u4yWDjfipFHQTTlxTBoSrVtdIBuC6ogBtL435g5EwgfMEvRwhS3gp/n5/5
aBY6spqcMF58BV/+vBSU+1ASrQZwjO8uYzjXLFeWGFvY1JMxYioKlnwIIcxUt2a9QRUcYtnja8/t
/VCu3uUt/PZjdRXHiEAnz/JKOl9Z7gqbcFtUTHJ26lvg0rAmR3FeZFLNVE4PRjCS6ZtWxu4sqyqB
Uf4bZt7OMeUg2jxmK2+dZTNzpC05ptOe7zdKQ7lrqrayhYAJPdDzm8/tEWElsroZagbXUfbpCf/D
EnNy0NAr6BGMflRbaOmVygVR8+YzfvN0lgjO7dR5gbk89HEGo08ERldgjq/uGg0Gtz2zDJPbzipq
ikGxNdu4FqJzJbxSFXBwVPcMyeDtf78dC4Bqh4Xzejdmi47+qs9e3diwN/PEWvtcx3FhcreSHqVx
YYHAUaJab3S+gRi5w9PJjoHzNRxZIG9ujKaIGwRHSjpvvCYaMqjaw1YdQL566lalmPn7iuoUhSYc
TKSGWYL6Xf3PfZVwmsMjgTKmACVKsXoL0PeiYimehD5tji6aX0CFRyIfQx4wCzu9ILr0MfNiFjeA
OMvEg1vOIHi9rS5PjPmyBZni4CDVYYmixR1ex/pH61E9Ss4hRnMbiCc0cdXpdhZ/rvzOh0O+t5Lh
E2CtQUYigbLcFXIOQpKhS61opFCZYJ3SdRTAMib4sx2nlGIMy2qS+AasD2Kpf9nurkQKXU0RV9LR
+H313UAD6pRaoSuLkNiGdCM15ozScuf9wfHdWHR0VKI1jwfPboHgLPB8/ZcI7y4wENiCRD/d6YNP
1F24ROHbAcYUeLxcYq2bDTY6Cjw+ZFMwg2wj3wJiXVsBb9jQvFmFOqmrw/itCA4CS86DhdIFKn7C
4x/7UxANhp85jiJ6zBeR+elAw842Ckxd+GFa4is5sbAMyYxNEvKaM5/G8DEuJj3/5b5xnlzN5MG1
MxyFME0BeOeAJz/D7YtkMZfWilAVfrnNb5x3UYhPxC3R4TJxSjUn8zJqAGLEwX5d91i7EdCxd3+z
3El5ttaNIunDO1R+ujMUJQo7TIo0X/Y4TrqZDGBf+IdjM7euML3WWTmW0SHzvwFymbHFArD9+3Yy
5jFXbf0XrwpJRyvcuJdrGcliyGaZeVtGNvqvmz1lOtqThCkKDGl3EGHRGpp7bVq6GgkC3Zju376L
pFTDocPKdB11tdc7HN4uhq0YeI05O9T3hLFYLfNukNjwKxxZNChdUan/GEptGza/gKp96QvaROts
8AxBod0oWNNUIuRiGVt6yYsVmJLadRvg6WkRRnnobH8k/s3d1uJVk9oxqkm7nomBeHrasOtN779g
JyCHHxGhGZdxt/l0Kmg4IYjz8pOnHmBoxFWHLLatCu7hgEmdsFPmG7glzBFiu8qajQPDA2kav4WK
JTbGqB9pFtKcFN0pMEKPE/gvjdRqdLugvwLXdSqFgjjCataDvvXPdXnTPXk+DxBZswBulq0deQgl
LtZD5T/ydLkJIeLmv/NaP6ty/kL70fdeyysdCMPSkA5hWLZv3CoJ+SiG5YFWKyhMWEGu+2HsQ33k
V6klNsrzllZ0Ok0JVqgav+uRsWbLSrBYVrRoHqy6wnK7TVX8FRN+LoVxoQh7sY2n8lYp4jjQ8g8K
NK3yJi5PEpomxi3nkuhJvZWajawwxuROUPSP4YHPrxRuPx/XA4MixELkbExDIEVl53A4Qov6ztLX
VyEuuygzbOLXEY1FGJzjppdT1JhTwPcLjMwBvA+D8dF9y5zIavyjusIx6qhAukqwLEaPARAniF41
395CgHdD5bz4dPXbQHbrkHHqVz8Uy0RG5WuP9M0xGxB7V73XuKVKYDX2u9pIZIq7o/2mNQVmTdji
+lmtEhqNiU4SzFxyUHYTXKjsrPXWqVNX2edzpR44xTIOfb4MozfNpvoqccHBbBSlR805Pu/GguAx
CBipujM7AdybItQ3bCSGqrvlC4zAdGhhImLErscqGwehjCQ5a6BXpwk/dEBzH3AZqm/xoy64kn9C
tOpOru9c2EWv/t9arTMvBCTSD0gza0mU97SHFdFC6nob0hNPcEswDkNL3Hy9LRO0UdnphYWQS46E
5i9/78v0IeAkAsJeWtcmNetreyaFFsaq5gjSuwxPi93A0ab1/GtHtlRM6cTKSuJCBER2/ZipsyxD
+TrgG+nH2rcrU7H55UiF0qhUdLuU0KDXgoZPVGE2wsgZiwMCOyIv+ufEBmKky2RWmsENEz4LcXK2
L5nXv+9HulZn0S+ySSzX0bjOg814hl723xtvF33xFcupqlr+pOCAyxxwZ49OK1GEBtKMFRJGLuH7
o06DT4aVvCgwy6FoS83Zig9vL6yERNm/D5kExPTpwgD2vAGzQu9Ln/dpYGEvxJot3DYdzPIQrOqz
uy+/sclmZC3pu5b14XYXaRsDRZo/kWy2TP9lcPplx4EjuzzCqcQc0EAMUiYRaR5TvcLRnmG0idnF
HcfTY8vovdF2FsK962Xf5ThNLw12hEXW61mMk2nBWwz4V9GZFu3bcTGlawwfADUEfg6orHLVyJqr
HR5Ea2jRdnthQh1QEDpmUERSSEBvEz8xTGHnNMt1rjMSFY839NoLvuXcH/cQH+9Q9+rz1X6Ixvbj
mAWZx2FRfS/royS8Ja9AuMUQikKfdpoYCVpmPC+/z6beuOOCYp8n+S6cU2wcstfKCwdYu1GLqt3S
3YMIMKqdj2U8PpUicxq5qiprMEk3l6/tsIuotLO332OFCDl4+HWXGu/4lDQOFn0r+MU4kEyFOntc
UWHfsQVLsYoBXhIkkw6EgMGCXvaVClAvJzLpe4C+TN9iZPgdZymDkz6IZ17/t9IGHwgoXLXsiRTB
jAQH8854tppuQycngfGFi5Rf58WcTSExKTlr1zlqCP2dIpN4XRGg+YgAMuxSqAFyRqXvKV7/bgPX
Sjb3d9kRp/Qo1hIFdiDKV19ULaLwVLzKegZPr0d/J7dNs0MYKMIXRDqeYpU6MWKCcstHhLKSnBD1
/+DL/cv5N/T3OpCh/o/SRhUw82Fm3pR4ko9JBPS9rnBQnhPcRbbu8TzJPFZC8aR15nHyzep/uAXD
Yw5+ltgHCf8uYhMQAoV9hhsWI3mofBhYmkQ0jo2iirlrOdLRjWJD8yKhFDCvgQQlVOFPe5GKmz5X
h4l3T0qsX/jECKIMnpWoPjTbERe46yJy4ro0jNESCg/pta6TT05bFq+Ilr0+noPMgYtG6Sq9b9tI
jWXkUwgbtjLqWlbnIBizXQi02DAseW+DdpY/MpOIXv2IgVNQnXxBUzLRwxUBn8IoGW166nlfkx47
hja7dUSDJpc2zrKT2yjNV8Qa7HTzYtWcU8yTG35iO1DncHckkG0tySKUHJS0FTE7+PUZ9cdvOpUq
zae4m/aYFDVCBOOpVYkYI95zYlQtc29j9cir+TyVISIbERkOIKwm/ZOKs9uUbX/Onip5GSNG0MQ1
SVgUXeE5oyYvKevDuZijsurdIVabgCbYd7ieXH8wgVBxuk16VfsAkSXGuVopTfbpLITq8vUyU1KO
B3i/+7xg6S0TZwSDIrTLUMkfuLhJubomYvpjVyDzSlf29k8DqD+sck3rQ5JzHrI5EjEqiCqceZXx
ciUJnf74Ioni4b74pw3vCiG3Id9MlOnbRKRgiHivJiax9TSfxTCyKDCXtmkt4ooUieN+P4CB3Cuw
7oP/A6NuJQVRkhZZH9T/rmj+smP+Ahlh1Y9rvKDjtpVgG92waUqea3s5zk3/CdbYEfmX3MDhjzXu
wlPdtYQ93QS90tgM772F9kkDH2BgvuDDDAM3xwyepHyFB3FlY8kxhJL6gWZqwIEBJfLQt5sgoTRt
PmMa6+sH1rguH2znpYcG/1eDLuvWMbshu8v8Nk+9oiVDwbTnsW30jQltZSFdnmLyTKZU8bzC6eG/
Zlj4TY75v3Wlj1fF+rm/jsWzXFeArGeFnDiLxIO/FsDKFL5ZBm3hF9Y//ZaSbwhkwR/ie0dQA97V
wxxRR3zwf6LkIOSRs2DrO4YFEginOZtrDuBx7pfU38kqAR8Xe1RU9WqrryvwCRfkoAkm6/zUAdnl
e4yhizFIeSJj9mnWuIS4IG9pZQkHzSHsll1rpPctzdWnQRVgWTOMlSw27Cigyjn2rnUrDSPWaMdp
sguYQE8gPzhsJU+i3JLMDjXpV+o5qwo7FefetBjVhrIq+MqVHjqQsr8TFVo6TKGJG18yZJxPaJh1
5mcmzCm63JkBP/3ZVTci9sQXvTQa8YwRaMn94NyOwctbfXBXBjyjCRXKQJHCDvsPzGM/F3FNndLv
eAQjYadtgis+lO2SMBS4dgMwEiN4uQnvNRZ/Csgm0ilXOakrM8IsBd8NvmAjQUoVmr7+FbT9zMpS
wn3f3XohIE1ayMzMwE6QCigE9Ct8qEX5V9yDsSVxOAh9BcSfzxziQCyKeuoDa9gjoSPq0gzDXuWa
usM0rFwjdOEV6Z2XyZ4/6RZg63b6TtQgi08mCbRxl9p8mpdll/PoD8eO1U7TdsUUmWmFqBKdZwZP
N9vCLJfZ6Ff9OIU20YQkHrR7fb+VBJgiA8b7ZwDCh5WV/Cn8ayGcpy6fZ2f3xLL4bdnhWM2laSnw
gS19zvhqdkeco7sE2Fj+Q5A7hvXCWZiNwcTf+z0DpJlvEBU9AP66t0PaL+bHiccW6EfNtzskLsNr
MuUk1/E2J+P0LQjRnwMv+qK3MymAVmYBY5cLi9zTJYd7W6U9U5bYoH0rfRDWCVBGOQMQdY01xUxM
nZuCpgtn9TjN+eKrx7HvuVZdnoPzykHjMDrZd0+iRZ8GcZlMijm4/s8WA/kPNYzrS7v55C0fPTHV
JSlx8oCt/IMk0nFJNnfCrkOg7VFlqupACrPIiqv/L4wavEw/Sl0s9vzETKJHixlZi+ZzWop0jsVS
3kQVsECW1gvAuTQeAN38uMr0fW9FpfacdUKV6L3Ao/fV36Oo95I0gpJOXDMs7N8phvc+Ih7pLUF9
/2hNq/ZIFPLfqBdig+hPm+/ixCiUAsnSP04ZdB3X0fG0N+yI7DI0daO25cfdmhQ8aWQ8k+ZT+z8F
NqJc9xR9CVj2hsrvUFF8ag3QCC8I6X0d1Pl3RJAxUK6Gr6jInaoWHiOjSEeCt1MikkaPE74jeNZF
axzM++QdaZAT8IM3njl9jngWxnZvq9KDdidTgBdFBVwemOT9rP08FL/0T0UI3O2WKu4A/3CHCwY+
dta32PdZ6/fFrgK7/QsHPF9MIZJrzRggkdwwXXFo66CHFS+BagzbOhMgNl+0X/HQHkOu8lo8a3/w
iPoeI+J5tBTWbPzt962Lm7J1p3sBgGaFIT0GkCIcdtb+fdSfeQiQ2qgvqtqcQCZHmWPw3Hkq+dbN
py0ddJN0Hy8j+8s69+abbaoI5fs1kAhRwwUgJI44S7A2HF8OvevqCb3znhdUofba9AgoxsaOtj8B
uR56Bv428IYG/VTwcndUGDN6V/CrNy8z836xCsoGFuDmeKRz7ghCyfXYkUPu+VlF7jeQg0CqZiSX
fZ7P652dB3DZLDE/bXxJo+nF2Mi1MBkcj/t7Dt+f59ihm0N2R6J7zjp0itGGpCS3wkw5vImaHPxO
uBYU6oRJV8NfvCBzb6jfJWfZqPGx5TOeejLUQ9MYt1anVXRy+ZzMS11qNFawdWdhwur2qxTutZVG
jUUUDVBZvOY5I/K4xNemwZyukqelY7j9dw9k2VD6gEWsP5NRHaLZm1aJs5FsVPrrV6nXjR3xjX7b
I4EzIgrPZpp3Yb7PEgHiH7sp8GWmDFZHzh371oh1QJzRDe3rWdoo/h70TF3QEXoWTWpUsFrw7aj+
SPUML+BBpX4Y6MHrUd3a1WNQLLoNziTcZa5U6Oh/UZtQbc+2REuTrJODRddNrGOziRI3l9RPjjRq
Wa1nNYWow4nsxwDL0eFIOUdgvPWX+iZC/pALa4RYswBKFHYOOd8h5CD+0QS5mckviC6DFdjFx/kY
eh8LAlCecQExM89OHylOd2+6XMM1wM29ezIafIzynY6eb/sUvC9ixFwegXuKSNSHGdr/s6+lsZzF
8iYsn28DDIkeIsJBBg8FGFJgLD2eGtoc64umOz0J1LgTI/c9QaCxfaeWrQNOj+5rj2a8CfAvSKCL
JEyZIiWvD8tXzzYI3j6uBYAUrxsKbrA4Sv2xF+4hBdGjE4OenXo6NPw3lt5/U7ABKQmkLOPFNQGk
E1VUWMAQGMu48DHS9qpz+Dw/ryjrGa6Eoa3UiJNb/0ROxWx6tadHIpjySB6F6y7qRgT5Ubcj3W5P
4BLrN6ssVde5Mu6qqVlVlk11hAh1SvubqdE/ofMjidPtVdAUrMAraiC8UBKFxaBMW+0PhAJLD5yG
lcD7JhBrlPIX41nlQvjMrUN2vMsyZlaJSJFbz81zO8KJgBgRNqzm6e3pNOWP/hAR9xhEJC2Fi0Yd
wWtecFw03aGl7sHnSkEBRYhtH/G3YPk6EpcvpRCBdUYyLcHfmY1+G+Ie5tYLvHW6aztXzsG4KKI6
sILxP+rHGyOlsaitOY923XqBxEWSZFZ40ixT+ewiQsAGzGj5Hi6TjF/Bil7KSuNzwj3y9w/Nl61g
lh68w2CQLEYBhT+MVhpPbuHZ9he9LSQ3gudYKzX3bxXzlPYddLifhhvlyLb8LVzUUs1o4eooD2Tq
Y2dhjWeIq5RibnMTX0tuOctqV+n0Y13aFEk7+IUXOjBeZG+VqjVcrq7EQRMqX4EmuPvmIrOn6i2f
jLyIpzxCSvlxLfMb+OmW0D33OVXsDjmXePQloEFfkIQ6TSw0OWvHwr5f9yKJlJ14gKFG5job/5ak
Z5MRzpxYnADkGnxWo0UygrH8x9q9WsyfHvvbZ8YlDr//unIyvba1RVUZ6LzHvSTstQoWf/KVkp/x
RZoGsrzmpRFYyNidfzYZiKFAnlI7XouKQjC41ofmPvPOKPAnGfk7yAX+w0F5DMhsIRc/or6HLLXB
+oylnjRVFO55yVI874dm4XP+/USLTAhMXR25q+rWh7tGV4nv9BcliOwXLXOVuDJwk94l+UigkfV3
a48anzlciUZ8U52DzXPFqyyi1Pyg1DqqeXgCKC7m0LylXV9sNKv1D+7u0lxUBD2NDzVj5TYdqv3Q
DwwkufbT+zs6LKhS56fCmjqbb3SrgMX1U8UgpbyKZ/wWJsrXtGqIYctVv7Qy/H4kyW3UHLQFIz31
P8kbuzE7a5NNbqMrWa7cBzF32XV3BELlIyxFPsSweVBGNyDK8SdmPoxuTec3U6Y/gumuwS+A+Ktn
JZpNGlKdVplVNL2wRff0Q+TQyhrSrWVJX9r1q24b+X5czY0D1HVau/0w1wvCxmdj5gzAG8TSru8/
C8PM6SG8uHw2XKsxekhdpguP4au0zqjKv2mzBp/TdJIvZhfVkMmBXL/nrQymTmOsXfvcPZLXKWfH
4B9bS51LnOLzP1pzpSZAOUXZiut9bMpjxmDZts9853mqSGbRKKfhp3V0DiXY5NabxQR+coEjQ3KJ
gN4sxOBzpjW1aFgie8OktL+5dbxi1ze//F48iDOw+BWWNfIVXylb1Sa5I14bI4S2X0OO2Zg3P5k8
dsscQVOwdjYaGtxNjJRevkVTIZI/35orXy8Lrlbs1Lomi/YJa2r3dejZy53JJR5NNAIs82PE9RkJ
dZXPkZiqsE33eH5fhGDjf2BjF0sfwTEYrf3RVGiEenPnV8mzqZMka35cv1K2x/MI+uRp5hUTiNS6
gAg/D0mx2mHcU3FIpkqWgdNeTJZrXW2yjzyyDI0vV7jgIdh+utwtJgDpjLHKS+JnIEEtTsb84tzo
dAvic5h1aBIO+sLbUPthQwjz9JIAgpOq96fCJPMRTGVWu1WM+eyeI4o4VB0XJdb5Nkn2hUXevJgW
ZNh/8IaCFPRRKcB5cqlKnSn79jxBjNcPOOyvF5fE6EbbbD/JMlZKj9b8IZO/f29ITRy3GRWjiNIN
IkcpiS/FDeAewLF8I6oKsWnStchHMH7opSKsRTOPKeO0txqAdcWaklIFSEbm3S5ik0nbF7X3Gyqr
Fs/f0E9Njkq+E1/hRwB2hcHA3rHLbpqjlg/oUJ1zHzF9vw+aoOKX8k0yD40C/YMXvtrQ01hRVBAC
Wjbpy6riLRszeQz2IKojnBIal2kSzHkYyDr0N6M0Wflxdbt+yc1a1wMyPvLXyXW8sn6YYE+JEKH2
7CF5pZ64ActiPhJamU7iSyMr29+wlq76XsL9AohsmfMgvlQPj6Ady6MiBUrtvftbHuRVLQyeAfOC
yNi+Sabw6JVuKHzuOU7yf5uC9Uh+JIg5gimhk6uwG9Y7up2NrehTPbWeeM0clP7DHBlZINqa+apC
bNQeNSbw2PtaOOhoMN7yp3//XakMSeET/6o7wu+rOeln6bi8Io2wmw1/e06jHtZVtTZpY79ciHON
0XOlKAChB0gU4Fzt+jMs4axpWh6XtMT1QdIp21fZckf4TTFepnYITWE9/3Xs12kBSAI6jTQgc6Zb
8/Z/QxuuvmG3SMpEE5OJKR7syn/2qW3Zh7HSFpkZxMuRni9QOawIDoPwYptSDQW2w+WJ4p08MF6f
9jBIxxapHoOKjGa6oM/AxSOI4oaCOKdaI7NF7s9PYf8g8Chb2Rof0489PPjhGSkA5hPWBFo8Xgsj
Kgru0XZ8XHM+Zpn7WqkNRaEh+EpMrANmCzH5DNiYNOCCvbdG/vETW7ifMAoFLvOdfTtk5Rt6ZInp
BFk2thIFMddb3AKIVx0UTByM701Vr4BUThgEGAupAi8kWdXdd+I3z3vaLEKfaqe/byU/dkN1FONR
wZF35cDv/uY0ijeeQTZFcbVBjWe/JqGgwtc+SQ9gmjMlD3mYHFbnEtHBwBhvYQkq4vV8+ElxItLi
0eHzL2g1KzE2BZaFvqXiobQ7HIWzeT9mU+jtvbOsDnGA4PNfxVc1jK5Ug7zFPqzrPVzkID6uM6GB
nPhpj33bzQcwbiloyWqnNBhG+jGxm8HbX7wl5GXDoiwEA1RtINiCGzVeuWwDYR2m2C7UkWSjan3H
Tm4b60IYTBC30cqU5Iv4Z3AYLB8FmZGespPGV05BQqEaBslXnrE0kGDVaewOsgZGzK9ahbgwMXzo
gVcbZJFxewaSfVkxZrNEwCIN39btv3CojwTjnbCtjYO9mEBxdk/OPP1FAklH//BEobfR3rKO3plk
DfH9aWPDXbe7aap8NqGxqDsSrQCO+Nfb086HFUFOoKJe8M0tJ3AV8pNKq5EYR+QVDA3Aa8w/e7Sm
dzsnfjctb1kutvzmwTV8XFdcEiFgCsJPKZ2BTVp9xNn3byo4S44dmIaZ2c8w3kHOR3SF/mNhQ9Jj
TEJK7OWhAoqImKJ9RXULgTrvvljDdLn7tZrs9L2ucmRd0jytK2bI2L3zD4JC5EwnXH6ujymNEuJD
tGK4VcBJUg7BymDbRs9vM+oJsAPRD7VrqN18YjeywVoxkdfjquF2Q+jaCWQdLdmnN7OegXsWJSlq
dtnNjgV3rtmJ5Md2IuZyLIZHUAiyQlHVjvrlqs2ig4Vn/9ATCuLr4QYQZpqNZ3atGVD4KJbm3qBe
aVt1OpaFvQrN77n5z1ue2wo27WHtDb6EpCsXCqFSesY7tnIk99V5Mf47pLi9MFz6CCs625S6r8D0
eq0/tEY/t+aqOAtK9ayNgtF6nX343evzodAmWQYH7i0V/VeMfIOgU+u5dwHL4/NqN/eE70CUviY9
yD6lxwecMd6KZnEyd6bJd9Qh+zJjEWKOvrAsUlDRlUmtqUy9FxTqpGFrfIir5lPoISoe3dEuoVrv
EIhtqe9rZXGgf5+iZyMk/ZWnpr+hHznKNgoYZIexIH2azb3/CxeLKO5TVUs1rX2QjlW31QyMNXwr
sqDj/ZGoshge/KQe1Tz8CsLFWwkjp8i0KuRYqLVcU/JBXx+VypdKsblgdglWSvy7q5eLDz593W7n
uTzZjA5yd4bFPCJAn3gZmqSNt0G8ZA+925hktGnbTCNE9pPA0s+X2TkisgYfsVq+6Bf256blMqNf
uQN/sGDML7o3GMzM7/gv6ohNt+N22eGPt/IeOmx1imH0oJj/3ckem4yeh7prk1HLDesjhfvcbjzH
1kZbwSIoh0QxGnnQBy7YiU7aGPZAuVka/IJIaaVKV9X7dS6jyVa36bw0qlN7R5Jy/7g8X6R6cXgJ
+ZXuvQRQVSLPyPbwPPDYXI2t0mwt23faiz16esqmyX8oEa0QBZohhq6O6ibunt8irZkNkSpQ3ec+
vU8mhiByA3vlAJEjBRlSUEDb8spqlSokaZapC0a2NQje1unwjxFFmBzxBk3kB/VjigZ3sxRs+k4X
n7VJyKsqRGv8Ntr7xMGmRNFC850/77+yuJJt6JqPe69r6zqsRytWtOdL+TwpPzCA4BIRtCAWHp9z
BRmKno+nNrMTHg9bR686XmCeJgGA/fh2E0FX3zxN8Z0BI4dmbW8TPbHiEghB0hAg3KGMvLJcfpzZ
tpKKbBJbS8oTh2va8BIJVUwKiTym+BzfGKQVzqo8PTuVUIHUbJPx74zedqrMnPoMoQOF3CtY3I5U
FZQJ7bWehH38LYGhJpxxgKy3PYwCKfzMUjZIMSauBkIpVq9C5zmfTSxD4aj2cyIX//QMIOV4BIvP
D7E/s4bD5gQjNNdPm4oL4RQnfTE9sJDGGe6H56Jb2H4ExIbYO76T6C54hvdUXYdO8UGWYJjioBVr
ZV46gydk3L9AuoOJrTJKbFzl7UJCNN0jydoTkdpc3/mak5i8mQa9swKyEJKorb1DqfH8AEdBzLzz
gp21My5fTe+afob+anLGXTM0aWRGHWff7lE5inJQa6ZusXAYpm+y98mgGtYsguzHVyJVj1CMWBS0
L4O/kJwAvq3CSUO4Jvfy6rvoHQMCRiy08rBU4SrS+TRUyHt93sUVh5lMtTnVo38FBLcZPzM118Zm
/Ra1np8hzI04B8mAZcDR3eofLd9ik14mobkLUOMV2R8+gpfbNX2/DTcam0TIGWe5tF2FncAvj9pf
NdTP/LswFVDpSfzePp61h6f4ouStYXleE6B0WCCGsE1iVKcc8ol+JEiOBLtBBsdZHREPEEP4OlnT
/FIJRimBUvoEU4X4XQ0fRcI995cASXm8mUjpn82NCGFVCYi/ED4CPbnT/opwbhIhXMPaGamivLrS
/bbsMx9+YI2UOOWIQ4MmW14ttgBPawgnAp9G23p0CpyjWq7r17ZT+XLn5BvngjA5XoypOhUpeHJZ
dNDOqRcLo58SV99Z9G3HDYDAIO8qChFUAOJU6+m1dfEss1vFHlf2uAdiJZe9X5R4+skJKniEAn+O
jNz5Y/oB8XBhn7R1y7g6WFy28u6/5C6DQf2XE/dpe2b1Lj5xDf6xl9a4fnNJ9EHvi9XEZcyBbJcz
+dV3xorJ2ivWVlqeOV43Tqcvoq3J5iUa1VQ8E8lnzlTTylWYJEb19k921MguMK8Jd/oPb0aj8oJz
aN4EPB0PFy5ENaLbZiqV+vZsgjJUfhTQuKilGucSH2dxOmWWUxdDOw47D5S/agYFShJI9myYJnKV
7cv0Wi2Rcd+uXhbLvAzGDGcF3yagj212R3zGSLQrM2XbKPPNCOiNmdeyHMMpvgAuw0yigFfTGgh3
O3yFm9Uhzh23hCJ6uuMboYVTaNCH94sz8t6dNagcX2J/Qg2EICqJGxCBPCAn5e8UCzAY3mIMU6FN
roclJRgicO1Ma8A5rWrG8RpC3Nv7vqJta7Cdrb4NBidkKMBiAbky3nnkqpOHm4trfDGq2L7IVRVy
BSctXnrdkjGVgn38DWSdIfgyZ6ZXcsiT/YbsWEf2pzBd/rqkHx5BnTE/hc0pL+yFSgpDoTVci9wQ
zwbQt2az4mQe7NSm93fQl1JvqFR9tQQxbP63t/i+UXjwNqfU40DNUrfLxEZXWfgdzhk4q/ccbKQF
jXf4z2tqd69/tf53bBzLP4SIja4s3SED9Qpea2mSmGug3gSsfu49C1M5AZHWQqIBoIZwk2wp53bJ
DS0PDoSR5xAS4QiWgKDjxqbCrw3rw1ddvq3Yb0K/sKNPkeyCAEacZdqdpUJ7I7gWJdCOjNm2bHmF
bgoGwpQWOXUYqSna4TOxko/+tn00QiCdyEU0RWSDKtMHhFAVn1g3PzyvkEUlbKYgXdu7cJq7ZYDh
9dQfjCQJXX12FDPBgDyNPjWZ1z0PsoqKIf5lo3yGRHoaq0bAUVLojCDjDjYlrIo7tXZj2fXtmqfT
5RzgsNdglvvHZ/qLsUnllDkKZotuowf317onGzGRDGTY3uOttmCLI79/NRTdtTVAcDaJg29v4IvF
hbTetbprEZnNp4U14+EatInZ9juTrnm2HzggCdx8q5NNN+z9VzdM44UAsckNK4nE28azwZpBziqN
RsqV3bLxjWjJHIsEPrGaYxrw7kCB9j0GvljYkObzee7rfBCZgn0uCrFPvdxCFmjCv30erw7ha6KF
aRw74PfmYlngwy9543fka8pK1J4QtOrr9/Boy8ZknwCR7QzIoyggKho17RcIGjo9pDPAht1sqtjn
T8tRsZrsTmtWsao8rwbIKQ5wkD0jWONv8IsXvedG/EqxJgNNT6MvVdpAlv9VI3pa72aHOa4y14KM
JGkxRfgxg/I6r0F88wIGVv9qV+qEPXcJjr9J8svuTt5eX/LRnHOpAS7JwveS5tqBLozxfaXnYFiD
srStpTvFqsojFvP8rmxM8HWx0nh3TUIOwm/+sL4oh5YXPIHbbWQMWtWOytfbi9d7WR4Ofgsf4tNU
aO+bcyUrLlf78FPJKZ+F9IFzALch0cQm7vNNeZEp6PAdCPT1RORiCJFCogZE88YhlswONl22Egyh
xCl5DYnMnMy2/8mGYOkkbweq53iJ1rWlqPHf9z9eO7C7ADQKVcXp7DrkLxNiPdeCEIDmpxo9VRdZ
k/RI43NL/Nu4/geX+fAAY0xdFh8BmyC4sQYOzj016DFPGB6VNb/4kVIpN9nzk55l24PLYWI0RV2z
FUX5XJO6WkLgS68/ZJJnDzEumwyrC+5Uxbpj26hDdp1qRBNCdXU0XNHbQropJnZFWH1u9urJSKxB
XzeMyyvYrZGYWIUrs/ZwzoPI1z1ZbDcngQ0suqJv7XgNPv2Elbp5CTHfaUN5U6JZ9N0kYmrpeQFq
5t+yZQ8tuHh4NwcTNYhtN7DPI1hmLQTQKW70pwPXD0gpjHLfy+0+3ueTu/HpnBSX0o7NQzOoQ/B+
NR288jrcchIWEqAp0BmiONuIZiEbjNGqReeL2u60GG95MN8YhoLOD3sn/6U2h9M4OKvXtvBO565X
pj8x6jjB8errTpMDjPiQYR4ZEPiebOW0GZOtdVjRzYSLopBU7XoLjTaXPxQhGxVXux2yTG0IqPRH
eeoAerbTxTb3gVX6DHG4rWwXteWlQdoronavJhdH7E6AZDhMbBY3UYTFdO8SKSuk9vHv2TM1xn8i
+jY4aO2079rV+GS1SXqwUfjbhKRnDM7PB7ieh21FyExpFPGLIYXM3iaq6ViS6uR8sYxMpv8uJHKr
UgX/ngb5T+tmUU4eAv02BfsYhb4kmquwqRRlDTndH9CrXM8fd60KnDXrhQO0Cf6RPmPtG/pvQInZ
GRWUrQ/NoDbdwpDU66KXBdlX1VIyo4bGCc1oDQL6GYoWlx1VG8uu6c368IBIv+j984wm5qMepaQS
0wLlmlvm0aJ0eh/xJN4lJ3CQfvhGXw77x4iP164BB53KlBXv+0GE06jTWoLDv4HwQVjhTBSbhUTJ
EwlmqnY61zK4tbjvy1IpclxS9qNqCxQQN0Nj5G7cuy2hxdTLYBoQIyNBucMgaB/P5w4brQsyZvvi
pbPl1TPG4saV/bIOrdtuSVmROLVgZT7vPBUNTncy5N5Jy9/qdb4pQ1GqvpPw326KnTEfiVGFlBFL
Z1YfZ1c1BIjrfysPvmkXek3xaDc3Q3eHx2EXqQayM01CRF+IwPrRuL2l5JKzTYtO5Rx9oZEQpINp
Db1itBNwrRvEU96iCGsNLdolS52P04NQ0QxN14Gl0YzNS4rsvg/psbayHZY8W4HVtIq9A01AkVAr
TvdAR7P+Kut7BKDqlsXY5SwDeOMeqd88ndYWMrx1Lgbzr4YnPO0F/Lonw+Jss139h7wIdOLriK2k
PcS3urfT1DvJkHq0w3kTxViMreoM8NqS3BZZtkEmxP/jc2+idQDoWN6Wa2LZHwOICRigvTowNAus
KPcmhjpgATOHINbBKi2VRfUAzUerQzcdL4TMfeHYW8l3M+kkcx1ZLOF0A2P21uWUAUMwn7U3+3e+
qU8uXtqyF8hN8H4fhSS5cy6rvlTzrDvGkEKjB1rR+rNPcxgEsrfwvZ08MgTuHI2L/KZ9gONIVKmz
xXzkPH+V1qnPfE9qh1pjVXEEa7nCDj9AqT1URQH1bRGpAT/ymbm7AJ+2P9L22DGohv15+nLq50k8
0Fcp7waWdz9o/0DfsV1C3ceIw2flZ++9wUFhCMeX/o5cTuPoY4+smpgwJbmadff15LebL2IgJVw5
nJdkwqWRxwTbRNxYXQ334PRJXbeGwS2RPf/FoD2aLQlvhdtT+0RzC3XMjF5Cd4b3sNCEz0R1kcSm
CVhB7Xgsyq+MAkSYIhDjx5ilfIUMJCYVzTOb+LJRzzjRnjXXRgoCG7L+7vjzGHEYYXumnmDNUrNn
3WOxOMV1QgKSrVP5bZFlqnV/hfpAbKbCCtTIPcM1BHSTSG6VLgUKFf75cqcrsD49+mQAQYETZ2mw
bqAt1f1Q1nVclfA/Ic2eAIeEB11gTJMDEjW9mjGk5FXu4e4TkGxJlt92BaFtZhj+qd3o8L0TMEQg
L2bSRi54KFxENtlr8CHxw+GkLmOFK1mEDWJE6a21Z8kXrND+DGBM+hlhFqeHvZ8mqQXkquvd0MV8
E6j5OHM8aif8rzgE43zXOZKNwvwGj7/dGs6a7Lq7N0kQVZww7dgkfBJis1uW3UQwvaBUzMBikBM+
mXNbLr1Fv4BZSFxFM4jhKmiaUc2TQkuNyrYBCkrhJr+WqgkPAzPzpNO2PLRDCFgy9yhe9TO09nwI
bDL4sl4i0e/Utl9bttoP/kT0wsL1sZdWx0zcrqDqvgQ2Pkl9QYt8ee5KLjNYrRpXK+/+qM0AYpE8
H/YJMrHfPLjXemeHcPSgl7XZwbfHuuyq3fDs4UiX29btm0n2M8efkAy3CR0jjHquINU7FXI2vzuU
eVAkDRQw0EvonTeNJQuSYcXgfZF6vMRFGmtxxBaJB3Fr5tQhC3MuXTuEevd3oAxJcjjqPCK7hZa4
1gNT2Ga0iGEpOTTi3byr/7e8sJ+GZI3sdsHCZJw65Cpj9H+dyb64O8OJ5EUqAR3GUuAFpftKkJxC
/+FQ4MFsGXURE5YRnYCV8Qp5QQzwDZov/Jo1UHTXNG+0ookgxmLVgPmgV1NIqhYcIFXgib2BOYR3
TSE7n/nACgPUxBIENLXuPNJuN4K9I6w0PK07Z/kwynx+CAnIsDJnVwA2RMELeyF/dj6Z4VwUvg6b
ipL5Xf7tKE3Epnc6MuGSoTfbDh+8gzE91o9SWlTNeBirYrrKqV+7JAnJh1EMmP2SWP5NmU/zDClv
6gcsyk6jYBa6nJ+LFanIZ7Kse14qQHBR1QzQ4BBvYkJOqXUAgS5wf7XzgMZavOCdTKKoZgh8gt5Y
gXG8Of+Nb6WeB/ofIPFHlMsYwZH7VR9GdFhRvVpNnfcVk2tSvCqgNhMpG+QvPW9gwy67oQsoeuRS
pugMZF9s5RM9rsQnWG3piVY8ET4H5OEAAfaMKfuex9YMI30pfZnMyec960LdpIMHxZ379JzlF17Y
/W74CVFuGbKc2vkkGh/bGE0dX9lg0WfBXPRkpmSQOLvtN6ccLBbhLxkeQcUHocH5VaG2VfKuaGP/
v6ceX+x477hnwi2kcmUd6dA7QWzKoB++AP3AyD3+M4JnSmB/6JW/xoHWyb0b4UeS+8D/4HR3LS7p
P2toxvubMLC+51v4KAUJw8pqYQH0dId1EpdmxeTOjNW+gB7gKYNT+IMRgiWhtbWLTIePa1OgxvAV
ttvmrPiH49D1A3twQxjbRWfeU1Orql91oKmFJZx79l0wSxY7XfuB3RSJdiC3LYXULh7wv5qzuZiB
6j5sMUAPK0U+fSCTNLiKALGJGaKXOISOLCZ6p36iMmVn9UcoqNMajbkRGFvhpXsk7sHFU1Oiz7dx
NoZUhp9s3xBIh2rkRpz/GI9fKhkV5oWNpgkS3V4p3Vvi/TbB8XVBnrbz7jLm0mJLtfFVlKZM+l3/
mBJVM9de37HqCwUUf4gIoUTzFqtmxE5XQDMT3TbSrcU40YIEporatclcuJ5oxBIumjTk+1cQG1Wk
6DkQn0FMIltRCdI1PADJhD3c2T+8FPraFFWVJnwsSpmZ8w1vbrsMCTbPubUbqFYX5u5J6/+K+p8f
QnnFtEwqd7Zmm+xJETyv5qmqVcF+TK9NFD/c6fLFrbbwRTXDhSeEhKUfwTEU+gAH+voREeBu+Cu0
b+uPL/gd/1gu8gkvHHHZmYUOZxjh1FQKcbkqzqyNVdEHbjIVfl1lKiwBMDLiNGMTo++JN+kPNtV+
cmpS5XwbzIA5HLKcOmDogv1z893Nq9I59dDU9z6kqmTSO7d96KhBm+vOtDWMebINz4P4Jq8UtJiL
RLr5yvvs2qdi9GRvMc3cTK6kLyPNR4wuxpGbID1/daLyYD/Nz74ZQm8wuQjFyPVFt9Nk6AOJWXP8
BVo0lFkzPBRkoAGdUqn12FJcyL0zk/BlFKrdUfQjg3nC6sVAfybkW9xo9pnKY3TDotXbiVTssz3n
s9IbP3jDwP3npRdizTIERidXa6VxW9dgIfsZ95Ceqm1NWFK085ICbD7r/dUYLoAjGKeDdzTkPEbc
sd+e8UPqSYRKo0DLqV6cRSAdR+O+RiCZIBLgGENC1SP77+FMbcUohRhjuxEvxGC3f3rbB/zcZa3C
F8O0O0srxa9HZtH0ix8SvJnad34jNvLIFWKh7PVzkGjaSsUHYilgikw+G8ZMY/LOEDrYDpoCjEab
c95vCWHOKYN0QeFFF0n0N0C/siyxRkFgQ/nq8nRoPEw7WnK8kcWrYX34AqAZpoGQAqrxpjiaA1tW
xQkzreDm5kpk9cSxxJbn28iQ9DBqh8oW326cvA1spN5G7vUnJi1TopPe53x+PpBvJ1dUUXViI+IJ
lCbjz/WrDkiEc6wV3qDYEz2x0oanLP2cvhoMjfO0wdLPV+qLFPWFQh4ZQQa32ikb3pItTRoFlReI
CsvuHgSD6Bqk0DKhY6qfQ+oiqm0wmNn6E0w8r24HZFU03+dHcEmQmy0eIEGUvzBdiWX+RBNhvks0
xbUfKTZAScecR24Yx1tn0Dt+kSqHMgdBwatYV9ZJ/vIrkCaYReg2YIVacW/T/xis70LdIW7Pjr5V
3SiCPl2bfFnGaN8gSpHYJNPHvHDlZPeMSK4ID9Q/1/kmvnxiVJV+QQL0KI5CsySymYcChR9MU3LN
PYGyi87bLrreuMBxD9CRxhHgATINChq0JbS1q2/tfybtS6ji5L1dD0E5hrpQAekbwY0gfYIBSpEY
FOJPEbY+qXPqHOKKcbdwS2Y3RdHOgP33FPmXRnJqP1vTJO/lgB57OaiPGN3OZMdHKcM5oSWMpjFb
BsWp838RE1tcXtL7L12jOrpoe7yP7dUINNerI3E4gql5EtOYuGI9Y3LCltHJk2+kEIloYZU3hmci
kwYg3yF3qS4Gw47KW05C81AyXmv3DqxHAIbgQq8NKTNT4S8KwFBTJcWq9JDjRXL3Jv1ldWEqecxp
NSom9II1gmgNd4at+/XnnM8cEUQAIp1/aBTd5vrZP17h7o9x9CDw6aspJ0k450Ihsi04sLAQUtve
RXH9lXf0tPiz21+kIZsQVKoTyQV23EzQtfgki2gBV7BygvrWpp/pcOCL7IVXPFzg7LwRqpxpPW0J
lUdGi3DbYjujv39Rh6Tw50y0Tdb0oSmuqjsBn1r4OoPtyG3DX3h7Fp+ipl9a3GPpRgEhyQJ3Y2wt
05hjuL6yY06gbWcjHs7VFnI9ippyAyurqTeF6zAVAS5FzES8IXUp/YGcAbe5z3WAzRs23uL+Yyzn
BeS7t913QwHwd2j8HsGlyLalVCu/CRdYTUSCKP4EnCZUl7MFpnn4LLwfyIbETTU+mGublUWvj630
Ad5byH9CctDrGBjOx+qcUWmbQmNldZoYNzM4i0wuYL5z5ftV2yMNXRQjlWtZ42jRher1bHAHYZSl
bKvbIZKPwzKzkyrGTJbomitcw18tTxH6O95YOY86ap2GpDKTtZRVto5lRCxEFWzrEt4v2lAHUDi9
tcozgSrgLmlSiKzRFsD8E1nylEYvJHQcC4+5Yi0mGpXKMLyPTRPFAbZ47uUi2uKZMRwWSquOO9dE
9IQTmV0hc9shQhr5myDz9yzm2M81hO+0DkkwRncIzCXmOh/6NWySXzuupCXF/6uFz8vwGdFbEGQu
F51Zigr6CdOrttuVya/L+vGHGMlufSeFG2nUBMl6Zrhj5N10lczu3yqVxTHyLCtJthXNZ6W7pfhM
uBWQKOvu4ynfP0FYQ66+hOSX+Fv85jnQpcpImoOVI/WK3TwGscpoFP1TmmzGD3NaNJFDXVyQ8p7i
JtEt88x86nt/lpTgICzEz0hgRG8jT5DDz8aNlUbf6EQVIKetk8NEdCUoJipJbG1h2CGi+u6Y7Hjt
GJ7lHdMbcNr1MBXlnzLp79+cXzlaC+vXhw3DTPv0qhqaeXkkvEoa5hfwOjgdlfFCqTuk+DfyAhwU
1CQZPsTOyekOGAfm/FDewCbja+IEP34nScSWnR5bDuCXJAiNP4Qi/uguuResbVrom9fh1NkjwI5P
WROoerp3M0qngIl6HSH8jH6Y1dOmdK925cMEM1luSuhHVG+viyp7tmuwqlIAxdVmNMV6YvoClWdU
FI0SJub1lSI3KAMdwEF8kOoQ3Uyauc4PVTkU9zrxvOQQnDP1a4wSd6RrCxSdzacP2HbIBPeYT80g
MsLRC4Ol5T5txefAD8ksVLR8Qzv5W/NRL5b3lL755QLDGEKOH+uvekdgvIEzE0oRRgIKwzzRookm
pB1Xch47YZ1rDBQ0vY0Mn9u0i/bAHWXEWMFBdEWBuB9Wo5fbPq4YyU8jhv8Yo+p2KU4cztxRTO8H
D92gZgBUgpGQ2IbRU/TGWf+8oytfWUIhakKdf6PiZ2GhEOL4dbHp6weKe4gEpXX4gawU95Im4HQG
3cHXza+EccPeXdV7EOF9C0reCicQRw1E5TCRCK0DRnHCBHXGWxenniT7XkBTeAYaZpMy/24cxM2R
spsgQlpvwRDwOW9YWvvNkaarRK88tSMWniNkr+HBA+5egNBKKWybzaxyjsQASLf103DFl80kAit0
h0LagvdXDfobjDwJ2RUonKGALDfcgPnxB/GDvWyra+E3P1eXzmaIxLVdW4xPuJMHK02JeNdmNGSa
sKR1PDP+efXdfRpzC8oHaLlj/FTkkJSe6gx9LxrBbw3rbdOAC+/4ysE9d8MMK7sE4i73fM9NO0v3
unGvVTzqNlOv7NTsQJkiYPsptkaDTCWJscn2607To6QdMDRr3MGZnyfQeVGMDwG4u6tWd4rp1nDJ
sDSbpxzrq9AXj95kUFyRwmDrDhWQ89ROGAAf+oU9B3W7O6+926XzaHen5d8il66fmO67XczM+tbO
A18fEYc3q8t1AO0CMQI89bWrhrzh5cr58CJWPXMKcWaVpLdZLepLIQMKnK/arpNT7NRZtpO0h9gt
dLEpIqxyijQPTcbCD8aD2c5bJFhXOnEKwct538IFQUWn6nwd/yJTRIZNQmOUdOG7P/3gvYWqfDAE
+nGppM6OYi5bOgCLN6Ys5yPwTV0dfscMMN/pqNdmTAf12mBgzcurB6Q8X2k77+rFi8vsg+rEMpSt
Nud43Sgi6REytdbb7M5ghgrjoUE3zemzlv+Xg5QoLg4g8Di53jk+dBvhP9i6n6+pL/vS9awgo6Xs
fEvZ7z58YA8ZD3RW+NZ6L0vmmKDkFnwg/WEsUxvxQPo+wTZwNIADh7v/mXU5Y5I2+JqiL5dH1/E6
ctDAds1JkS198oT+jKvB0aleeBqv+dunYNEvXXJxWGJQFRi7MZkkuP/GeVuCEz8sqXwSa6J1vwTj
92Tpecx7961/5QebcqP/ndU6AntpzfBX3L5xcLzC3vOzBn1LMk6qhbOt2ZIaeWSy5PDFPuxPosJx
S1Rt+/X2LlU+ISYnppXFkBx0k6GN9rFreLB9F5oUZbzmk3W24PVlGAfgbDSkcGvLskBY516JqdBZ
l6YLuZ9jYrORi5jivrLFTQy37qOiRWPjqL7FqAFAs3BOKEX8vGtA2qrcAoei2pbRPmaUFZno8ZAx
WYtNt50cXWGtPZBHwJnab0M8roTxb4etX4pGdXsJsImAMA1rk3VK32+ZV+mYGhb0xwYJ97txSnJ1
n+3Zp43WdQvjnxyV0DWt+3OewpRxRQPZFQlWvsHkxAGOhsfgRT+a8+5HaSsogcir/z91MEsvVRra
z89Pb6pXDB5yFTCnAQpLDq/HCmx3IRd178ZcUqqiycHc6ScUTEbpb1+stp9Ckq8u1rqGwggkL3D/
hR3n4E5a1dIUHyzzVjUpvGyVGHxaOng7W/+xrryD5aNPEFOIu6/rwGWp892HBAbZamTygTkkThze
FoeVTyKo3cL5byDobYH/Z4HhlL0i1/j7LqWK4yYLVUs4GUPvmFDMf1CknL4F2Y3L6v6yoh54VjZF
VZs/gHwxvcWr78XCjnJhYzPJ63HN/qOXJUDtYrdKHF7Dx7Eo4bAX+0V9GnL0BisCoJ/WP/u2ZxQd
gc+XIlDIKKbk+sgu7zzI+vnvXjT1oGwlht+V2GIpGeUxTvsYFkO4wZaWF+qWlZeH1fGcQeucP029
dwHiXR+s/phGF88aYaMLefUDiPiNv5aN67zwiHb6n2aXlwf6mdS54sNf5S68ydX20bmc9BwJAxsh
rVc+kCE9HDpZelu39XxQSw21afddXQOzBG+ucPm+AoaurfGZ+J92hrS4+Go6MP4IY1ATy2Otc+8R
ouaE0Rl1lg5Llu2/WMGrJqXxLJOcau6ayJCTZck2K4xTtLNzChXgkzAzJNk03POzkbX9xU744/xL
mW5vCsbZRkF3o9CkwKgfi0Sk4jkUmnibbVMB1dOVkhDzMG7jzGRvzK5HOt6AF21N5c0UI5O6en8U
o3fFDf+hSoAHQme39tGd08hBjWUBr+4SNICcnhIqRPPmQDwq1F7e3eNh5keztLw1b3Q6tCRa6TL8
1fDWqda7mEQ554tAILqOud3djwEGDiah8rB1SP9V1c9Ij/L7PRa6Eri01ZhRsv5U/oDrM8WNF26C
CRyerBGEvz7Ed/N8jAwW2cNr3anwM6aJb5Rrr4oaZ9ZIs352DUkvYz67fa+q4QRbaNpxeNvYhXBv
iWfHlLLA3/m54c+kKwpi+0/J+yebmKXcRzaQFR9hVHAlAy/ZvJ3OMtzJImYPLMX7ZhZs2tbnXrev
84EdrwNYAt+hcn8ujeL6yDc3DBfRLaNRonrSHwZSlTiXcfCNOgkK9ht6ZKoHUqbeyQ+9xi71fsM7
BRN41KRuQJqFhfudzEPNhkSJPoG7ZkHXJ5VpJnYZ7ERecBgJsWtyXb/hUJD9bJRH4rnhCtqzf165
ybEEQeLZCS2HsdIHZ5kixdyRLFPORTF/3Vm7FYRMJfNQDjxchqAmkB27y0whDziChSTFh5VXzRYj
yLVNokGQWkMlGsQVsSDQA+LZioTcMojUMnsuPGBc5gdbWdRVS5yYrQ0tFWMyL/16FRgHB0btTN5+
g6cpglETCN0wHKplBZ3x3OknlbmqCCWecVeKnHBw0/uKzHTUJYqWZnlsKt0pGfa2FznOGGZiPnU4
zKTgUgmtKPX1FxhdTYjxfyrno2IDq+IPDpU1D81s0B0ZE7wfgVXwIH4qxMP8d3MPekUa7NvNu3gP
KlZLA2p1XNEEymZT5KW30PKbGkecXgA86WjmZRPROLUTAoBTQEPsZMuXSa5qJqmKeqGrZgib/tdQ
0dEy6Fq2QEPH2HnQj9GsuIegNNUIFyVXkr28BBYKceXuQlFfdMJB7IeiACQ+5bb1tp2D/wYpP9pM
imxcGByqE/r98nAkmAUMEMhPlVJLzjQsLkCMoVMu2FxcrhBdM2vqjPhAfCEPpA9HFFxH1kkcdOuZ
BAr+RK/bPd8r/aRpnxWYbWpqn2E1jgyao8slwLgxanan5priWvt3R+69jOY18H0PCaxLI+lOCnhN
3NQUeLmsp7msIqlWimglvtr8YTplsAjc+//+qOEgLb5Cefs9SZOlsF2qTSiH9veT63v4JA45Rxbo
qDL32tqzy77NNmzaLXhKzHpYG3+rvCiOMyhHIPHcgvBFJ2yG2FBAdL1b4J39AP0O81+lqsMEaGU0
agxWz199+6MgtctbEvCbHd2m4PmhpA/GIk3zCbI68/6FvtM6lBZ+OVdc8lVVZwAR+gXGgsLQmxbi
Q6G0KYbS/aCJ+nBJDmuEfWsYYZ3PcL/RyE1WPPIrWMKfh4ZljhyBRg7sCpBifbskyt/YvYL8Rt+X
ayBxNHvBp8qJdinQ+ej9PtaQjTw2d2vOQhJ23fnR+b71QvXCtpMDULKrqkGNT699E1JjNL7zm3+A
WnwXYNyvE4VKoYk2psPKGCfkhxc0oSqqEW8tQ4d3JFvbmNs7aMhxAbD4LkwS4KhyPnf+kEchnFPl
JOd10UaKgv3gNDOlBNMvM/0GszvWbd2U3XZxEuv1v+hNps0XUCV89nZQxsgWShVgt5vH8aDbZKol
VMUMidTRtNxWev7V6VKDj7cZcEHA9Mmosa/uX6LVaaK4Hl2020lBYMkty6krt+E1BHqDKCKKou+D
hb7mBFm/KdSTSYWB9GENkbtK+mvoe+BhDB4Xnl+ooxXvaxvjwW3TtS/JU0560vxB1dRmSLBlvKhk
e9gcHYispy/rBbFOy3fNFZUcRLDte35qsbUR45ewgXU0EaXtp8Sw01AXiyiaexxdkz07qvq0dtAW
MYCgYOmtjQyRO8xEkWHfABonxwWGBjhvG2VdSjF1042DyVJjeTcPode7tU0QmwZPn3H/dTR9Z7Io
yBlhKoI/7f1sCm6QvccPeP6FewRC6WFWJxSbcIEcqmiUlM/qvgPPaMHLwFESDNWrWN5Jv9ekPEW6
Xk2JpzOkhncqBiY9yq8xn8DL9Sq/qEEGurawPosB3pLIthnw/L5xS/GG99BsK051QMW26Ivy24md
K/Kx3+IVrpeSooXhPrIzy7ZZ/GKrEccs2rYSWEI9f/DbzXYg9L/+e9TyDTpIAlyrn6xgLeHO8VUi
UU6qjQJJz78dHDUjyaAnTu+AanWKcKifSToMxS4Mug53wBWDydefH/T2xpNDZajs6mogDZn1wvch
T2ZGvCnGN6zrKCTiaw5JPtjUaxsbycoS3p7GXqBLpqAWRgX8bzvZ2QFuKXf9loBURi31L3aR4nZL
ZMoyG4RjWz8nUDjmWFdrXMiRTG9g+H/ZR1NK5tVCfOddAgKnTufqXGQLp0MpprlUTqrxPxuljpt9
D2LBEhzz7CF+kQ/5XOW/hWxoA4g13+w/DtNllDrlQ4Be0Jbluzu6zX3ywxFmGSb3SBK+uIfwvxr6
Vg3PdeEAQ052n1xCwXp4se8EnHpWtIf/VOpr5/DQ2cnJRYMRA+k5mEnm2HlAYD9a+lBIupWMo7Hh
Ku8ZE4KivRC+IrXoUJGnCCOKmhfMgep3+V/ZVLSW0dyvVLx3rSsQw32sqeAqMz9SuugNtxIo0qAL
zLTqlVd0MUczk4ZD3eixLX+U4A+vSK7g8U2661Y0c0SObCrFZe5wGBOnCY1vjDUA7CZhyWC+ZmAq
KDXc4RFLKAf/5wymjE9/oIiQWPShqoc/hbm0vyrON65k7xoRbrSzFA6KdBj3FhpeCHFxbDzQndBq
PuXLinSiL3C4lQfeeWollUiXJMnjEddaregIAMhKDx1fiUVPExPHf8+6H6e4ByhgYMgYPFliHlDl
chUGVeeLrJdlKohl/0D0IFGHPPLlKppmOkHA1KpuVjTpWEk3cMyAKNwvQA4Li3hDE9yeniVr+RpH
sdXXvAc6XzjJRGQhlt+9kaBy2Zoqm8tMuuNtUdR5UNNsaKX3GwVxR+9RkLB+7U02gDZsp6OfFtYK
T+RMGjBLn5AAFdAOgEQ/mq7XcvQmNH/ksiQG4iR6nWwidwFbC85WLr/WpTQBQKHqOD3dxpMpCA1L
LMMvAm11kuAfjMFopiIK9fs5XRevE3ZqBMVPGT4PYXGuvggTUfaangMC3JIks7y6dV8E5CdBBUEa
pG9J1PihlZRH1d0mPRLksR7Yks98+klpDNnaqrXsbPDGeh6PBQPzUEyfFcuHCfU7vS0om/IqVSsK
OnM368ww3So821kWX5Zng6EulwCm1YB0I+C5DOMG+MhA2g76nIlBCYdD+qnMRe8v7rovYmUaU3Gz
LHAv5XLU3xKmO/5x1p9r0ZmCu37x7t5xNKs54vMXzHX5zZXyzb0jHcPkf/hkc6LTVJGp6Vvm4PKi
kuJd2dENHXbQfkmdHtPYEjfhJQYwgQZGtAE5keGrLXigkAlSbnpPkoCIGnQWQk8dnC5CIJ/sw8UI
FGDPAP2qojgGjdQ23TbZv3ejRmaBbD7PBnKhQ9wuHWyzWvphp0o5GOxJ0i3RRhi0oQ+WCjem9MHC
o76/IBAimbNEirHuMkkSXLGHB4s6G82D21sCOiDf30DAxeHyakboYhYFbsaKoDIX8yfzfPiu+tOV
GmGvYC8J3kK6TWaZHYNcpCqt0a6HjkbvPcwO99NfXuW1TCmyOQ1HqGFww9aCUd0r6DoZfoF7ikd2
ty+p0AD2FQCiTKtUorx44fAuc2yw2+/2Ltdx+45I+577Gil4dQg3SF+eFVlQtEIISvPGnuXdwtfh
tUh5FlWnvX7dBDb07GWgYEQPJWUB2KNKGSiPwQwzhEX/u3zs2tOYp+PzeKWavzZjblQBZ6jSDYCO
vVbXO0h2DZgf2Qhu4ASFLMQDLvQJlaYbXR8sMD3WV0Q0enghpLinzk90UOqg9KOvxSmFxYNRccHf
410xiUqdE9bt7LqNpOi3+sVOdWILn4A0ugHuHo5TZnCZhShwq0Cpcn7uxlp31O3obv5sQpgofGyt
VmeF7TOmYlOb7GpOyI4B5bVXoZFdhKR6kR/iK+OuIVEzDMbueU/fPR1TAmwA1KZuYVcQRbjHOYXJ
UxH6qp9PZxSMkHfK5jjqrOz/D3P4Wf8+Z8j+69yexlVUIzND5ciUOvVqZ/MDt+WwGAPQVedti094
7eBRwT62lkcDgZnyQ+xT4FjLD3gZLXDMIM9iwS5e3YIZqmlCl/nw/mAMS4wMCTPHHjrUeDCNRiDL
0iI/NRfESKRgN6xDbfWjopr7sBMSHqw7sf1tDnp1QkZ3sb29i1r9N0Zk7Lb7ldBShWeMS/XqguNU
8hschERTjRJCsnzU3tHjQiUuNS3a/ddyNEZu10bqKlual6+6zEu6RcFzxXq2YmJoy7VQ5PuW1t3B
A3iS8pK24F906cJUstP481jDKa4/pJLgzQ4nNILfuD0vMWT6QAHpqmRbhWx3PgtMld6hfar18jGL
22x2tO4+0vYej1RnUFlrdbZn9g/Gm8q/QwC8gxkHmtjKCAEnN4bwyHCzrPiV3wmoSwN6XXDNc/0p
dmj/QS9kZPu4D1NWHCaph752zxg5lKBRM49xtNnizwxK/cIwElmW1vi7Y5SSbC/D/XNFduoZRQ3q
vg4lVK3wtWQ6T/SS/Y10DI5ObYN1xBDVTssBcNFlT8Jo+t5xhMEcoJFoj754CKv7AS4wNblPfcHT
Qj5yELa2zrfRXDNAlug5aQvL3eDHXftLCUYFPgFit5Wr/4ZMzjW5WxzPo0t7xvEYaCV5pNX2esry
AVOnBkHcQByQi2+txWx0+V+/BMcEBuVp9ohvPA8FVtuZjeOeimpfBCUyXKZc0393/jX8yZ8pAGVb
iXPcjZ2HyHSZyUMOUGquWWHTLMtmMMghdSYkGPaQOg668Z1wBr0wQ/G1WuGmQzDaXU+YEDHBMgjG
MooZpFMSLVjhrM5yy8dWDmE/CEGt9O6Iqu0OpgW/CtBLNo1F3YbStk6O+ZUyhd4TEe8nPlfKuVQ3
UVC1y+sWPBD3XniqW+bJgToApGK2FIN0ZUNIil0KqgpChUVSIu+PTwZClETfkUZYA2yLDgjL53CF
XPQmzSM5YWqeUFCgLjVsqzBHaHorOHhE8P0ki0ditXILfI26Pyt0PP8po+dg12xta2ne2+it8RwV
Jcm7bAofQfwSA5X0Y6IFLQoH3Ab09K6T2xRI529cU00I/FyXzIMckb3tNf1RBNj6IWwES8ShOAzL
/TyjX8lJ3OE1MrMq0AQyKHNOWGU++g6LnYWreQ8hOwtf9RqBJmhieqyRyGfMCB/5561gCos7RrPX
+u0W2Hzjqnj8Fjrqg2yQDCHGA7cY3nlwLeLNJ05TIRIm6vhD61co4+zU5TzdMJvTODxdBTzjWwDQ
r1Z62MLZ4BEmjjETFQfZOq33bP6xQQSlKyfGT1tuq164svrE3hA0ZTlCeK9oYcEFxD4aJS1mnirf
rP/Xo1Tnq56btVbJZTaBVIImllHSER/2fofAxTSaB/qfeA/E3z4VpqL1C4O1Mb/Woo7AiV/FZzNL
cFlsOvJYoadZoVbOBmVljj7bEKaVKhiqhHo9/Ys7c3n8RY9K8P6b1cXPqEBhcgRXmip+I3UJ/JOu
TSGBgqH7xwaR8gSPRqDkto6MUCh81PonZQcQ3BYeolwgyUwrDComcQD/DQDOiINbbwxODXxQrYXb
YcC/P3+aeFX9DT31eNzJ+dC1bZSVC3yIHNwxZT3C8GCw67c6kem04QJGWUGOPbbVBxlKzfa3L50i
f9MW9hyHYJzlsH+e/AUM/6Buo2B7E97nSg1Yjom/+hv21thjg076LNXeicXvff057o4MUi8X6xzN
aYBBLKWXCsb/FxoRF5SuzU2GZC8w8tWzhshgtsnS6coWv/229tScZHXJurAA8Oo5Q/00L7pdOJq9
xqeJD3ku+cxGB/246TY82kffJayreTFe4qpgcJiOV2RkW/dh9iRgWpm7GiROV5ww/r7io3wWmWsL
UYq3+dExqA3mT/KAbgCyc3HACEJ3vTJ9ynhM8+9woZmvMiHjUuYF2K14dVY86OGUmsQ2Ydh6hRTb
a/LvgpkvMXDQ3WH9KUQzu0MLBuTDjSRUEEXIKSPr/HmMhOi6nl4kszeU1gCr5O9TokbD90FEop+9
sswSFOFIu/r7Dpq8xXqsuvl3rmz4fqqjRHdx/Dm3bawOlUKLMnKX/T6aN2TIA8maXNGdE+k2d8xk
4x38h1jRIXi0ABaxWD3iAkj2lXi8LeQVgJL1/HOpqQx2FEA68lZmAjKHrJJ4dYg2hx3UCRw2dUx3
QPAdtXSGLRgFUA+Lv28zCB3uHgoFqpWHUjloYRq7vVI9DvtVldRTbv1AmkOygSX0RYNwsUEAXpDt
3GEM30pkOdw20bFSPUZnppFqbWxHfMP3MmigUnHRDBvq5wELrQ6leaHQbKaFgR7dvC2Z6WNpqK+W
AB3/n9m+nt0zqsAhPPkBS1BSmG4K//g9/N2dzODFe3bqDo3aKnM7lGMag8JsWLW8AiVzH4879qNm
iOVXCuQBpjFyclLVtCeunRCoHWJ00UPJHiS4Uel+qG7vRDV2uZsbnRZe1ZcgVMNW3cJ6EHLLY0E3
ZAoC6WKUVhEqtH9zydabujpOTywgY5PqJ3BWUnkcXnxLn4ZQGfNuXfw8h8JNDcQPAMiccgnBtteF
hRjFhQy4Hj0XXDEhGrkKbt25Dl80UnunWN7bhuvWTzjgHJ0x/UNzswc9Qb41fRq7LNehGAWTiV2b
477fvjWxYFVBuHznGZ+S+SgVwsNP/RaZpj0VRiHto7Uz5s4VFfc4OUQv+TnI/OI7Dgc7VVyk8nLC
bL2W2RCMqdum1e1W2UHVBb17QxWd4lIX3pTM0ZoQqVBX1wVG6HzhYf6C1+404r6QoDCoRXvuWDXD
NNG1fx1iGg5Le9VOMB69PhlE18mMQL06knFksn5qvXWGk9D77Y3BPI6c/dIdBH6pE+IriJD5N7dK
hJfn6qo0bTdTSxkTXTaL3FkZZ58XdgZdxm2sCet2InCSMJPgKJZ4nx3PKaKAeQWRxcwpBr5lhkVf
M6uoiYcMP0xHTxqRsVAWJWtdL2BwygPBLsxYkmCWXkT+bdbBDKmz9xLH/+KoxdrVyD7p48gfinI8
z1S0V/4tcL3B8w9mW/SIG4Z8UwRbGnmfF2EGfQ3M35D8Hi/41M4hYtB1QqZX0KXGA/gRhgTRYsIs
gwhd8tjEq41cloWPaZNsr+g9MgQA7SJQbzbnhrstAkcZFzY2REXN5fkfxkZuc1ei8R9Rxo5gLnN5
rO5BZ34Dh2xWqQAxUrWkOpYzlp5A3eLlhsuYNMo2HcQVo1JFEW55KBtCQj4nraXjKBjYo8kNKm9s
t+6MCoNsNB0kyj3zeI3w+LXRqVbGJSpd9TsWLdEzrjYBLBrpri8F2ybANnkijgFDnOJhFRyjrdHy
V+9bZS98XLyFMP1Tr7FW/anxOfLXEZYoKmWI0w0vjX882bYQ1D708ce1lANbkiX2BY5RiZWHaLxW
uFSMney8ZZqlxZut9323VsfTi36wpIS2W3gdTLOT14uHZ+mv1uAhvuL4OB+V1G074tm5kYxSBkYi
WP1U4DBco9gj/ZNX0ZHG4+G3wc/3T7bouX3C54r8enGmCvlcdguh1MNU/eCO5EofK456YK3ouIUt
OZT/N8Zfk7UmQtq8lAFbIAig+QUd94AsRKZWIfvqN3omtvuWU8Ckh0QCPACwkGHtSUEdm4XnXEYB
dZdKsQiRJ2DjCFZObkk8DDtm7gjt+g2Ad/tWJGacpDnTqR2WnJp07MwOlUz9F705UPKs8ClZ5IRL
7UZlWYnvXFHqgj76SMleJyaZqFCYG/XMknOX+T+uD6g2JbF6md/jJUwFco+GMCmhhG8VSzcLygL8
xVFLaggzfF2gR8WHYGPPzDsGa1ti8DrG7g+YKGQ47LopiLtBBoD8F8RqUc096l3xjEeLuPbrrBSt
46uomvArDPhB7Xaz/g268OKTV/vpOOtmFBZ6Uj0Vbor9AK2bM8P+3HNJxVQDjJfl7EyxpsshjZBX
pdNX2fa9kt31GX/GE6zhKkZHMtGD68WddOrcCWKgXQEnQnJxAfhEbMROjqA4P0/BwC628mT4b6+T
V0XQaUHdBIuGHxt0xS8drPXq5Jx7oXfEL91vBWR4E62vo+COA6YuQJaE8H7QUUFzhQC9K+5FurqJ
70USRsg/gtoSNrYY36/iyrBWhLOYFog33jCQp7ALe0B5V3uw7gGntO0SPIB6m5tLRfLL4Wo4+A4G
XAmlVR2XmUAY+n90Cp148cYpo5lRHI0pI37fYXciKGQhxXkCte5u9mOkQtpxnMJHpnfPgdBGLFiE
LlR2BPAhkGa/hGGZBOCTh5mp6OJZbZL6TEhg1CPTMzzH24elGJMw2cav4ECDTg42q/a0ebrFfo34
UuUy18SzFD0zG0zir0P8BwIRofPI0td03w7vaOSyVjN4o/8/rMsL1JMvDcFwIdmb5+iB65XkzRDq
RtR5/Ckay/gQ3JS3FirmCJcui6wVGs9mEdJSeNzNYcZbegr58kStqDeIXpZpMA2Bu1jGwA4X8PLK
qh4EbZvXa2lRjWEA4khtohJf4NnhftA4jt2Jac4bqzEDcfuDB/6h29u4/ReDrV8zKoBTKCsq3749
CaKyB7VawTBBrEPYfBilS40j2P4FcrRVclXnQR1XMlW8NR+He7iU4DnKsx3Ecz1vcVugKIbV1J2q
S8BOhoWiFM5WZkRUkMOFC/Ybx/fzb66cOpkBnCeHE5WbEDDidcISiZ5MEZ66B4msmP4G6MLf0ajb
ymjtIRi/6/BRIijojv6nei2TzkRhm7adBC5CpJ+Qjn2ghdk1NGxAt6GcDkl/CDO8hS8EYwP73dbh
gvMDMkDRO47kFi6m3V5noLkojBDevYAPpa/CoZibctL18ffTUYUbEay+3FAAMHRes4wFGHR7Z0Lr
i1siI61V+Z64aaOzMZ044d5f9L6iOnMKCZ7iXBhh5246q+VzQCDMZsoGrwntPPxHhjIhtsPtCyV7
ABXxOIBCfkwi18b47W+tLxHnonK7fj9BV+HPh5bM9+ZQ62o1A5HevkTg2+qNY7cqSfbIwht57dC2
Se6IL7Xmx71SzEYewbOi7rLgyanfLi3LEO+nUtVm0elTTv+b/B20g8jCGTuu1rtL3q+4yy1OPUPi
4DgwgWwAK5AgikYenm/boEv0N2w753jFLJQjHBHLe4mRxyMH/awCARnXfuwj9tZuMvUnmx9YON/X
KNU4tDA+r/6/cnShHy5p8gl/JFUez17k05Tt2jVWhCvTUsJ+Z3kurWs1gp7ptUeDHNJnL0/6PUXG
hu8rmG1iNGdJ+7/z7lDuNafmasG5lH0pfkNVe2N1r/IlLGNIR9E+DvIl8aNkHTrLxwpvgA+hweAV
J4oc/+Rcxgwq5fVTPL0iP59GDbBUqTSw94FyBvnI7tY4oL0BRdAUhDB5Ar5DnjkcHjAn6xkOReAk
4GUShxBNRfsX11ebBOisz35qSZ47H0dfqAkYlo4VwIvORBw9t/GTVzSYYq+F6VbdAv8A8Gqpyyzp
gd6rSFHbhadsfDZHRaUnlIxjSdm6/bn1qrFXmux9fderiuv2DetrRseuNKFQR665h92x4eVgK/lF
h3EH9Nn0UWlFVLCDnsARenC2nl2qs6kGHmWPhs52DTuucpwGBKiBVcw8LFQkGw4foFNuUBqytmP5
j66PQQs4aU1ag0DWpH7S/nlBLhaCPKsxQQ4jCYZSaKUyGEh+f3Fb7l9fJseH9jvcJrxCpgR2zBvO
v0dwU1jTbZSJY/4h1TGeicZMTtsi/0NkegjaTfsFpQyf/XQp/6LmiYrLMgTwdPG1XyZ49MhRQRBI
LMmfcw/0PZ8lTDZpCd/z97JgwAT3zXfRrIjAiNxExufe+Phbg7W5unP4kE1O/OnfBqns6dQmneb6
e8965zw75eJpebysE+QMaNruHGE3HrhDZwBCCm9ztUFn2qxLubkGTdPf5tqtGa3uwlfAQiaXOmvv
aKixVDN2fe0SlGgwe46V3rv/xw6mbt9JrP1SZZzVNHHrQY7MO3TBOY9qV/7j7W21VWnJttLEGnTe
1UqWdy/SCeOHUoljxuJndFq2MYUDozJzziNq6C5+1h6CGLB1EXdvlRXpJW+YrSytUxQTDZSOgh8K
Yjkxu5REpE3w0XqF3Co+iMg975+1/l08toz/Gz27ZV1dnysTwFxoyAsWv+sgrxbFBh9eCX9Iut9h
LeLsjQOLvJoQLfSZ0pyPuiJmgk34Ny0yKwHdz7gh2/5rzuTt5AsA+iB2pner9VSdNlnjfzxxrz65
InelJEokMUlB3zS0/R0heeKDdGTeSUGeI57DU3k4qrHXMAbqsA9M0qqZsE8jHKjXe+/+QqOEChgB
dvlepTvSy1bZDw50Oq4bYw/fmUofXvTXIy3c2uS0AxBS3a/G+DFL+QXT+9envjJua9wGCEyKdQHR
qF49IoO2bYXsTee8ZdM1JC/N/IUc0xEf2kdJB61U2mhHJb8zpSORe4ooeU5Gp5Dnr6BADR+SZGm9
vlXdhUiSK79Keqym8E5xNK5j7i3YAXaD1wNaAjWTUhtGblfQaE/F1b3bzW2AnxQwCPo2kC+GSOtc
VgIAOqmW74/dpPtIK6e2SVD8S+KBMUdKWcgPScMWcyB8fLwD3AuIz6E4AbBxrgw7SPFND95XL6Ky
2nL6CD+RB1Luze48wvvZ7WWqY4+5KNnoFUew1xGq6IT5eSPUSzDX18sYV48zUllgHlOfOQT89u7c
dL27X1CCiVbcfbYM/+Ll7VU6CWrPB1/7e5TD6GrnCsa2DcWA1YQFtnjYYphT4r/WGHGPqJnyN8V2
J+4lVTCmESXrevQyHjIPeudt3ubbVjffVay/C/VAiOc7mr64Byu8ia5U8QL9UsPgYLqNy1mfTesH
pA2hwXLyjbozKtzPXp0JdRLT6p/pzJ3OB0z7i9iMUm/SCa2GobyfXavldpCR+Uq4vbOhYMgA/uZT
oh9QtnNZdeGQpJBfXlzO0rNCuTarxvvCQWx4a8Si+pjAcmRx6pn54QViwEInG63Scnn8O5MgPOYC
805r66lNDNQFpqgTHOtofdVsBYsZCKfVMh93HfP04da0kVC3qq1zTqEX+0/frDSEg6dEMWIrWfdS
uYqCywP+QR6YPPBImCz7D+zQQsVH3mXcRS+yXEV4GoVS7h3j2PfqywaiwKPD5O1SnMufWECNgyLq
WU8QfWOsd4KaPwvqhTeFy3td6E/bB0DWC6pKLOicyRiMTxdoygNwL1Amu0054ZwyqSjo5OWFq4iX
Ts7jT1EexTY+Dx1xNXgUBWxxjFrsa7zqrRRlSI2aNiLDw9IdFoS/vhHOCnhfD69TmEndZm0h0DTC
5im4LitqSwn/s6XIou7LCAw2PwnBbglnPGrNbciwyrA/xordkx5L1PdqDrR8lQBwOaKQzD6UBD0+
Ey5KWoF5rnx5jwwFs7OF/gHP56zp5fSlfoDVGYtqAMA3oOI+yxJkp1ULqpsYtQKwx8FMMK95gwtf
VsncobI9sdvk/x9i+ytdxYIa8nG1kNlaVM8y6ykPpiUIPIleVJ07f1nNMv902pBQSI4T+2m4s0BJ
vIZWFvxHBxsPKj66AHF+gT0NsNqGccr1BPsfsHwAa4KvrllE7F2mGY/l1zoN+3cc6ha13JkuIoNe
o1rYpCytdisYjYhSKMlz3fQ28QerkH3cYY7h3NkG07rW4qKFEduFHl5PJiCQQQgUxu/DK58YBh85
EHJDGWCPUv5xquqHBSpt/ks0NZP5HZ2lvfA+yf3zxRREdrxvELHYZGSK0bpZURlGcqixwzry6YnD
3VxS8sJ64S3CX7mPai1qZvN0lkKFxKcR13YuLZ4se/ytxUg0UpECrhjrD4lqNMqv4sGWHdaDRnIi
cA9Vmpz+ahwG9znXCuACdHhUMgJ4kdJs8Vj+BvtIS6QHO+hmDsqfO3ld+p5rlF/adxdmP7Lyc493
c8XhZyRggxIPyzkWqi0rCRvQPdeCBUFcExfPPhoXjR0a4wsAr2DUl+nR3vczI0JXNgC5z6TqnXdD
hL6PPs+OwDCvfrE1OJD0EYa4pvho2JfLmvGbEas+7iyKEdj6pN0iTcDuft2dy482JWFntI6tV1hZ
KBNrf5F0w7rmbPWMSu9lVTnRlXkSdnFf6mf+iEl3ly4JDp4NyUSxgjoIEqPfPa4ROgGG8K7iLG5J
ysEirfjqSAUJBArG5BTYzUknzUxUskd2oJ0xWMl59RaW8QnJBE2Nl1qGw4yTtijuu3Qi91xnRsKy
NFj0AraiSUxu9zH8icnOuVYFL3Esw7G5dznz0kaoSI+ghMDusrNtcqW0kq1auCuqMXnxhwpUbcVZ
Qbh+n57FodDrsv1tGQ7bnT96yjHGyR/KgaC+I3m8xPOqKDm4U1hMvfECSr9Qa8Vj+/mKZDTpVSyD
MP3Fx+fioP+lNx98aWAUpJrKNmqXkNZAG1aruCcFPZW3tzMcenUHUM0LJ+WZIuC6DGhj283UVeKI
Az+t92FsDLtdnEvYpJRn/yo+hPya1jLLJze4sUg0hJagJdQ351HFgOW8P++P+vFuYugBZD0YTr3L
VJAPm9lwMD0yVtgZaJpcfIwuJ7h4SP2WU+YTg3tKDwitxvn+RuS5WI3VBbaWlcbdK4BrWRngjzb+
QqcEc3iU7UmOruKeGgKCW9Z383co7IqlAOLiFFJ13iYkr3KHdrVcCApccxYPsvf28rDdbyHhqV0f
i0C69cZbZ4vxyabh5bR9fRNW+OHycw7+xk7bRtP6h5Qs6eqCRhCeavLTIMP/xH5wSRqzEyXxRw7S
uQLqaZUkcVKdXeQE2/ClonDIdq4Om36Q3qhbrw+LMy9llhhfAVM1yf5+xyB0fNXiKqjNLXJvusAU
F3CYrHIM1+xm5kxeNkyLoXnY3oRrApuK06UiXhkipRsu/yZMf7lCMAXUinIur1vf8cb3+1HJj2ZL
lsW+fwLUGe4fp/q40+eHNcbQEMniB6HQxMz/89kQ6fU3IR6D3IH0WV/BdCQfQsR0Xp962Odeft/j
ocj8BUHpW69+Q73QMucoEL1TMjWPhmbK+qmjhNOsz9Zieag/yc8PO8Mhu+DlzHpTd2eyQ6hGDOQL
wS26sWyxJNMFzd8wqzLR9mTdjPvBPIFGxV/P/Tczarm43FBrqIk8NwKptTuZmz6VwXAi9/WRmWEQ
BmHZFdYLb3V2CcBFFJZK7QHQQlBcmtKyowFeCvOYSI9K9BmSQMGzGc8cZfiCNnUCVUgStOSn9eWW
KBpWErIHD7CztsHiN3fFOWmnDcbCs1P2XTtgcDdQcNeG1okBQUcgHQOFZM0txkKg02IOvYrK69Ie
Gf/ZMVIOMMdNpp9BeRKxN7WqKNaGnzpw0uiQPnRZH/m9n8vSoGomGyLPuULqVUhFer+H1lqtaGXx
hjOOJl2qYZVsENb/84ztMZEmnm6J8fBY4nQakaH5til5yDHfGytUVPwBQXimyzWvIOkYP9L7lNqG
7wjxhTsZzr4sSNt5Qxb3iBjPAwjt721jJHVMV+7YIFWSdvWLlLKWx8bhh+Ygt6ZxZLC/sJ+bY8G1
KcIagqxRNMoDhcpeVyI7323vClWB/bymIzGmntCrK6thhBcqMy62Ut5MQI6+uujteJtvCCxQ42wz
fV0PFGuwmeFxQzSLGzENR+1mT8Vzl9K1dmqbpMOMBLm2WZ3ssj2UbKkqgPXEDavgSsyavf9YDZD5
NJfDxi+GFJUO4t+JWoXJ6xIFh8KebO8nf021e9SjdoSD8iKaKeUmbjDcjCatExEYdfMPiiSnxz5B
CpAwT3qnKPHTMpKrVKAa/dglz6kMOyLUydnLybG2FOxw0NMrX3qB2couMf01jItWAf5jNeemZ8oD
dTV2xdYnnLA0EYR0j+7y784MrLR5SyvHnD4ihbJirSPxMgOhpfKVXN7XCStTytHcyRTNQbfb/oYZ
u4NKwJHBT6JIg3+QoG4CSTrh8TGHV/t6rt3WVUSAbHv+QfL8eUj6teuA/MwDof7TXUoGAjVzEp9W
2TdVT51XL1Kj0Ne1AKpoUhFDcKmKlD1ViqE3fnMF/myEjGKWbYIMY8iZhJrrtnl2FEkogDx4TE35
KtvvK4IbmqgQq43+SvRz+y+e9iNBBWHUR1BwrCUw4hxJUUg+TW7Rbzvyh3H9Cj2WAdai0twESs7L
2YIlSkBuQjfWk51Ju0bRxYnNGf7t4rTsGeaYHozVTYCxzxdTPs953aCskZ3EW0QqCtWTJtkZJ8Yq
KHsBEJvPNqySIKULOG5TbVffVqbjNbcGWrZm4LNitMaYHXTVY0S5nxey6TytQhCu8YdgtL2N2wps
4SvROwSCj/E6c7t+moBQ/VmObGXx82vAz5EQCzaTdxfAqYg+VmCiczOZT4wWg9L6L8ctG963RP6C
/CWaX1Mvtg9ECyLi1bte9c+z6NXcqY1IUnyXUGXJ2r253reTUTU3pBpTlXhIBNbpQfvPy3LNj124
6oEXi3eZSoQHgbhHbxllJi8JwqT5EEjWJu/1nQa3ink1+BhdKunN9ZoSBT9CtzZLoG8+NeAaHUwm
/v0Mc/F8XtK3J/ToL9fgLrMqFnSKswizw1eNGcuMyvKH3uSpK6duH7R0GXM91oJ2eK9dYD1lvwXG
AOEoqSUea+m8sqT78U/3J8zeAJWTK6GOqzEDk5hz/yblt6tipTnH/UHoyOgeyzdjVzbxRKzN98gc
mvcvQc4WDFnsGdKUOVOWCL+FzxZOj4M2Om7ztKOlR9ZHD+X93st+h5O9nlOfP88U0c8Rbl98+yLW
OpgAiSuNBtLRJkX4kRzqJaObEiwnHj1mTrBhMvs2GdFL1tbE7z2jHFpqXN5zQ2zx47CAdejECJvQ
EzzepEHpn4h4ZTtOOZsO1Ea5nOEK7QXDsQrcRSm1xi2rRgj/53DcjvTQ9nnaGW5nqRddZx4Q1aiS
WFxU3vaiFmaRNolzMTVQCTGQUgo8qGJmwMbUP8D2Jj/+ORyJEltrlhV4tExDyJGT9G/9DgJpJm3M
zZDfoMC4lHJulYhl4o0X6v7leN23UaTRyi6A8oQqRppiCxPb1PmLwHCoSEdFBTadG7pFwTjkOgp8
qyARs/+8GXnXRK2+zP/XVMRxUtfKiIxnUOR7dbB/ii5Jx8KZ+pgMDdpZeQ0LzaF1n9C4/QIZNb53
z9rzt/nI/lJHhyjFyCpuRni4z8W5heqSjKsUyEGqrTi1sjojF6IQkUe8TslxgqcC449DTEzHtDHi
naHsu7fkJkeXTvgRiG1f1OM2qwBz85/6gZs1ui88dtRf8KeT3+u68Tkhn7dp6HrPa2dfHQgdduDB
1D+N4z7iuQib5lanWHSsniV/nRx7PnlK+3+Lyr5nQ1oIuX3a61ZXs2OG93vvJ18bx3zr5aNGN3Vb
hdnI+qNywotLGtaxHsa234KPcMzAJtB84EqmypQiUeVcI+68yLXM1fa0h6iVP/qPgfi7I8NQuKTP
6jcDx0bFHdmqc0szLT2FAkPKXrUoXzG6FKGdDGa6aifoflK297DSOt+rycIJusJnPEuHdS5IUlbJ
U1S9rhY1trxqF5Zyds7i6mTO5jMf1oOtlMe+qO2ID0bcfR+6oXT4IeH2df7Fm64GIFSkCNIKx/Dn
bD46SPzE2kUl1kwU/VJI8MH8BOpPLn0Ftbluw9C8sZ4NbfnR73ucj0laSppcEKtJYD3aJqTDma6S
buzFugIN15Z3+iCgO6dmMkO55497wTv6DEkJwu+l5e3ubQWaC1b4Iiz2fM87VkPxv+pwwrLw0+od
Mjd68CfGpdsz2/Tx/h4GkQDjaGaxqDY0TrfQxSkrsFOYL3961dltunLkZ6HLVkDIsZ80BiGhfs/A
0f8M3onKHpNgYW9g/JShJk6CnsQFCCbxNYaJxhkk/8yAlmUddugxplm4zPCCsJo2Nu1tWNQfxc03
UDYzKzs8fKuTfSRcJnEKiHO/vbcDyIQLqZDS2mzXJa+DVcRtCM6iaZPXDtr4WsMFX3Z6x4M8cEAW
2SFdyU6LJCJb6T11tHNub+ts34DKZ3oO/SQQ+0O+BUMZOJOilEBgCFhsGQ9ChT81PcLkPjTmgVRs
OWu2MY1lApENFEVFwhq7susVvaTk/mrvJOkrR7DtfNB0Wee+hoM60mfLR6JZ2xbLpwl0J5D/+IRU
89uRxn6o9GcMSG9QWYKg7Wa+uOFqhXAOoO/mmrTvK9rGUdSTolm2zfqv7oz5evKuEafihz2+CMth
WlqqGDfI67tJauhkLg8yapLGtG9fbaojt/PS7FZw694OeLWmjaExgcb52zoS1g2b6XbRBrhchwb3
yCVZXkQ0eleTTzw2lNGNYIDV5jY87ytJEygjpGN9u3lczAkzVM+kfZ6NGCMdIofWQsE6n9DTrI0a
L59Wy0DKEoyIT6Hr/WCP+nbX7QTViEwlF8aZTKnkndle0+c1Bf8QU5PE3jueYYtyzBGiI+dutNih
/+3o4fn4zSgS/kU2+Kzs0++LMUgnVS8UZIyUchyTi2wjT+iYFkNPpl3RqLkDILL9tb2LgC4EzgbF
Y3G+9lgLrZZ+Vh3581veTbnCMbxBxh6In32YkN7Aq+NjBgCrpWgAtRS0Ig9mRM8vSU/R3MoIHekF
Mgf9nPIQ/E0NLAnyozCzi4dPK3duGkPpHNqa46+Ubg0OOMVWvMNe2AMAOe3fzbsdSoUO/ZOIPT+o
9nwoHrHwJqkFw03oXhAVWvC7AuyJaxkoWdpe0x3Wfx32r6sVTG+ppqylNreBCChuQkMjOaha+83H
Vz0DzZA2Gc3/670WjxO48qu1UoYJ4EWaK+9v3YtQNzTi91Bjq/RlUr5OhmrMPp2B74Gf2lPovWGH
pRau1MDFG8JQ5Qv+QY6vqXv3yvFtY3McdJIbqbeQCwW7jiNKKSM8nRVzaP8euoWD/xTU5vzvhClE
PVzukZjt906IkRZSw1DMUCGn+N8AlZr6ApUgg7UstJ8+9zCgKnUZbcaRY1DIgz1gqaUTFopxOxzD
riLjsE53DgMOpe/OdDJPMIMCa8k9Lnq9cXJ1Oo1p8sBYzN5lk0vAQ4DNvxui1uXBx3cx9xPM3CX6
SL7+gKqIz2TjYmzcfI/8nxZq73JEtgH8x7Vw8hXmqlytfrjgFGM+HfmwwXFDFF9P/ImaKQm+rYEn
FqzH5rgUBf/qi5QrN+d1Ls2dwM83EfGTenqMVQq2fZvHrHstqCFWit7z/NitnevpTPSpTHsPH8JO
FU9kO0zcA5JWWW5cu2qc2oGlGgGGpdS5CgDOL9LZT23OZbNKrDXoTRjcfSOWh1MAMpMWPmX+OyV+
Y1KLFaClIi9nAX70bJc7cAzfjvB7iFFWpPKk4jPBUtQZ/we32h+ly6vxz2cm5RR0izPSOX5TtYZS
zaSclg0FQvKCAQ1lfeyf2vCbcBLyUWGBnXMJquwxFBwauNAHgePPldJXOiJzmlPg1M/SWnK9mkJ6
aazahyGsoTaBzza5Ujw7lVI5GJiF3Z/BYvEg6tD4VthkoSteZhfDlDSPLh7sviB3wA3ukxq8RqlR
IY9A7bw9W8yeIgj7j97Z01Wx0SVUxRITqju2wENuMW2EMrFSsgDZfEvt3ZS190OSi7zHhK17XJio
md6mM4ZFhNOY2nnd10ixWfQCVEzIvkVK90VL95IglpsHk5vLXNqoyxaGmD7NURvw6Z1E+nAfIi5O
aqCTu0iKj6s2tU3rpqHbagVfOwmQHZVpZI9Ru4z88/OViLvQhfeg+grcUleJfktsW/Naxl+9+mbb
f+NOJTdDMnDU5wu+956QVWvmIal9JHp8/L5i/5nJUK+T+STtlnAA8DFxAvDGkq35nuRlH4gGmO6w
s+U/IpLsENFevumLOkojb/ZAUWZLisSlcMFvbZKtyEddtft7MxSRWZH1myTLCOrcBXfKtEJckaK+
WH1ZwysRcZns1TxaZNjf+zXjgI8OW2FzZk4SyZ+v1/pXvYtASbJ0M5Hi0us+BqHnrVVMx8De2Avz
HE+RRhvWydQDbhvo91DNQvxY8m0XDQ8oXyRD6ClYM6Gr7SQZ+02liPFdfs4mft+UmMYA86EdZ+n9
F5X91RHlkYp79XjDpmMZSZDzatllixTsMvBNF8ovgabMIWGR19FLyDdFmaXZ04zlBd4gaIYUazIT
EPEal90oVhqa+aKnGmjbLnTo01gSg4r+Cq/OzGtj/QvkFjm/5zgLDjnZT7YSYvyUgqBxMLCyLNQa
bEld/HSu4sSblem6uzvHrkBfF4LcIwXpGZlM7fMSE9Ri4dYURiNbfeksik8UC/pviAPQzxZoIUks
X5VWglCT1Hvd48FGe4Zs8JM4YmURMC+4sBZ3qEhbcUsgFOEFfNsDoKK5J/z3wIgGYtvEFx9s+hBQ
hzq5FWw3rgHEHlnPd/HBqv0/SeKHVnPABHiwwYY+gEluCnaoga7hzRCqDqREnnqw51yMBb/1w2Y0
UsWF1JZfDN0LaNBCG3QQ+EF1QHRMupDwGwrKkkLm3rSywd0tg+EBBSFGEXgOn7B0mf2QgxuB2g9b
Qvlj4cO8UUOW/dzUeCw+lTqulQqmJ73io14/sK513/5JG9qdZo4ouIFgdekocxtYcXVsAg4CBxkA
qT2ISW5/1p4ci22ujYx9dVZcwK1nwSdw8ujoRxhjwElPXXcUjWSQ5/jbZUxi1zIJv9v2b35JA2z1
fGiDQMU3H40/DhVn7UBHK1KEe5z4iIyGZLD/NMldhMXt4DtDOtzf3cRZa7Iv1qn1hfIpwiE2M+OY
tWSx4ggJHk8ibPx5HQIaR6jW95HH6IuoYul0R/dXfQfJez12staqce7+Be4UtxPISuZk/RWwVVZJ
iKs+oDnCQpf3heKLSOuj6bDMOZX/Xoxt5L4FTVs7xpcpbh3dt/PkIneIQlsmFvYo6+wuP0YuPq5J
UBF7O3A57WYboG6/mV7Qa9JStjDGymWyePNjjpaqjevcze82xSN9UwjJniFN0SeiVUiF930SSR81
mWo6itz+UMT3mKRJJJ+kI7x4r7SMOTNBHhg59RN7VBQr1ogU3xX1UdsciCoT08RaA+1rmqRuQryL
4wOkrwrFZ5jWL+R3UYJ2o6cNpcTyYDpvBEexJVdQE9tTuO3nCqQKOOZAQr1PHgjKaiqFeKS7uGcD
o4ARn3CRqQTzKz8AVmZXO5/DkAJkotSvgAWgY/ojFzY8sRnGOf5nj9Dyn+yY6khX0L8yJCbi7FqI
pyb/jIHjkKT3Kya/v+esYfBHkz06lGzuMHzaHTaIhlvahthaJa/ITjgRdN0pFiuMghbWlqK+G3yk
1lp638AcrCr+SpcbYzWLiZhiPge18UVJMm0Je8wyPd+nntzjbGXdWpjH2ch86TO4+KHCW5Ux0ldO
Pxdxm0Igbyn1vMbG+NLoVX1GohsaGSaoULBTUHOH/eqapOMUUKTNFuQodlk4cjZidzO3Zc7JVnsT
U7vSMryiJ1IgO1pjzNFPfSMo+OWezU7TkgpbxVm6fN2zN94X5XhLmBwJR/eAC4lI/fSssMF8R13G
HdjP6Chy0onXGNXc6f3yG7pxGE5ensdTE0WetP6xYur+JwMAjvQkNiig3fkyM246TXwjk9PVVGzG
8Wnm1ZJZBcsO4Q3ff5zBortlOPf6eCEl4mDYb1/OmOeXSjkY4bFYXeBCk4Mo7Vr/CfxR2SHA1ycP
vxDZQinh97La54MdYVMgw1wnMaztJmo1QWIgHKnBvhsLZi+dPzMkDJD4X3b6uIf6ZWNm7dUzARnb
6CvGtcVqmgG+TRTx5feIGJUI30fO/oKIzCrBFm592nL2jUkDcN2OClm6FRXZEAa2UUoQJ8WUTdkD
slANmqSKx6Qfw3ef5rjBfPwR2ePrF4q7TucoDhYmSii2d43ieLfxPO/YN4t4OMvR1g8j3n79e/QN
Xc0RaiBpApQuZ9rRPTFHzEh/vJz228ZCgjrQ9ivQeBmyD1XOotdv6kXnTgARWa09C4DM0ND4ffVd
gZ+CyKRYeT3BFKMRuE1cabxoL/Q1S+KK0K65kyx6wOGXQOcussPdfGYhxce1t1GYNf5uMqYqb3Yp
+vnd7iR3o9dZ0niegrbYTYQi5q9LPX10124tC/GN+ibj2Naev09Dpdz8FzQhVyfKbmmlOg3Y85lL
GX1Gfn60RnHzVTRkwRuiyvGSgg0O/JD6nYhxqubx/d2zZqkcURe6bWrD3Hr9giGFGGFdWXrAZVVx
fxyaT/I+HR3qlaDVSToke3hpIZ0paqCC2bGxLXJSewuzs6q9iCXFswdeALiLbaMQq8h31v1nzuaU
O4qSOpuJvAtJij250x2ZQtwgB5ggWwMPwTGqxdYARDWFgPlVqihY+XzZNynGVEEGbeO9KzUNaykM
8k0BoSBOnggnkM9W5jdlHIyos5q3hmwH8IYlugXUIVWNZEVAkXcZWf+6Bb1pJR9jpCuSVvcYPi3+
Nh8RMqYtSlFFxUiBd/cH3JQWZ6lUU7QaPlMliSnO2BQfX7TBYi8Lyq3i4aV1ZafBcq+nDLp87TL9
nLuLzXjFVXqbMwcDyVpEXBpR0JXlgbkgnDufmHtHmaeqUjwGQuclI6fgbe4WNC63Z0ZjOc5BJxt6
c9Xt3+OeSTla73pXH8E6L6VT9SE/1gvQwdphY0NRJL3KgBMOXJLPBxr8yET2mcLVOzGVQoPas9wt
tGuPRXwPQNFxyV0u6eBMtO1GqYPFaSsBtdiwCT5wyjaxFspENMhLHie+3eV6N53zcIjw+PfhTxrT
cxsNYonOi93qt+dPDE2VrqumhwPvXnABB9RamVBei1gwOkqlKHE8PiGqcEGT6aqjHfD+FjA4fDH0
9FNcfu+1c9zqLNFJ/M3yK1i4grKGJD4wlBvdsOuZT3LNtMxZKyYgT2KjAabu50srCbBT38W60yn5
D1dDLnm3kC7f12kI0sp4WsEo+7MchY2fVqESSMEIAfNSDhs+/zSRFAcJDMsYNqCZpbowjZR5V504
G/doLlREp6BqDb4lUASeWwPNQE5Mj7DyjN6A5IEjLT1VDrqjkUdvzmuoZXstg9k6kd0lshNJDQGD
LytdPbn4KXE2tw0Dgk7q/c1bSQLslOrYOQsNzo18ZVB9Q1ZfQZ1KKExFT6O3mWe00yH5iSJsD+gU
GKMoS8wNCUDuHCX5Rzcusol5pBCdgg+mC40+uiE/WuzNvu4Dy/WdSXCnnleZcUw8JAviAtwd/DJF
xwIcUjj/ftPVkvK1ohVjFmMgtnGDrvNSszY5wa4C0BBD7EUECNOyolBpS/wcUABzwm5ZDxdVaoTU
a0fkwdJmocidcEH1NKeo8DaG4aGR2Ts55Moh6cgyKe0qVstOYsTMyX4BuoCYlF0BoP5LMCry7L/l
kgl0BgNMtigMEGKelB5DcEbRyarwyQL8ZomuiAr3BaFdz5ngz3/62uLL6VRbXK3ymCpmmYQyxSJw
2ieiaQONME4tqks7tydn12TiLCLP3E+wHrQiDGzHIaoWh8jKOPx6DN4Xm1lA1PYNOqO1AmGPsKmE
NtoNtjB5zyPRroVlioU0mr2UBZDoKiJJT7ETOzIr7QW9dvfn8YPOnvMggWvfhmDZd8AzU6FxtB1A
F7pFZhEKE0J5g7zZ4Yv7h4SWeSPNpPSkIK1CgW8Dy04szea7H9sAyLuwmuift3wJEFbifF9dDAuA
F35/PzF4bU1ZV3WZPxjYjwWuOBPNxEztvAWeyWhUI7qvXsh7NpwQUvyQmNapZ4he1KU0CjtzBzte
Q39dfs6iLA/pM5HAYBWughJzGOLk0gtyjxDcnXIQDemLZT2IDwyAbmz7rlSSVonu3Qhcgh0J6JEc
v2dt4XsKNkHZg+bI2b+vBTkRYZUPRkkIsax6rhKn11vSYud+R6mYq5z+XIbY6+eGxQlqDyHIIXzs
zaLI17ftDjnPgHuPpNf2RtpStWmZw8+7k38VQaHBXdwWhrEa21KRWRxKc5YxUZQnLmPuFITVd48O
h+o4bKUFbiCJKNRuCYZnV8/ATCAyUchAT4M432sn6qy4gfcdM9ghCIMPfHEGWe7C/Drv4d3vDkHI
muZ7FBl+sXlkNJP+kT6C3wbQ3nt1331FAu8Yfnzixl5l8LpQdpuBnWHW9q6oNKY1ZTznJl1hAXhx
Tk18Z3XZ7DNZjyu55Lb+aXgdJXkKOS/Su5Be/ltgW92lz9LhSKN7SC0S4B5nCnBgjpCuGe15ZTtr
cTF6o002rDs09IFU3LtZ/VJWTdDa/RJI+EsXXyU/I0TirAoaSoH/Vttx9mVnYT5zFnQbEDTn5lhG
YQEIVX+1v6v09h99vJ/modWzbXk0kmO1iT+3/jHF5rQS/eGQ0KMcRnb+Qfms3jSjn8hM7vAXo/8m
tvi0i+e1BQpQw7UZMlsE1fgErE5LKwp6XJ91dNg0z/JrXPa7peeA7BsAYUbDdRtGCY2fEziXuL7H
/CSdEPDjjb0GKtrQGP6Ao78DspgXoycvITbSrJbC35yFWQ5KSDX4Keg2dC0JgjV1bEY7+/TtlPBy
H5pGGr8kv36+/j1WSokN9VMVsZI1jhVe3E3qpM5DX8KHdTE380tIvaYYU0cLq4q2HTmJeq5qIEt+
5NSheQDIHdQ6eur7iMZQw0RFVSXwBrBO7m+n7I2aFUN9wJtw9YV6bp4PEpfaOKbkaksIUJ0w1zfz
k7aJFgqWSHeD9LaPWL7KpiZMhzJN1ykzDwu7s2FIDAPaAmbZz9KMHbBup0hLctHwIiIl9QrVU0G7
IXONxon1LbqUAfLsvYe7+8tpMhsDycoyIwB+rvjTdq69lJ/Ks181Tn4cQ89dzi71NqNe8SSMo8QS
TCTHHlICxiUg+/EpbhXmdOm2Nb35vLjaSZqlzSIJIl0Hv91r2TEie5zZn+lxCZ15O+9ogiNjMRg1
Z/VNnj77gOW4+faCTWoz8oR/djx9XOS+8MDLQnOwMEMRefDDuq+Vrx72u9c6+DBuktYsGJdTd+eI
4+GSDT/nqVPDlT696ThN/CUcD8jXQMIf2uV+XKgZiPkgIXJjqOZS0QydrR71meTznyS40VtfuBZ1
h9nLN6rHOdNlYyR9lh4tCk9owB81G1nYJ2sP05Oi772aGlGi6a2CyqQibzDclCOAPAA8zGphbA0F
k9a9eKY9bpk2UQhclwW671Mw7YMzTsMFv6irep+7ex3XLDsn0ksNDMvO1F/CQIEpEwqRidZuZnWq
k/3sg82Iff9pf9EOzLnQqPzNZ7ib3ERoLuKz6r2sKGXhs9skfBP5ZwrLoKKDGnNfQX9NZfP8CpVq
Gqcxw04eca1vIr7koAbRKlDoCVA80WrCkxYvTRSLz33+oyCaIod6lCdFPyi17vGAXGvlhjxSp6Y4
RdcCQhsmhCkoIczaW7ARr3Y9xHFpwzOpvLmMsP4SXymWPIYItXw6jgFVK9aVIqb3fRHA3IJzjCwA
CQ5p4onmEt98lbjN09xlxDXT2aEtnOUoR64U2JczNUbDOAzyM28YiCnKp13dMGJnr1+8lZ338N7C
0+zJP5DEdZtbg9C2pPYEEJNgHgRj79gvuWcL4J5GUAihPPTr/LA+8sGSXxB3jWNw7OOsZji5Ua79
63QyFlCeqGFLu9dP+KlpP8IZxu6bwOXP2mm2pyYg4NBFo6T9oh134xIEJ/0z6mOf49qAfa013L2o
eObx5aEY95m6ooY9BbOt4TsNuQN52BdywP1RBJaBSyV8NcJIZwPSsx8GbFBeoFczruydPurpsaN9
u1ZVx6UTJ4Ss7Kia/gsYFQhrXWNHEYYIKTDpkr4+NUA6d+hpok/2v+Jyg4WBkWqTEA5LxgnIgjhy
aTY762WFVs4Dbhq6ypQSmEsttn1RQXEtVtNTREMShhsjDZIMtMkjVVn6VJo3aAvOfXNSrc/oWwuS
XzREesYhkRtht3dMuW/OeeymtP/WoLgauQozvRFCpf5aNSfw+QH3kltxMrHCV9+vdAVtZQu965hY
sOu1jAMPE4Rs9puKmMtOvvmuhWCGwNDmxEd8ufF8hC6qm/2qrjSjm5WymUov/9xegjZVHgCURS37
tuZqkxYKQh57fnS8LQnRBueGPIJWIMDdXHEDLGMK09LRXuRpku1P5AJ+k0L2EJiDCAde+Md5R0Ra
EeccsYbqo8YX4Z+IywRaBM2bO1QcJ6AJ7wkoj+yj8xQsqajL4dfI9QAZ3B9Udz7ckbvMNVcAiSiT
ETAxBVamcCm3NisMmHIbfycDw07OLgJ7GKFbelHwG5w2W7PH1owVnsgUjjm/P2rUpLmKJm7oik+/
N0mYAq4b8GREpbJ8ZPy9JE1PL3scaJX63s1d/Tox7Gi8LztNPDBwEpAkaiTn+b2/VZq4pVYG1ycy
Eq0z/nzddkS3/tOw13TjGxrWX350VcoUs5sNTXzadOvFFnmndRJ4IUbWExtSUKeHy7fM/m9+NQeZ
QjayTHUjwocLTEM80VGGwVMUIfbD+acLs68O23PBIAQE0hD35aRJfvA+1X3qUGrH8Y8129KvXzmc
u/p9mv+QWFnvBK7HoyYkQuHbtJ3IbO1bqDu1rPYwHkwGuJs1i16syGsQjhf6x/AroirYPMPsE3X6
rnrvqqcxK5OdCSqwQoooIboGA2f1si8g6f0AhmPwUlxgNOZ35AQV/g88NarZkm8I/p8Ru2FsqJiF
fiM+tpiXsRh1UhVC5Rlq8+FZ+zyUQQ1PzDSP1IvoZ1DsbePvDK3egKCaby0+Onv5O3eUJsZdTzZc
Qr3573CmGtQdU59Fx9YMvEAKw39cvycLpUVlQQ8lNNWpg/OJNJL2+FbwsNLgHhKZeRnjHRdmbMoW
xxdWg26R4GlCCYjy7bRGsgOGzcuiYCvQxeK47k+wWOeumiSLWXV+4iYLkTsN2H2EyEZwPS2bySML
FH7qyF4EiB53B72VVFYCzikg6HtNAexhOMIApoGeTT9ZN3pAYuJpMIpw4Hbwmyh+KQIwEZaVyhMR
DGw2e2K3YViXW67u1cQKZwqVqVBHlNioi0k5IK//2d0y2Nt7ktocXpwRh1jhnqfs85fwGdLcEgBH
LG4tPVycn/nnyJ8Sv11gNdh/fcMKYjxrBB+JWg1NSK6XGlB816G/QlR+XGpLXNNSuRX3zHcIQAhJ
4kxxocZIB2Kwv5YuAgaYp41z+81krWGjuWc/UbBp2v1hzw7oUlepErXSAD1FFowl9xp05ii8qayp
dCEJWFiuWHp9o708UtM/YBrOKbqgvC5nH3qthCazb9W0PKNOR8/UHMaOslQGlxGCD7qk6j0RPXTi
Ykf5xoAqdmwXSMH4zOVC1VZqRHRCGcEKJTnY1gau6tOpf8xGnKTJ//6P9SXQZkIlx6FG/ju4ALvm
VIekX59SQk4RU9Xi1ROe+TCdOIZUOVWEGIQjUw8CmX2sz0Sb1eUBMpNlZ8lPN9QjmonAqT2ApfD+
iikzlFDxl2t2JVMnMRt8Ing9KuqnC9+Wsge1uNPm/MD1lVCVr1slfTWniXYZYR4Ev1xFsD7F9SzO
K3GDaNCdjvkxCL067/sEU3WZhaP+xl3Stqn4MZ6vKv1DYkdzoRi77n7ScIRa8IrjIdpYf9n3e3JD
7DtImcHcIR8cKu7kecGONC06QsOYdI6WKydSnY1436Uk4gzIzscCOIGY3iFCBb9ZJyPn1WcQDX0F
i9NchATCYAYcXXvt4Evg/ryuEKw+hlWqkGnIwx0fmW/LJyOmp2XBRCi8eAEGcxwyjok6pToDS2EI
A4DElTNKTg2SlczRvyL5Xs5DOh0ZgmX/KwoPd+gwIUNZ4VFf3FStfcrLeN+YAM9kyCN9k9vzjuVt
eQYk9+wpqJiJDv+PmRzsV5uJWSwxGXa8WXhf4MX1DcwETc3cvLKADJz2Ef52RxXBv1kDxymr0cNg
tnU+jd1aOxMWgIuJ8H7mnbisuqVwZk2+bojZp4+QNEb6OurDx1ZtXAER4jyxrOEOn8KcZmeUuNAU
yDnkkRXO9hmDo7BL1McZR77y6SkX5eNY2Whxw7GNpS0K+vHdkMj0eVh0ViaItmUekpUMnDJVMK+M
MTyeaea0gVHHqMGg/22AzxAgZZFk7pnvXjWyk040KXtDVSeCEWf7yAmOOJA+2l4XwbmCtRLpWN/k
4KwWhU90MAXo70lVzTHjX18Cu9ddkyloKWW8khxfXN2wYSX3ACzqtopZzmhdhtQxFpSpyNO09DYo
LH8ZEQH+ChYOCkLSmDPxkm4D1e2402dkNc8I+EtB7A9RQ/DxZOJOm3i+ef7DkXV8sON3vCU6WNcT
B3zvpIVcckmelIlm+snozhy6AgT8vvY2jDnfg+oRHE7ui0M+s+B4IKUd2Q/Avbv4qRkC0PH4FeH8
NlwwQq2ObjXOO76oEpFoC/0eu4V+X58KnGdySCxF3QZBeNL3CfMzbuENWa9178B/eiZhr3AgfBbW
T4PEO72OVSwDWEu/mSFUJtqxPTfJh1IMej/4L5XjQ7vJkgnclQsAqEkxwdP1OBT2+7dK3ZcXbKfE
U7TYVP/u2haUwiBL33RaP53ghwW0L1Mfzwj5MEMFxPqHsgwBKzx2Ps7KJHlY8xSiKij9E9DjxrlD
XXQHFESayvB2eDY+Iqw7sebyW7skXeyUQbhPq/f9+UkBdQkIZpWp82lzhqbxtnuXGKbF9OssiNuM
tF0lit8qJoCrrzxlDh/G4blyg8GqHwoxdJAYJiwam50kXoDjOPIkzsqhetFdmv37HY5tuc6Dmi8v
Hb7YUxUmQJ++CJUaA5cFjO62glssDqf807QCWTOllVEdvZGh8K5JscvlgacsWdp5Pl5iGMaRzogF
/yWfbpLgTce5Ok6orE1W6GTu7iPsRBxOcrVb+O3d30o7TP9p7RkkN7UjyiWp+aCafKx4Gaa6o+vr
gJxGKW/Y/aVkJKi7BzvpU93O5GDUp3GLXDNHBmIvJlCn7w9n+2fQn4P4gV/4vb38d6eLBUMNojox
lQgGGlZY82oc7pSG82YJbkbuci9H6RtKDItbMIQxfjSX5IKyRL1dAVOHC7h2P+Cd6vvNO38dCA7T
+I7rNF6pnrrGUIUSmpG7P4dD5ZHRlRyY9aOvEbqANto8j/OWZdzAIU+LRsevD8RYffVhbBRjdFlV
nBzyluwVSMsEVrys57mcP1wBvaFPatZw7q2yu1J1cRKGlwwfuSIBInLCuPAzFxaAVHbX1hzGmxM2
l/dBeOkSJ5Uj6X6jpguK1PPFzJW4Ofm5NiTmoZGUYfwjfWOxn3OGVg4qCNHpavlmppbZRH+uwqRh
HCfJ8n0ur3ZN9WNBn6gajiBkAaIlRYRtfvMmuYFySKawhFPBCyapQCVvI/NtlIl4I9+JtlXuVxJ6
Dzv1migCGK8HK1nPff3/8J25PGSGl57Z7EmkdcNgCiNDet9orOu5takPl89KlSc0ZGq9iBqwKAYu
qR1BsOed4ZyudyLZNXvitQqv6ybw3+4VoLgc59wbh4SsMLQ6OuUQRH46Vo0Jsbu4u7DtS01fqWJ4
zLrUqYKFjf1IBlU/oF4YwKjNEFqzOQzd2CNbm7KGULkPyJoc3utdUJNr//KclzDkExDp1nBcZkA0
75gEOkWKhm0OIzShrqkHe4N6L6S89IcEzPQ6wkOzeVrK50jXLWJ2udiX7rJCeLU3tqV6ti3iHiMi
bHJ3XERq3jsxfbrIi5yFBMRqAFyWP5Vlgq38Qe5cyu6x0vEDdYj45TZlkW1IlORO2ZD9Ztz2IHzV
tjR0wbhBAVTfW3OIP9v3hPtfihrPn6nG2+Z/HLHdSrJZ/C7ZG+NIhvGSyZhzxrVS32MZ0xHQEOwj
aZvMn8lzt2oz1Q9Dr/z7KQHAdaY28Drdolw2v87DLnhux4y6gR5dcMycrO8AcKbNzUPXrFshq5s4
Yaw+C0eOCEggaka0i1j61q1Ein8fdTt9+Ze3E+Soaa2IfVpl3Rwp1BQTE96fd4GuYaofxUHMH1zw
YPyZr+gkB7k80PUZLkS20wgc0QsxoDv+EjUKiP3L8JK4w0LU+y9RZonODjJ637/eTo5fRiymZeo8
vDEFIFYrMklIKny35sag2C6F8dzVeBwrzR278eBaP7lQxhoSjtRukG/msr9ltNdUh7vm/1soqNiE
34NCRE6Rs59WiFySHPVLl85/aE83h4NUu1J4o4dyZ139pNXs1nVF1oveeDHdEwOndcxdz4BhNYYo
IGJevAIYaZIRqegZBAChtSNwrLwP3O45O5+68jooDReZFINClfeiYmVM4OPM/FFhGWoWj4X18cpQ
//JZ8pUjt12hJb7U/qb1+svoegRiriWoGP8kDuK1Vy7nMjqGJqD2i9SauQPdm1uP/byjJv8DwsKe
Ehyf/CiLKEBwFMfIVoasvizLRis6ou4zO65LIZcChSh3FPQijEmagHiuaiRNj4QHMCrfTnMtFm9K
jHWnSqzK6Y0OiqdwgW6b+TTK+brimqeIwQzTHGVNvwl8GB9t8EMryFCZQfGLekFAW6IjAq1+81Ho
VJiFE//aUqEvOWaEkJUASrvfLkV/44f7VC5+BjKAhXqKK5OiQP1T+0QZu2OvXv+dHMLGKDhtlAZf
YnQQpHZiq0sOHO2ysh/CA2M4sQpeZbJ7jxEJHLboCvMBItrryu4XR3NaUpbCFfh3WAdjVV335ZXZ
E6+azUCPK98OgWtpKBTcfsXzITyPu3uDmXLb9MVXoEZS4pJqK4yX0iJUQ0jQWIcvCQsJnsN/dV2z
U0iGWmn+OZ7N9ZhfvbJZKPKP0eiy746poSV+Tx+9E49zGo8MfUvW6OG0rBK67xKN/Dgu07SFIIyp
AJ61nzdIacqQC62Q9OVlVcPhIitGWYKZ72VsAtX4vg80uZahReHuePsOXKv+Cody1E1M811y0XDe
l14nuH48Pf1Akg5oUIg7TZCMovAPiSTz1pxzbuOhLg7NmbsI7o0PFVYS5taJhlk/KUz9T2h6FjI0
Ti37GwhV2tASIOIC96tpx6chXuLImkQ2nlbbXlIfk6xrvydE8k8Ombjlx7YEJ07bG6dtTcS/bCmE
DH0FpQZo7FgarnjW30DChTIuc8KgsgC86W5xXTHv30GPgErO5jtIA4D7neR4i4paZDi8DSiJzod6
OKZMpuep7X+z9YWoUxnhXAQxKJq5InH/UzZP/Nyo5d26EwGkKSUqhYJ44zuxRi2PdMDzleVRn47n
aIedeTu1GCRGu2cVU6JjhfRrAMBWJTsQp1WFYwkjKYdx0lzcBzGGGv2UCLP3FD97swRaNH5MLsOy
mudG4NPG4txNVUtV9/Xk4CQBQNRIw+DQ47rffh2sefbYR6XUGPWfOgubl7x4aiF9PQ/4k43frD0k
ay8VMEMJlwl4STZzak0HIlgVUosUptvafUSiHdzY3mqyhZQJP6Iq9L58qGPoMdL9c+qW0bsirw5B
EVLLGbBgNug8R0ShD5BDV3cuPQUXQsCzoAmty5GgizkUnrSVyef3LoqRqW+TYOKBjKU7dTUCfc7r
iBEu2yY7H3q4zy3UKDsx+g0+vu0VMNwznReCId8QQsaGiyQ5G370ZpxKxj4v1lIssJcYPTTTJz3+
qtZkHnurweTWxp4TBzau+4uwIEP0nZWiR7aVHR4LG7keiN2DHKFkcG0H6ytPh3VBOcPKzHZ70F8S
hWZlS6TghxewJjKtFkzhfHSYCHTWVb2rvG4z4Dvs2htDc4o/r5s1X5smRcrTcd+tEwFjo1u5VJsy
vOtR74TpuO86vpVioYysfvi1UbGCUCcDrXFFDRPYN85A4hAK1uEvnwWmavsQgCkK3tbNs14xgl3d
mG1GHZL/5J20iL2Fo1sTIJOjMQ0Wn3jQmQMcIMrjZdlNiaoloDbXaUjbrfI78Dy6jZzti+Wz8V1N
Q8fqkBEPC05q99+i+OFr+gj68PG7/8FSkNDrnszu2Rsb6Ta8onz/N8S/+lV4USgeWx4ZX4D5m0eZ
711bwLff/N19rOo3Pf7LVVfEYLSpKOx1CEOi2/D4POHfNH+sV4oiEwm6TSDd4XrKsNIsWrBQOpDJ
rfo3iF/3AjFl3yDOuSaYUgWwQz2qMWYYFK6Kp+FIq/UEz1hFri0SMPJS/avtZIymFJuuQP6uoeYu
hb6CACV+tgCpAUvk4Jhf90IKpH8gVQAvAR6rxQMAuzexy1qfOOhdm9NY8ZFTHoO5Ha/GQsYyuCvu
KLJX4eWHrWDR1praJbqaN4xrOB1hlZzDWsLjSunELHBM0U+3zCY0Erpi9qtviYp2TnqqzDjY0+wq
xFXB2x9X03fmfv5NarFHOEQXHF1hG7kZWjuC7HcbKQPbGmiPfu6/dxg9OS8YuA0GG/dEy+yaa/o9
gOK8/sryDSY5+t7bFGX8xG1awITMfy/fFPPxbzKYwcnvB5mxAfZ8sSsMMq7B/6nv91Wrt9HwYDAb
mgce906STFlV61xLDy6KsSBiagEE8A1SktpPC06V7GzOCP58mqL0JHi4fR+SBo/Mn8jtYrHoc33o
r8lIzHzJOqLjjuLZtLxeWdnPgHCja+Z7dDs8uJcuSx3VP+Y0UpruJlkB9zqvL2fHaJ1yBMd7xbkc
WIEgHSLU6ybbeYMqzgTGNy5rqVwnDU50vIUedz3GhLAq91QMrtFotNKmpiiwRBZrZ5A9byh4Tr82
Vy3LF3Rw2Bswdm0nbMZOXLqYY5ZqZjN3xmv8X0YBAUcodDYmvMFr1sqQ7uAI0rqlivYeSWPBhU2z
VjtSIdFnU+TNHLW99WYjdLWbQcpR7ygXTqPgY1t/iO9DfrIGOCgYjjQTA+pfdw+1HVAOFv8PishE
jkHhmtkOMfYhL+Q198eOMZytJcJ5udqX1dEmUCvXkzwFCAQH4fW7Bxn7E7rbWAw/4DDnRXyU8qIo
5OwL1wB68mLtzInqs77yfzJkbg10nruy4KIZT48b/I7uho4MrJLUBAuB8oOpP7348GDg16kT6OSC
18TJ1omND+cKzZ6xmRslmg6ZaYcOWBTD2t8TWzn3uaxhHhSWH30yeWl6DJR6XM440fRsStE+Q5vv
C5C8wzFEGDjxSHKnVC+1aOfddPd2/uq4v7Ot3x1ZaQEJjyEZSZOIXw9d2BscE9wrMz77rZDxTELV
oLgYo52bN0ipH0NP0xxEs5BqosjidYhpowhTrc5IGSr9Y5F+UXFDq+Cv5pxYGNLAOCOFNCZPm507
i1iDagdOgYUVnQCknuFzC75U3mc/9bs8mvW+02Zpr95GUYR/oyiuwL67tnT8ytLWlBuNSx6Z5i9V
ghNzCKFJ5sB7833OpWWkW6c82z33z0CVKcrpof2NliosvqeFoR5N/2LMgyZpv/ltZAWizTfMq28v
p0190DIj91uPTX+6SFtcgyj4aEg1KvxXKhXI/fBBsgcQcOJURO8l7sfeI6Udqq8YOp7A0Auk4/Pu
WZm5ZCIzYenRHhOclkWLxyIDOtmbeEneRVeBmqrbbWRnw1r0D0MyeU0g8mozVSbccdCTasNZ9fIN
WRePV+t4ZVQLRl7/ccJJ646nd7f5q3x36gmMrVvqTOjD3zswmgYe5YQXdzJI3UpPZeVeGi84tKln
dToPj4Fi8MphUQVxhETlGClswbpa5xS/3m3Xr23oX3m+TSZz/OF4LoAJNoVZ+bYpCI+O49zK0Qzs
TnoechmlspE61LX9nh5lwX8NVMLh64p8ptGSzQ0IuCRKydU1Mv5L7gBfL6gMKTOw7pSDUci0gPar
1S4HfnfzKNT3nmh0FgZgzJ3gXjkbybhzDV5Ymykiozntr/bOTkjDpiJEv8r02/THyrpCET6DwCn+
9FoyHRYpA85y9wbHCStxHUQK26Ye4v64iVMGGuGNs/brv9/yR/9GkxxaoJwXV9jeYO1LIqugF/tg
+wlNiPAcNB/iu6cCwsPVnfsKL/ZqNApoiyCz6uwRQoki0p7mEFQzHzFh4GlLM4sy6NjHxtRRla2q
h+T04k+eUjnlcM8tw8t6sfhuhY9Qv8aHCtnFXOGDpzmdbG1JFPSSsA0mxjX1mpwd4QEKan3f5ezm
xdq+LnvUD3o5uAzszdM1/fPx4kBvtDtn92hej3fjtOKFDbDJxsdxAtJhPyw6CBRmhJ34mS3q/aV0
FZ0Keh8l4vvMNXAZkWFi8owtQ0sp/E2fkod0fRicFDEUka8EavE3WbV7pDC0xv2P0NQOoHQrcm3z
WHGuldNQ8Zs8XxWw7Ba5cWtVnZP7knWPeR/UE884Nyu66ekgCb4Rnp5O1OheekobFAC4GAQy9a6k
RUl2szC8soTMbKD3VRa9Ri8+pThj2uG/hqIB0cds37MIgxSaCmuTkIfTktES8GEgyTI6IeSHejqi
BDsdwbGgsaOxf6yQfFl7UC+TnPWhSxnJgtMqwQJu01xoLB63R8JyDnlnzpQP0JlnM4OiF1f+roSV
GZ2xYjyANGDBbwSvs1NjGoJYmlOCBT28caSGb2XcQstf7phN6n4oKCz1gRpLtJGRKJycayONyCLi
AUO2Rw7LoHY3JHd8Btzc4TWoZbIeNXSGEyDs3/BbmZzy7TXXsJe8M2eqZxrQMrr11EMRQXlBwzYq
w15ilpyxl9mReuggqumGmdrxBPKd1m6ZJ+8KRJvTRMnYpukm2zpuaA8xfHsDk0YqWTelyfZuOK1I
Zla26EdywZx+D4rBLGWIpTDONxbNOSCwREsIVvUk5iszTWIJzlPgN/977KYFycRKJdvNQxb2lgtu
SKGFAoDeCbXTUx+ZSaU9AQSfD9I4AllW5dOMX1Qjj1ajWX8rKQVqrGku/Q6giUjufmcIUJwGMC7x
BrLAXUGSJdoL6XSIW2C1DyDFoTMy72c/EHCzelO6Innflw7FhwTCen9InTHUqlzeSDSwTcELI7US
N2YoJp5B5xej5C+/GwtuYin5JOi4VYKJfaFth7G2poyiIn5c2Ys+iu7nAt/DgJLFDI2x82Yq7La/
+rbxZgHUaKkWKfaI4FuixcQhiUtK+ur4l6UZdWJkXjOtbh3AUENQ7rlSgM2/wL1J22ITWSK84RDa
KXl7GcHHLVwboyR/PSEN1XBZ0ztNvqxIUAbwZXzvX9yPByG2e2j0lEi3VqUC/JyNmwHX3kJ7z6Cp
LbNlur4AVhLXkfOj+lsbdGwkgqIEwku/I9J4Jxq33yNdLZXc3mwjQjNjqEbZznrzwVhdPtPev/Sb
SzCLtZ99QEFjWr6+z4YYmuZHS4KB1cIUax0itYxlTvcFQnR1d2yvBCiQ6OjyiRObRVCKHLxUT5Qv
x0Fbn80HIopxBWgEyzA526RNR54QuAxBYO1PyHjsHzsSfF1EB9Ov6BE7o0ezPxV2g+xioqaJfzVF
1a2AR6MdxXOUjtC0LUDws7zQm95cF9o3VkdIIGaNHh1gaq9WsTSXTaUramIabHjDrJWHrpz7C1t0
1UuLSDKVcsabR3TE5oWkBZO/Z85SsDlR+pwrI7c2cX2OfJRoDZg924S2hfD9ycp91oF6bXdXDN7i
vVmIdOYtsWpGI9NtcK7rizW+Hm1aOzQamiSMgyX0ck7XvfdbewLCadtuABPwlY6EmUYGpzkfHbZ5
iuyuvZVU2ed4QIUVqkEFrquqzC8goV696gc2tq+HjWWrV81G9oB/PNIlG6u6lvB1shuUUeQDEfmG
QeHWF0/DjUguUANnl2931nS9cxMEQlO7RC6JlL2QN4sfsmXcA493Un+7zblVVwBsD+yXoU1chGFJ
URb3tiNaa83Bj4JXFDI0Fo64NsLoFwhz1CzZp7Nvr0SuijEK57Ebm9U3wQTD2Kbp84d/eUNBqU/h
pfAR7eJYvob6ruSXCJNgs6umWQiVZ0TVOcTmJtq24toVp9BvEV8lTOlvpywkUHqnzdW57YLPxNMQ
eRgWvLfRYM2dgfLVX+f7iIHqXsg30QECQHSEHFa2TBcDgNFkeevqJeg900O9fZ33z6+cS4tYNbTG
OoDz7qzpPYJ3ODfTX5mK4sWtC1MnBYNMscFU5FgcwPdI01rNYpAkbwOeSt2AvL80xM2iAzG5uK6M
v2I7ynawcVDy0RCs6dHCaNzLcPYC0BHywm7cE92kkIr7r/9gTe7/AbVZCFwymKkPYOS20cnRirWI
MOERVffMy/fIZDHxo7TNetWuWzL0rYMagUQAwPBL/+7KVw/yvlUrh39wxBidl0TMGeBexSycWEkC
MXIBmFfGbvaGdW2d/bZTpu/zuATV4vFGFKVBvRgq/tAffLu14Ilb4cJT4Lhm+MRMvVzHD3QYzvHr
dGOSakmeLXv3aRQwKb/gkeziY57xhNaYwjMnowrCU/C9O17P/4h3SRQ4VnwO6l5yBO1o/b8/pyXc
o6PCJMHrnD31HpEfVjtcgb2GClf+YtQiTJt77ksQpwm30htqhjnWTST0KaZLWW/di3wyCo/N+td3
2Dkf/iMenX7MSJVXdi6AuJPVLwTarrz9r6nP1lNW9Yfe4HT0qIMfnSpNV0FL2e6asid9l6phB1XH
439MvZG3w0NZmS+9/Vy2nw3n/9uLcri3HC+7pAVyaZzTgsnLQIdPV4pSbNd29mSBHcR7ZkUx7Wym
V5Rrf1cMJgNBBDhDbHTkoDQsHc/W02MSwEuuE8FhznQHePTpAPx1u9pxqVA0+p4bTackyXqzHNNo
fZG4rLa/MaEosHpYAC7Ofc0pTo1p/2UCVBmuZHQ8fyBYTQx0kC/zx23lfWOj7NaF4Lb6gHo2d1Lw
Snn045uyFkfhDkfsZQi9B1D4UVYRuDltiOg6nrkVLqD63loVoBC5Jar2EKtRexH8dYNbp1iYgrbs
qDxvSXT6eZdvNPs3aFTh8RDcFMH41njFnDDcFugSs034wL4n4w7RzLNca7VipHR5ieQjdT/tyWoP
OZV9KDRHfKU96QmICEYKLdS7kExxXbGIZAinJSuW3fKoKUYOt83xleT45xz4T6w2qhhyR8724AE+
gtlNBVhsokgJ5IEvkxIXfyegQ3JT+dg7lY+8oeZdlR6rdfVXma+vRhN0PgNvTK59eDuTxYp+5u6N
l9ovWQ1tsHqS6/+LjacnRn6Zls4Pdf4GbuahzDb3ZvMAGWQjie8fbNW2XZUFOiBgRD7oL4HijkLG
MIEWRIW/acYVlV2xGiOO4CUELRjySTq5Dh4xzxklUdK7XJds+HutOtaq9zhQtDUQHQuIDuxJkCBU
51fR7QPVkv3/uvag+A4WoDt3SonWl9FFUBUgUGynlV8wWb9yciWKPTH2hUA0yUzCmqgSfFKgUyg2
/3w07ho+CV7H2CZrgYJkUAcr0Lsrbvws3IPAhe98kGD+tBBnGMyzAHtv0j5yu3KBqFBm4kjKXd0V
Jv2FLwPOWDKPbxbnJMuOy8BPEJve6CEodMqATGpzKcqzir8Qj5elB/FY7WGlIlYs0sMMpfsvR4PK
3uepfTpqZIlYNCP0Mv+WM5nXmI2H2BFFk55y02tp0khCu/TTqij1QEFFZVY7lz1pvzYdcH/Ufuvg
fSZhgU7bMczrlM0742Z+5g2Ue+PhXOkS3BRVZKbvbBKSoQJgASwqvLG/S2N7goERg0Kjuc6onP4e
SlfCZlzwUU5jVCykRS0Z81WGNI/WTd22NZp6iPEY5F1GUiTuRtQBUe75TrcmQiN/Xu45CUjnlkTQ
svABmj0UJ+qVGJoihsuPjWO9WiUeH1QG8OFG4KvYlvE8zYQdydg5MvE8j9IyfQ3AUrJ3VteHdGZU
26vXeuui40JZC9V7pvMsWBLbd+ZYXYNLthmpjS5729YOpyfuGl5GyhFdhhJwt7E9iLaXjkUoOTp2
AQsQkT7MLRM1eoDEEeQ6rfenbcl7fZvTzMeQRrtLKm7FKVaWstdtl4bnbJb6KNcp+6n05FEUoJ0J
+zBM1BPwoypZKOcmbe7h9GaRP7lz+ekTnULsYfFoTVhyWNywBdKTB0tBorP491vSIhzaIDHoapa+
gZpaMhE8HoHdH35eeBYIJiXp0PyjTsnsx6ZtpUEmwhj5jiU/gnIKJS4xSOEl2+/paxRpC6s+Izji
NLpCzqm28a0t2r/IZvru4UIeBJhEcLlSdjMotJj4oNggCeEQQA0QQzga2PCv2s1cL2aGt7skfLu6
Mr4412FNR7DjDlJkQV4V3XQV8Jz/dGS4xmVsHcQiA3mH4MkEd4MUNrVHQ8ywsYeKZ0WlosTo0EH0
6Ujvvs+RPgnYYuT1MMPqoqB/5dTrRsChabjyszdvEc9og8tZpIlQn3P4gnTEDB3pJjQ0jwy2YelC
aDxH88jb2Ffs7GIIgKWzYsFKNzWe8/lyy7C7bYS2qCm43kRtn3I2+UaHI/bI9pa64wTQoyYSeHvn
2GKU9sfu1ZMSIIhTMsnDZZbxRkNCnFn6GgUMS7NU2QQUNUTv1UzJHTzEPx2HLopalbzqpw53j7/C
rXwC4vjrVHbf+EmUWnx4mNCSHeNzaRU94pD333H+iLL8LmKvw8x2PU+uNzLpAT5sx+GFwy4xPcAZ
1BzvsdRj8vef/30Gi2v9Ov7tknA3HiEPhdsn/Uyl4K4+4OLkkOtJHiTGajxnnAJXYd7/LauZnbuv
4pec1WF4W6PyYeybGLVFk6lVT5toIu/mXNbA0rwRIfmUOJ11CNpunXyDGiJ6VrxydYuIGbxGFylz
b52WbWh4yvrhsdmn3KxcRZ3Zw+0Nicx0Tavwrs3aPmU3XlN3c+G/dBEqi2RafmrvAOKi5qQ2gheL
pKiyWJvNU9Vpv6yYr0ysxNn9YilswDwvRFjH5MkIi2lQJXo+GbdvwswvatR9G/Y1K3nW+vKT39/0
nVUmd/n8oWGTzbdmXZK1IwCAlOAYJKmI9bqHHNPPixKn4XuqKX6Gkbwj4fl/Q8hjB+Z2rAZjmyTZ
ZTd8WbkEeMkPZoXcdwumL9sglqn1wj7FipYl0dtiTrmpoW964Q9zD3jdzQkHJdkFmq3XNp150ua0
MlM29emP6wibLOSGt9QMlhNBS9ipROlMM+OJTrgmQxWdecypENiYqW53xcQC0sIJdABDDTnkg0Ec
foKqH9Wq5OEB40EjSstIibfucmD2oFEFldHWjd79dzEoyuXO4uX7KvmvZzJ0Z9lEOX1tOImqLeEd
V2mc02ZqFPKJz4vT0p5bZyjMfI+bIYVc1bVF02dameZOiHm3BWI8UIp9nS0/HSJYlumY6RRwVUPE
0KM7itj19u3826MBq+tXrITbAAs6CJqWuFXSXVC8NmzMqPNxX1jmQqCGv39ZtwqveD5js8co2Qt/
/cvcqvirDrY+0X1Szcl9uA1gojRoIfu7H1g3y1L4+E7rZlShGcJUmEWRo5CAXv7j3Neaq0YI2ZmD
5Jk/RMNaXeoL9hvRE+4aFBr0TqKvAwAho0ziT9nXHNn4vUqFA4buSx8SJffBSRqXLajgsvXklW1H
MYZSC/1QSTmY8FxdwVZnSxpaArQcAIk8ohtURvA0tBlLKMbcWjMh4N+hLiadjGutGSdxnXURCpij
tVzutBoZBG9G5BAcWVNS1humjjZIKReB8cRM7fCUW7u/K8vu6O5bVOIreBREpjNbR8OK5iHe9GTX
J8vfjc1fRuOgHcRTsEDQNWvkYgv4fLPDNbP2TNc99UUwnZmIZuPil5Rww20UB0KEYV1ua9tsiOuK
I7poWRYdR65BVDM4Bmt6wv3WYNYcsEFVtNeLepNFN8WO/oEcBFlQyDBQrLuQV+au71gtvACrRRzF
sngzVwDndxEcG9UJgctYGb8WwA5qJGfyW32Tamq5Vb4DL65VViqwal3yrG9hYmUGBFYudSDHa5Vi
CZ0drU2g6FhD8EkILejiH+wm24la7wlR0yTmRTiNPECSxV0uKsqaA/lYcwc/JHHPxKJEhxTOA1Jz
5+/12+Q9QfD3Mk6Zb04zjMdAb0Bu1OVaZ+bb7/85C+pa8OvyDuhQf2viCuRU+RFG2bAwMIp8t/nF
CuXBPmvZWe1N49UGEbVt+kSWgMO8OPsMbrFHD8j9BeQVJHM5n8Y0914qk2WHw6q1A75PsHz9k2W9
7Tzen87tBOb3Odr6p/pm7m2drslyelQPCe+M/GY9R967hawcfFiudxbokfd2GznjeRvReFEg9Hxh
dWjpWkk/AO0RqV16BpwlN8ngD0BuL1eilQnJ4XFnIioZWoOtO5OqJqDGMb7S0awxpK9o+blFKqeZ
td46DVCTfev5SDJOe49pSxpmpvBHzYYazqNpV/FURnDjx4xfC8Urd7X4PYNHZmbyefYE26aysUST
/vrTGJ/irdcdy4hNX5NXxvOZ8mBVfV3tJENgDyDdwf19KTnBsmaRZEJk2Mx2FzdjhQrazJTlye3f
ZfneSZMz/8QWRADNWUcgz8PId0PKnojLC3Jf2VXuITLX7eqwzoSViPclLMSGaXISRYjm7ge/6f94
1U5JsrFlXoyxb86gXxnCc6rl33batuTC/AVvWXyQPq+3bwTUhI4BK6SiRhExdt17ojtGWWCLehtr
qEy27uY8+poLy0awmWtyTi0brNm2ikLG4ZUVO1vwn+yV8YVLQ355wlxgkQ7MlJJClIzqgdDnUx1K
4yT9gRWULcpySL0eWY1u/nlMUjeA1c69E12AiYUhdE31Wk9FLzoCv8xCg3v9rWVpBdlU2Z69d3gg
NJXn/0eHTy4XEp6jIh9Cw5kDdmvMrdTmn7BiSmTP/e1G/CTUDH72BJNx0yp2GxWYTpjtiHBbpYIC
fOmNa14/+mj6igxgGj++Z1PEUZQ3OvGN3kKZuVf/bO9LzCFYSkMVf0JEed0EO9ju8lJJgZpF98G9
QO35cyw7awGr+nYCtvHVdxJIwivXemcDPisAwNGxDOyKzmvYj4iF7yidTXrxAeVph3gEEq2q1QWD
rvzrC4AxIecGpHfgX1DVNy2P/a6PqAQ7IqGdkx+RTemmpL351j+4VnkCkXP69uChZ82UKk4d7eXD
twbvtHGt26bJ8EsIkHzd7IPdYvjmakd1ocKShdoq5j30D4sBQBgitGV4BhhQT0LhI6rtXVBZf1qt
flbqVpTuZwdtRpP8KpOYetekdK9pl0ytdI4PZAvSd1OfWJgZaMECIccmTcydgHS4iZkLPhXSBSAs
dXeq7+Dus4HDx3cGXm31aBoL9kTwc8tKOFXfiq0+Njk/GYHW8GCTpaWto10N5wiIzLIeV1MOjbJs
IxSMmuBP26WqmJQ2bklKVLeELycH5MiyXCxAvnwhiIrSA7s6lMMoz7lBjSdNrHA9M2syAZoTlVsx
p+KsKTDAMTKbhecHNeiC+dJYUkv6E3iZHxNKIjO9zNByS1VaWFJrePTS29hWEZshX6BDcbXEiU94
YipYJOqzOFFhF0jsZOUvu3JFbo5S2sFRwPzzhx7jJJJpAKaaIQUoD0RJIcWSv9SyQNglGOiyODbi
YmStMTMs/GFyxJinV00Fh1hWp/Ym7f8busJx632LAtRrVUm6CHXYxPNAjB2+weRAkjxHE9jaLXE1
CnvFl7CJT/5UmRz3PX83MUYd8H32bVgAPylzSHQDFeO/XKqj3UFnKSlRzguN3Qp795/eJuvNBcgw
JQQ5frgTWt2wxApvVW2vo4gXAX7DI/sEjyTzVuCZ5VjRD75IMatFWkVQn5iKgVQiy4/OAJyH9NT9
y9vQ77+oh5nVvZDIBbcRz81a2Z36P6GnMhJkZfP+H7vYeHiMvLuAzdC0T/7N//rtQ/soNheHwVz6
OwkfIm0OFH22fukdvel1FVSO55L3ZZ2zpmbfkAUE6F8utc/i+l1o3vWvLDzbJZ2PBMAh8PfBztat
HJdi5BMnSU2VZ4paCBLjGDuzv3PyD+CUTtdoXnR6+SAn/m/kdYsMBTtbKkqlYiIeo0KeXh9AHB2H
Zuf5kth1poGiicOP9XBn3m/KivNKB5LGMklJdt+1bE05QsXw8dxs9uAd2ePK1aTUe4A+uorN+c1R
ojd4smJkUL9bApE0VxmMkZy4EVWpAWalZA4sF7BCO1fln+Fz+Wc5Ni8+TratfU6DygEehq1iYgxu
xzIpbk1I1jHLfrQdtep5VYQ1xiG0mDaZwwTbhp2aVqAlQpxE7AdwfAbTWjsSPL/KsiqrM5zRFm+a
WkL4HI5Asg8NgFjYJQ+InuSpgjMMkkus/GUk23LM9X8CYrymQXx6MQWMZHv3/0OxgZmBGzFoOf42
ldoqg3YEywB5/X99ELll/cCph3ddExtpIraMFki4ffYHCg0UVGe48Nu+6BrlQcUEAh/8iykX75Re
oDoQVMyKBhzwvkrHHR2uBZ8Z6BvT+ed4XnxghIhMV2iRBcWAC1eOcF4zAsiHt2uyDL+9f9eNoWsb
dIKf2Lcsqe7onuym/pW1Dn2zcIzTOwLqNVC8XoyCBGAsRuvz5xRgSgmDu8SFObObTgft0jqGCU5y
uPpZU7zlycbzGAJAyZfHSz0eFYQZymV3T5NJJLL3ffByt1yoFTua3Gmo8bpNrUiM56tawTm7AavK
vQu4sVgXSnZzVzLCFfpbIsHhdily72WE3frRUN7u2ynuG1CwscBoNGcGf+USG3koJT6V0+W1oS/L
nEzsISdVngZHIDpPrqcDqpBOPGrMl7UjuAQb2aDV95Vnv3t6GJNA0lZxqKPTa3dKE1+staMXU6uj
JlgnAeQhWrUhyp3M/aMYi+aGRslYFEJ9439kbQWF5h1XuCw2whAsfKE1kPIwislKCsZkq0qgm6vE
g3XKbp/0ldU0+MU5b9hjOop6b30m9VM3AT0CyaKqd3bq1UJrE2Yv99PnKCzgaCm23SnNSgi7jKEa
iMWoYq0gL4GlBdHWyPrD1x6/ZiIKjF8c7GlfECFI3fjAIogHIIUyCapVqz0plLkuKBmTWDsXEcbj
P91AuYYy9gsmmSfRCpZyCWi/WqB7ifYAPDit5lJoxw9FNHg27234x3oLSH3n0lJOmqKv6VHqI0db
WIb9B5gqCaBs8bZ+B5vj8OJnAsc//CehXZLaL3Ez4B4LaF0IrMTbAv5IfMirx/6lyYgRYoCYS3mS
mU/pjU6mresfAemDqyd2kemfG0apznRyMWNxa2XEX13YVld2sVyW9xbjUKzIHHyBkM1b0KysvQ5U
UgwVov21QchuVFYJBy2CHbztGUlRyu1kT3QcqvL9YkRyq7wKZmvWq2Un9M2lN0hdPekJKRVoX6uQ
PKTEfNMRxA2nEgPQrB8VDX95/WBe9/iAiOeyy0Rfe4MNqmy7zhwDzIYLlag1rknkWCnI8eSS7YAi
HpGeLCzegn2Jlf+f1+7ysNjaejC/mmFLdDpQydYFouOHrwooIRrwmRs/MfUHt6Hj+9mc1YRvxlsR
vAFE0shzLw7ENG0iJAnJnER5wToXuXy7Lb3c9dppvClUkXmcLEH32nqLwD8CGBPpHj+c7aIGDX/W
Q/OT3AriHZWbHXZFW9RPVnGlq0EDI9jqa9BkybT5U+cuL8DW9USwsXzHcnP0PA+VT23Ssn5QQINn
M0gZn2xGVFlHX24JICuj/IxIiHiDHho3v8kUHWwS5iKLXECIs8izXUXLaule1ti8wpcl2N+cW0Xt
hT7xEWdRJtKfbetGdKZv8k5qMxfQm1DzlCCv8HBfarPtM8V+BTUb+SGq+x0RuoBC95mvYUhU7qsI
NrrYOgu6Gf7QDT4BvnaXj5AYDMsT3vCDlC3Im4HVrX9TyHZl9tv1DdGOemSngaFywzLil6jzXMnw
3FahYWQ1brw+out/HFF9pJaVkxDbHh/fW9dXGK6Pu0+wuHxn5bqc1F6f4xDmW/43QEu9cQv0QGYh
xZmXx4xpPinZ6BAjxGn0Z51+bc9EK1waNL6dYbHxv/6fHHJCyvJGcZdCxiF6je1N/P1fUWkWkrSi
kc5VbzBJHT+XCXwJJo17wdStTlmfmCG9ew/SBCgjhppfpF7Mq+mOdt0o/Ptwo+yOTBx8KSmIi3RW
47bcZtNPgaJvEI2l6fjKoHCy2Md6W3k09iNVNxlh+q64qC1J/fYtVhyG9/NSL589U/ThaSw0PnKk
FRWB7fgeqUHT7B/qUjtBJsQU+2ghkhYU4lcSLrRdqksTM+SzNUAjGc23nyWVgJLK+QHNsuFRkJIe
W4fFD5PvRKzAxgTCbmpmqkSXqL356xzKt592WeJHducwOlb3HMrvV/Szg8jnW0MXRg393SHRNTnd
AaOi7xTlsijdnog48jGaASBQvKToQatABhI6TXIB8vpxIsWUVMvJke3CLYaW+YyoYJ6i16IsO3Xy
H/AZC16sC4SwTOCqUyyckqNAVFnKys0wzy27OG6ykQcE3hLn2IVX8uktbcyu+bhLWI9AsMXJ+GbF
CJonjsW5s6LIAlUlzZZiSJoUe3qw3mQATTkDbW48sG2F8X1xiUzW9NsSrVvkRU+uE4dA2X16uWgr
XXtZSbBkW3bl2nNQoWesZxRcfhyb+ghToFSuPAxBblyDoehtZRRfckFNtBwknKmbXIwWrfv0fdlx
vhXllmvQ3MQq5Px8///XqirQVY1PlLRATVaarov1CJaU42YLc4/7MkMMRUOJ/v76w5mtD1ZOZlPV
JwyAL9LI3clIhMNgZOvFnm7K6lMR/kh5JlpECUgXDPqBmmS21p/6urkCGt8x5ECpqCj9Pz3EaNlH
j+3RTbLTNUajNp/WipLB/ex4nY0e0jDKS8HY2ifqzTVej8ydog/unnVLei1Lb56TrL39SPaQyA9O
CxIub7yy59UPzRTAxKhrRt9YXTqC+FZ1/C4ATEih7852Vh0gfsrwVAH6IlHRLHZr2NYVE+SvCn+j
7lsYM7DDxn4mbdHsql1NQot+MqO8wRcXhOx6PBztf9Ik1GiNiHhqhuDwegEZjfjBPk0QFPxnt/mW
FV1JJcoQKWrGc0aly07tiztIcI5HJng4049QUlEZ35h36NZawPeNiOsmZUanpzaxlMU8ZM0cKwTc
D56JwOfznq+zJgsS2NJuufb19MyP+9j0wJe60i8Gjy/iZ3nB1CaH5nFbUvgi5MI4WlGioqVmUNs3
fG95coFZU3X1lv0CtAVB5U9QJs1DLhh1KCvbHLSpt4Zxj2VK33C40jDsYm99/0Q/9NSaWRGQKRSG
/cxWU+bFVSmn0P0oKq55RvwaCZvTYX5U7FMdJLNj3Jaj79VINb6DipCh6HGu3XFk/4D7It/S0Nq5
o37618I5t2rqbyOyrDAU6R2GPaNpgLtaO1tLa4mYX1MWGwB2Z09nOX3BQOEyDXdoBKc4pxeu0msu
MGfeHBiH8OCf9p5FIubFQ/cXewd7R68aGFnDr5G3DI0CZhbJqJLZaKthXxpwYJr3oCX1Sx5IA9eh
yZs+KJzDkdrTlIpDTjcAczjGpTyuotsIO47saJPtrSCuLFpI7uAUR+/1sSruVyWeJhmnDNLO6Zcy
oT9TQYEMMefiIGXHyo115JZ0w1uu3uKNN/hItVhF+/r8HEa/gECAW3gfFCRZkfUGVp3PVkAFkhTy
4zZ7U8HUvQlQBhlnOxQG5x49DSIA9pm+uoCZYfUGtvJNX51glQPiRnvOV74xypbmKrDaTkjiicfs
ogihtNuSoRwdg3iJcphjZz1IGDPSJirXWa4G+h44GGeMu2f5tNHtKk/fd4pPPOKMG8vKAT97HsgL
3F/0oD7viSi22EIO5xdjq/GlFP/tPyFlPAqCiqVlzJoj3PFZ4NeQui2pEn5j3GrsxuohZ1iJFoJ9
sWS8x/ZzjpGZuATdiOjCg5zO+uUevkTRgyA0bKEwkya4LPNeOoQ/zraRJOR1EXzzO0VdCEX9XX88
jS7yB9vnO0lMolgfhdpSdZmPX+5aCDgs8HbPpgJ29jRG+h3zA8t2GwxXC3xMRy/+VQSW92DOTXZC
ozmQ02RlbcfZbQ3I0WlvffOUkKIu9qyXWxLvIOGXpdYZj1tAQ7whN3KJKEO7porp61rwDl4EncJK
MbnUTWGid6Q5a/O+NKNMX+d4gj42ZjsIWGufDZi8QV8EnApy6p/M9lDuGXRPEP7ys6oK/mbcVGWW
mKr6Rw/lDDedtaP0qqyzc1Gyz7Ug/LBiT9vBKYwCKu6J2DJCXdrJwetlkWLo5gwhBNi0A8aGS5Yu
TAMZ71GDPCDUr53VAImmmMQa6gYXr1nFVFKb+6ZbPE/KVIuRU3Vkd6hNff0WUNwBIXxLbtudlx84
gESzQbLnL5pWJgKycpYrXKJm5UXD/0WsSnLOmxgx52QZv9CsQDUlr0KKnm+XkDJqlEbbd1HqfTVy
Fyx29gJAtCXjl055lZY7Y+xLc2UgjBi2GszgpBsyF3pwjSDN0Iaioid/h34unMgSjVAde/oz2e8P
kdIzsIOVQN33rpJRuADLYNBhvxjwPAJRojoYI3BjI5eH7UcSgH1cW/ZBD/688soDsc7RImhvj7+h
mkxcLCcQzWU5xfCXp7OY/TYCcxDSFVZnebTx7WaQBTRi96krOufjpGJdiDg0hXHUtRP//gWEKxnL
8tc0PPuPhILDr/8gzmlmkXJWUN1ayuueNRDAxrhqtFn6SAc+8R/Q/+tICcw2tkF8rHhTibgtaKko
N1/IKdYmN8/zBUjQH/g6sGwqYdBDjB9sSLzZC1pcIn6J7i0QVj6Df9HuDprzfAm8KO9apLCJdHu3
PPaiD05G+RY+C73bBSDk97JtUTZPgmQgkaHsACD2hDyceTTASxPlYdFkQr3WTC/4RJh9jv51vGtU
lYRZl3mB6qolD/onY0sHaHj3wwK7M+UH5THCOaN10P9/Xiu9uhoL6IWhXVo9kEF8nvNMH9iU18qJ
gZb/4xY0f4CAEvow8A1+eer+g7UK/jdwmIbh1XStzyaiCK6IWnjsAD76XWBn5xRa5dKEt/zNiPHf
1NlGI6csh0NAEBRQJIT6j4sWItjTaiIjEiykJCaJ5L5L1onBvsMVfbjtZBRDQnjW6y20pyZUFLU3
HW/2lk3cj93BtlHgbg9U3fafgiPK9yB/CwpNhcS/v+uXrzsMuWKTb9crGNj5cdST/fxJbBnHEQ7e
6DHryo45P4HSpZouYz0GY4KtV+rT7Gw3l248fTMY6mM5WBqT75Bi2l73Rx7Y2mMBMJIwQ2gjZyBj
7+ML1wAVuZFBcMmC31KqOvv6w7NKannLEw+bReSN3gbAzV6TxQ+vWytKrFjNi02Y53+4I1G/RBQo
dPK7bHKZ6ZW5Ic2s3e0J9MOObu0yWPJdlE0PdPA47FPl5WfUr5masZFmi1dEL5FX3XIMCgU0EoeU
WwZP19/wXK0alGpkP/fe9rPY7Q5xRxzMTCgtJAalNk34ojeDyhxs0MTdFh6xVGIpGGZVnZH2DvI/
Brb4UuB53G4z8l1ZQGiSyvC4f2X1PqxrHppM9EUcS9U7X0q46z/8Hf5vl0tPitTgJBI+MeNZs3NM
btTviB9lG/LfEwzE/KANoSTW4AHfSPGet/fianWkrAzBJ6NmCrPn5c04gnnVx0wLjqCowJYdXW4W
ZcGkSzhHzlqs/SeaOR2cQJY+uPXBZnMWe2OItpCowuU/oInlOXV7ASzx6hcwOrFn/RYpVyExduvl
jlaP02IDh/ybK0l0tDyBWZn3ldLbXrgsr3ZoufM1G3LKsQ/+ec62cMSuNMMUKMFH1KF4PcNgDlTJ
oi5oQrkh5LrCPKPpU/noUTmshid3woSN/a6MZHes+moxkSs75KqiAxeB4zcyIkE2F5YSR0l8SUmG
s77jujEMczGlNGofHW4MPwkfjs8g6CAcgYVX3pjCC3wsw9MklnPC6iemZnWwI2clWCAQwUHMkrlI
xH+Q3oHoIScfkRn1doeZjjqk/5y0aWfojWnZ2ATZCRvNZuDLqo/kjXq1oJYZkbj2chTyXzriGgaM
N6ouVDlMYBbS7B47PQ/xjRymigmLU+glrelmxF6ayZ545rssoenm38r6WkxVBNDS+zf1ZD6DZGGD
L0iKHChR+Plxh6HUX8yB6odVdw20xzlx3odZbuEMCotCm8hT032kII1KS/Xwnip48YbgGI5DHfoF
84wyIdl2K/BH3cKoRzi3Y1GjDL6ZagcTkL74j+lmHlDJNRMIXRem6eyp8Mm4oEaHx045pt6QKk4C
FPWvrLtqM8EJxEvvRA0tZ+cBQCo7nOuXKbe1ND35qDdr8jIU0WzPjJPcyQU8diGtu5n9pZt+6Cfm
fX8xHeRQomoncHBHUoZpTF9BKtsmqxnuV4JiKzsyy/i51Cbx7uRX7P6+LS48vlxZ1gHNjaSCHVXy
SzA/DTr1PSpgQV3gsi6DNr9jmlDRdyegh8A7lAovfHYZKarfdliU+SbrbJAowEoRPMAvZPXuFA8e
qL5otPQVjvDSMTgfrN0Q43BIKtboxSdVeVyVaYQVhucXmSTynattOpe7tFwEt4iV34UMgxRO8pgb
hdD3OujVhvASpprgjg4AZXBrnq70NF+iGRjJOnq5c/Bma6zUm5IPO0nnzHxm9GI5V+7zM98tUxUT
PQcuIJ2jEABI/3hYfJrpx1lLF6+GvKo2ELAuCM1eED8Ty0lwOJdlpqhA7D+YBucR0zARSaJQyyaz
1gk/jjnlbEblVFhQB3ZQ7UhUVA4O0jS7q9ni2SbRJP1BG/CvGLMMiLrE7l3EfvVuCM3VC+Oe6tjv
TweLiTbJmBPIb7wIE6emwmVr5uQy8TyU8mlgg0r+SaAUPPi961Wcj5YrR6oeXBHdpTeMGmkeIDyR
jsYgKHTAathg7SykDoG44tXwtUJoJhVMvqtuLgQ9RCx1wp6V5LqWcWeXvB+adc8w01WejaDLR7o5
UKScGTNtKB7waWyt0Ku0MwVasyIlzdSIU9qa6miMrx/PS5hBt4URAx+yEPdCvmbF5mKibUAwZocw
yjjLpKpHWYtBsg7YYxse3hzzRRQvAdQk+I6n8LUya22zTVX7O4I/7NemfyRQ9rH/VV4e8aXmN8u3
kDepemTKtNREyHpmVeSeHe4/ulc8I2SjlUVK5ASb8U52SdFHZH3p6owNnoMh0y02ONFtrRA9gFG6
fAlXHMElUYvsOErfNvzlPUcvT/wMvP3FuqPg0EWde1EaWC+MRfBigrFl+1965qC2VV3GcWEQcJXR
2nm4yDj4URp162eX8+1o9DRKKsxfyXlD3Nh8CuLXPA7SqOB4EX2RvIGOGNuAyC7/xBtmYDFeM/RY
omlpKy7g29d3nbh2KKNbUiFeqfXXZda44n2bXrnwqp9AYizy2h74QktyUGNyOhkR7M+YMWatpeCX
5T1lCrRXMwkuw70B8QclFqGr740Hhx6QmZMKVu7pfMxp6T/zAGVL/CtFKI7+RxbmS7LtFJwh47Vm
plkz0GTpKwJ1QRYJN4m9fQKyr+sKLsOA31aHZQTuo+yFTFfNEgJo4uJogkQFHXGr0qMm61khT+2j
spNtRkllnvYAzO+GNU9nD63o8dTfQm+2pC40ZXeiLOzJ+UySxGHOkdNNdsBawjTJzrn8kqVkY8zo
A6qWd+FZofc0a8MHT83OXEJoAC8P23L3lj3b+nz3Fmq/tVE+rfEf+adaPCdKbhpwx72PraekvBH6
NwpDZp1DOXpYU7bgqwHnPKCf1fn7diB40HKvlgUEzDByeGSZQNDWFAZ1GWtNY9yj+6fLiYkjn4ed
CCwdP0D7sM5OtW8I1tertuUvqncREEOsrbhY43lXcWZPHChML2oHLoqg5kzDGafpxhkJnZsOGVE4
k4QDe+o297zvfccySRZKiOt3nH9GAb8AHlr1WlxVt1ckuoUoPV7SD2lMfyO5qWGLtAehSOLKelT1
0cdDEMQlf7/Q/9HsbMilO9VCAv7lThbZMTHqUyPmZYHEL//aVQxJd8bocXqVLBEy54ZJKJzyEQg1
kzXqxhuOpZ7gDnfCLLcpBIKc3Zqh1b2lmSptT79gwy1NESRInPV56pOPhJBJS22soFG4t4OGfXbQ
o4L6COozCbKEyTOGO/ds9F7tRQdI1AMUhNpCfPTfYAN7ZRUx8/yBFgve9s0jZWUhuQV3GxCh/BkG
2Mlb0hR93juANfM00zS5W2pD7mBvyuewSMvrh3llpZRVxtkV9mgUeeIuNKEF6fiYMVfZjo29W1dw
tezpxMro5kHWmy+YlKyCRxGyWlA+Egd+G+hyr21HuukpXY+SFzVVcucA17TJ1MWtEQl2Hh6N8R66
ztL5SGZX+QB4LyutLEh70eG3IYgPTP3QjVmi/QpvCC1udx9BRJSE0C0e8fjvIsn2YHzo5/u1TSDr
5qaovDbnq/9K6ng7q8CHzpYyh+qfekgr7hedTTfweFIyghJNlGAKCh2OXqbfWr7njrG4etVTB5j0
oEqbKqmCJYg3EKShPEU5c/BZ1kOGoQuifS7IWjVNa8Lm2fX8RsnTW1RUJfWVqp5OF6AfyvLe1oap
HgGBmFWxf4bSZPDF6zLr4x4iU0xNbu7fw6G4CwnBegOZJTCUvqvqwfU08cF0ydY+rqlP1n2MV+GS
XpGlB92PpLYnR7rl/GF41arKcQBzFgrKrOQ9THi8OjtApq2AaBIbqzkEnkWSwsvPa7NhIehqNi1H
zUe2maiBbjAA6bq659VsrDRAZewpxelslA9JCiSB/7CeN3ctAN2EO9GuQX3kAoI6MxPL6L7VsZuB
aUYYH29H6j7bv8UBqn4wXTojzo24GWGt92//ZQFs57hhMOi0LmyrpUxSuGseCJRxhhf7wPPKD+Bg
Blw7Q01hOCePwJKnfK2zCVlAMI0N86KBYoZ8rkxgFBevjFm5iEyTs572R6kKei1YTjFa/3RJDFlQ
NYuKFsMe9Bw5mCTVm3P1K+EqTsMr8vYU/fdqfGauRNEhyxe6NNJuhC+QbL1dMiG2hR2Q39e9I+hg
21uGVb7nGMgllY5i+oPzE2UxCeKsw4gFBmTovJF015YT2NZG1SUtKpe7eqJ9fpItRJIgAm9qrUNV
gwpKgEWnoRZRDjSltL4phZiYJaoezN7UqmPWeZQDq80QY3wJVl/BZubMzJoqaJi66NBqkq/+wIj9
jOfjkM6ADrJyrlL19UtpUy9G2AyyUcEdMAGO7rNbmzz9nx7bFi6F3IOS5J6U3vTlIfUWwG4TM4qd
ERKiZ0uoC8LfgsVdE6c4f3Lxg3prDWPrR3NQWuaKuRRYWC6JU3RZE2CivtqnT/RUQeN+4dwmnyJW
3YziPDfn+a2RHveeHuRwYV8uH4JvilAJy3d/ltK51/tGV/+6iGehW2KXCRytZqacphEJtiqa4ngM
74m/sjWmQflQpFMk9de1I6yexxrYqN/9YyrquWKAnpN0+AmkqPijMgIANDAnpjaswRfySmvfcutO
d6GqYCxI39z2SJGRnoasQII4UMHLF2SV67qv83dXEAcJGQiGH1H5zHzckgyUxXZVr5QptnYLaSEu
4s1laZNJox8N159wBHyTOP8pyMKY411gHjrSh9gMite2ck4SUNQNrF6T9gvVsvwkghsqGxXCTlB7
ur//Y9mm3uMXMTXtAe2hJO769f1EhK1itMc9W3UTOHKBx1KlgQ3ysHTIcHRi+nCwncOgzItd40L7
78E2Hc4b2CY3Frbr4cJdoY61ulhejN1aFtTm7scUC2NGvnACupkcch22ZFbNicoqdtKrEzWPHde5
uOBfbEVkniOycFPaj/aT+CQWc+Kb6FqvHMElSJpl2D/uzeUDEaWsRa3rwfPJrzk4lPPXSCe0bgbV
UBa1sKe1z5hnf3UyYctdkFJe9z36j4wuCUmGMRC7XeuMFOE9hWPp5WGS0M0fq1YpOgWxOTsNMbXM
ap/wLMSu8dT5Pn0dia++s2iXA7n7y5DzYhUvKdVr7mrYIUNcpl4hLssqfGD7md9svVAi2nET2T+s
oSwaRrrMQswxv7aSGREW8QJt2cDSFzprOocOf6KtETS3satR7+d/dnMqCvQ9j0pClStT2lflRxRT
NVRhEujtSsfFzbXSbegy6N5mrSuRapAtvUCaZIXBQIr7axsx15dEH2+Q1xKMsdMMSR3MiR+f8L2u
AjPYtQ6CcAtSauzVjl6HmZlyWzObE/2T/skinSy8OwSF88r/uqRvh2fIAMeyqg1KFWB0FVwqndv9
AE2DNs5bksil0w70VmIedfgYk+qYxYheaUuu0fKB3WrUZ5fvChan7meCrgMlvbkOZPrBFEBYbULc
YCZv1wkoDBZBBdOo7Wcw7Gh8HssWKZruB96R81mo9C/fQx68okefhEAnGs4Uqm0d1eIu70yYetrW
4CzICsFtsXM/MWIzAg8rw5akXljp8NXUbPH4jUKdg5MWAq04XmYaDFBGGFAQWUqTf6hH8wgv027L
RQHh5HnSDz2z10tG9BTuAKZ4v1nqS+20Vya6G6TcwXkaN024AocFpQ7NJn2BawTUcEWQcUcFEMsH
nCCNAj8K3VwuCP9O4EcqRHdRl3FnzJIx4JSSM158RNv0RxmtVY0xXysdqxRjjomLkHaUm3QkMIRj
33sdryf7B9ZNpYE0A8Pn1qq8TywAMQN50A4sx46gA+BD0SKqTJITZJqsnAfY89HFe4m9PRasY1St
03LimnOHKjRkDnZWn4CAM78btM2BJ+LJJ5ammQlypizYmxJS+0psaRHrV+LaU9YZXVvliO/8THCD
yQhK3SWs5oRhgfrpjhhKb/Xp+hG0lka8rPr4lJpQaIEaXVJR6ViK5iDlEWnFjdqu83PUQqm1YuZa
2M2WH3UFfeAhQ7aOrewDvQqoQu9BID0C2dbTOAQIMxVc8VFqBRLBaFDFPNq8wZHqghOhXtOYjWrG
Ds5uvzHSxxCuV8j5AyzuShqzHVGa535akFaXB/PSt2HwHAIZzWuQztBSreCfTD7gi7sZd57/frzf
sMGXa8O+39yQWIiZqAOHRuqwLLXwSgA3HqxYVa39ZpMUACZ6UFlhWCZLcdmeKi2E9jWwexMPBS+L
GOTvuYphqZnsOaC+o/iViw67z8EjVj3XeLx3HcMB4UxYPVyuheGrA8DzR4PKCGIaUarvmAogoaNg
yGZK4/4EZYPqc6tXHMETFyo577LUv5QmfQvnNLlVOOrNiqHXQRoIMFBuao2mzSf1k/lua+Nuq3cf
MoXHfsoDCRgaVPEdC2nPWjL2cyaUUgjto/4Od0hpu28PNTgYoiMsI1qMM5q6VfHGBqpSxB8VP5jS
Xz7Li9J1ZRMJ/dkfn2ci+Yxy+Ia/HhJXPOObPXIHEEsGomamwV7XW6CMXx+F6Of3f8FY/0ihxzkQ
4R9PFfMQgv6TcUe5weXD35H5WJqMD8s38Q02cvFVJKWAn+/Mhp/0aKzyxmh0dU+cszPixu+zyu6g
NmJxLMwLKKF0Op4iX6pp/zVWNcO9V6u0/dj3VG3owta/MmEFJvhclHip1eDSTt2hpskERiRSViQH
80Ku9YSk8NT1MAlBU0VaK6jiI+ppcAM4ZDNSNUEf1n5pdBnngnpJDiGDCj89v9+PdupVBD2fhPw3
IhaMZ7Xlm4KXoBXb5AU57jgjLxTB+J4jgIyYOJxqd3K9fLsIDi9QRmA6T/Do+yxumE6c7QO4tpgn
6EyXEiuzG9grL3I7ywYIB2FyaOquRU3Zqzv5AQ1tfGWGk93bSmj2Z+gaFww98GBpjjARNqoi83Kg
relJpbw827Syp+Hd9Aw5yHZjVeQEFacVXjOD1b36+4bQuoVkDREg5+kBh0427y3Rs6es1CY93W4w
kISFBv0JQ+GCcBIIphTfshNnhjYttlH4ML62Pf1wW50XoelboHbQPKtXMK/QAhFLimFnCDGVt9XD
Ogq+/oenajvY+qp2dAfJ7d61enfODCzN+uAZwLNzQni/Z2zHw3Rgst5DbbIPKu2bOHWWJi4417Lg
9oUIyHV77HZDYErdx2nmAX99Tlh7OB+Ryg8BjM3rgqq8gW4iG3oZq2/hrQwOMHNjqU+f0lv1YBDJ
MWA3e7l02XMFiAHTzjDxN/48bOpXwCfmuX9t4gCCYPF8xWU2ekUja+QdrvzgCyJugz9SnLDsZxXz
vGJN3TbZYbK042Ym6BZ/u74ojthrYPChQEL6rsd0eXvIgspHwtXVoG6BTEnt0X3AbWfgOQiVVryD
DzR/nLmGiyNxHOXIfjU4qPmOlRwTpvMmUXSE7U4Zly2fXrMyX+3kKjawvolqGJmzDRsUQCRvZ1tw
h4llqfLvAWNmNrE9RX1F1+Y6Io5vHX97TKWYbjwHZA22VkgjFl/R3P2Q2v1ex4GuwBMAG9jMH0RV
nPnY2ade5wUVNIZC+MWAsAeXH0nMfrtawjcpZtfatnhT19pjnH7eGeMfF0ZOf9JT9H3H0dtwX6q5
I4OT8BVILHxFtk5+O/Nd3n9Jm8Edl7BESgXfuGcNCHtanVIxjUwZrrTteT7+Fb6L2o6FzSo91dNt
hh3T0dXZu87dvExaVA3G5UvayM9SHSeoBgw2RxumbRw+Onj48PJ9c6tksrI5+1l4FMEv6BK2DyAa
P48Em1lVpZ6GI5Ama9ddhzJ8mGTOVt/EJ86aHFt4QGEaGxWC6F7mqdllzFGXaFuXW4DCgYY3Zo8G
qPAazuIm+bhwa/hpi7uHxudMWiLuJcHtSbDzoovmydfGHT8IgivRTzSWeg4Q5kvuO+CQSxuzkxsv
7TRMc4ZQudQIFX6G22MsDn4UMi6QkzNwgjMK+qqxGCd376iN1P//i98j2wyrZIB66uDEZ4ep9InA
yoOluB0xRLtXVhREYc8YlSJUSdwdYWAqtxMwgLInpzFyiRR0JhyasvVIPwHdwi/4axfjIQVPOyUe
9YciB6b6y9iQSyCiT5AB1wEetdOwjhjs9aRMkU81jaAOZad8LFBPbnnH2ePytTySY2z0rPUrl9LY
74HjNjMkBAVDQ04CaOSGcSuNqmGAlpchKQthHzKk4sOpU7GTYFj1ZUWpFe2zdRp02zXDsRPP0Vpz
v+Lr0MDSY+sKLjwt6O9gzI/RSjQ5VUeUTL1fgvgqxyiLCTyuxFBUMuD/vsybY1eB+WtgbcmlulgX
4mbtuJF4pWYY1br6lrNwCuXWrYHvGcy0QgmY+hYsh4rYIlnAWNqoZuFqkUZd8Si0NpHyI4uesWJY
dhvCFyuYLhzPdM9LdSDpnKAHvfY1xXZAxFS5s4mPxPNj40C5hfHMDEhqQNvAaUsf/RzJo5TOb6Pr
Us7G6R5oNiXLA8AoXdVxR1dLBKlKLdC1+eny5eMPx/CXmPwX9/HpaOsyRqr0lT/RQTL2psvu+vVW
HOpRnTA9ZUrt7/zNekbqjlFYh/scWkaSnBsvDMICtJIZcWbEYToz88Zrh/4/g7ZSmS4pXwORsuNc
IRAVyKQ52oGs1+DQW4nAOm4MxSXAlV6iKOIYFd9l19ozy18Nt46d/Bg19AhLZjZoPjFSn73y/56G
M48m+6+Ox40R9FSDO4BIJ7pVm1cOBWKATOBRS/ocVbdr+XqTRM+5gt6Pd33GD70jWGixHj4b6bcO
Hdbx1cDql305pwNnMer9QnzXXvUvrgrPPVuo0YOitgPdfePiqdkpvpgfyVRmgVgOiuymSiGwV1lp
GudEVOy9URYgmzgRlicgxV8QuB30vdHJIABY4faRpxnvX1ZaicFPzWiZZFiu/cIQS3bkdz/lAU6k
ADgZ1FK0xQdjPwNTmfIBjXe7QDQgWriFbnQku467nNpVNgVjrzS/VXYbcwxHT4p6TAPwMkhA0hwL
x9NMvPC+vKNjdCPaFI8sNgQ2L2Mp2PBz/+KCAwGvcq1q/uGTquvLitYVScmDKd4tWoZhReF+AxQ6
E5VzT144/NGAFa2jB1zDg+tXkvdF0k772sNaJnUd2CniFnXIsZ1jfyGk36npe13FYSEzhDHVWeRD
e4ZEBw5qHCAQzq3yISkqdRcXbbJxSHuAnEvJpitxSgAFH2BWaxJ4o5EIGeGS6PmzEo94laPOESy4
H+a24chIFcuS1Bw44F3wMyphTGn+PUssDtIjQKMyULZqdw56BO3qaNZvwmugaNz/tc3L6qd1mHgv
kaSozV+JhoyUBr6ErgE9Rlw4ruFQ8p4RUIzfARo2UVOPG4/Crv21Xjk9XamMAlGjxMLTme82CfPM
IUKwqO37ExucrYnLM2ADxX9ejg9Ix6Krxzki0vqmWDXFfft1DKbjL1Mj575u+dBs4yqa8fRRVPtc
LFiFIoDmFqkyUDNYdcfALlpoPkMUUZPaMgEDEuJy7E6A4h2k+1GY52NQeRvI9yUWf+7iYzg/p7HO
JIaAKzpXovbnhOFxL2hUweoZL7dNb2WmW54YCyOxeQwhiJe78hdD2suJfZfCX3XhT3jgIZoaRbsE
pB3e2qGsfreIU2GCPid5r7J/g++YOHirhbKxMPS9DMRrbUKanmSLwBmEOlWsxrZSS1dJHx/TGyeU
y3uaa/9fzKmAv71mIq8J4DhptUB4egNRT77rwTBAnSBPdn50UGKGxNUI5tA7rHrU6poV3hgxzre6
noKK03+KSRZ2TIXv1qlZ733l/ngegMg5+z9xxpO/qtSF7JVZGDg7GpjNBaYILoa8RF5bUECzKZVI
NP9TgEd4EpCNx+tVLXvRH7Ukii7kALsJ9cbQfQ5eVB/ajoYfKZ/ziS+PqWh7C3f81FUm/gDd9ah1
5Yn7rUF4KHEmveLLELY7gXrlEDjCXVEijJZoQ0p9mKzDRP0/KO+HDeXIosccXT/xg4ZwBTezLstF
YSLbxwz/zqEycgEIp/JzRTB8cIjzjvdpvh69isYcLR4ewpISQ8iUoHmX5XMPbZWDp5+XFbcHhIzK
wMdUIF5tmOmADQQLmvetXO+6P98AOkMVshviGPzyzE0GXszY2LfGh+GiCzjytYPpRA9u8RCz9snO
nLkxvsr8uHe0dKRyMuY+spm2Ej6PDKHxbpsl9bZIyBiMTxPTioznMrZUL0nGzaFBjbu8fAa3233o
8HfQ93gw0lezPmR85wOrDafDBWWCtgK0oLFMuWKXOWuhLEt4C1c4oHo7klVqRvciUqrUEerJdDld
m+IN+Vhbiff9yLmHSRN/14PIMTthGz75GclR7Bq03oRc6FYM3zQzXc+Zue6tFSCThsBLACjkzOK7
Y/sQKTejdCJKjmawaQ/OQyKwWQXbysMW7NgAd20VHhHN06DU57Lr1zdHB+B369hiIAwHgUZOeMbM
pn1OdONxg0O7nZotywNByGvHXdiPIqhn9Yt2O2T7UToQk61h/BcuP/EixuK474YZtBLzusZmwJvZ
GjeP/Sn8XDEbME4Cudt8dTbnzpbt3k4b7vF+f6gGI78td0mlj6IAT17WAf3/QFCTBTTL7ynH2v+a
uLK10kVzR6FPzEAkIvgZ00qNZUNXofdVJaiLCF5Qhp6O5UfPrvkg9M/WrFSVC3tuMoI7uM4gZ0h6
cMSEso4SFP4mbPEYuoPe3bit6NSok7TQyaXoS75IB4U9dy2jkeiKU9LhH/yvp5OTPtTiM0CJb+8w
acfTY/PuTJDl5dYIzmQeDrNG3wsKMZq0m++8stdJtVjoZbfZQw3SKfnS7AqvtvJmw8WpraNBuxTY
dYob6ZspR5XrclKLNPrKFDBl3CMsoHuiTwGGLcudLe8yE6f+30SllCS39XAPYuJe87jGTlZEAx4E
u+w9ig/88f9xLw/pBjEM7yWpLR4F6x/22urC1yMTluaM04LzeU6Ey8usrLTzXqQJKBXnbLnFgFm1
e0cmsSBi5zRFcRMnL8BtZz4hfMe+IKORtkVDvBhjLzT/HgiPFzUCzgfE470lpP4G02eQV8wPfSBY
hYoXQ/Ugc8hKkpY8JhEOg0VElXfADlDqU8AYMhg7CY79bIoa4irg2yTElJG6YKL4X/6pzn4sLzYt
34FkvCSPrV71QGG5KxvsalGN/GlVf0yS7GrU+vwH/btem7QFgDtW7GlR0nLG8mgqH6f7e4bavtEr
9Z/7FbfRu9kxUtMcCapFy0husH+L48NwgS2IDue8iijTuMtmQd8zYExdpKRPedop/rFREEbG2lAn
qkaN3buXrDnEzJo1SC9ZCy6gVxmKO7hU7vJjlwowcvHblStcCkCDAzr6oM9rRq5JCU7tOuB8wxz3
ZlF+wFDAtHketfEO4mwq5HHMTJ0hRPMqM2po3jfW+NP2IP91MJokygcWZVX6vKDSiWu8cCSSfQN+
DdcvHlVXAqazIiqkfkdqzfJm3OYcM95Uy9gGuIVBckL1JaAMr4NCbZjn1cQhhQx2KYGP97oQJj5S
wVe7wu4pbEac0pao/fB4zVtVW2NNPJc08fwJ9iaVn6+CcucCCkA08FnOCtiGIyHApAswdvH4Liy1
AAWuVYhwxlg2S0P5bkKhFxxBYXAx6rpUcKNrubklUzUuqLfw6ojNBRHiOs3i9/5FVf1W9Nm8dSNT
BWj4I+Zgy+LhjM4KoHgQ3clq9wexXbXOmn5GT6sm+q+BwDd8iQ7Trf2y3CsCT8o6UYqmwoPcWpl6
kjJ8JYhCEVvgmZjIobEgWKOnl8iuLad0IpXyD0TxRkYHCynlY0jAUq0QveerAwVljDz/Xv052lQ7
s3ks3qmTDElsPuN2WNZNixiwdGerMsUqDaDDA34Ii5YuIty7jOONVRJa1fcuX8E2m1SRDgzCKak7
hJ7cVsEG7YxTlEukUcjo4AMKfiucA90Z9pqzwOXOy1UofzyM36ck3Nuaa7ZKeRqJPODEQIIm5lqA
PEZ9rcw2iMAJOvmrRrBmUy4zkTBZe7RPf/DL69+LSLqAydAfwQPuCrgL9PBkmO5GIhH8bk5jFtFA
oP2AnV0OKXK9II9YmEdF4onBsHFB+GFpBe2BIbNFFMAJiIXO7pQI2x5rzOwT6pJZg3ZQilWKbU/i
nU9jKVbKDEjt47gzWyfY6R/0hrJc070f0vih2BLdwvnQlmmTdNxcxAQaIST21QlveryThrhMbIeg
VKUNgPxg19qAqfiDfMMb47ExBSF6uqQdhs9R0jj50K1vDkPcZu7Bmk3WhOJsInxrUjw3U4YeILw2
mB/tSQzT7QT3e7d4jkwhNAUjvPyiR5oDWJUGV4rec9/1hxkOQHgQTRqNfmrXwDYMXqmAIMs+0u1N
LWErYhBUjuMGtg1NVXZilRiT+bMW0BkyjjTglulhxLsZFyTGq4rMfxKfXwH/8+D22ufBbsa02ZoK
ApCOisTW5ZTTqhJeiqV0lTn81fX0BbCtW7Elf2YDK9rEOUGiqXGH8Xmi+7VsqbETJaE6cWLkF6DC
QIgJ8PurEaXdka3DQGeDgHAUbJKpSKCpPP1Cq4nUzEp8jI9epj01ztY5Y+0jSMviV2c3iPIStjmS
4Cm7R5dE0d4LdO+AnOBQ6+2czkD9CFv2IXWg+HF9/ZbJqt64siMteMfFJ9yLBXHSUpGO+U0IwhVG
Bx4BQ7RKOB0+ck+khOzsCcV4ZxmRHUxxu8hcEtplkEk4RVMqkDty9rmcfUImjJ7/Mm35aJlCnfNX
tjfUTZwMOQhGmeHGPQnqY53ON7gVjmWpUOszqAxj6cb9Q724DmLSQEynvvx1osE9TnhEYNBnrsyr
Yy9M/9C1HbBdBRpvckHAHBHQ5stHrreknkMneeT1RQPrtHrJLSDpNaoh4ZcE9Y1pXvZ3jlq/mgWa
woUsGZbar9v5rUnFqKHTTY1Hk1jEO8v8k9oHQqrlkLga68Mfop95VZJ9DOfM3LTOgx+TT0yTg4YL
MXbT82ejhouOlYz3Agptoq7Qw8sWZsVcWgLbLIKlzWotbhuo5S6giExsP5M26dFliqoYxyY+6Cga
hDYM1tzQpuBWO8P9BCGcMPmsa9hpbGKNAl0cIH08AqlwZCsRVAbjtAXpZ2nrqHeAOkMvDywcfkaq
10s+oB/AfBz7V8le6n+Nw2S0Gy+u9p7NHze31aLdk/iFCZAXoVo0DEukNBhXsouEDk5kcTH8AYDK
qbk98qTdpZ+B3UHw1POj8U5fNRZCufyjiA4P1HdBu9RDE08csCvrojLzPWv+QkYEykmR6uPL4gmt
wHDAY4pMGJ9XLhdQv67AovG/tcuLBpx1jUsbWxg1G6SBGdIgpBh+ngztSHNYl3ww2kcEWH1JHNka
MuZiy/Yurs5NpNmU7qG8H9C5n3hMEaqOSykGFnp7ttovsZvRr/o5fxIyzTK5DTprOkJs3JwCRpV9
cJK1v3PoKpQOi/IjOxX85itdFBzf9p5SOQwLfoxvOKVhdzdojM5pXUDgJ9fetCi3HaOU6k/XcPh+
e0LJCB3JBT8ecOXqS3vNlrU0WPwdn/ZelHA4M61RnXKYnRzk8r2iQEJGHoFG3oSs6eZbAQ7FzjRW
ljLyZBmgiFiLSDXx5ACNbEH+z7mcUz4LcdxQqKfOY9ei+jylIVFyVCaErhTq4y0ljT+RvovXt9BL
IYvzdiPP1vPsBKGqJKfYe9dQuRMpLg3BJ77wBXRiTqsPfHTT9GIOaR2igwIsU1J9oHL8/bUS/Cpy
cuk5dkLa5/T2zk4AYUMSVy1JG0sosJtda0q/qmPi/XWsNdIrGIUZeNjPwI5+4vrUCU6cM91V/TBk
tKgyyr3jm8Co1ehEGa0yZVy9JtCJpbiag/jqlwtzUNbIUQuQLjRauFHsxwYjAdfAx/mq7fmmxJlP
Ff2lWwk+rId1Ey2/t+k3QvkjH3Dm5AQoBfJUMIZ+cuC2HCdvyssjWCKOSTEGqOGM79x9c7dRgDNb
ydsBuP2RAgk8Zr1r5a98h+2K6FtyA1FshwmQ+Qky2NxByt9eQ7sNHEzsP171JkP3sBLHHhr7rxPr
+qz9Be+gt4xgfTl/fBoyZAln1i5GZJq9Mtf7hPV6Bv94jWXurFx7UTrkrczPDx9164GDyBe2tvDW
ZcRyEquM+wzF59mXOFOpAl92/FY3J5z8bGAglBtjwbgEQyhfPtf8VbXpw9SgAiOzlYsFXLeptT1y
jIKct2iwSFIhFt1g6RKJxYvASvpmPYec3qXEHM31X2syaonJzTuxcbwbegoXjp+K34LI8WTNTRj0
8uxOUPnSQ2QMyoXZ0vKRs4BWmhoXBMYG+ItFCntoEMJtfx/mtxYxWf+gIC3d45ZjlvgWPKKxYDJ/
Gv5bGXZ415Xe36PFSVz4Pf6/GWYGWN/ekt2eVfU8kdUzaPJCAWXUXy3MLQC3PFau886zPkdpFLRP
hbdxFO+2KoIFFl3pXo6xzOxg0xXdrCogI8JZF2r7r7qcw589VULW06P04V7r8XydsXTnX/tqIp4T
uR7QW/Xtt7vGJZ6k73vSiLDbgCD2DMBG3WY1OtXodzYn/N3C4QdNvjn/EOfgssY3K/DkzXBiveqH
YGZudXvzZiUuRxUuZ37qbSbKviIfCe3CL7IcI+WcqIpo/G6U12i+LC/LMiExIOy8/Ws344WJ0lD4
KX3AIUa9Hyomls6w29PZbEGAxXUGDCQh95HIS4waRc+b1kTqspR12nZjUpUWRycQuMv9BRhntSVV
XE/rBU/+RtS+prEvL9DjaAzjt3qC4BYPJBJ2mZ1mZqn1ursjcvpCOaV7kM1D02bjkdmYBZjiPNje
8KuOX6z8XWkufRWtrstUEur1fuBfUZuV3hJQuChGi9sYxEm4H8m7lvrp9q81xf4BPKoLiYYRqJt/
JE3JsNVHQNX0KE/46ftRYG3JitGZJQb8tBoP6OYCnrLd9Otv+gSonQQsoDeNJMjVMP3S+P7H/7W2
hh4k+HSyXJJhFv7lPp4XdqzphHZxfkgYSpE9fXWK0SZhYdmP2x+ixZxtRurrzm+MKcvl/9T80U+Q
sVn5Zvzpviw8jP1xg/4DUj7ZiYN830M9aQuZPuge1fjq3eFet3GY6dUHgiUhRO75PMubTOMwRH6L
LVLoYG2ta9y6S54wFTg2PF14AXYEkH6ceWiqLcsXp4gvIt5vZ5TDzIxzNwa5sLgYl1SoIQHJf+ZE
Rc+qkQrshhAebcWZDKBeW0iqYXJNyfs0ztbh/AuplWkOIV9mRa0QKEaWMCGtY9mCzedSSxhqv8XG
REoIVVYc4G/GGQsYhui5Zy7cc8iVqJZh26fONYxywT0VXAInTyjqa7zBYN91/rZ0HNiR5CtwTma9
nnrZApTZ+evU3vXauzRygyWmeVO7isLC0zt3GhG8EoKQOWELsg9/szkD2TQWQTYLCKmqGFuuTT9O
Msq3k0upyfyYQf954FZK7Mmsx8TB0s+3wc2y96LwOXu4SBCRQKIN6WIyIo00pJdzeut34Nq/zo5q
xOgB8ybsK426jT33nwU1sDNkp2xsfncEEO3r9XEwdwpJF/SWMOf2g0KdB6FF/uUt0G+Sx6khrBjn
TVvK6aVDPdFzzAxnR6YPFJiRteO+m17C18hCm/TnvSo5uxAn9kLvLQcdyz/pWTjdGQtuYnsslglF
b0ZDejam0ay1hrDqckCoEX3T8w0GFOPJe70vwJXS0gAJStUZM8GX4zZ0+y/8SkM5EXAXanwybMei
rzb2ulV50mS/NJ36kre3WN3+Okxq4womsNhSIAQTAJ2b06EsFcWbVn4p0zc6HO3alVi8nw03DNad
qA/xoHZ6wTQB17AfiMBx8eAd/G2jroJsX3RO4GquyepbdkvrIBF24AvlMuI/pRso2qLg/oiPCKRj
cqtW4cWa5aKvPPozlwTFHltblaVHIc3eO3TdWSKMXSIQY2NwGUjqG0qoGMYm0Mf8Exa9gUZz5B1u
OvDGvfTXuJ3n2RkUrnwXws5RYMFYuESo0PZB1Ae56+9hOaAYaB+X6Ti8Yte0fSbNId/0StWpxXOy
5w9mWJyOoYhO+JO1Gw2IPOmuA+FokFUB/QzHO3DuXKEKU0+iF8eK4egNnX8ITyLgnZhpMnGRMII8
hXvY7b0hKxSCVEfQ6XVkQCxK+88DptbS6dQkuL7chkJEjpDpOwPqRoA7QakWvXKVSkqgjMMkLENq
PPiU+hTzhnw2aNXKL9CMguArRtjbbzP6GqKbAfOkx2m4UyTBfsio4m1Va46uJ8eVx2PbmLrka/ZY
DS5Nj8NP7pKmkwmF3ZxUuy3TDqucAPzFo6AS9ead0DPvawDsQu8dK/oVWmWsE8D6u58ufqS/O6PG
mfitV3C129wyS7VKSZy3S5RryRhuUF4khYZHmsADTN6/NcivkYViFoTXhfxa4k/QLpLBWzcLpY7z
sj3L/vQOydEJza4JaJqKF+ebKhM18AxtIU8lXEethd4PfOUr7YXH7Voc3wOyURXMOrjthu83ZZom
F7vMzNYnNUZdhP+scOBkrSF3qiRpH/Dy2EHQ/v9iYoXiBgEHcEnq39XJJ8N95DHuMia4qIOhMTnw
7mHGoAPNbM+dVSQFo0ZtKZfPEhNVYQrjmddFvjK2WEqsKsDbVQ3ybi3iTwwtsWBXVHra/+1grVTK
8+Jy4NKwRd0avwx761G9XBjh1f3FtvTLDwgDCwHG5otQWTxVQXyVcOldwEbKGvGqTlUq20JeoIDs
USa8KTQCWiblajnTaem8bwzV8K3uXq4MzvHSh1xMJSTCRekQkM2hEeqSRVq1j1wn2a6igNxGTImE
J3NuXThz85DwNPNCn48VN63m1sjnhM1rcUqND+Px/XPcVzaQiN4QjC85UGQ0rQO7Vj9kQeJjVUIh
qF9pDRMuK/q1mLJjXy/L0ddfXbDweR+z8a2+8J/cy/c1c8vqx5tJyEu5fidrw4NltXrgz5h5mAFC
VmPLyiN4M6NszC/+VTgkjTJhZRELv2vEWGu6hr6EsAwifukAO0cCorGAyFeB0FbNRUiMxkW2pvIO
8jBmcUocd1WtEwuZEVZAt3DuNLTrSBRCbs1/Hg1v6HdgIxxafMhgweFy/7CfWAur044lNDE0Vlh9
zSbfRbeaCHjHdhXtRLJPUI/vf+2EyCXDPTJPaD4nwKwcogmZcCqTIBJGCyg4Cf6PNlxizkYS0BxM
lb83C+5sQ49/WL2x9AGNPpY3bu1uZzLqVIcEw58s4c6BbocPEPzmVCpWKAoO8YtSKgaoZxE76EeX
e9oAOGXiw877gAa3n8llGHr0PYhmPNw+tvIM8w7eyC+rjoVzBETEmanIlssTNle0JKPcxqg30Ige
bPyur+pm6ZrUf3BG9JG6FYfWO/njEWQvWYHUOXjjNrJsqwKdumrE7809NY8ggDBABRXM5p5U3rXv
VkgkcRLmt+27E/t6Gf+t6gC1mWm20vYspibs4rZu3dfbqoP38efGHGORDDf9xa5FLklmEMFDOjqv
DtrWT9F126+2NCySeP4UcDfp96zrdEMwvdnDaoW55V2Da7VXMulYysBSggWrnj96qoefIG7Ut0Rj
DmUl6xQ+ltRhx0wAnDH+1yzXgXnB7hXJ7dRtHnxkMFJN3AFhiNc9LdQZgTIQDxzRSajJMR+hkRm4
S4gCntI9a2CA43xrSeqnpCtnya8i0TTfJekBfC2HKci1llpdXiB2q3st0ATNkFo2sWg5iYCmva/n
swkoiXoQUSpOWCnpmaRvHyxEmQNLF+9xogEHqycxMT/Y6BZ9N26AHXQ59eac6anJm2ZxiYTyLq8A
wLYqrvjuTy18sdR/k4rybkVX2GzxsyksaAo/ZQACTDRGPGPXkKSBx20xp8WAUmf96cxetI8pvdVe
ODMi+IFUg+Af3wPU7gDdcr0gZcaWripicKQbhxpuiOWnCNoF13eSPDvUh6HX77LiU0qo6uPPt7oz
x2A405oaSAJueAvBaeJ+ti/Ih0WvNCgL9DmF8LZTdcn1AmBvundwdTiH3Zref2kYW3sZXSP6y58p
TcIRUvdq6im8lPLCh0JOU6+EADYH9QIK8JcWk0XGX8xZ7YddtFXpT7D4TSn/D2u8+SWgBOOPs0ls
7rXz7I8g3P2qJGnmg6XjunPF0NIYjU2qY+bCfAdzcWOc68q7IFnwKVY4plyJHGtJEDTR2853ylri
cW0wfwLlf1RB3cb/MDHZtvHypw50YKGSrMeajUpwolgRGb5R/X1sHxycRL8dmBobILDCQ4gq0D9c
ShmtOOYLgF0oIpaHt1qamhnkukNWdyBKigIfmDibmCK1v52AnH2p83tFvqsS040qqgp3B5BvWQGX
B2kCm0h0m6H87DYWmxTNZ8mBDpuAlO3PgNIIaIGkTtGii19hSrIJvLc5VnKVeVubDTkjjJ3dMcDD
fWtqohrfvY96bjTDABAUrvFLq/S+uSCujY24l+emHeFvJI6xD2I0EBCcRvbgMwiZPC+623LqJzwq
ZnSJdh0BDLfxqIIH4k7wj8nH5zAnpCC2oD1WcO+tMlo9Yil5o2rjqLGAZMGIa+ypQpqIFUKnGItk
QI3pNpIPq97si5NFJrR+wggydibU9ewI66dc+HunWrFg38DssGLgBCsvzrts2MVpiY/S6Tdh7AuN
nnx1pEH14WhY/gE5iMXv2FCoaRxeSwKlJO/hBXqBsjffvHam1r0JahENAP8acvBRs/pGogaDCQcH
U0usOEURKBl3yBAVl5I51n34cjEdzBZn3eXaV25Jt/ZBSkUNj8eMdOft2LS2pT5Voe5Sw8Q5+x9h
rq+orCHl7MDKsN1GEK2PRgod8bGizkA+uIS1z4nIWkDP44t0t99h2WChqnYw89fgLRmIwg4fnS6A
Bb4LOePhrpWn5xg5eymG0wiGofDPa4zuaIA+HIXWgFfHG3bQOoQmVe6rgC3s8UAPVAush2cZ6iyH
L1PlAl/3Jx7UptKDNO7caCzatBWTxbRaHGU+KEnLBr3BBSFwMgV+1D05v9tNM5uhF3I5Ial8dLKd
Mw/9yfmrEtqSqhf/MBAqPxrBtjqBToHzS2T1mzfhgRzchLb9vFYrDybq+S2wAfrSe+E5ew5Ya48D
q6SL2qbsDjANG9+9UeZ3RSCWn5pssJs9Ynv/JgKZef+WdVpmUwESTrY4ypeojuwzfca6TQEfwhrU
Yg7YdrXClU5IJRkLnGmT8BvnFeKtYUyNiKr/wimU+J7EWgCu4MdFDacinyPWC2qxcxKDEh63X0jk
yjVUnv11CnfNoh9e5uqEq3WMQ6ju8N5UiZm/L0w7UCkwg5mjmT4wYYKRcKpdapfWLH5EeBu9cPtP
qyXmxYm3fU3aZ3iGWl6SmS4tMaX0+fV5L45AytA9Y1p4pCdwPshGODCTzg0mX5rrr/IXyqo0Y3Fb
JaFHfHB6kRWkAeQDWISUAgj/aPvbolMbwHwPIS79Hila8QM1dpyXhAFXwYwg4oRH7T7FTaeYHUza
+lN9eGHh89y6LieMyFn6I0xmzvGEGRCD5h0zWUeTf1dsnFIQFLPgOqDyOrc1H6zlZLDBKR5ucgel
VHHZdzr2BbOqvRFJk/3LR+iekj53AGz7JD0yly90b8pBSE1maASj5/5npipKl/Y6XcSgft0PfIqU
ovqIKAHc9xBsRA6vvYyV7ec3dVP1jg9oYmf0pUB6S5k1dGKAQyA3C55rsqaf0jc36KIy6jgQIHsr
dnyIWK6nTMqMmyElUPByMoQA7uxbg/nSCZ/HxXDC1AXmGCjwwCCfw51ABN6XftAkXR90+N1TA6f/
zbL0aWMkmBl6Pl3jmfdLKXVVEykF8Yhv7k12a48QDrKbPBpMNO7WVhBLbyZsr1/9T4KJzX9gFrcj
eT7FSNWiUs9PJCc5IZH1TotuEHyX10ShawA3LqMi+vaCGO1UcShiyi2wND9cqG4Ac7h7fHEzqYxZ
eiB7fUhNp2dkux0J2Slp9av8vHju+I5i8N7crr8QLnoaYtuz2g92kV/2HiD+pnPx1XEiPmCTfLqj
ZLAkzl06J0njv3b0uXpJ5DGoYzRY+5n9SUemwK08t6/T9/cs4orlBHBTJRGtI/MR0Qbkk3kbWXmZ
glkPXUZrk/QK7pi4x9fhxVwxG6YVdsKlnI48/c5AEUSs0qcR7E8s1CUPK6m5eTaTACz1MoR9QPl9
C8UL2Uu60yJg43oV9cN8cy9HhjZAsj9TcxSL7Pt8PV3GLnalf/GpCRU+Eqx3oH6jfvAqVNtHumGH
ruAyOnyvajsuMMYjb/Q9ySxP2XKEVaDpQy05qLxv3ngw1CAkcbDjhOFYr4XK5S8R802C/KC4btBi
nccAtUneaznxWjbIQ04WyYIOzBz7XdO16zNSXN4gXBVFTap2aGGRl1Wx/qy2o/ZvKTyiUuaJafHw
qEr3TK9B5YkbHAeVfAIQ+rXg0qqbMbO4vtJlUFoP8xp1cjt+Uo1guZ/cExFDvkL8jSz/kZWefdPj
LFXA193Ta11XCJz0aStMSaD2PCsoHVykTwHhMg7AdvMc1//zRHPe0Z3OGEwYs5lCh7I0rdyBzGGN
fj9m5tLnk03CuYYFk60hFOHISyOLGWkfYQED/0cehOJYxSP2Z6NyUSGV4RVO+haw6rD7Vyg07P5+
Qyxuj3Yl7AO0MjJA6GrH1JusaIaYW2l7M1qfT0yM28ATYnsgLiqpb8K0DMpXLPEJELKuKYg9yUQJ
CSiPgUrKsvuECDKwywQbeKGKZgDLGvkBIheIPzjtAYrPnTbw7KGLuE08rZHEN22tLvs3cs4MQFi0
7cwfIi591n0JhgW/gUWtgh95cvlXI7jzSlc0tt42eg4VX8ff/QGESA/Roamp7zG8x/waQoBHVze4
bcu2m1/iaQfQyWI7XxylGpxZz1LAr0/L/7dkdJGj1Chl7nAw5V+JSKRwdV54mVfQ75LMuBSW4E7E
UrVK71oc42kRUngA55DcxDOFOMphNMZBBO9ZmnzweAKg68eyxKhWjY/BZW2JoGCBHk/TBh9wZ2Qy
BhZ5nn5bfj4poSjstrnNKshzY3uA3Nw25cCCG19rHMfFYgTzqRdQVtmV/Nv4NrdnwFtjnW9ZAVrD
IrY8IM3iniEr6E99rg0Pb5vRLZVSve380rQwuX6K13QbLjghZ/ZJVcJPGA4aNIKpe4uCUIiBRX8s
VG2PKUc09AaozhXDNocGjyPW6r/oc9L1nGrNLS4ylyKGbFa/tb7tax91uHVUcSkNvKFZfKkFSlCR
mBtTSIUSaUgq3Hha/b4QimTMmnCuWuwCHS/piw8FcUkuryspt2Vd2dkMzvHVO/mIrx+q85Qlwacs
VA5EqPpqti4akwOAU6uVVY2JuHXNL/+ODGHAVPpX5pODp5yertBlSkIHyxPqtDv7xHWDljlgBM5B
QOvddqL12N838LKq8epZuSdeNrH0/zrNRz5KBZszGtfsYJ76dDk9mGczHhcmwS7r6a+03cKGZ/PT
VyzKpO65nZyDADIbhEpTzaWwkbNmPE88GocguVNs1NNItw4HHXlfYLVD4LQc5dnGkMvqIbVe4Cf6
lor+Y1ghsqfmK59FG6SxLm3146lDYLvAVFmWkihkLhMoMCyX6Yp4MRqpAqo4mdeYzb9v3dNls4VK
ci8zfVS3Mo8vjBppumGmgir0BkbwVfkAN0wgGRP5u4mnDLtKlhgTw8LSxTzlqOYlQrwIdyIP/8oB
YrcbaSKrs719uKUCY9Xc5EcLUmEzNgjb+oF78YxjnppkxY8m1bofxr4mOCv9uiHaODjda1AiM81x
Wellf2/JS8wQYKMvgaEru8mtN4dR79qg8RyBxO7UEJB62g9ruJFR9pwZF7z2P7ghiP+XBoks5daa
T1G7N7OWC9SrelxYzAaLmuJghPPaW4+5lrCxK6jpDplHq5P9BjT1rjs5v+Nj71WzqCq1B9AfndFY
L9ORSpSKYP/nWn+jmyKMP+OfRTwqFsq035Ycl0bMa6JARbcQW0R5T8Mq9CFM6vPryq6czP3ne0FC
SrnbkG4Jz+PPpB1kxk2maiN0gKZOWbowQK6Fk5hUoiEpTumzrs06iZVyDle6AWuDJn1keFjpAiOu
9PoFWWDwP57Sukgg6wCNCbnfu/DZvUAYpbJxPVlV/nrdIKcLRStx3o4sSp9nqH3Z/ZwbV+dqcfIR
jN2mq2k4SC+1tfsR0EzcR2S2wedP+0mFganbtmnnY+i62vZwt2F+Px6h9Ww/UP4zII+XWzl9w9P+
24Fi8afBfKjagyG85CzM1ZSuOVTxT46O3KgP0hj1tguvdRDjOmlifDokJybuh0JWPIi2DOSMe4er
pe2rWYGp2pAm1biaAEvF4QsoWFfF/HAAnY2q8lyEnoh95rZDCxot/fMGqnx9oPRtfpnPv7E35sic
eFpA0Hf/j3czRDCUlIf7ev2gf6hBfmXoHXjRMeWfhycT1GxIlA0z+thrghAJZemoDNJyWSa3NQqR
GdzBnXIQAdhiehd3cPeeBRsmtPBsJTCrOaNh90+ZTfQPXVtsk+O9emrbVvJAsfSN1up0IsKxDUmz
FlsIRFC890x3JvojUYp41XTD6FuADmBvdYEOE3BIEEdwaj+zkqSghfnQjHcPI7JQM9ht9W9fvou4
UXXC34eAUt5Rqi9j05Zvv8xC0ZKOQn+580+ZdX+t7JB4+hC428lAw+SHrGCNczJC+R4Ue31tVH9w
BHFSR9uVkUul/HVZSi8pevw5tBqHWa8LFw8RZmqFVXpyqpETbpWVzv2WmANOl0g5aHIhTQ77VwEH
tJER5d/HaZAMW8JYgI4XjOe37jAeA4V3+Bj23hUOJvEBIqqBm7SgmPq1G1bZFCQL/7oN/40OY5Qf
U7LL+3gBKy+Mpv63agwiCt8iqwoxm3MQSwKlFnqN/6gbG4ojRlVwFAdgQYnkIIDxgRJDhG1GAoTd
0i8TpCf5e/tflr/DWEKRjDCfd4Ldhv7gLh3h3V316vqIJVeIuLYNPy8hc1Za6LdSXmmjqyGJSlsk
XTMQLxaTaRNHENzbiU0j8KnTBHJQnjYOftmO+Sbbxlb9BFrzaLIffjnRFrwU8WulQx71prGZKGCK
Q6X/dLvJbM8htaSJpi2k+CH78cAU346E1l6HtjTM9rtc6DbfHGOsF3yhEdiKbQE4FwzZF++f/zBD
t7G56vHI2O3ugZtBEHJh7A0vZFPe+fvhBPM8SbyAYhmvIDKCI9EzaufJmDqmKJkrO31vvuXVr+zm
h/H3wfDzsH6JaE6882xwfhyUDdpkzfaO4sRGV9x6KjUcuDvh0QSZiLQ0X5LZ44QGskugXtdo0PKG
vAF2aL2hG3N2jLvd0FBg0GuRfvPoXPDOL2bH4QEnJt12+VBCGmjiqSlYzKkr9zWhVM757R0MhfDH
i5eBvf5hnnCjUoYf7XBHYPaHCJiq446djXpe8GEbR2XErn2EkydBE8kQU3kjpdSdGoGOW3fjGxJx
PCifqJnOnQRezp6l0MM3nD89uDyHaSqUQZjscsmjTMQBihhyZrYm0JOTCupMT0/6oJIv5+wumS+k
q+H+PCOPPxDjSkuWY8uesAvixGWkQf80a1mG9+LlEWzB9lZITINoxy8Wdfg86sKQe8uv03l0Ou07
c6E6OgmEawRaTsNkElvCPXKamCsS5nk1QWUWJQSEuFluCfNz2lTVb/7WWgnlPxLruSiyBdfuJwuI
gTwc+mysN9hZ/Fdm7u4MZpDyQxFrQ51m/buK2ogo6qydnym8/Bda6x0SwAz/h7knmEuMtybo943/
VFvszqkBark2ljGH1uwU4VitCSKH7O2WZwzm+H1D+kuVvK5cjhGP4fdZSY66QBKkgTUThQqYRvdW
n29bM0/ONUt4dXFt5H/oEc/AW+RUcBG6du8q8Du1Pxa6+rD8M17SsBVlGY+dcEQ3412rQVLePy9T
cQvUQVF0DISH9GMB5zgSpQZWofAWId6HcgrFSjLIolHMk9wIY9povDrTLYhE/eYshSJIt8SV7mGz
3/7fNi4ubpJYm/QB7XQ4h4L9OJpWl9QUAXf3yZYGwLp3PVrqZ8LeHYB2OMM4IxX6efCH+wFVLU9Q
cJPIy/UY9bz7gzFwBkcYfGO/tLQj1pEa4z6vYYVvUPh9s30slnYYaqLAK34MBSAjl7dWnLj6vCxP
XgcCbnv8Vx/cGLJsTvxbY28PGCUBuabGPijuzw/WuD3cKPO5oWMEQjoUy1DgGALX5MSm9Oblgko+
Y/nq4EKhufDbtKs/kjXE4uQjCctH1ukndZbITay5/HM1s6WwcwUcCspaUWpeCXbA7ht0dRWBDPls
bGFKdta5oiPBfvqaKiMkJD1SQBEdCIJ1BRcs2Rsg5i0QhCJ56DESP8UhbqfkMqX5Y5PLNZn3Dk4n
9bz/FhWmElLZWfTvdMOLGfWJJW6oBkamU65slvgpoU/v1VzQAv5vsR+er+9Qt0bJNjdTlMlmkdFd
AuY11za2fkxMwBYxqO59Y3YoQjuMD9AITsxhwYcQFMO/J+nUwlhjFPa3eA4ZV2yHt+lYCEMVUUFZ
k1sqrSUhLykRRmpRkDNahXzsfI0bj0HBqVkyLmVHRP9bTLdU4THd45b2lFRSdFHVrmKUq+k4w8/P
9r1+kwBqYjeZKHdqu4UQvg5sa822QcmR/I7zY/8TIJHLGwnnaqc6IlasvzCsqtOD34Dg+LbzyTBD
VDqdjYeR+LNbb6rcdXCToaEe2FAm7HrlTr/XZe7tiMIfk4h2iLP/QZ+kCcFlhgmIttXEHp35k2tH
5HmE9HvH8YDou5FI0OK38dldIppop1NWFlo0E5ZI1Vg/Xso8WnXT7VWiDL5I7GJanFqg5qoNNTWW
A9BulDHsbkKpMUwTRWcdXNh1Lhe8Uhn9R8MnqpBBJj8q8hKwATfs0cickOSFGyN4mLcIGvuF8UfJ
Pjv2G3KnaqYpFGr2FMveOfhIemIHrGag1QxNzmA9NyoYivjHkAlq5/z/cjCk9Sicpsuhikek5TtD
VQ6pBTxROFEHZ1AGPEwJBvsHTB0dEgvRXp2tcyEEiH/Pzi+EaCk+e1ZzS9IrZvAYa1rOK7W6p+Gb
fI0OMhtWyMAb2chdLKUP/+i4piouCm4dwCLGH99qhpBlff7/nbm7BCDDhYeKBmRErD4Om1MrtzhZ
vGtlE2jggm+juSJCF1eP2VuoQqCf3s1N1rQxenKyv8k8xQU+xgNHENZoCPVoxeCSh2H2+gOM4owh
lGAP0+IccU35k5OX0lKHkOt+yuVVzLcg3iHERclCo7QQXslBGY9LKKmZ3lt2b3SaUbQB1f9LkQ5p
hM6ofKOg0mYTJZzwejlb0FhLeeq7Shlm3lfTGsQbwkKdTttqmevojq3Y/vRL2fRdvW5D8Ce1olr4
UIsKRGQp+Q7DXf4EFKL1iuQWA/b6R+kaM9djerF52AYag3ZvKRtNKfOINnfXRxCo4h8ZrwdWjWRQ
obNn/+Xmabyus5xfSgX2zZ7Kn637LrXhkdKmBp9g5SetFuzGSt9FIAys9VB2rCB9exinA3c6TRjl
NUdvtzIC+u/JaZ23ovz0U64mtIsSMQo/b17DfuitF1PHFu+tBkYkRq02ZQ9PdATm9kMwnuKtlQb+
0u6lo3zCh/AkT22YYixSKHdyhUQzaEjtMdCwkJmv7hWiBsdu95SX9qNv6iR5U+OAbKTudZNeuP2+
HFdqn5fHawEtSuVQH7cVZV9ZsyoaSr0YQabeAogAcqtyfBzxoFj9wF6qKDAlP5kAVepJ88ADd9zu
dswwPr7MeK7d+nRCh5SrYn8P72QqvriztKcHZ7OTEw+ZknABZybHUw6UYW4LaKoTD3A7yUFTpH1R
J18Cth2Q3EVrWdkGs37zA92au14cetUZbl1O/HG8ma2odBZrE3WkyPM78mjZrZUDgIvQ3JktWarm
dAl8VdIu3K/kEQMx/Wxaoisa29dCvLIXX/mqOJwANEGqZCwCC8IURI/G4f6Ga5QehgwaecI3gpze
wgBkwJiafmVMp0bFEVD+BCbON4rVUmlBuwJ8jLUVy8/oSCK5Rvi+qMJXUVCFHxKCBazjLKb34pfz
xltW9O59zWCJmXPdiwLjCQ+1tEIA0IsCceFdTMuB9phMUHIy3Y0eYixzDCbrY8OGeqZi5M7LnUP1
LdMG1616u1JzBGGe2NtOVuA0sNqBSbu+b1XGivrURt1xOZL18eJfoA/hVCR5tPuYUGzPL8VZ34Do
48E6diC9OEJvWJRegEmvL4Jmwj/strgc+vnZ8imWEqq3Tk4QSSunrzAObpJhlQR194IedrC1yY0T
b5C+JC71lKEMZihwyYXBeJb/k4j6/KqCndy/qRXj7BzaL6vPR0gudWv3LncyTKJUozcBaOBfu83I
n4Q0hb41sIyuUMhhGHlOFAQPlJOfspDobO9uN26KxwUt3OULCffNUtmNdk39dcCGYnctKWRwWLcN
y7hzjOvG0fhi5/5oIAsEVwN3vCUkaPrxfeBlbmSImstnjJ7+MVcGCZ0CpO2AGRoi0be/VGu2ZKCT
DRXf9hgMmVB1dfkDmnq8sJc0o3Rwl3GAyokggRunxASL0WIdFrbUH2QCNMvTKECeUaHyeNeUIR06
dqXwF7NSsvGB+qWGcpdg5ZRvPrjZslP5IbozdFmMhcuXnSuqwuNkrQS0pEpK4pTb8sxkIdjQ1S0+
uFyNE/YcHOI6yWtqgsxKngunKvlOc/NKaN4Kuyd0GRnJhrchQadMu7qccTN4+pozxsEgfPScb4QB
kATutypNgfZMJ5aKacIc0uLsen651rK/acsy9StAuJg8KDPXkCIOHyAczdu/igadLYnZ/OroNhQS
pIEVmEw2lz0K8CQXFsZvQK6bfnXYAZsyKTXiw4RevZBeTKp224TBBgf0dgE0X8vdoQrXn5XiNj+c
zDSElZoSG1qE/ikN2D+SsIm6CZlSs+VRXK+sjMCC/5JRHNNT+hJrk3/vKihKM0Y2gQXQmH4wYZTR
xpDt9FmiY6pYWEmRuMe4ugge5rsDx6EYoiQPQUtDJNHGasgRC3vahlVHiF/q4BtSRhRu07VwHJze
wfT8DpU6o26YXmmDStFnPgRcAFn3egNiIdwZUCo5TZY0KOTFMFvJBk8SmG9XkQNv6yt0E8W8DtIo
i+xBGIsFfG6cWg6BDc99YPz9/Vc7depSw/uzRCjlgy/r+C1/w2C5lgq6UND4HPJfsSJB0b2xpYqA
ZivpdCOQRvvW3s/sHF2wlLVOJ3YiJ0sT5Z8Cr0m+7lLKEUrhlqxH0KXnh7lbXwixsPlueA+aMFav
aJvcTmR9JFpO4/t6QTylJlQMyxEGj2xGM4RYxwpCSv2GW7rONwPKGzMynlDU98k93EXtZNpODb9v
xqHkIuuk21RNWdCjxLa9A0mENhorDOM4FMxtgZGqwKWaR7N0QNAnHGlp7V0MaqBJXjQH5P0WJ32w
n/4Axet1OA5ZiTZofi5z/O0eSXxpNrcPL3uKgNWd5rWFofM3BF5mzeJv5JQoWj2hZ9alFg/B4oDc
DubtOAnoApWbOeMZSFPlvHsCdQh27dZKhkziPZCK/4btsxhNqA74ddPmskv+zvr8cKjPhIMfNsrO
GM/mNg8Qb0D6WJIGGVtn3FTx3nPVz5ZQ/m22xLkGdnRJ+oRfzWY2dqCGAVWX14v95zjJjXfEoFvj
laGb7TIKSU/ESbAVXu8d4nYG+wYEax+2lzsTKGqdtt4Rd2xGrwXDBmDqIERPr0uwjhHFJLFbuzpk
qk5CtAI+fqxJ0obxKmtO9Rs9ahI4ce6+rB5Ta5Q0qcijizHtMnW2s5gmJA6frKMwVAlUHaS4Q+TX
mfzyXQBX4i6Ry+z8tHuSopbPnLdAC84y2QmU7vvt7bDMQskt1aa693VWT9isMoKf1F98K0mvMzip
77I/frUgSB1XeNwqqVABj2g7vz8EaFtC4AfgChPsx5Cv8uLTpyaJ8ZD/fcgi9qNTrHlOWhVZlm+R
p5USEVjD+uEbIUnSZnZ0HOaEkYUMTPzUoRFDne2gYbAW4/4RVGMdL9WnXPIKVIFOV7j07CI8NM7o
vClrgNQvHK7nJFmpG9xJy0eIPI0GmdJQ5kxRmOoA6v5jErH/8lDnK72KBb5ScXcJb+v+lRteoGEY
OvNgTf4bZQFtH1dbKLGEAVPP4PZuAQE0Wo52C6KGazMn8IizdsMw0T6MOpyN8cx4l8AEL4sgbPwT
Jh+vObbysCuIaIyJbmHYBWydjD8P3/RGO9qJ/g+/rti/DJIWayO1gPZ8HYg7WyoU/ibnYLRHqovf
TKTiIxp9U/qw2v1oNFJralslCRjFsygXRYNjgfJ4KReEMBnL+tEM9ZmBwKDFIrWsLvaT6FUOlep5
h1oSrCU5/nwbRTSfZk0dtk+TqYeAMkpuLlvOHp3g/5PNBPRV6Mj3ZPOLyLOVpNmMzpo1L69DXGkW
Av69KMoMe7Oy/NudxXPZb1sBa3P9Zbr9WjWh2p3IBnsPBFd9VLZlcxBm/EikmV4ltrMguFnreIjq
Nn3umPy2GA3oNLKFGnoIqH+f3qOQXYCD7n7V7xK29nGtLsQcGBQiWkaXY3TzfHos/9wa8DMyUJJy
AfGp6TSBVpx8UCNDVU9L4FWlvClmtp/bw/Ev+/rCS9KBz4FVvtcNwi/HvFqYFIbBQhXRLlx2FxG7
GF5iecDcGjtAoM3GT//5VzqaUljv5okv7mQan05vqBv8sKe8puwlnQ/yvzXQf6yCKfwOlYZ/7KQZ
9TWe1gQpJFUDHC9L6zItIIrIWVv1s0yfHnhs/n40lODWQw2gQTp7ekfXJ1olVp+kB9IPKOexFOT+
EfkMR9fCxCegUTF156yGmeWmLOEcGFvtNgftpNfTdSu0impugQPJRmgxsZc4NGanHeOeRY9ONx21
MV4q8wBRd6uyQsB30GrZJmD6y40jIzRRhKapoPvSelBD/raODj0SDekBBjAAI85RwCpxn5wt5dN2
/wnTZqNRi0cUCTrY2raD5VUJ9jYdCjWrEtNnyhqGefaYi/Q95Txgmpm3kS2orLGL66MRHSm2TYHo
tqomcReEWTn04JLP9o5tMJdS6sgXxg+Bnrj7uLMZ9gNpOip8Kp39jaOT8337w6Vt4Y1jYfWzpPqM
969W0J3dIjCx5/iuOSVR3O8sqlTG/0PV9ZzPGdHbvQ/SFHO9PZZV7adw4hrPGJi7C4MQTTjYckrR
YQnQVv1zSUF382qr1EeAr4Frg1SEKQrnmdDlfYILu3ayQFWePBYmoYI7D4VOVXGB1Kp7qQ8Be85o
Z2uSO9yCZUN0hX/C3GvDc7Hs3ik3WZKuSWZaSlBAR+TuOVVIbtrW0cweHEkAaXi+oUjG1ulg3SA+
wLcCD8uH5qiQ6DHTRzc2ff2XOCzWl+Wx9h5ON+/WUqBiEzEJGHIA+f6nN+i1zyxlIxFxmgck1oR2
q/Dv5P/mNQPwbETwkV57/XE+2YxJqmSZe10XZGMmxCr9oKenBgfJquLew+MS2wWnKCC6aG3oEN69
yHnO+RBvFSLso2e3SskeGTdzRdsLPITvYlGcuW2Dp5kpN6xB9zVafjxiDe5tIPuxUv6Pum8jADLL
eLY2MaqkLhsr5NvoT20NJCyjL3ApZtpgWp1Mp5UMDnI8X41kZsqh/rMfHbX+0YkcgexkZ7CiwNIj
AVpInsZG39atVX3pDaj6la173R84+93jEtIiPCyF6iSZgQUWxO1KL8MiQB1PW5XYhgqmViMlNKyj
UvJWF9wAS74B+WZRsLLfOQlv7tlMz8fCtZxOm0E4ArPaKfze5o7B3MvcyXU/mQWKScr+pMhXLP54
9q/pqeQfzms5y6+/LPeYB8HY7p555ew3TeTYBjNMKoB44r/9SypsKQuMHvYBybQfB/Rbxcv1XLMS
CTPlFemt1kw1l6A+2kySoFartdzKpyPZrvAvBdgGrFSD2U4Pv6mt5qX0nyUaRXgMQvvz0wpTkTaY
GT+8DPQ3SGfu/gdO/s4w5u0yIcnEFvnWaQIDaFgjpUOwbzTsDNSQ7SJVSjEPGdBELnna9o5+MOUC
DSTPl8eXnIjlSa0uAZRLBKWpRKk/DyBTXojTRYLr8nG+4nK+jdBheHGLMP4Vk8iVOpCwxkIIE4/V
EMRJM5tdKDwh2ufNKvh2KY08BHL8tUQOYdLRgZIFwlJd9IgAj1A7kB9bzwAfWXoguCuw7aF/jHS4
23MNi/1S5HhStonFoSuu5cNKDOA8bXlGaj9fP8MP+X60pFFceeyRSosZXacFBoFyvaxULAoaNLVi
fLjbWNdcGNs+sS4dD77fePCZxihTmHGmu7fLRWHBsNIHTVd54Y+DVbE1aYskTeszqRl5lcUm7T/B
rVBU23owYFerJ7OjwSiG6nMVhKO+5Ot69STY5gmmYIvgPfeEUfAGH8TmAToDwVld8nQ9/kLiFdmT
EKQ+SjMqD2Mmq+zfe0wP9n0msdlIIwtJD1zkH6EZiq13afQONIBjWrrpSC1NRhosDM9Dc6R9SDS1
qvL3tIz+v3rDhe+/dFYY3IRDV8rGugWmFkF0L3NU5+wCEPZ+sSPR9w41aTafF3ZuBl+nV4GWzkrN
+IqGBL6g5HLdwVYyDwpTfRaO3sRSGy+9uQ6fUOf+kYWe5/2LkYnHVhyfFvHm6XJEgQDefaCgZmnp
R4w4xires2sQorbdz5pO5/H9wzNqKAfEvt1Og/dsiuouC6YRLtoEpdkAIh2yRV+WBDjpnzi9/T4M
joFX1E9Q/s80mP4/WzN9GkmG2mMB9viCHZCqh3S9tUnHMY1H4Kb1zmmPcK/Q/cg3vpwp0KLCxEUE
LViuWfwgAeEmL7GrhNIbZu8m1vm0MU8G03GPgwC/DVb3w7oBoJyGbW4ZqT17C1cVkOspGuQocFlv
Ou4mlGS3M7+9TRr5ppQJ2WwfuqXxn+PPsb0tMJ6KQYN7f5Q2Il8npU3hOwwPwnt/5T4K5Lsjrwdd
1JpzjBhyjM5H6JGPQuc/yC83IaZ+Nte036DowkLnXAql+vvqcnNCqv7H0Z+67bF25buMez0uUXqp
BLAGv+/Tb5AujBkKCVRi4486amDfJhfRv43ScxH5s6VQwoL1/Tb0qBblPuJcm/mg30wPdD6vqMOp
UqMLRC9OuShzhaoJIPBOg3xztQ6LZxdaGteZd8Nm4YbEIJv7DXifJI5FNofg3mHdEgpZwnJz48Tp
1GXSb1m8RVB4+8nxGuWG/z1qhTBnmz46Xj4syDBBJgYl4m1yxuOroQ3Ssl82hWgxUkWAvgeFlgyB
9Y0/Uual29cjKo5cLWkUQmUKBO9/L/r2ipxbEOXhu5EvhDiDhF5AJDV6+5TKEbufCo05PKNYcXiv
6vzJcoi4bnVkPz5kJLBuG5KmGwcDeNWe9AH8TilTVWPNk0LXLJV276YAKL3DDjLMYcMrlqxbV7J1
cP+R3E0zVvzvUpM3rdpDntAXAZPF3O7rbxSDovAzEpuJZTXcDvDQ4bJ4B2DC2Hi5Z6/ldVRFF7m/
KjfKxRvpcioth8/Kzr1AC9WdsfK2OwLdY/BWG2K+veKWal44TQkUnHhOuHIRevnBcYTD+PbLk7BT
2a/NY5uQjpNL6dfVnlhmw+XcCQPSC/yH2vcGKEAQqPjNlDgJJ0V3LjuLSiyDhVPe1ndaCU9NV7NS
TgxeLvOBAVcH+C0ZOha872sk+U+pdc+kNzSdCWerihyGYx/uKmYrBrERr4SpjMUeUirp8Lg/0uHN
xH7NXuKEiIGk9I7xHs1I1DTTwbXU6k4njX+GIRvKiSVirweQQrxLLMfKmmbJlaW3Qz2KAyEPa8VL
d8JmuKaHFupn9zIsHPUwHr8gAUoNBoTUeb4K7n+FWPz6JOOkEDC93yXTbKSaboHe5rVLXgLTLv0g
thKC24d+k11O76/RirfmMiuSIvmJ0Djw4sSXBKByd0Y8kr78oR+3jEh+Ym7LoVc0LiKnZuCfJIUS
Q8J5GeiafL72ph6TR/OTyWsPsuZk7IHr1Kytg/7BIELYn9O8CRdI53an7Hljv/YtErQsbidSF0fN
JfuHRyxUutWiAdX1V5zhii4b6ifVvDiaZ3I6vHQl0hu8kBx1XMRAihRopyefjRISXAsC842jJu9a
L2MgLZmzmSkxsWKnqeWt+rMRBauVq1FPwnL6N2uPugXUBqXYql7J+Rhlw65onGP+RseXP7xMhnnt
u9Fm5cFX+jj1pcMCEvQYsXYA4RjvSaToXqWlcc1Imx/56di8YVCfS8AXnNrNseivwZBFa5jk5Kgz
HfC/totCR+fWj2mmRpoe4cI+pLiursSoptpFaXRJ7dqeIg9v1/3u6dfPBD2eEGwLgyWQo+DHPPv3
CPlteTau6/DfTGUV0K8AaIRJYgDq9kP5e25lag3XBO3oBEk5c8+/xQt7ct5rufMAEUUXqhL3QZm7
m1voEYradHuul26GlKdg3fLwG00i0KTsy5ytR067ktxX18wDQHiIOiPHmKz9g1TUw5jRWtLfMg/9
RY+YXQ92lFN5sp1/32EgJPKVm8AhkiVn2VGggrWsxorQTsRCp6ttO5ZEwO4UXYMnsRPK8Z1/W/M9
OjJGzkqX6+4BuJzGBNkKQouSwj09Kg5iWtO/gcK1Nc6jHGKr8a3arZl20xkL8SdD3U3zQhKSLxAL
IQOefhL81ufHqQsPYjbp8NBRw1qEV0yX7enXeFjdPqRGf19gcXbal8caHjEIZw6Tza1bAZw49awt
8nr9rNwS5OXtvsD5kEpG78ect28gg/vKg35bq1YpUVH1T/88tdBTsh72vFhzn4EZ8149zcxRsCyZ
Dor4/0uV1VmqTV1Oqcsy475kOHH0xSFrYlylv0lzDK7hUauQmilQQkFfo6r5jf6tdpIO5r3TpQ2X
GPCvxnfvjtQKTyXKd5XOgwyE1JOHTnJpNMSzRIbECSw51os70Fs2zpQCqmtqSsbM3RVEickuGNFM
9TvpMM8UoYmcI1CGJ/DMFP3q2ZHR+7MIPzBOgLhDDM1RJfiNzmHXl9kjROpvKG5i4g+U6T1XKBoo
pLV1URmvYn6ibQzRFxpQdyfHyOAd4mEq6P5Dpi7NTVL7FVzZlWbJYV5mHkQt0xccZS7fmKcYc1+U
rqkyqvHKsctZce+rucWb/xuLFdMskg1KPa7W2NTN8LCXbkg/l1qy/1YsKtnpVBb44ILw9khAI62e
SyrnSOpiizcfu/v34cfjz3jF8A2+W1ry9JbPUAvmTgMGDIAsWaUCBfXM8r0Uu/Od8cYoDk3glboY
TRlreM3nUjKf5QMC3u6uMM9KTJpqnH7xzK77cjuBKI4ZWBh1qV9uG3+BA4+XGyfHZZ0xyoCOOHet
3gR9ohtn0aBj+qTwRs31Kzx0gmUiV3nt9V/ifBtiOkiMjwTRFiILgDX8p8ZW9QNFiUOzfVbPe+cu
t/jIm8Ttnd3H8R50tMLKWtx/LbNUVep3UQt139JBXz32QIFM7IIh9Xgrq/paGLqV71cs1snU+GIw
6aDfP3DGWMqYmii54wL8Hd5UhFR3bUptBCpZzyOhrBhWzUotATzhZ38zxjnvrG6xIjEKlia7ctqF
59o4zEl5ksj3cDCNAep3GVbRNBQbPsUFqQuufsRMAh2mD2X5DdXwsxOmBVECbDN5Jn4FVUTPNvan
dZz4aRLMP0xFXLTngK8nI8ikeAnRC2I1zVfY17HZltfb3UGOIKo8Qe2HNZaaDDJEudHiyj/ULv7C
q6efKBpsGVZ7dvCmvHzoRfdToA60km/G1oWgNGR3j4FhxSk8OqGvsbNtWr7lCHqcrGHuDFALswJP
iMqhx/wKrXhEu9hmTqWx4fzMsaCqWM91L4iTuqdCeqjbuQDLw6To5D0te0fxSG5yioPABQqsuRvk
tyLllyi9W1YdIYHSGjBAgchDyPhIjB1BaQH48dBTZU8fBrspLdIIxhm8bC0mVKjW0P9l5PEOg1QW
NvDWbKSgK81Fs5N5i054+kdI6kbweG+/l4p/IAGOCLxz+Ts4K7iqELp5GP+n20W4SpWpc68Enzaq
DukrkjxolYG5+4R8E4ifrXFJ6X2zUmiwIlMgNrloteaCzpKz8sifITEjAFjmCjE+73RfVqFf62hS
lVa3J0vXaW10O1QBcBzLrQJYg4xVZ3TPyqsQz0Q95V5DYx7JCJv6PUaRCT12L2/B3zYBJQU4Rm80
t8COGYCaGfnpT7uqsLMzoroEqyjBpr9yA72jn0Zv0he3w5l8DGK5Axx5ysKd753DEqbF2xZOUldd
3uqKG9KbUZ8LFUvarXgGd0bFGPFTdAq1gsMRfMMximtOioxuC5WfvbvWIdPXQXcWsWv6+eijZ9rC
o36o3qRHYp5SGAMCsRUU1viz1To/SlPDx7FmeRUEyN0EX+Lq/YSYH9x8uH36YjFZc6KlzMYUay6f
zrKdWw2mo3YZjtmyH3HpOlFh0HMFE3Ld9pJu0m3vg67PTI5wZgsBLFEaV+of9QV0/WGU5L0XJs/J
20V9sGFBMGCGv2Go7ugmBxEQwI2xwClj1sYANcxpwciSvsCRsOS8kd6gVoV5zlYMmnoHRUf47egI
V2gPlEBHi+5b6o6LAHPN84VL2hL+1V6voeac1xaKe+9kG8bhB6QOSIXmJV6ODYVLLqNbSSVGFzVq
sLxMOVC5HXFt+BUHQGxLNDReGQw4peEBovHX+HZOm49aQQMYohRSGG78b2GeKCR5e0+rFHXm142I
Y1YmjsgGQOrO8RLfX7HDgYqLX4yFKGb6GO8zzfQRE8u0KEQ9k3o8/OWgKCqSNB6Ln9SWVeTiatax
lYk37Oo+zqydUD6EIzfp544FjTnOJno8iPZiYYxA+x5lmpqTphV8n5nuQsNE/qc3wWzTX2bh4a8X
lIQP7DP4Qg1VJ0dHjgVakPx6usyPZ1N3tXz4jzXQcp0p+7gDRcYP40VNsRTuNYMhqKkQ7KkuYglO
j4qKo6vdcjB3kkcChQTNi04sM78SZsJV1O9ZhK1JdQlyqlSWsi6FGPqa0tvtZCoOEouyT0kRDL6E
KjL68qksUnBlgXjx8oxc+gk87ZFUUgysJw/T58vbt9V20PXsuV6rxHDMSH+8GVv+SVYrGAFAMohk
NHRKYk0sbIUtS/ZZYiFje1fWxX13XiueKJmtL0UtGmEn+CQ4zH0OuL2dWp2DDVj7tSIZLvJDX9Pw
QydxWU6jm6sdrbvUjWcn2s4H56B/gFpDmDweWKbDcX2aDKDUFKDNyGh3NHHJsF78DRVSeTlVJ7jY
O/tsQKIMiV+qHUvRGTwx2Yvz3aLQ0T35A1VU8yVnpvGMWi1cRqgAGCrD6IMqz5OVkEx3H5roB6ND
iE1TdTcpF5hPIEdsVNgFEnJP05ZyK7OFgXO502bmZX0LQZgGPyswr9WUUV6eQ1a4d0aXjOEAMM0G
5Hd2lReBsnvYeE6UEHHA3E8H0BJ/6UpTu3itzMKz+mxRoL1K1vi/Mm+AoodnWVa62P1ckGitan0S
6ZmZyuomJ2A4y5XR40KVTh6fsNazqrBme9sn64vtIInJilMyjGSQ6LLZBh6O4S0S6mKYug59bd2G
rkFrjMfiGYVZc26CdtotsS04VCi95srKx2hGcBm+8Ib/HgCWMnRG2SOyqTy5usMf1Du+RNZFwv4V
/ESIUEITIsHa0xHgTJeB7wS/byNSrEQjpexkzfx6hHYmz0F5yll85faTDXqnA0abEuCKtkKq18ah
XjD48qJ0TqPIWAnFgkwRfGIkFtbxLJJ9vGjBu/iop6nKgVkAyaZKpS23qyPeiqfwFKXlUC+AD6DD
i0iSPJfmIkz24im9V0Pj9bQpn5rhuDBTOGb2sqtkqhGI3Z/O7RydbTUGes2TtP1iuaIPPV5sa2lw
ASmf3fKWSlZg0s7RLwcgYyGSAf0oGpPi+Tz9mtw2nJmNgR560dbucqLAC2gJaSdknywr3CVrmsJM
srORylpVztphg17f/vVI8BkhZH6GjpAVU4Zos8USAgYEQYeqXPogW3DvTK2BoxHjJ3cQ9kZoC037
XLUy2uP3iLpFeAoK/asq2x0X0VcObk9WMUDB03WWv4taSu473Ovt1PO1PmmDKAfws9PDYrJ9bouq
yv0LwahcDgrcEufpCi8BFxs2drw1M00KhVF/24ZscUmz0bEiZaOHXkdlBXQfLcWL67r8B/taTHyN
9r2ue/NxdicCA6oLEQrp1y2/29BX/6uOKj2BSaHmfm/1oC4nGDgo9MzpMQCY2fNgAxiC6XcxI6Q+
go+lR8NFuKVcsYFakJhYE4Cnboqi+9A2rbJZT2jDy3WNqa737zXNR21s9uFlhTHDCaRxaZaP0eDD
70DDa0FXQB6dwVE3gc5dEFnueVVEhdOrEWk7gW8MDznkpL1OjIb+uMlI9FskpGrvzszxIpY0NaAK
z+tQpBLV8lwKB8ooY6yfhjmnz0labb65mdnFNuiTtAY0rHUcv2OtEY8JgVt+hhBShs5Y6DlbO7lh
2m8vMFLBPrx39rmo0Q+6v0oIFkJdyEAZp6IH7MmVBzI7z1lF0hOHe+uWMtsX2ACJ1AufpM3ceFjR
cBVbLLV7/haPOs+d2wvmZrxvoztkaYw1Rw586vsWraErVdg2MX8hj68Onvnk/hlWoAft0AMtHorb
wrIGTtyQKUx0C0/SvLYaaqsFiPPS+d/IFq/h8729tv3QXftg0olPZE8HK+ZTdfc8x33ldQtnxr1e
lkZsIV/J8U4wvDv9tiHMvuHDzC0zVC6XTh7W/1qU7qY5vn5RfP/jROndtaFHMY52hXSIRtk03j4u
bPSE7VqFsLqxrjNixzgcnrA2OZ+nwblQx8aMId1yfgFJxedJClWT0VCTNGu/Ll/TE/7ms3ETIViZ
vukYo6ZmZBZpCqAeqAxDBR+LUaRvtd5j9DcLRpZ0NdKIrLjfVdiod6qqBZOJEWqmoBZqEP3gnVo8
wTPaEUby3Yara4VFsSdbKdreS0Xvwx5+sQzTvshaCX3IrU1IoV/IZF4glYTyMIvmLlnliL6AaaRK
M2V9W0Zjj3tpZwAk0ArNOlJy59mppN7CR3OEtyYG9w2TaHaEfhARbE3ihAmW3zYal9R//pv7waVq
Z1xULjiQ9HiXfTA7vFUP9nSCaCCP0hEtYfd8S90b8ckwnhtsTw7lAhC9LPlSmcLprNvI0JW7uKfQ
rcjxbfkZJARaqKxcSPWhU5Dube60f/ebKxOOFhkevxEZEoUfr4lYhnftKrUGn3IDVm/OqM+diC3W
qoWjvZtese0NJ6CkyABYWdclM7qcxzMeLwkhxdVIrKoUowXMx36maGe6y9vFaYt9YvJG+sb7tQLq
7R1pv1Qa+PC6jsn6XLYhmRse9EfNPX2YWpZ11BFSd0fQpVr9sF5wdSMgv/olqexO2df/nZimZbwL
IxjEbSlMtSe9pjtF65xKm+41vl4RDSqhM0hvEiDmQXM9pzGwQ+Wy2BulDxGUDcN4m1V7b3P7lQ4R
dGfEpeCENCvHoAwg1PLQIwiSYFSVqnVA3PEi+pfolrvoZf67GSKYIWSnl1CgNK9Msh2OCGscJrLw
i+OUg/eLnMtKRPQupjHe/vFAA/ZlSsspIrVDnPXk5SuK3k2EjBMWaAT0poRqex2fzzuOuek3w9I8
HPCGSF6gKXCieqcTsYZKoRvHGjy1IW45RYAPMOI6TL/5uiizhQr1roxT7joEhFUFrJaDK+nNhP7G
7uaYmPD3xVXWWHCyWQ7cXATFSEV8955p+ycZU42dbTm8DMvwVPcxCjgy7NOCpyD9HIIFtTw7otea
knmfqcaslAlqX9CBX4j4URgLDtYh9MqZe3DKPUy/MUfTnzsPBcYKxJIFP/tuDFpkcruEIkKeleSU
yMYg8GQDuHhD4rA29iRg/LbwyhgFmFbbk2hhi0nCpPu0WqqMuNjDVOHTOtobt2VfCIRfH2ofxxWC
tICnc8YiBtIVlV57inVzAOmpim4V/OaqeAYdW/HoDOnXlg/hawU46uYeIX/8dY+NS7XPwg5veNtE
j0YT6ijavQSc6CDVfCoF7ah6b49/bbJuxi8yOc8BuTipcu9g/kLXiJ2v7T8GWsrvhOqKtn1BlFH+
1QeKDU7QjuSZniwRfUN6wiIVqYY4AvtDVAnnXK1t+GnRpy0mPPwVJGgx4bFjiC9Vu9TTvPuRMGDD
vvg+XlTsDK2WNudg5fgTfvg5+DRshgl34m3XL+M+GaM9yPbuNEm67LxcsbLuVBFg2BQOTlWq3vxr
Sz4aAT9crMHt68zCdXB8pEdfWAJ4V0NhSNgcLF3XV6EoKAXsaLXRwbJCopE+Q1ohsUwb7V/vBz17
IWNSsFIwkS+7qUEhgWcTl3k4qxIBe6e+MweNDWdXFvP88K1Ax/SqcJGKxcy5plbLe4nW+5eeZe/S
rPGIvrIn/ofKfH6Hnngzsei830RKJBvV8ki2eGROD43y377NtipiS3L4tkqTgvfTpuuOhgt+8Bs3
PhSFIP0T3S+Begyd9cQsPSkVRy8UrXskr3zOYXrBGATXXk378XGvPknZHZkKpeFZ58ctkwTW5n+T
aecRTLBUfz26v1IsDHQ4M9HdrMJvRTz9vtT3pYOwwig1S5ZeQVkz/qlQV4A1GBmLTaXc965i/1BS
iLx4dsW1OROy507I3DeHiovcjzw4z5WhTXaaLycvzLY6l0+l2tlxhAGjdna48xP/YlpDMKsypaeF
RQsOEE1KkFkH0XOppEDVhtyOIyOatZwudXNISqzn60JjQotAUwUHjESq/6pdWb7KzAq5KsZkyxyV
yhlfkE2fUXli9NQKdXGFDwYhwCtlwnOS9hcxTkEOqnaHpPmXEe0S37hGEPs0f/QYWyuple1IzI3x
dzaYb37aflXmjRcJNNXxgyT0ZfJVYYJQwWWl26SsMoXA7ulDJJx2fnny/zU863PCOg+/FvvqMLeB
BV6Unh+ciCXxJ11L2j9q3qh2X5TN4fdF1F3DHXXRJzkNqCBmrkHH+f3pa/vs0OJKccGitP9HJ2RJ
HUtM/xEGyYdNHY3LvuQEnYSknLJtXKOKupApfxgx8T6IFswyJkdJWqC5vcXqqRsPLZsO1C+xkMqu
WTE6niypvzLwySsQdIoNFj7UQWgoCxL4MKtfEzs8LmsFECe4m7fKn2UjsArTkRaPTAtvNEC2yQWU
6qh0Yk5fbhBj1QGp0EpP5aV/L3Hrbbxp0lfLK990v5CvPit0/HcZC1vjNUC4S4xjxpoK7jl6D7R+
Z3bsy7cN59f3M+AbzLW6kl4+iXShbeFxZDro6QSFUvuTVDPyvBDx7fAEA/FxJ+V361uAvzEXKGj+
lSj6GEhK7+2mkol9Qy9P2J4AHYaVrc6zNDokqWntk+1yM+RpzFm0s5SEIcByOl+M9lCzy9/wS6L2
ZD4Omnp1ZiUnELrL76PSZN54b6B6bjIg+sMkBXtxXm0N+fgOcdBaw06wzP+S1ZcWWYwVIA4f9rqe
+zz2xebNFY4eFaY9Xv09usyyK2ovdJC/P41oDQlketaakuI/ZPI7lI8mGU7De7r8pRlc8ephKyy7
ZopPnb3LcHNXc2dOa6WQVDXULuzdhbJh27NGqVgq3oFN1E3BD/vUcmn3v51Ri3dfCw4Cij6sn/i6
xwJ1r3tydf1KD7AYIw6ejShJD9BAcPkYM6Oieelr8dAz/0bMZFFv9iMc4cuovkuuNZCWAIFDPqES
zv/Bh4ubSVGBDNuUCMy7twbpy/z1I1T8opc0ZpuVySFS0ndtvzPQXWNyfmXHB5vWjbTgYicJq8I2
kgOKPNgW9wIYftvRCmsgPVhJtiykc4GXjFbKnnxPevoacRMoczYj4vf2FFR8BnrAVoZyzxNQV9Dl
faQQ1PPigOTKyVF/aP22rVauehAX0kbO/hRxzVULJ4jxpwTh6RJuVLzqFdW4w7eoUfb7LcwOt4wd
prErJROVG5IKGMznNSbv5S83wHyM95WVyiJR/fGzZ6Tu+jMMQ1ED1R9UZWVU9syNWm6efn/6foAu
zqxh7WQ5ImGrmb2IZuVjqV/WUwCn9rtfd4uxh+lb4qQeLyFQpCtlbNxBWtE0dFF7G1uk6uzC+gWd
L3u5ayyg2W/q/Yr6DfV9g2ejGPbPgFYqDJ0gVyyx2zq5Su0Zw0nThtY6Ihb7RosuZbQIl5U7HoFD
zBK74X/DF9vNhN/jesCqkqa5iDeKoNByzw3ZsXtg5Pl5w36GfldX8wsxVLprKxAyItQdkg/7MXZd
+T7Mk6GM0J54C9NZZO+CsgVqOYQgBXZJ2iA2R//74Hh/4m1BYxErvIDMh8fAdjkjwHzPNzttRXP1
TdwNohJkD834muEXz+7ryb8VNS0T2AJLnfitjw2A4rt1OUl+luq9jByD6cc4NXirIL8kV1iYOr3y
GmuCoBi7HlYaPDNw13yZCPE9JCpFimL3AjwVYDu9rPvfzlchdc+IeLxVBa2Iszz01CdEVGcMqpov
Oht0yaSd741YeuI0SZZFaopytVUzmvaUrVQFIPyzAt8A5+BN/GvtcwUAHCwWUZfMYX/bQ3V8rw72
kAmNxgcywsl3ptg1Ra7dQLEaIf5DdHl+SrFCWfuFudZmDsTP09pDgFd6JyClX18S8fHAqsc/V43N
jOnc5LY7jcxsxQkENryKMvDuR/lQLYFCXXdIuhtvFAFg7msZ2AjQ2T3co5k4c7Rw04V3tNW1eATj
/6j+JK/rYMMKHKclXYLvlXgQQkV7bWYTkEzwBpkGU5pmuNWzS7SyLXT+T8I4ZplmihNIRQXoycrm
MncWEyEu3MV6/t6cMAhZd6yvyy/Bbodu5BYnW9N0ZS9XLCrsOvg7+vxfGCkI9nFh79A4/We4X8OQ
hwJn3XIbnLNkruFTsMm8fzwHwZm7mpTNzdiG61oCSHVvPAJC34YpWf2i7lLLOb2hsLQUy7JZVuF+
gHc0wWJLWKmxQPJGzsT3EFmFSW7HXsmjnmCg9K8z8vMWVEiwyxgKR7LLwuH6kth1NUL7Bhg6blkm
MlBkNLtTxC00ti5CHagrasOhyzZDVq9pSZlRCYuVCeggUgQWorTuyAbgcX4lLKoGvnzdwoy3/L8X
yPZXeyg+xQIW8a2Gwl1NNYOH1Leez2tWXtdoGLXLFrxa62L6w2wEjy2S0Ux99mv18pnQbUyeWtPr
3/EUqmYWAYdpGiW0ZPvLZ3OCq1pKi9RLDgYEvlB7OH77E0NuhuNPd+5Xx5ieyq2FWchxilzDAC++
VAb059IB6g1ZyfbbG47BcqR1miSwEzT5JzwK1rNtZgiDoq38sBuleX5SCRA4jBSkqeCridNpr84f
E5xZJmmAj+toWuYNRHt3Qcubp/dfbaE4trswxu72arxfqbJd2mbKGyqyEV8QL5NCimiFV7tkY8fw
IQZPkkOzWHph8cuACL0k7Fd4nkD7mX0plxz+rwTa6WJMVDLcdEEz6DAgf3JE+aFnsHCEH2PAMoYf
jDISiXHLyOMe9iP+5/gcfYW6zr17rYG+mlzI/G+hJXb8boVvzDCTLI5QC9aDPv3jNGj6w4BJ2O62
3q8fmv9IvsB152osMAKcHejSnLi1k5NwV3RgcZiA5F41/PTZlv/RCKbPEvyv1ZsELCpUidkGLAfO
fCfhtCQ/UWp3qEKQejOgnnjPqL94DquaEWhVnb2+6nt5YziAedD3Kemce0fSE1RsR0oOHsK6Ee+W
XIX2SRDkH7oSyBGp4XF6MUsvRRKVcG360dUDBW3EJYU9pwnqpIoVJhmSiYjndp/QyjFl9R5O8S9O
Ew8pjJwhDsYxOwtTt0CDFsJLATdZIDVRFEShDOLTa8cF8jaIZ8QKZpMqxHbHvqvRqU0XColarNI1
Gpp8FWkTL3U58SRpBTdgUuKn9x+7eNBhVpSZzyXK2JzRgvg15UgMz/v5CToRglzIyYyxI0HWr3F8
Y99ygRWpwXUJm/28E53OVKiKe/g4J9cxRAKyMb5b4+owKhSTufBAJ+dVMku1nzit6F7d9Qgqkqt5
JyUQ+4ixuftPiSoGaginD+CSt5O7/2HNW4xuZtDYiwhXqtpcQFY7gKbJMCJkv/EJsO7MKAZMoySs
ps2HCtN16zD8Q5c0rrRECp07X/CAlC0AlabDuDfTBiKbqYwUUTztEF2uEbnfGJ/iNjFchZMe6HGq
tOmpaV3T/4MHN2d0f3WnXdg4mHsgDtL4NzW2kPpj3hgdSy3LV4/fD81h98CzToSxia6Ymhc99ExY
Z+KRG24kl1yP28ooSRwhT0tekud/L5kzBlrdKgSghJ4vxL+ZaR4AFgVG1+sfU4B/jjdxP92X/ofu
AHjunKwopk6b0+/8LAMxtKn2LdeZTdS8KigPeDO7pE8CcA0aNEm3sASnvbOjfgJxAm63ebnAhNsU
sB8WN+2hWxoCBr8FutrDwU1mdYM8KhsRon2PVulV59ILRl9oHDCSYblnURMNbSvd2q2bEwxBls5U
fo46op20F9vUKqbQDLJOdHr/i/YuszWHvRnpXE1kSV5RGOM5kzRm5Vj/bQL1Coc3drD4NuafCVuG
GD6ldfvClO9x/Z9YfHDsaIK7hNVswHHsE7PdxBDyPHPWxXRofMeJ+O1XAzf7ttDnCA5W9EWaf3p2
oVrYPqbOoFQUfm7kN7GcLiooeBcWePynkM4Gn+PCUevQOfcHsBlLj9cyRH++q02bx6szzQJSy+5c
HyAKGSKqsvnWW1Gt74cqAsTZhJFucy2CLLzi3rrkPDltIUOGXNDcEQHP6qo0uwfeVgHkKLr/DD5+
0rwC1OvUI5eGxeEtvDBsWFhYSpxCSjtT1AoXL2hg0o88g960ro9vBr4hAiCoe5q8Bth86UmBnmIV
z14tbpoEhBZN/y2n4CeaY1WiHEQqoLvbEp2yzevImmrXT0F4Nq2s/ATDSqRNSJQChxBATMxctWBm
bUTGsTlKLdShqLIVkYkqagS4d2akwQEbAeqC6W35zZ04JxVy57iPRhb86U6IUPuCdsWPWtgYjU0U
0qQtbg+C0ZztwKyOXPW9aQqzibAyEXruIjvVVFIo14Mf7NslJHxYoctpfXde8KnT97XTVNxeY6BV
7NtuSSzXLhk3ruUBCx9/j1YnZMoTJPe7R7bS5YODZbnUZP7ZfbUiXeQ4ABXvldE7t/15gkuOgIIC
7vTbj14K3B347f0iuzdT6670tgNZvx/wkWgJcol8M0NN2LZl8dCrbkG+/f7D16gJLrCcogoyYiqt
RTC7kqB9y4LMgNLFKkYqqnJ6pU5cgT5LTDWJmUYHJYGV4he5K4Sn4m+Gp1YH5d5kJqour4tWfdpk
4ltdmRxQfxAkqkIEHTYhAP5tw+77jx2GjDh1xNZusxGFaoJuqZBHO3ufjFayHsYcjUnG7NtAhnjk
+9IL2gYJibHhCpkskyWzRyd0fT3k0VnqhTN5yAuzMytiYsLwhrWsOP7SGSZ/OI+rG5f77VDYLqq+
DaM77hw7Am98zTaLWAYiuoESwwk7FI4hAutthV0QX5AHOYrCMRScPsLn5S0VjilsNrYTxVpxLLQ+
w3fwe+4o1hWT1CdzwyhnHMT8miij9JUsOcU2y1JHzZkBrTP4/KV2T7YtOIb2dcBx+F7Sjpc2q0WR
xHVxk+HMyqBmzzdo7sPnSPRVPBxwmWe91P2D/axviYrqc5fywlhUdAk1aPDoJPOzKPqeOcJGAeCP
Nyo34npZa68dlAj94XggZ0anOOgMT1ngYHs2JgLg/XIYX3JYPiPtchtdvlMY33Mu0FX/Cm/8WoxM
0fpjGdCm3F8v5oMOTSyiezCjYp/GQXitkM26JuZA27Ctbd/ogB0s/u3o2DuL/XlwinabTwdrhrcQ
nh3bEVYo4IVdwUvuQbJk4fWmGEUpQAwYRTuU0oyylUPp050znMPrXoI2Xt/f5aJCssmtvTKFVRDW
ErWhCEgFWw+L0fR/k55XEv5mgwUt3Az7ZSj4yXzuSxBNfbsYgP/Df5zMHUWmzBpqn+Tzf+AU91UG
5c3jypB/V2kjBva53PqFqcwe1e91wp0mID+rRcgDxmYks6jFdn2GTGw06fIGZHYKLRuKzq3+Nvj7
KmbbFH2mndVCpOZDm1vNviUHW0lvl5pVARiuVBfykwRhftuOGK6ogJiiT7Wjxe63LM6qwkAZ9rhM
Nokg2oOvCp02LOHn6S97d7d6FdRg3R/OfJ1oXnKAeFMtY+iZFElDeFEE+TdwMrBrxourOwVAcvwg
mUnEhRw3RpbZ2v8xDQwIphyEpdxShmAL6pWIr4qRWxLgqKi03usbizZSqoPszjA7a71wzqHr8wyC
ZldEre5PuooI8J844LyjBkFAfnWW6YAcrnRAI7a6VZLPvXsyjDVIcBXP+dSS83zy+1WFFk6niDJJ
gT+5wCB4T8mKMyUl9wzPYtTm3uZOxyATgXtb/Vaoj2SVCDNgvxM6rmLdhAwxAhGsKZNTchA+yCW7
osk5jb2u3LZ9kq7g0xOH4ZvA5cG5mFYRIIVjTTLnD73pxzpS34A+BoCx1ncNesjSH0ES126/pafU
0De4eOSHPqVwReddC8o3SS3qQc1/5IhfvlPeK13kx2XuFC9z7EsolHHiTQIyUO3+l+Iar+XeAKWr
NtlP7dkLPGcXww5AedhR9inbBDN0uCtAH70zm79Lxy6pnDUsFoe3GDOZAzIxgzD25x87IEfzSMES
MS4UMWa+/RZ2U+ATmCMIhWLZsDWC55F0SSFtGzRF6zak/C/m7izcjDoWm0tHvvsoJE/Vy81Lw+h5
CF7/dD68diovdpxi3hke2VjmKydH83ZzVza35P2mrdW3qKgcueb4/pZPN4EqVcpc1KxQy4Fk9Ym0
ynwq7I26YeKJr7IqV/hAk57grwHHQMnoYlvlVXMc3/ujvFbRxejJsfa1XPhGP9Nbj5wYH3pga2i7
GmOYLqTJ3wRvwVGipSTJl7co1AafHcyjFXd0f5+hFwBtFKHoyNkgWVNorDnWMXSwjs2dUz0/SmmG
PpxZpNI+NHxQiWITWKf/xC08LHkDgk4jNVlpQCQtawMCgb3/hPmsMYe40ipXv3FtcmAcxXvjdgHS
HG4ZgcrUEDY2YbTjn8RBJdLTf4kDob/r24muMPyGjm2kw8YUC7BKhLoFXIcNQFmxCEZC+YR6qOIL
ZrsFA5jQuBWsAH3QTqzn8UzfX2zUc7qOqQRt6kvauQ7B/ScMec12QsQwtfPDhcE/9eDYE6jjLr6D
7J6jS3JhCwW98XRNE/qBh7ffE0ceUEWoNncAQkOTmy/rxpygWCXCCLI+Kb42Fz0fw0sYklGNZnTU
UL/SQtC97++CfzQFmu90ZK9SDKeAwlo2GaoVThbsD82qgw7LqRxQXcHqs3HOMOV9jCpyLavcOiSw
FdoPOuEIP6DcKQ93rdl2xgapMh/juGuy8sISwBSbyig5Js58L7M32HIJkuhVLrF8WjzZg+frQOtd
OjGJiDg9UKwMQ/RpsTn/PZTx3risr7+GzGfwr5ujQXlgrMR3uoGeq/LIzCrYGggwLbj2MO7aQn3O
sTbDnyNGPlK7+LXtkxaLYay/fYSLgki4XhEIRLONQ7iycB4R1kB47FdS2Gs7+/gIfI0+FoMGLYHR
s3RELrbA2zMy+ESkK00eSVpJwI5H7WraB6+GVC1mldlCCwRzyiSZihoY3N50AQPJ56JlIhzTIrZZ
oDxchh8TqK08ItVw69qDHhZN6tjrMWbt8NnDSlvblFLWbgH4GOwaM+5qzBnOacumS7LSLsNO8/vW
nJueRLdQzNJK6PmTekol7/SDBCrq1rfOg/jyl9fC2Z1rN4+IGZA20roOOsLkaTh57lcPwv8rtJWZ
urvkQIlPRmVrVF7hHwyZtzlXtke0sWdJy8HFbpYejfX808a6uGg8rviVzHzt2PvyNW7vbgwnflwq
6hiocouYr4QUCf1fSkg0YCpZIhvP2qFcGKEXfQQEvVU/ctRD5ANd0eEoHPUE9jI7cNB4ROUdhfA8
THq2UrAwVjWUAV5irMzaw0S2j8RuYG3FGDzmAFpdiZd+2JMkaNXLNW6+QdwUj7PigznkyCejIT+7
H8KKNPI1pT18BSG8dhNkK5vrlUJpjjOMN4yZ+AtO7B7xKWxIDkYVFrUsDvuQX+ZcF5kjM9g/Bq9K
RjdVFOlOIri81V+X39Tp/ZnooBEGDf5x/FDBwL5O7Fd0+coLMtM7jqFCxQwLUzhdfYj7hD4a6P0J
LjdS7NfXCOoPzMM1jfKZZTqkkmxOEUvZoUquupnv/EtC/KDiXMnWpnq8n7ZNo7VTNvmDwIgiNgWz
yqGJFTLsXlVyKIKVorImkwQsIYbuKLpOZjcP9AvqLr5vMceYYNCRLZvXDT9Wjy/aQGmAfgRSdIUg
TPEflpjGwM5fDWXyDm3EUMd3PTFoYLV4sCEMRkqLtumez5vhBO6q6NFCCBVeH1inOS6d7dLXG6uK
c84GGeeiZQ3ed5ZDIy6AFuQ56/SrEciwwJ8YFM/kSXu73NB5LHUG7VXe2WMHcR2a9c5ncvYPxgz9
Dj7u0wpCd3xpYlUh4b420h8sloIYwqPwkn9z9zXgdIrJw6EcvXLWBZ10MtNjQrW3BnreNvV72+7v
1RfHMBQwudp0q4PT0ivlZIgbe9EzwQz35+Xas5k9unJHwV+BAXCqaVYDJpNX3I8BNHF3NK1gf1Oi
0OnxWpTBy3SRf1Crc62CzZG0If7CYdto3ziRanPhd4oMRzsoWp5ZLAl1bHyTU6CXRjwytr4eNUHV
97TG3Rsh5AFV1oxnBgACjzIzInwhrebJiF5ADbHKYv+RSoNjSDBqkTpxP2qvXJaI9QgT2SDAUNlf
kpwHYCdFIEIc4TuhgDy4EuDT+gB8JgAgG697HeQOdPcZN4bTUghAPwsg3vA7nGx7OEtFQ5P/3YyJ
uI/G68LVvVQyrknrSTpSOZOojDpGQYojh8b3x0guLBGA2DS0h450LDT7pFdIFiZKnkvkK92qmO1K
TXPSyZuDlAh5yfH/x6NqBl++my9DwT2TKtU7zwgNXJ9MSQQ6vav5IloN3LDh582+3ESlvQxJo3WK
Wt3F1q3cn8slN8M9T81YroMJZFCPk960viHaohRwkis/toHikvRR6nZ76HlA16m7qL2xttSOcr2q
zctyt1rm3PWHDWeYEP8eZwJbCiNGD1resf59zYFtQwKmaguqi5/ddIyP/Y0MpnCoBV/8czWYhJGf
v1oenDPd98xmKy79pHhvUVX312IXoE/InF/JoJaf2aAOH3oUfiSSDVWeVgXaYuzFJA9wIHieDu+c
+P/t5CIUacuT3wE3mgpg5/FoKeA1Fs+UOPu3lJrYlO/y4OeOFAzwRn9riDlXzORPxhz3zFV/zCb5
EXdy0ymPcdKMdM6GxuWPmMgKgVU7Q68ji0BUynk4LxHoQDEejsfVmPXVqxd3F0CoK4SxCBAhsgDR
wkM34KbqDLm/8/nokGB24i/+LZNmiVTDv745qUa32iCbvpztwq1ehfZnMqsA3Dyr8SEKoh5+h7H0
Bdx6Sx3ZEPJ3W7zT0ZdoRuAwMwyR7hhepzVdqJCnA3d4dTkCEREowXxMCn7Ax91X88DltguswgOf
BEnq0vM/jbLe1Y+43AH8xj4du9iDhyolmgE/sNi707Ykp9aZE5idGlXTmQwVudiasE4VGhpDg6MB
WJo3HJ++ASO/aS9fbYwq2g0mzkTUSAxHU+N7zv6ey6CirWkOVX6PIFxFCfS/FAoecQlSU7Fqiuz7
6l6F+UK1kRRDfiluArFjZtPxsF1pdQ/2eIl6bklKhNhGAgkaCRvU8CaDbq87Pwe+b1+spZJOccXx
aCt/iGz2eEfArgRpDvy6cG1HumCmZEtygLyIK26hT2gw4iJF0BaZtb6OTiJiMRXzPL2Njy2/yEXo
Ei0b0ltqEOMJ8q1NHThgt4BL4HdVVrbFYm9roeN7uEFZVD/g4Xv7lWo6QQMlsRSA2JByeTCyia/r
KJvJEdlLMHIjE50yYf5jS+Vuph2PU1hH+nAhAr6f7V49Tn1jfcGKsC3O2dJaT1esbEPV5N1E9ZRT
3xtQysp55DjGo6lRjWoE29FoRtTOi0V6QiNpGfzouFXZPrjOgqGAod/Q3B/YH2W/kQOOksU71d0d
vZL2b2LxQ4AUkLnYwYRIB+VWRZTr/OFRn93kbo/6v1Ba0EWMgATN+YauEY9nzRMR61ubEjH8Oeqk
7u2o52xDCeIOHCgy/DOkuGlSiDb5IclHC0HQNgnAzCKWjVtm8Bb4qn2MTlyPhbdXX9zcZKWmdBnr
BemJrXW3FcOsruesOcCkl1/9bZXzEHIOZMzR1S4pR8P26w2DwlWf3umbNlPXd136IvzPzT/vaaem
ov8/PGM+qlV7ABLcnBnluNp9CPix73Kzop4iaEcV6sZWTCFdOb1wD4irjnkh1Ne5ZSe8KczSxEPU
gqh1g3JdL90Ha97StOxI6tDZPWoQcCMdEfmndhieslfO1AQeY3UF72u+74bwVVXKs9lz80+v+H3S
s26JFgvclOZkdnLKHiyU0zTue/uX9tOo4g+xzf6Z81SIwqdDDNqwog+/tiEyBoaGm8P8/3duxk/i
01Ra5LSXCA28osFojdFyKlPZeYtnGNI+Nn3GRAlpcdKLl6P4OqPrkCpubn6Vkt9wmbdQ9PIEAqTF
CzBnurSdwM4B0r4YwPP18sAJOTaY0yQ2AkxDN+VqSXssbZro7sOkud+FFe3zyqA7+Zgmh/gZ7tKb
vHnDPuxpcsbszrz7KJEo52i8bb145TEGZonSC1MRZqns0lvXzPkECq6Ax1psYdNULzpRONp0V5VC
CXLbTbcJHY25xvO3uttlL56fjPimUIETBiVfAdprCbtiuqFEqXnWPYFbzqElF7pYgl/sqDM0o2TB
p+dZtUg4o0/IqFxP8hN7hBR9y2FqU6BQ++uMPaiWbDkEx8mk15KhuviJ5nsN2DQ29nw7KqnfHB3n
w3eKZGCT663qn2/xkNwPs+Y+InORisD8qv+WhXAl81fWk5ym1jmBvhoISqnHmZ2fVH1f28G6/vie
FSn7cNDCCQ4rDQhQNWUCOBPrAxfChGhbW66O03XzBBinq9ElAENhE1v2FB3iRFy0LnGE1yyyUkYf
8Pna8OlyGtUYB22F4rl5I0o9kdmFMLPE1LaMS+TZbYGwKywTtvVnEECJhBO2bgZeUEKRPoOVNONG
KSnwSK+EHW76syaX5ihMV0whJ2/2uo1t+BqU1JRo/zAadgejF8UWsGnDVP2H0AjwHIPgnKp1Nq4I
UQtZmMSe+7UNAUsbOVkNhCLjk/+FjdpLyY82WxRgpRPVPUDOdtNBZ7FYl149P/CMtbh/wHragLY3
ubUl5V9J7c/xmRPeaB6qvz0SZ52IB2tSTGcyXeYUM4McGBcqb+3pAVJJbfwOC6jmWFqadfPsa4Cd
A4vH0xL8xNX3zhWvrk6K/7qpZYt2oMBTbBdTUpDCvDZhYb2FRqPC0kaj7nBJQ/aSGAi0eC2MybFg
RoGqZdSuS1I0hBBpOVi7iVJVNZqfrJecSA5B1MMUgYH6u7+CFcLgUvY4h25wBZjdoteahYNH+xA9
ezUzUq1ajxd6TZJX1MvRqhQyQ1Qs6j7MjO1gGJCHMqsKBprwh8UvxE8lfnuSSecyb7djp7LxPZXa
0ByF88ivvlKhS0g5vh36OWZdIbQAUBN68eJnSdOyT8OfqkOLQA72REwUrCQvDX9KNksuA9P6MSiJ
tZ/vxIb5fy5y5lMbDb3R+yugwK8JbTMPZ9yK8OWOaN6182fqRnST+WB3alR5MyBCBxDsjk+4DTOc
zdsnKHuVZEy4ZTCfgBGCMTlxfIW2WPe895dNm/iQxYk14quyHEfglZGuM/gtWCVt+M69Y61pqmK6
JJV+APRBNdjbBMhf+KVGbCxS1p5PPP636X+w1vl5YExUi9wYNhyVOu5kgkWyLrsNezTtG0GiaUaJ
PLVIXxnS6tIkUlZn+pW0tFIDGWsLItu67UTTkmSoj0EhfBxUJ9giJ4UZyNSqi5Ovrw50WkoiwkIS
a92V36P2P5Q/P3tVQNjHyrnWrsgwFIwbk8pxmrh7VRduCDcwECT9ly41aOypf3ksO+QyVxoxjH0G
cKNgcJYypZ/mArvP6Ws8xgGQTc3uHypbZNlvJKNQeLm7g4g/ILDAXm9bJvGmomy7QGLD+tfmwEPj
A9gwcU+v8Oh7LnpmtiXl5L2EHcjzK52WRoyJyS4ekd67Vd/K0MqcvslIaPuqOJtj5ggFJzQS9HJ7
29baFy9XYVRx5jEGMI9zuHA9kxVbHkXYieb7bJQ6vFAajt885CL7JoS+GZmw6bvtp/bE2vrt/Qsg
Az6mVgw/XJtCMAFtfGqlgChjcVBQXpvx7lyc4ilvxhLV7NBZBtL6geh1fQjV4zZkE2/7EqWU3njP
vD+LT1SDbw7pEWiqmNQMjNj4V+2W5vB4eJCcmvtCTdcyclgYJKQBPQxnMPbB7Qf9pBslgwlEr3B9
FtUPjS1ib5NK6ED3Jrgh3ahxdS6XY0ORxFy0jbE2DTkbUe4AWF1THvcwEI2JC4rNd2XLFiJoBy02
y9csiUN2izxAsEhLCkQYpsU+R2TrhnnZJcW7bepYPlnJ7sHpKQHr2+Jwq3LpZMSD7OU5eLSvloFL
ik/+2tO3iHkiW2NxDO1Yd1OAOCMjHqsnabnrLaRWoshKY1Xwut/RuQU2n/6xG3bEvohgnPVtkmmT
aNTqI/OUDDT0lacstlNscKNwvOhiZYEZV7KwJD5PHguihQqbeTQaI6ykBlZE5v9wTegqun7kTsvm
68BM4/Vpfg0lxeGlKhCdQ8WuowZ+OSHRxeTVZI/NZybSfkJXGLsLHNy6afAwM85fd9w1SedRRQib
jHV7kQroqGNrVQYGjpdCp6IXGljZ0WwgJvv04dZDIRKOBbbZuXVft9M/rkt0+YN4PoS37KipPkUZ
TvPXK36a2OQtb01sTm54+Anlv0Pzr55n9zM09hokGeO9kGusUxpGvU8h924XmkKCAou/iB3dJDwe
sBSciGG1HqBWYrYi8oEi7FwAWW0IHXtJ3tYuz7L5vGwVbaj60ziE4epiDqFKx4nVumXvM2MKFUep
Y4kvErDc8+Hfb8oWRhtMZZfYWA5/cyEqy8X1KiQhDp5o4IjRwXvzxeSuWEambsCdTU6Xf0ynA6DU
fQoJuH75h1vQjoPhWFdMX8ejxQ1EEDPeMjlOGf2NW5d56/qsuENJBt5kAB2ZV/53jAIueo+FlQOJ
IQUFDwValf0nUMc0koWi1ovUZs+agMSX3Pe4aQ2y+yRShu58yjZw/TGBSjqCHGbQwyEAcgjczy0F
tD/wzpwIE7CuRTyWipK95971mH1tm6cOJeV0GwCM02XdjiMvRcfFEAl6sa9fMQx8l3wFf2pUWWo7
FCpKZqQAdoyOBLJc7Aums3rd8TVb28tOsV7V9rXajQJX5/QgpgECI3XsBXGu0xduFcFx55teYbWV
31fc+Ti0VKL2Iu2K6l5p/N59e2IeV3nJoBS6QtvQvgcQXkG7YvsiMq36V9ug3A5U7QlQGyBPEEbR
ZQ+iaR8/jGNZNOTf+QzJx36ufmyNcZvYP2M0ebhmpDU9UrT7PGAVaffCiiCPt4HypSwNaGKw1Hcx
xezVno4dvwLtJ0P5jFQDwO4GpxyxZ+BbZTLyqn1CfCiEJ51feV8+Ntx8VYQH0lPSR61xmnGOp7WE
fe+9DI6T5SdHlaC2NTg58dpJLMoYDPkGb8iu0yMhIkC4ED14IGIqepOGPlHMa/AFwef9Ukw5xuex
JKSXLSMVhGht9J64rvP98bo9+XXvU3wLow6KjHZ2zaPepr3tP0KuCgs09Hxk9vcPx1MQ4k/FSOoW
klUA/vrAVQgv+CzHhSLqb2pYdyw3ruFERZlrpb5+kQGlyyUWJfICrgmFJtXYOu9+jBCPryREmfil
EQd6BGYfXXjq5WfRAnKTvLF05g6jkmODVPkEgb8/ZP10MhmwD2+Z2qWj8/FnYXbK22aHnRpxh+3K
8KnxSMvaLhSMEfWS1U1OvRX1eHX5v/yX6rK1bMpJ7aYyysyCXr9s4A71WcAthZkvXf7JsOmQ2cwF
parlyocEj9F7x1YqYnxxayl+oEqXZ8K7b1aZgCuNcjUYxjjUfLmOiX2OBx37K/ChNchZP7X4jmFB
8qii28H96WA7ETvF0b5gFk+hmMtCc1/Vu5Eg1f3Qj3mmPotjp2McfjWZlVtJd6Yx4piA6rik2Jyg
UhUAl7DLnPZEGgZTjdiWScUWJBNQha0tpV7r4Ds5zwv1bapQBx99alcgGEAWaZWKJ0gFNEUEVEvC
j2cvDGACas+Xxg6MIqWh6Be6WZjE9CawsIPSIsNPCL7ENPtWJAQl3EbjxwHalqyvcrPKfNlulIj5
IwH6zc3yz6tgIrVpZHixNbsb8XPjx+UCbEHF+2vIFSIH6W0piWkj1zRZ8V35bbzYtZFe9yaYI7C4
Zuk9uLjyrMVceYvt1Jr44A/745KdqUhUBRakxgj98ZddPivxay5DKH41NSsRlyEjI3KdeE1IyAu8
RZhuDe6UIODyDJJVT1irWus+HOX7qrSomAazpvMSNI4RVqjryIjBDBkB/4OQULNU8/inwca8ljSL
hKIauhrRnHVi4+GUzZc/7N+UQ+iFvlGzAc6Qy6UzKevu8mA00MGGuvVe66LuB3yxzcZLtpZAUcj2
1+j5GC7jGu5OHby+L/dIxdyR7cewnraEZW5Li54lO56y4wbV0tbURFX1x4H0SvDx6zmvfDATm+th
1SbJmO4SKQ+J1qrp52YdwvpxjOZB+F0h+WTJb5qimqgcRpiUhhlgk7VJAO70unOxK1WAe4iIdCLM
OA1VROX7mLmeIRyeQoVnutgTjGCKy2UUmbMLLF00UX1HvjbTGJZ3zfGzmptqi8+280rgLiu1Z3BK
BcMw5buvR4qW9EP1mxjpt4n4KSwWN8430/fplleXBhzk+g+sDVXhaSP+SFJ7C201oo5fbX7JI/CZ
V1LDiqdpcWfEAW08tXhCv02fChxk4taQlV6syEnOEnKhNuw0B7qW8qKTNQeUmY0ZtpDoGmQfEhEe
OFhY6dFo4zaaIrkwGrc4ucIYCPGd7FoKwHg609IY4/sDUOpbdyn1wz38r0TfEVx726brh+exFaiL
RILTpnUZUfTTi/577J/xJOS8/KoxFgD+Jw+2w5Z9hUDFvt0nk/ewpvHvYRx0cmGkXg87DeDZ6//t
tJC4wSLi8lBhsFIs+jkdse+7TR5QTGN91WHpKn0vxX6eu0qelFt0uJ3w6YT6Cawa1Gymb46YjK1r
erh6/Su3ulc3TQAvit8IKVsxxm5b+S6WluDPRvBF0ZkxuJPmUJya4KGWiYzjGpjrqlMb9swV/2p/
eSO/9ii2serkV1Yn2LEdPJFXo1kgy1iA8jcpTzKDCbDBOnDbKQNZvnwzWOklQTpllzOIPXdPUkvV
mUNDzoxnV1UYmp6CA9MhSk+m8b/w1ntaoT3lEkqzp1KtlLLULqqiYqd4Syz7lZvLZVHvMOvYKLA4
k1LAmXJQ2lo5NE6b7Z9W/0AC0SQhwhXdXc+4v+C2u4N7wAhJxrrnugCI6JiwtqP4FS/V9bbf7D9I
ZIV2JvqiwoitwsO0TkSOOAW8M/qAo0s7B0D48FB2QrpbszkR9w+tcZQlZ6+CrY6yzyotLDqFL4KL
aoW1pelLhraghKOpzdpRjPgjk622r/tVLz4kRuRr0laJtw6wD7vstUKeCt8Q034crgJnO5WnnA4B
U+gsFhZ1j5b+dYa7MmvWhD9rBUPnsZqX9eVknitjD4r8DZPsjjqmp73TZ1uoZ6ozWmAr57uZnEQD
qEI2PinqcHFyoXv5PxkYD1vrKM7G8GzxTBXMR6BaVUk4eHomPcugua0EBIL5drntiJLQOlyDU15i
G5KfEcV+SKBTMpsBtt2QW4pGhIXD5yNcajA4BFvs/1Ltiu6OU6NuxgmCpVLZ0y/Dn2XJTOYw9a75
7cNnvrCnJecRTusmaDOYpzzFzzsLXsM15IfBSH0p6db7N0WLw31Z/ht+/P+PYtIIlvt2D35Lo93S
cFqpjiyYyIqKAsaY7hx+SmW60GN9arrDaZHEiYdn4AfwstgUeq4vJEet7incsvrCKjb0A2qRRJIg
9nSmu6QVzfNZ/S21FNP2JXPLAFhYKTpwdRPY38H0qfB78RZksHL1YL1G8dyoBdwBj5Yd5re6CQBB
CBmVWNCB4uoYprgduUo5UhwgAxupkof3Hr4j6FuOnZWh8aK9uflefADO6NNkahz5G+iOAtBThGc0
AuqFSpiLa7lQuw210euzvVfwP3ID+tvqj0kWZuZltCIDPgqHCXF8UMTSQUS6XSH2PpXIT2coaft8
V/MT//Zf8oAQZE/quqfEJv4DfvRrcmsuMBiui8k42Qhfhxv68ByJn+pswoB26351PwZ3tnhyZ+46
x46U4ktrWCcyo29EsZ5LuRxO+7x6zEzMaK0RGb0CgSdkrgslF4FU+ipH06w0hFRZzwGO3Ya5wtXK
qaInsCkoMHusOGJW4wxp3ueiilR/YMP/lrrmVmaEh7uymBFB86rrYWjiu6ly1kdBK+6jnvZYWW0u
VVTDlDnWd1uLiF33sLoCblz9ogurZLyPIO9DI8fAH9WHDO1LoBSc5T+EvRWIM1nhQFAeA4Tt0pkn
roDxgGL2DZHlPP31j7V4AO9sP9ajjNK68256irT219hfqOV59g00Dc1eggjpfhp+cNiEU7mLWOb0
smlrne7jymUL9cXh0qr91fOn7ydVdhv8JpbAgZ0TmYw5rwPH2BQr4KrbpAQjvIyHZMCjGiQFWYco
aVHzko6988H7FJwIP/Gy3FRAckHOMEFlrNyRE5n37xVXoSnBD5kxreETar7+yd+KRVhHqS/tDKoL
KpIbkfdLc8K/fBDoNCR6Y08lzNw4/PTecWltdxD/x+aX0486aPJEPQrXcd2hiXx4soGurNzu1dXB
6IyZUdNUxNggblO4WMyLvQcQvrO2uEZ9FHIs/CnXNzdNS8tDVdqRcoq4Gpegy1YFuIKW7jgBwtoY
6Pzg97I3av3JmBwTOYfONA96ocjp+nerbC8+7E62fc4l2ErCSJdSNu/pFrDs4lW26lmpJLwFqOIj
tDDjeVaZJP1FenWITZUYqDButb5OK+749TMm4uDeeFCa7dzbAqHkDmEHaMAwCn212qWIG57RXlra
G/plYVJVqY0oueCSlUqLWbx+L6rddVZSkZqbm+y0jf6wkUARK9UNVdKikJ9dHeOvlGVd5vGwb+tl
8dlFh7IRjsY2pcoMqRTwbsExpYXfok3tz/nDVeNjapTEn7HdGAXL215GluCj4FXFZN4S/2zOWIOX
Oq/S3zpEYrAXGw+p/NnfPE679Wsup0qh7v5xmeIRR+8ld6uSNJkjlklhsY+IbuOFVEW/xxWr0PFl
hSUW2g7Sgy9Qbxhy0EVONy4+kseGTa4dXyK8L4QvR1K/J9hhm7WTDnX+faBdBhhyl8ZlXIVH4M2p
Fx2aVUH5OABcn05WGa2O5l8SXfPAnNpFY6y47QGQBrWRgws833R/0nzhFxbYby7UnfwVe4JRePNN
Xosu5A2abNu9VH3cbv+CEJP0gBpZL7p+N1pXALF8Ktl3M/bIWlNUbU4gtBm3nprhtlFOgsXdOqqT
IDvsWuRGtGmwXjTi6h+7JCEyWdRoKXLUXEWUwtDuHq1z9uUwH40HGJUCRNdPBTigmIo8yqLEItMU
mjhtVNP+DMYefJ/AQqYlSru1WlDN9dqYJv5lFMp60JldnuQgdnWh4C5cYsu1T5A3+YuwGzYa7SHs
YX2ji7bhem0DOk3Mkac2I86GuJGl+LmM52i+8J+wbHnoeAt41hPAEw5bSkUkzt03cMYf0qPIMu11
kyf7/BNwT61YWuqCxLSnU3D3gY/fQWiTY3FezRiMsCIXfcI48xDfpDzzHXZHrTbPJgxTvkoQSvA8
dbSc4RmC8cJsSFZ0bdKxegrc+H1UtuswuSrS0+02Woi6HCL9LZwcCVtKconLrMll0xJ1fQgUPg4d
VYYoUfVoNVAOU5aldJf3NW3vnZNtRhKPwl1dAs58492PeZ4gKbHs/9FohKRHFBhG2y7Gs0O2enzA
JjU/u0JEw8xcVWVbUH3hRcUkf6Z4J1POMTdbywiK7ibbVE3J6udyDsQS5jdElzLgq6GSp1xBj+wH
MMHMc/GmlkruiF7vKzyt+FjDW2qLxJXrRKnstQvnKmMxQUS5TNmduiCAAGoKMwcNFKo+mWUa3AUz
oUp0yq2mD7p3i1h4RA88UhXVO6R6Ci5bTIm4aoJ5Lfq9triktGtLy3wzNRpmFAoNO6TCz8xhhfqD
OILDNORK7nEJ2XIqP++/3LMgkgdBCw+udN4bTpJ3K1+kyCinJs/kHMSaVFOYSEegeBjOpakfLEvA
fz3Ux7mBuP1YjQSj6ScyM1JtnTSKOwFzHwNbkfEKtFjQdMBh1UQulR/vaN6DKXATiEk/F1bPWYqg
j6BsAUXOvEFw8/+OATuw0jgPGMeTJeCxv+V04RlZOUttaVwDe472W6RTE/IW9/EkugZxa0KH2yCW
7jqED6yGFBhZpe0RqaSAjyb2guzD5R95FQSwO7lYGCV1WD5Wroq/omu6soGxGts48/fi3O7zFORe
ll5reTVQxdpk/FywNrSxWk7saCr4cOxxbzg+hLGJr6VhAzk5nLFaFX3FfxtqK02PVDVB4DaWyncD
mXKpF8G0HY6Z6RVKjOsmJABlrtTDQO8rSR7E2f4g1Hf72Xrs66Hk/KKycjuIiC7VMSUIyfrOTtRh
AazNzmqt4HvjdHUi8Y+BOyVmY0BCd4Qik9JRot1G6VXPEimVEJvTJ5069y7V//rQgSrVZjanNsNv
H2sgwLaw5zImJy3e6THkeaWsZ00qQ2uO4BPaLPtvsZSU7XLPJ9smK8Y16UmhRCNlEzktOY9rXa2g
faoFE0bVbSObPLydRlX2N0NRhoTeoc9IE28ErOubUnU1fzUWHyj1aaqdnlwZ7grnCObe2cvpCd3t
uQraloAEGEwQLPB1fY3YieTnEnVF0B9R8qddBPQc1qWvK3NAO/ov4ZdCshTsQGXvPwFBH4DGjs3H
IhcbjiMndOTIjLVe+kKEyzSdi/im563b93thLfPeaNngZxesfl/HYpeRiIsDzvLGuXOnyDiwSoR+
6W/jyXG/9I+y6C1OCWiMYqcWSEr4j+qkeoiAhF1ZUva5xilO8YipezVSpjYQ6M7ZlI4ENS0HC+Mg
UPFPYd7gukjPywf+ilMxHLKv1HSNKCLBdypzWvxNdK9x51+/nj7x/Ix4A+oKXiY6f1ioNjtjVlNT
BO40H4FSGDzNMJz67fKA/Ud85G91gXVZ0LZfrHEAwJaR6nLtycrNvI4R6KteCA0arznVl7SyxG38
z0SIdmHBfBH4YWdqLHNKiVBSzrVjlzVAtTx0S9TTlap/+dGvLCuDZ9N9yh/Wki/nlwr4FDQma8al
kgyVNTaWsthMyvIvFEnsr21cQ0kH81SkXSO2vtGpfmw2VFO1fbcztDr0RLg0H6HAaZ1GTGANfb+u
pKd6ODnHRHJ18T4QgR+Xec7d4EyTdMBfswfGDvgKC+FdNETpETsIXP5BTBxwipUMUMP3SntUehlf
WoTYPk2LzaBff7Sbu+UhTWZZYiOZvdAcstH4eoYKrgv7oR/MRgfMHoq787ScPjHawvUmD7q6ThtF
hLw2qmWEDXEKHvTeMJb/FVSoUhHDJ7qNjr4v53F6J/qfvz92g2PSEFOrQbFpzfirleu9wM1lc0iP
DeqUPsqrZBtVNptdKDmALYh1foedu2U+iS9Muixg+Oz/1HAdRBiO8W/a2z5te6+W4+JjUk/gyB+x
DtIU837TN42orbp/O1kzQNJXBS9wZJ+Zd5LZlVGgPJsn19l+n0icLBZPtSvEwQhrCSc2S7Y0qW1L
sRCSXy2KMomY8tNx6tcWHsSwCE2vh1ZTl4g0PIMALZp3MbKvSPqabFhMBKY6RoyJh2upVPuvqeB0
Pvu2vE0U5nhG5rHLj95FScBqjQKl04cEnuMfIQkfIVGGCHmZ7W1FomiXfUxpOjTbR8PIiPuQBclC
Oyn9ZrzuyZ0cSDrKvXQLE04S6fxvtMdzwtzmT29veCqzTe/T5LGvZ0/8GjjMaZNE+wn8IFFM5I/j
PhlSqpcvs44p+EQn0XYVNr6PTDlCGpHhn+nNMdFhP5RAU0b5LEcZf6Ff8RBtopUsjnpG7YKKpEJt
VVquUbWNXyPzgcz29yenTZ5ZsJAwWk/ttfa7vgr/OV5nLaiiVcDmGy/PzRW72JubwO37blNnw6N8
9263CgRGyOs48l2Bdwl1BeYlcCiAfbVkbnSBTZ84fZz43TYAX/fb5nw+IfgjfFA/UehPhCn7vgKJ
5mXN5Hr526qedwco+ea1eqSes47ZdIP+zS3Ns9SpF3d/r0Old0KgQlx8npYG5QB6DxMXWP7iHdWA
sL5WuFPa9Ugb7KH6Xw1DF2wY96VBO2CzH2WAqncWqjoCbOSyMjZaonRGnyYGKkJB/aOEiTvpGy98
eFpvZspLFQt6C0Np5hjpXf6eATZvQL63k1yCVfwJ7H6IDY6RMzaddGuhwRVBkN93XRisUmYyV5Yx
WIib1tJXtOIyBP7Lmw/zuNqwtJPy11afqRt4bqKuLNaKYxl06kDoK0Hj4UAySYslPMfP0JHeBn1V
dsfKfBKMwAQWq7S6bgypf9yKlC/SdGA8YpO3D9mHYPQlCd56nc/iPRC/GvD810CKF6UlYxfI0qXf
oIkOGQ1QRHRQhAoD3Ss6EcYFaHdIZ7DlU98DMODybGsnGZfGFLTaU848r2EYHdp1Eb93xdHCH9D+
WR9VauWsLukjM69iVNTqDU5kYjoQoNducLFzFq7esRDTXj6JsUPjWlascbKQzITRTqpddv3mU++E
YhiXlmNjdIlnTQc2dwCUrztFPj3ZuKc41ABzHql94n2Gw4CPzcEndqgxxjc+gwm66IjGWTj4/Wt3
m1CHCrEMPJYUP2BpNuvOCH/lUoJsMtYDZqLxQad+nXWQNnWRLbrIChwPrNbDs7336tHy/fcV+ge5
iPrzUPzUZFpt0r3sWq6u+M/vxkRmkLxdyOsnFXIDUYbgwdljIvYhqT7MA5WgmUErrGWxxCg/O3vb
X97G0ITKv9qQpqYXZ17Ch+OuVXmRQNlsCUBj0jybpug8EmakC2Gz7XLxAZM8SCQqHaNWfS8l5JKe
L/lAXxWdGYkKDJ3XR7z0tfOCphzzND8fc7F3wy8Me1AlaOKVELyAILhBoMwczaFqEgRgAvy5TUDL
ecB8pDVVj65d+0Pd2ApPDDB5YRLLULIW4npux2jYNJoRSOlkehgRj/jHAY2fjoF4J0ieGawcR7c2
9cleYk68Qyn60vbXoywd0FiUlX9CUM3uH3udAHsf20Fhl1epXFzfUM7LACagtb9/ILtaJLcHIvXq
n89CfiQCZLbzBbwrQFd1ysawHkpwvf3kc8v9XjioWZJWMnW9ynslt8jq/Efpzkq8t4l9XxHeM2s4
XtrQIrTPYogbQPOFHhC02c7XD0zINduNUi8nxCfsZ5j+1rBpZ7xScinjfISIkNHckndqwrW2RMjw
XVXrbEUUpYxs7hx/lX+zkumNLWtbPs/ti9k/1DyAj7UhO4M+d86E+r36AmVKgWu9ymFAGP2f9H97
UxjQnRwXfeiSfhbIHSCG799R6ATSuucGKg/Qgj39279ZDhvVe5BV4f/NxFofvMfLwlxz672Sjb60
sci1tVjQbYE6oojxKTdyaN2G/mh/xqulnzcxBaPvppMxAagxGteQNgyrApMsQFDT5JGYgoLlWD0o
7jDkjYg9fls+1YuGwlwk6iPmeRS0hQVZVXyGdA93OzRjWnCi0J+w4pq3TiX0lFCQalhIytBmK2C2
YXarqSuYObOB7eFi6e32/Pvg++sdjPsKiNTpbFY3Q9wXAsE0UuQOj6fgEk13qeSgLWdOn8ujQNk2
ULE2ZWJMNfNfsJInDE2nnS4DYWsZjIMMWigaoqiYYtiUwSxrYJMxbBj2kJigOn0NgynuriIE6Rps
91woHxeVHfhlrfbDuYqb1BzSupQVxwQ8Zk7pSrF+XA+k2h5XudMLyUguS+Pi9uKTCU24Dg3yTpRb
N/rsCzDEYCHVur+e4DwFq54d63mI/eiKhLUOpPCq8NmSlLGkuAcAdDoOkuvkqcg9Q01f/MGctoxf
6W3gC67yOK+p5hboPhDuO5Rajx2SZdbwWs7YpjF1D/jKLle4pPILf8k93q7XnXmRGLpoKhEQHlSn
IJRfkf4vRaax9qZzCfBSzYyqJQwRhT4Qmnpax7vPIut0gMmBeI5WB5nocPK4XFVZUsQhzT2geLwt
LRLgSxCmxzHcj5Z5JX4FocL6yM4Bf1GKnBfN2jCh2Ua81TRPcVzh40er93VL7eTIIY/IMcizqvM2
vPCryhSWmZAak1TGIJcMKCwf1a/1Ua1c8U48f0ioiXhNb7jDRHsmhCnwV33zr7d6ykxkJn1LKirP
TGp755ca09/SshPIRAWaD6oHFuCvAqq1TGISHcBOCrHbSnE3Lc1HR5u1pRGvtg+KBm7PoR+kZ4Yu
PfL5KDSRwwtb3zIDfxsoEttSMV4ibs0wx3UJYLKNpRXbpo3bSpuQtvnTbZdoMwfwooiVgvKwmwtl
VZy5yq0ozfeVzLR++b/4t5kSbDlHYZZOOmyRWtVhMW93kTneNAu4UJmuK8CZv0BKrZEoTlXRz5pU
zeS/dELFioEwb6391QTHR4rhadP+W0eGaePtHXXWblMSq45tncsTHwyd6Kb0xDsxhtlXm8Gd/vYX
+x0jy+qFk6UgDSW20lfRwl0c7s3KGhridsNy5p7OsyAKA/F5NdW9DIjcQUsREPCGTFT4zk5Z3Ce0
v5L3XXhuU8JfW6da9bCa4VdYe21YrpUnaSa81gevxdNY89cpgaTfHCfne00CLa4TODlk99WQDJC5
dCyBjkUb77MRErP4AFkXGASk9yYkD0sLHP3fA+CsdZesfdjhmROmXK5lny3GUvT0sLi5LlC6jApB
ruYuGrWNESlxwyK8jEjMG0qBkyY7jeI21CmZXzkBfy+Q7gBh7EoDU59tU/HviAeGfyp0jaTBMt8u
ZKx1/mqPsegwQNtsl8qfn42fxESHiD+JFuVytXeo+iW4QAno3PSIcYHbjtBYvVewEBq6AX0ghAIR
KIQlqJbHHobKQQ1MhtnFsKrmTfQxhNHUmWr3vh/Z8CXUEUvaBTPqnRZDTjADFNJX6vOGZqeScfOz
z5UoRE9WxVVd6ZeODr5lRG8x2PR7JPon9pMgHYvIpkWSCGTxnx4ubgp/Esvg7taMMVBjnvXOWQ53
/Q+QK6MHzjm3fWVaL3u2I7eqz7hasmhwdB44YDV1ve9EhbC1UGbFU6//LENwz3yNCC/J0F3m/TkA
nJDQ5UT4D5L1Ns66D9TYQYfp8joS+6WBCpJKkbN18Mn6seu64SJsZ/GeKZlamQ9p/DmYSSYWLzXq
hhgQa3GM5I3pb7hAh0+Lcz5+Q7P8iRFVzQGWpaKGmtKrYbtBwLl9zms8rxQEAf85V9Sl7GJudbxr
UKu/z6YTRHqt4Cq2uC8vtRqCQvaZgwiO2bPWzW4RORQITkSsJA6zWS1tIuOHwY+jtKrEVOMeVcwg
YV9VnHTDZQXtzJ3S00UDf3rFlmgRCDbJj5Qb84dY0i02687M2Pdds/sqL0LsOebIHK1TSw4qk3vR
B+pMMAUVm4ZZx/6AbWB3QyljYFN1w5bDwNbyE+K+AuoSEWtZJIr07k2AVvwARaEWXnY/X6Ei71pe
EZVM2T0NWEvD7L2WZuTgGQud9l+oY4TzdK5eVFxF/FiiIiWI6rt4p5pkjsWU/MF0KqL7vmcuxgoB
TStdBr7HAZgnjdWLVxvQizgsjfPlhTCObQ3/WPBapUYtcC/SFm9UtRjFZq7jiiu7NgC/jkNNaF7m
Aja765nS0yLxzqMIl5QS5Wd1qLaOr65xM4ap9N+hbHjBDZNSRuZf7N+G43O3S1HQU7fbjsjOhVNq
l4myaet8d38qnZucdalDfF6DSyOSDTpm3Sbck4AZFN/1nlTMGnIaGujq+K28ZYsjIVIF348nE+8b
SZl0rb5zPvhTSmJaTNwl3+84jA913wJ0AWD8WZ5ICt2vrGkpg7PZRtD3hrJC/s31O+CH2ND0xkUD
moBn6TMqReNok9i/Lz+/8R6iTKT80GKRWS9/r4iPZUzZIceKEzxD5KfszZ+NaPoWjVUTOslokcYi
kv8iI+e6YazNXpyKMAlOD6B+XjmyyRpDVTUqd+WvXDHAf7JTKMTdtNiJdudodfV427che42tOJGN
dhVPeUpB5gydwQI50qfUZFqh5ZwnzmvnnKfjWq9O+avBwC99sdjEpwDDLTk9ANDUZrP4uNce1Swx
H23kPrG63NMRMFrXAfi/XOi7Ay9ElL6pQlsU4HiYEinfbgeJvCH0HVrC6rpZgkE93IJSG8+zcbxw
jkS0KXn/7dDzn9APJIjefHznmZguh8ifEXfinRfL1KO1/ptJU07yv9eouQEK8pzwa9qLpPM7QZnY
1ZeVfpMlKImuGoohjx354HMpIy4W7eq6yUOszxH2udZCHYIrFaB4fAMZNNjout11zNrdReQDloki
YV655+LjvcI7Hz+DHN7bZdn/7W6VjWVCgTXUScZKfIGbd+T4iFNccIi9zwVYOnshrWRUgaqrCwrx
o+8ZH0yiP3NqRXfIx6Z/TUsQspGPnCoQV86snG4me6tAWnvSarq0Xen+RjtpwPA+GgUWvtBoP9K2
fsIrEkOalvdiMdcPhvq8zYDcS49JpYrC+9+p789ttTCAuk0hnOAruptetqkdGnUBCRUVBx1/wiep
BxCkSX0PDqRFEpNRfKRtVbkfcXYFvgKkc4BKQYQCnFYheMki0g9iPU1CETHspzBraQbQsTXrERxx
UK5VS0lVYjzarTQmHCkIuwx6WlTN48rloVyonk5aGG7XGMqSksl0jQ2UOrYe1IeeEh9gsCiGEnjv
RQYjeTevLgSAgWKo3+DY+YIuoRJmUOi6lcn9VE4Gxaz1IgRjypEBvcXyxo1+hQNplZh4rfjjAX7S
Gk/t0TNhP2VHQvsKvUj2qseADjUt4F0DCj02AK+9SZt57eYhi9XtRU5/8rBkdVmuulJLjcUJAZZy
2G+TZJFjGfK7kZOHal58wDMvhIhtcdIrVX4A8qK91bEj9VTTFmailQLpDQRp+jZKF7a+LeZa5lRh
7/YZdMzuoh3GRkIMtblIVhGz5RAEXjVGPyLwb5dS+MYdONJ8rbqrLVP+Os3bQLo7IdKLy0PDNvxU
eXjwDW7Hh54uIFId8MUFDluq2JscmVzv/zqPEdX397DN775RtiCmHL772T4XLVYQ7w2z1iB7S9ul
OmJgnVls11uZEjVDC16BQxdM4hrYCsfNMMRF7sZTc7tXWRDj8vbgHFIuJiruBeVzG5TSfWOl0rOA
RvnOd6JyiX/yu8SdUPy8j8GSAuTygtp0gaFv8/1chKXLjbrNHWoLnLfH3WY5tKCRSTtWkH3q3Ku3
tjnnW1Nzkp3MOHW1s+M403uuSEvDEZt/zhzl39cjh13tbx5ERJ1Rrtw/wU2+vrSxk5jaHGYAi2eq
4ICASrOGNheX83AzBo8MqOD8zx8dEiFSpn7h/KtiFbSVslOwE18bE8eBCZjTbsxftskpM5ollfvQ
sMQjL+IAAKRG3LlGhCmg9P/S/uPmjNQ6iEHveT4ld3a2kU1QXbEQJW/qmAyk/fmc6IYZVSA0CCIt
+ay5XVshNd7w4EVpmWZjQF1JwAFfgT/au1XkjlaKqJFUitjGKfhcp2+5c9hpCrH9U8mDUoCPoxub
zc16k4ayqMNbJ1koaRo8d4dQhZjI67HGlvTlRaI8E5/bfUBVN+zTEiniQkMbgxL3KmnPrT778Z7F
bRGMpeuRKrz6sCRQJckCkR3dDjSmtL/uDJIHlDfnhYnddSSWn+1qDe6fFJcqrjzaJgG5UcdgokNr
Pa/idy/Khns0aGTTO7Srgz3lZ5MWsoB36BPYhw/OYNQxC0lXwgfb0FS0cBVrcBRrG6zs4YDIgKjm
klvUPxQY+vnKxGiBWU1AHSbRbWpfDk/hbljne/NXJehWPQB7cpAvuZiexJgCNVTQvS6XtebVNKYc
f91sVlV7AxQXu+Fo/auxy6xIikisIlRxnfW0maKEOgxPq7FqWa5f5F7b/T6tYN+sAK63is2R+ILQ
faRcJuW43cPOKuJygDq7UOz6xTPrpthgiwdrdE5he/IrhwD6TL0fIc80EeGiFWdXqPQKSw95TUZD
u8o/W0lkaKy5ome7z3WvgHRtY6+r6UsczUsIISnZpBty6BhXG1nuSVil2yXpR3Tx3qbViSrcnoLl
tgeN8lodSF6vyFDBwIzgoDMfwREmZ2d0iclV6u1yLXm7MINyMG3Fc0F0M+loS0vXhc403tPOV8Cu
71c2C2JwxYu6AbduYUfSJDzS6PnG/qAzXxQsb5FAlLcUkmmQkstMpRYUeDe/CTd+TxsINGfRTU1o
oS9aQJ6HyARDrdcKQWJwaLN0NKAjsEY4BeLFVkYSiuGlGddhMsaa14rABVY76hDqGxWZmwZ+SMIO
xVh89WVVyNYJMmFiYEievhNH9r+B+8ZY+2B950fT9EmUDTVuXpph7qkeO/4UI0nmOaQ/QFB4ERZD
fp2G9ynShRFDVfFy7HBGr8Yi+rXEb/twEuRMgztuxvpyN0kNSwb+Td/gA1NjFwYgFMLlTpRU63MG
lM5tdniiy5HCm+AGGwhynDXs4cEV2akvX+TlfZAhqwNGm9q6qtWRK7EjhOhixCjaO7hWxrsrd6ZW
xBsHSSjL6TW+zIuRuATqULxR1AmbhYVuXq1SBVh8RSr2Ne6So6LSrMYpRklA2mmJaLVTVfe9AIGE
FveyP/sCKZckzvt6p46nXE41rM/G8CufSSod1TPpkzPVg4xCjsGz2AhvN63qUAYEIWMPqCzucUTq
lm3Aryxm13jmsaplWyn5sCZtWJI309OjUzZ4AYP7j52XXBQw8W3iOG0/bsDUPdG7T0AIIA9lwQys
0MLIbILhX1GO3U9T+9isBr6Tdv3XrxwpydM2TdHHfj2f0mCrv/8CDWn9FgLwO6jJQTG58tQmUhVn
WysaJ2x0XTmbwaC8bEoHxyHMUaXHdaTgzxszTqQUnpdGizMj7XI5i+Ix0hyDjy/mWW76UuDnDlVN
l+AhIPKRk3g9kegdXq14R838g2y96hraDwaaOzE/svJqX7o3RJI5ajvdkU7tO+Jy/rYF0vSzfqdt
55ZbTQC+n33gn/SzxABk0pajml0ff4km2nT2mtE2Z9B7nyWJ5BcnBP7fsa+g07/uuVX0tqIN91kO
+mxvuIXTEWsgKVIWxDGC7FNQKg87NV/B6f7I62aTCVpLfvqiPEyV6a+hpu6BkDqloVPvUYUaValW
Ax9HDUqoc3Lle/Ii02/BFSdWtack5/Uul0EGKK4PxoPWNfXIt8DEDZv0SHoURQMFPhSQZFWgylWY
bq0kgEUGDxQOvoYBKG2foTc91iPtbF84fCJrgHtmakPgqLOXjOO/6I68YMjNgUTeBnEXHWTJcVYd
H7n+KkWSUb+d8cbg/NV150llz1V31l6aUWAN4Vcb6o9OMl6PBF0G92ENNVBOQDMGuEy4Xl3hEtbi
tJg0m6oeNd8XdBhJnJ1uJqHtjt/2VnQT7sbeL+3ubVgLTcDu8xmMXxx/OkxeeJu9JGZqcXMJChxD
G9Jj6TJKC05+so11h8jkF3xOy73wTpotVxktrmdXAv/tTJm9gi2dxY8kQZw3LTr3zYVXwl21U0eD
Ie5soDgtB+2WL0oXBQLGVAZx1b2pVfmSqQKmd01vnxVTiJ6v0dwuh+5xWOv/kwrqtbTMtpU2ywpe
PePlzeCER6pPORcMl7vIIx9vrofG65aeIh8lAjyXFDbtrbEofuV0G4BJpCHeWcAZWLZg6vwOrR/6
n42G+2wnHMqIe9dIWR3osWZASOq5EFIe56W+RNXkB+HeY1I9vH4GlhYH5lMAXfwxOE7mMMX5docx
1i8KVvrRd5glAPZ37SOYGyXedqhIyC7Stm7I1tyuzwNtoi4iihVlXWH7XwnTmqOQzRdDq7yOewxa
6SbjZZnt3mMEqJeWZ9Qgi6Gl3c13Wvw4lWJW6F5/FuWr4L8cHediRGuUMH4JMU+mgEgLPTqtD+kw
7oKvijYUbmQBAs9N/QaG9VgAWxS7GzTiZMSfnt1VTt6blhpZ9TX5koUCSrraUlZkm1jHTE/hH9jv
GPhEjPsI3KVbmiywdFN7xAeSihreGKSIA9YibfmCRGLLrRGvA0rpvM31Keg04tCeC3iFKxAXCqhN
K9RpaIA41xNUIu4XEpERJx7pl/+AHQ5betmw+GZzpawpUCSzdJ7UTinjHMS7bZ0p54n1FjQ2gEyj
4pqiJDyqmLHgNmr6NIb3KiD7n0Rsv0B2boheRVHOj1kOfUEvtxd30haI05p6wMzCwDv91mnCg5o8
pyXhRlFXM8fEtzmP7PMYFNPXh7CBLynnxdZGKTb/AfHlOJ36QpaH40bvflNjmopdth27x1y9H4NJ
dXrwwlwv3ZqljNk5fZHdeQZxIYUCNctCXJUhCxHgvJNxnL6qMRygzJHzPkMNgaI3kKqliJhRD1+r
HoPx3uXAzDizFtdUZzp0GqrOFiyA5GNDBFxl9ywIIb4mIAdr7fu0M5pMHZSWRiu5Av2/v+mrmupN
tka4Xi6++WpE2NEkdN42So62k45kYTVnJApYvh+Je8cu/INBqjpLvxbzv2II8fh5SfKRgDJSzVAg
TG//oiYYyjOSRWLMrcmwlEQosWlt4yfPfWCdGhCNRVilue3mPEQSkfvg3A+zC4JOz4Qbw7hOITPM
AC2zkmOopvDG85SNjlED0ffXZINj+/8VhhhSHADFpdyPRDNmvn7Z745RPV/p3H3+s86fm24Rto/7
wAKyL/d0CdspB80L+NouTJfaHR/N71M1TvW/2W5wagipge/+o6ceXemPLe98CX7LcQXNo9kp3GNf
tOOLzy5B2d7kk1K5K9pmtKPGRBTi23LXx7N3myeAKLvDG7jG17TZG4HMSswPQqBXMX3hiktCIrZG
xOQz25yWl3SKyMlvNvSp8rNRy4uUg0rZHWrKF31cHW08hXeaDf2mzHIasvpF3XPXOLVaneXg0z6k
zgQvuZablHJHRVortHjS1aXoqhOlOrLJzK2mwPFgcZ/Nli7dy2OsEAIwzWE/RpjlOUaczMcb7nZN
O6t9uAUtNPU9zNTj5a1l5XpICbRvGbeR4ASC7wqlakK0zraDLvyR/C8qRihwFFO/AbQxIJYWig+I
9JL1VsshGMlVaLUZpJ5Ax3wXYFQfj2DE51K36vnyuyXVReDW4QNXPHO+Bez4/0KtP3wecffg5btU
7egjCDyIQb0zgHG47OzIHCVBlQMJV26Hx+ObO2A2LRHAoIRurxLCwyuVuNHpUk4uWx2fb76RJQ5Y
ihOHx0LtMNEZaoSEDiyORItC219lAwj+0MKKVFoP+KpkRCABUQj58EXDoCb1Kw8oPK3xFDviT0uU
ycz9jUPwiKf44Wxwtvjd8jEQVS7gaKP25wmFOtoe2SV54TV8K+n2jKEujyR3+K0vhS0Xcn6hXdvP
U0E8r1o15cIemjKGxmc7fXxQjYlUtTEZwFFIQNF2J6pcFeoo83VKJKYsYJFrcZbNOGjK1bmGYXEO
z8RawjZEQrmfUxm59hewCvcwDldwrYQYRFbgKpfl/wonffkRyqRW9b400UHONoZyRs/voRdsv0/l
+42Wu7HeQ6HUTryW4LtFjHHn8z2norSBfzq/wzn6K50MpZJ/4h+q4vV9/ZXckq2fQY/qmO0auxCG
RzZaKMy9Jl/SV8ZmelE9QoYVS27fwtriEfrAWXwb4II8sJuTpv4xlRdzlVk4iaDTIhRZEsQyC/79
qMPjrOyE6FJWhrij4+mYvOPnX2aGp/g43Rc7baIcXf5ZRZAYX6ftNb84vcVm2i8efDUMD8lw5Mvq
MjA+KpNyMBycBQ4xlwP+WfQrmMYBr3n6DHOHrZYXNJDK2NxC1ciyd9lHPUBrkPBf3TeAg3sLWHmu
boSunEqyJ4QtRUW6fFujuvD5uXiAAbkxRQorsQfrhrm//o3jzFSE9qfncZfy8vEaeWA6QsBd0hQp
k04lZPrp/Wlf87GQr8zh7Tv0STxt9wb6KYe3t99rRM1h/ouqu/Q/s7mnfokLWvFIyLnc4BVjVDeg
puNQLvls+f1kU6oEIUQPWly7RVMgxGx3lS0cM5hgjSlaifn8x/tUvTOTNqINv38HZwQ4Lo6sU42o
S5uD32WsLi0seA3Z0e3RY1PIO5MiT2tb9IPx0fuDkd3autczyAjJ3XQEtb44RWYhaYhQSJ41udIF
eBRqQUO7VpSzeROBncvyz59ZXZyRzUUOEhtI17+0TdixpNU4ewTcNIyChk3JkYG713AHYpMnGkjP
1BDneaEpeQ0zxng5tr8zMa/76g0WFQr346znrgDXSKR644RpD8F836fdNkLnkFHnHJ9Y4RIUWu+s
5uXvTBe5YoFI0A57G0WR6O8n5pizk6zsDMxMkreZ5qCzmXK5Z/7aZyHW6DuDQka7DqFYqIHfpB+t
7yo7oxR2RmREghZClzYg+uy2gnAXYx53jPf7NsbAMP3P2crMct3Sfit7URYevmKX6XEpC12B84jX
FQLzAXt9WkM9fFBnGIfZWPJGgtGAH8Ff0Ry0uLbv8RGHFdD0kN+lAMbT1BRQ7BpiIK6UFB10L23+
A+PtmdMpfVJJIrhIwmbQi14oz8wSv/YUh9hH2TH98vq2s/XCR5NRGa0z6nj56+JTaKKYdmRT1QGn
Tls0/dK9cTuemHdasllGm4FKNwwJk9sfBoNareqx7FP77SB7ToHvQLB++1AskTNgZ1A45TARnn5q
47zvAU1NWfpB+CQ3/a9tClDeOkU2AVi8LTpAx8wUcIJd5BXZwZuYDlhI/bEyLSEwVAyl+Ls8c1An
08loSsgTM93NHbV7yzXJ5CYzyn+WlwmrDxLHgwWpRZldr7b6TBUfGa02sFwwpx1EAI5DhoMONQIA
cFHNvm5EBgu0X2ubm53RjFVN9/wkWKIbfkibTihDf88y7RGwphk0B/0ZpoIfyLLSGaBKwITLvZGM
9oHVyQiiV5IPxbQC75u95QQfSCHAucFgmleYDIBhiA5+7IaNswL8aujD3kCHcFKekgpoc9yEiKYq
/5q57roHlvctUQFnNIPe2rA6ZK8aE497EEXpWfYQzYCyVUGstjchgaaeDydTugp5PHPYCBL5pBAE
3azcYe7DpWol2HIgXrREXv+4xrXapOGCnL8N1xkgcr0sHk+onPkplDjj/pPb3Tp56K3wVWgtCbqi
fA7bB4rCA9AnbXk6idVWYFGoc5OFhWLjhzW/QUxt/6OH5iBFPmu9FYPvgmB5LovyV+IUZjsmGW8R
FsfVlU0L+PUk9SaG1fhB7hDFBIxt0vWSaR4WPl69qCsT3hc6KxbdGamxbmteZkaPjIwn0OVszds2
IX5HEHF6bNlXw+BFdPZoqGcu1wiAnIj6mwDH0sHgZourUFWTZK0ds/QS85bw8HZuc1vhUEQ7dKRI
ys57lddnOoRPBemy4LNaAsMpzK8MZdolmGSrS0EsgMMyHo68vqP/jpjLlCgGgpAvgcjOsrPG5Ds6
luN3Mqdg4T7iZJWkOxlxHMspRMnsc9PoS8MLpSWOjwtvk8TWIsn9ft+peRRVTnB2buPvCM/RxfE/
1EFqujtam2C1nhACZwGhPBI1F8fNtSpKBDxocpYC0OaRU0uodBEvOCpHQ4XEDrNCM8ki5zK70apN
Tbo8/s0xscZgrhNzXO1CxkhCMrzyXGF5Nl7Ptljq7xgGnu3nvqS7q0QBjHxuUGi4ASg290lRllZF
Jh2sDuG66VUfRnpMn7XzIIpqTEOxZAHfevCyszJuhKyrFdKEClpt3paUed65Fa/plsv9Euf0aTW3
5l6qDKn5yjvS45hmO61RwX+eU2JK2k56/JGL8EC0WWNPf2T55nBtv94sAcVYSOQk22rU/k3k4e/I
fQmVT6pZD/A/E/vfqEI6ZdaC64J1SIFndr14eNArICvtNOk+F6Qr/RM9tefpnCZCFTtX7yccWZKo
tirjmyQCRyIP7pWxH+Aqg95+1LBIHwm0cE2XmHMkvyEp/QGqlT5wsRMd3m+2fPrcA0Yj/JBbeDsa
jXLKDwy9MIwKhiakTdYlYSS6UIq2jRSfwgsPi0dJqEtowbwUSISIawjrYxH0JDL3dOry85fqPbfg
wVURgVo1fwuFQyXxuQxzl85E5YjBXYE+DSLSmIrOZq2ptee6OF7DLAdCbnfIkLitXCAKomasZePz
Ov3YzWxxLGleB3fOyrLkXAl/OEtY9jc58tCwpdcu0R0ABE0hpldLt8mzrHhZAnQotesMRybnFTDV
sqT8p8yqNoBQ70e8/h0SXS+/XuJR6Zw8cXO/Uxly/koTTpGZADz58HebFLUscYfxZHfWv2WvAdgW
RtiiNKsquCUDkjP+XnI2iNDgUPKZWyQUmvm7qkQc0DfR5StRn7/Fz2MTV6BCmeGgysn2PUnqG8ZO
xXBrbuV2MwtIGq5sLT70F55hwUBB/Nf7cTgSCKFlUNe5CI91Xg/e1wWFE97LhbbM1hFejhkK4dxa
7f2eBeXqcTPTFhnsJyx9rKcmDrXbUWQXcyQmbIBEdNsX/XJIpOhSQFafUiHolFaSV593Xk8w0nxT
ci/QhOuy8TlBZ9KsDHyZGkAOmGC2KfszWtTUwyS6tYrxXcfGf2wiuJEw+/4NL2qteca0ETt+i00+
C07S5AlelOjWsu7/dPMQTryy9lyM2G7leoS6Nux/KqJx2xLmbOG7vLV4SGXH6If47dWhFy3q0JxC
5J880sKAGmhM/6ByfEbC5BSXfh5/lUoOMoaQbqI8ItKSLSPXYvZFPiNW1QAFeBg1y7o3XoVEYrjH
4D/ufiyUq1xTNWgyVa07STM4kWnKCoVYMLW73WpIcpN71cjn+hEv+waagcVPzl4761Qcwaiuai9J
qm5WBaAtG+T33f7pzP8VrIZJfWsjbZ58cQq5FiVewi92W0tBS2P4zuDYW2eJpR4m12sutlHaOYPq
jkrak35wQVpHHtrDzg8X3xVOWF6zm4lV2fRjns1k6aLv/mN0D343NKY/1C3s++R2yaO3d4xCgTc/
LMj904bdQJsyhAzGdMZsEh8ZTr5yCXFBqNbSFHW54yxlyrkZ03rpXHvhnv1fnPDBB8Px+sZwtRlC
otqQt7q755Hb8Cm6SPAWByNRgSAIDibVQlkn7O8z75/+aX8U1b09V3AL8iPKutGujDnP8j3UBNj6
Gxsr2SfI/28vmnnkhg0Yne+wmecx29gPB/igHNgD9pRN95XviMf4RJ5soNjzFl+Yr2La9af0Ig4V
J/qJkbc3sIlzFUGR5Xzg/FDRPuYl1JQq3+u2luiZtyojpfSbuZep3vcfcW1FkAnUB5nBIvL0OLDc
QmMDX3p9mooorZGLSCKDOA69KKpGLzlF4tm27w0qA295mSsyaLLbOvQdHkOL058Fp3Ko/Fs+lgfu
sW2jScxB/s0AUQfOIyzvMJ3tJD433pox+oq+YhFkeYIumG3nkP3EWlasOaTVel8B2KUZgEzC0mYT
9O7pjLNma1o98NyltaUqfDIT1cCnwL4PLRSlIG/ZQYY0KldndkfRUtic3+WrrjSXD3DqEkGGQYMC
IpjAAfFVgMRtkoWsImA/I4Tdw4UKKCl9iI/lCoxCdXlNcrnyzb8Ad1v830O4qprzR5uP7X+DKIad
QFhkeyUK00LVW5RVuNEbvVca5gHULqkDOvhuFo5bd5ldfkRbx+4Iai6rRWfgkHnMQds7nyfqFlqd
So2gnedB/FTutQYH9RM2RALFeR4mBRNw8ssTrqT2CRMvxVfFyvw9n3kU3e411LfkDTHNiEG+COle
VeAwtSBbVhKjUGQ0e7ms6Ca/0wpRKSWs8T8G94j+NLtM30OgbhYjkHguuMdWScSdUlYIHu0p6t0W
qOG0EL7/f3I4uks5+ti1LvlL0Y6b2r04sC4+AbxbvFR6Hc7GJAhbr5vEgaIX7al/HMtaBcc7lLjA
sBQC+MHIvJjx4QQx1Bzh1TJFy7Mz6Kq734bgFtXW3y9RzMEsiEpLSM7uOmvZxycKof7aDxjUsZSx
AseBiccywtmp+GVGPp9Xs0kdiFB06hFbZJAMZhwMlBB5fIdorQk7asqXaIsTs1PEUFw/pmfqx5kx
YxwvQfPS49ybYp60Jg13a0bGZNGoXBDUdwf5qU/5xDbVu+UM/HkCHtWud21bHMKYplprzKgBnbzQ
11IcaE4FKyM6fd6Qxmq/91fT2/VnGvbNUS/76Hwp0xlCNR86M9UQfSJWVFcaM51wATBwsFZl2lej
tD1WIWdav9sxUjQGH+3VUetNPGEdBxz+R3Z43EKZ/6+XCNUZuthBbey4h3QVTnngZmPMU744AGkC
JAnNA/h5c9v9jPaHDqFuVCVBgHLGp0AJSd2hrxZgja0d9SQNPRzGRH7Bx2I8cbn9uh2F6ZIZhCBt
XkhEVAVOM2mAwEiZB2owECIAszopPpeFsMVKz+WagJZfzMpv2jBMBDlxItidsfln/vQNnQmljY/c
WcQVbdzoUc9oXb2itywLqJi4X5+BrqBwAlTniMW2ixwLsHZ/C9lG+1fHaeJMH9eQbyf920Dh37tA
9g1PCSPqHJhaN9G4usE0J1DoHVVNZC0PB0UemLlQxtiUCd+79lpDoDam8WstnMuspYV09Fek3E18
9fZ+Sj8VIdrgaOM6BNEy/+iptndYWpDvBGX+HGY6cvyXdWYu1e17TvWieVni0MP0eTVOTg8S+2Ee
6hhP66odXaKBNkxwhWX2Au1Lie9YEdL8jO4UEhzqIOqATdf0u96vhynyDO5T6RZzVm7/ZBWhcU45
BnCMj0PaaOnFOrWNmElmcIynkXErd+tq/KuLLn3y4vwx/4tDYf24nKQayMvG36m7r6+Qt8C8YWkB
IujqgZlAw2yGl28DxP42XNM+LGBZHl0PIon2nrz0ZvKEJPo01qFiTGVlYiYl79MgOkZTteSAI+th
eLrk4wqbe66NYhC3+Si9z+z+onM/guERt6cYNF5nPIcEqick8Ran21ZPbsNr4j1oH/9GYRCAe5dB
ciSWiKrvmhHSvDqjkXbEr0ShBWNX8yEEyCDi29DUezJ7ptYI7xJQE9XI3T6ka48r0TBXss1KUAhj
Rd4vPlZ6pV53MLjtc+r0OkYgeSrqz0j7eN3hg8sT0iS/DYdkzMVeLBWK734Otf8sPejxHARuV8+j
o4Cwku9IXQNhSNMZdN6u9Ngo9s+lSWfi27ifGANGWZS+b3CzLO78mi297mVcXvq8g6eG8MtGJONu
v8VEJi5ZKH8h/+njO2k8iFyY6lYLB3vIK9KRHYtZBpqOiWkuX9MqHHLBzwtDHAhpJRTeyapQRGUb
VgUp+g7k82Dm2eV/x0id44chNkzobFffHL2vunrIaIlhx7SUOZQyPjvWw2P7bTFGslWMtymo1UTv
qcpptE7PwJMPYTh3RSGaiH5QuoG9LTYadDkNMymGUlsFCifSTNUrRwd9ASkLXknqf1Wtptk7kan8
Lk6A55U3aTlGjmuC/qMa/tAyXoLUye55T9Zh8ht2dVWV9MD6D5lX7uWvoErsKvZbEVW7WUJE8KeK
ENIxK+AdTbe4VuOrJDoUpokgp7h/F8vYnJiaF5PbWTqIh9r6J+dPx65NebLTS6u4F6lFLZC2uPG3
dobNSIJxombn37V+NMrE6d1bjNWHf5xUAX8Luq5t27tFlOffGN5vqpcMGip3WV7VcHo8bq1VgFGn
25BHKyBRsv/sHU1uxrZ3ifuBabPwMhJWJwdKLtpkPZtwBtZ7SArBUCw7Yw6+Osx6iRHstf7kY0Rh
VN5iE0oelVKJ1hwsPCL7V4TnI/xOndzyUDR+ZQ3Z3qy4BXvUe7Z+cn6/7wGIDs1/iw/NxYesxSan
BNKB2ckOsunoODXbCgfnuq5LoWvFKoyZtrfsPGVIiGJBGcjcNjrsChUVdWkn38/e+nKu5X5kkUBa
AVUcGrkGXl8iZC/4C5yBh+A862bibD0kudjIYoDqgAcEC0TSHooDOrqIwJZoRmdDSPmVhmt6ZMXD
NNMxSpPa9aYb+ZDLgv5tfoQ7GHzMwLfOJfSf52YlmxuLam+rMjb9tbx21IcYWmi2/0WEkLp8ljxa
WkZUryeVSlY5yz87YjhDIO7UpAAr9AqQNBphFq+zIK9mw/p36ARuQQetP8G/By4j5jMnc9ZQWKZZ
r8M5u8KL3e3xEEuVA8UvM4DlvNt0IBGjQRgAgDlTEP5942j7ijL9ShEvCbJoHE9cPBf977d6dEs0
Lowxn4ClxMyaz03fsa+f9tslJpphATc72gY0zzRV2MW/vzGX7KRgb9EJsclqI4u8iaucXohF9wfm
ilc+NImsJQExtam8mfZsI3vQ8IPsBRR/KHdiM0wcw0ZOBWLydllkgmoXrhyM57FgIrEhZ3QmuT5i
Gsu++sxwS6cZbP4V6LEK1k57iquWo+u6R3gKSKI3AmPb8Vlk0b/SnaCTizz5yw4/CXIsv9ZEdgTN
QpkEzEn5Jb2/M6rW+Z7ilN2b369hT2ndFQbqlZaxlEQBNm1a1o+4xIDsF/++SPhX8eRxfzCliVfY
zL9NsqQ1Mhg52ibbYU6dEztD4OhxCGXJHXng7GiXHNcQeA57fWSrsu0SXmlkBR92ucmrhZuvOCfn
+qrZfIJn1sn6MFYapZaSciJ6C+bn3uunSvlIO33G7ZDgfBeBPQeaoNfxt62iSu9zmmQ5IVQAkxFD
LapkQdXweOhLpisVM0Jz/K+BEwrvdHag13fM18z7CVnBFhTGbiRjm3m0lvijfjuh/ggMYPkcnNuB
3n0+yyw/ugJjJLTDer0DVTzPz+BQFypPj5DRcQFa8emgMqRDRaA/c28iuU+Ib0uZ68f84MQobNGC
EDe5hS9UYOJADmM9Zzqw/vhzP3wyTq1pgI8lvCKjdNdqPYi9O9XIVhKAxmtarA3OinVpKwtoUcVL
VCKwL1HwzsYheLWDJiAWVjzOG47YyWs+kCiQX2WXazyzQNIWzfc1F5pZz0Dbmc06bA9kTK/87Mma
2d5UDLUnbedTe+TZ+lkYLFxh+GtrwMNrFS6FpbGe4lfc3qyI7MQDDDIQOxkwg1j/hihJXXIZ2CFc
sip2LAoztvmteh1Wy85RIUURx3Ads5tQ6LSMbq1ntzWUWPVaViDTCu2IyZLC9qtmokN0mLbE770v
6Re78ElC8gR7BkPiN35TsrTeHvfiAhs+3HgnmGQDSE7JbLEJ5LVwyGMWfexF0POo3bGXT+cdpM1I
AwxWyVlxjJpE6Cs/J9247+S0HQOEytVQP6sB6UTvGsjJ+3H2glnCFZwM4xbgRarbFQ6v936XUeR9
2eczUF2lvYTCVKibmgiLDtEv+1FyrdRKbG79OwkfsTHg+1AMPTcWcNxNlubugh/oGCdUpUFntndb
IAGYrt7XjBSfC1uaNv/MJM5oyNVMvt4oF0vxwBzwotUAGsAj3y+olfVqb01YrjGgBe2uU3aa0W8J
PH7WQTfStSEia+IaQE6G/ZcCCUUG9WhYqxsuSBKBnv8ZPL7Pn2QAyL4VFAl65/odIYZhX0yUlkg8
2oc4+82mx0Rpc/vlX1U9Q9cRqaxo0IGsgYde/pSey5sX+rBqvX6E1rDNA4ZNB0yJAo+gNycNzSVB
bdUA1cbEA48Q/ktVXIZSesFBx8rqR0Nm/jAUf+F/q/pjNVp9ryBEG6/3xyDfZ0Q/gXbLXr7OKNa3
gCU+/t6zWovEvpSkhgqFvYYP7nOWxQEavJSyykv7f8rFActJLfzejTR5iV3jxU8TbLfs5Aa9CROg
wCkZLDZQIefB5bAWK6vCD3gP3fxamHXUSEMXPtHNDL3H9NyBGDd4JAsG508hve68E7thQLfOlsXa
G9+5Va0lqf2RXY5u2Sjow1SVuZ4z3+fPd+b7+O5wu5xGuXHBUT3Kj9VFkPQ/9XDOyQxWSjZip3uQ
NUtHvXG1doOOsVfuRPrOxrsoRxnSZ/A3bLDsShjizudgaJOPMrJKJ5eVSyO0OuXTeBsWkToJtU9V
v3DKaS4dnvzlfga7iyTXyvG8Cu1EN08Z+nAGcCFjyAx+lCzAaXShQy1WHp3/BpCqRoorTJR6KUri
QCqPPnYzHJjTCcAnma0vj4zXTRmdaeZSfiAW9mCR2J596xVIvA8Fy7iRA3pd5OYbnKnjLN4JcIxa
MBHItRc8RCkLWF3wjbbxTshYWS2r9SYqkL9QTzoCa1A8sG4z6n3f5gSDwC7XXIXN2YNUjlVN5GZj
B6BmDUjS2HPCdyAuOKNsXK2RAA5QnoBwXKhEJ+BnwZtOMhs7qcZhQMO83VUJOeSyhf/FcnLy1+kz
nkZUQlzpScFeTI+hP1jpGp3xKqEzJd5gq72lT/G4Pa29XjOm3MZEWVEUE/YzFvbO92brRPXoPxu3
3qAXM0KLB52ax6IRrU5k6buvnU/+FcgqPi4YKeO3FlLlG0GU28/S6qLbjsjDlxsRT0O4+uN20+YQ
Wju26V3gLfdoncSEfE9cx7U+StlOCSnYTnDWcRp41MC0dJXPB5ED6wzj2um8dBSim+Dm4jhTFzAa
RoCI/KqdqDQH3rdikzEToybm7KLj/htWmtcK78XvIHhA7C3/j7hqknd4bvnToZ9gp/wXcYDFFS+p
jVe1zd64+IUdXvq1CNHPVv+UQ+DXs3sISzAX/A0DCkcU8APcsYQJNdWUQuhDCIm2hHopRG6aS6ey
rTRGhIc1proTVNJDpM/L7Ghw2knHOCSZWU3XqQdb4VPp22AS0ir+1+FKuCU+uL9X7CdHKOrvga6h
5k69+Dq+E6/1Hr9vwZy9vAm55DsXDLE5shp86EubEqcNwURNSahIa+Cnuk8Xo/kbst2abVp6OATc
LvL2peataAHpwQ7xySObD7xk95fTgeeoBmxbpkGg0K3iUWeuUWrQqVUEqmLo+AY5jNU+ZsDu3Pyu
v2uwRT0yRcSKUqGaqKu+bX49K/HFnYBhqp8KQEw4W0CQ/YMPvuWKLsYUwskN/kGmnN1kKSOIN0ts
bVhaXUe1pPKl4W7G4Sp02g8FMWNTf9NPOtF5XOjgF9G+2kXJYCx402Tg5wJWP04uTNuPRkGww4My
DKXSbBvQavQa1KreSJRzq8fVO73im7PA5YL6eh7KyfxkkKUuyKBflKtNisRicJZjxcS/7IpNTbrp
7fSdeOMZ2px2TmSExS9xwDa+9rABEtBSdwzkmIhA3wyhpi/enFwltKnTH4ELxyj3MAjB/IVELiUd
Gk+TVxYFf4nzZZckmbBWoVZ99Rp4DlAZ/yoRLht9Jx+TjY4M+iwzSx9dkT8JCcnnXn5Fuc4KznN4
RyWkqkqLfhHfofWyRBOXW5P+Jy5rCIm1GU5mGpJaG1WhLDxxWel3onM9QJKY9pJRUJgUX0Bw6CX+
Ggct+vnfdh5sLaOIzt1cnjIcvvqnLrV2owiddC7ZucuguK9rEGyFuiFjnTZsovFkxsjraxP2i/7v
m8eGCJ21XUKFfB2QVMKgVDM0zLUC6rQMONrM99PRrcy9zNuQ5muYXxt1JEsv13y8dIodaJL4zy2U
vbbUQg1UA5uWboyleqKHTXzU5zZS4yONIEhBiMicxDaPmTtDeXZ4qxVFqBt/Xb42nGF/q5LS25XG
w2rwIktrPIgpeVZuwEb32u4DH+TvtDxrpBp7nP11Tlw2i5fyXhCn21O2yuJaxbSQIh6TPRHKDVQl
ePwA3xtxx903O6hZKZzXUpHPwnhPzqMVViw/cp6lnkVRsSAWWTDbpe+UnOjh9OvLvafGX2luCv0x
SGsURQARdWwKfkpHFp9k3nKARNfB89Xi/F40crZTTx/H5UYvtDd9hpw/XxoOpGBjDs99soE8YxBb
s7bgwko00jPoFMeYGtQU5PS64mnyllq+QPtOsKIP69IKWkChziZIKZyc1bg1M+QlXMpITn8mISCT
/EzglT0Yc2kRNb5galS8Z+LmoUbftfxfpfpMWhTFOQTwRdUok4xEUHYC99/0ipXmgbI4Zaga8BOX
4h8aNM/QZTIHT3rHA5rDDaDifhI62N9z+Tu71bKHfxhyTbB6uxsxie8SOEyX83CRIHX/1e/g6LwZ
Y1WiPeG5qwVB97nCkKgQaFc07bxBgxiP768uATdjxXLVOhKaiSkMC45fOTg7ZH0MzxtuuH+fJ/Ge
phyxIPkrcQgfG0NSz07/cdxsg/oiGPxYXndMnTcq13L0hNsGBE2iFtvuhkNjYyECK/p6xCe1O1Od
qQsHWTq5JviWOTYu/NOwCBwBkdM064DlWeIZQIULaRpKl8urP0cldGa6ZStcA22qFvG33FY7ibRn
/NYGT3FixLWP+wU8unnIr2BRozUY0W+KdeluAwxRAJYYA8dEFNOLPeNyUwoPRQQ5a/jw9Phxp6Dz
pP9LXZHWqED5702S3ksxCia0BcPWb42P2ZcvKMGYOT+ZI8hOPnIjyK9PmOO0PIVCrCRfcUqk58yv
NSFjQaYNZW9T6Bo4FtgIhElmmxqB/rCiz4avExMQ6eHBeJQVcR2vRa0ZDjIh5mJ5kHhjAcv2IXaO
bsNpz+OeLCOfG37UY8cKDcP3c/5tiHJFeSYQFc6e4n0YBoMLwe1+gutQrA2pKKna3g1D75u4xH5m
IPoCVHq6sYBwdfMq/wtkb95VvLiycCQXSlbXWoAalydWOt3E8g7nlk1da13H29A2LMY1ZjrhyhrC
zJjQEo7qYHoRKdwKZK0a9/8FXs6adF5hbDmZL/dfReM5Tdzjj5nZq+7y6OU5BRG2j4u7Gi4VaDI0
mmc8XyZYX3VX8X988hhEjmb/75rckOERId+jyv8WzglHDmnyRMFSkTtlSWvfGouen1jSG2OQiKwa
xfiqcIt22ccFVEONiIKS2kCr33UTTcsJqz0tZTt99wXJX8fK1yueymvYf1NXW8qB0i9BfchGBD2Y
de6Kqpa8CZcEA4ap1D3KoQZmEzKw8qwkPEpX9sSy/NRpT7vdiAnuYsyPJblqs2qlR/P5uQtqVLPc
JuGg98lDdo5lkf5E2oUp0PdNonj2Jt+XMfpr3f9OVo9AK0uyiie9NuTk88uSqPXul9nHf+GfUmLF
5rsnHlF259x8KqTkBUu+viCWlNRq6URd13FIVpbqaD6h6JX//dSes7Vc9obN3TaFhpg14loltSm1
5gPV8FgjazSs0JDgoWlSOWg9b1E5QlZ8wyD6rlWUYbVsbZ9by6PTg3BBR3GEILg+6XZ3xGdU3ecs
XZUmi16CN4CwjV888dg3rqZ4uoHamS9YNCWLYq/RSfWkNcepQ4OoRSTNY7lq7bj3eK10jiWkgFfz
p7J2nf37fuQjr1YrCWDneQAB6VKDLs7K9dqB8XMXeGS/S+dtQNIEfdT0c8A2HUqozpiBICWqiPBS
J1Ifi7CauqJic70ICZCNb7hCtYvlslWr4hz0rnNuNV+MD8/EV8c21J88y/niTku4b1sM4kJt87TX
CDiUxKGA9mO1lBTlji5iNekMMXfIC8jhfb/NGde362mJaKp/RplR40+yji0nKlKo9JaHtdr7I3us
UFWUzI3JH9j9sRTaQNLIJC7Mc2YLWKIfOhfrhy4ZuV405lTmNn0Eh3rAsPaWuKKhA4dAbgRweIOq
DH73quKQfu21WsC4GxTh2ibwJTYIx6rQA4CHZMplQBpmS2bAPfReKToItKyAsJHkfIzECAANS2xa
LaG89MtnfGdMwPFKKCdp5v9k9I9th+DGGxCVwIF7kS6nK9GqD5jMz/gXWPV/92zpd1IOuaXmttw5
58d1BQgtdkMcmBAkOzrV5zlBvw6TjkL+JnFz/rQyX6sh5t91oOp4AUl5x396pVlHtwqWm7bm7BVs
reG/ete2XD/prCEQJU9PP38B54UZdFh87Gc2TGNXLkp9wkr2wiOFQGxWYD2sf5r5t8pHT3a9xE2y
jerX/9z2TBgHgB7pZKxhXocgHLKVPpw1h9ILv3M1CyaJmslBw0r4U4aAZqM42rRlGQFKswmUl1uj
0P5/XcMRdyxPn8TUrS75+SJgbO5tv7sFT78X/iQrpVnJYYzvpEQ+WAC8QSJpUYc+F1WTEYeS3tof
NLsk144wTFO1A5n78v/MaXJHSnprNn86IKlMtdkf0DcD148WjrSZ0W3UEZb+DuUTyG0FWIWHYnFQ
is8R1rmosWGyuXBQ7RaYfwXfG1PhgqHO4c1+GsYLYXsvsVtGwjLfKEFbugQZKLyCR6nbEVTojk60
h7Z1aPO5KwUeRFadDC/4CeVyFYjll8icXxqLa5r7VqTIbtR4btgWZ0wo+GBLOrvpZQzpR4eDOeJq
vHLSjGUBqE5UvncftoGDjW1Xq9CZA73Iz+4oL1WHFx2giVIBC5/ScVHAexBxOJoKhbH2REj+QLl/
zL+/OQB47AEM6H2xo8FxfZE1n3EBStPVzpIzoidW1sryuzSyDhdzTeAona0UDf5lQCQwt6KDbQph
2EZG1QHuOwwF3oIWApAntuNFHBcDcqmfUg+IgSpI3l17uWDCSH6jpTlx4YYUZ5gWYIfD02eujNRv
pnsveFHP/czBKSRZ8RuyeBGbi4fMTj0ExM6wtCwkbLhVhFUlBMsjpkMOqL/QYjkRg/zb8Ks/Fh3O
Hab2AC1i9zxmcK2VtP/GfskaruKD9p6rmCrZf4FypS9zEbFC8pOTbbVIkXSe8sYSB40niVndLNqk
4LbvxmKA/yIiw1bz059+HqxRbvF38KQF2tw9SLIjhxbAxeppi4+gwt64nve8KKua96P7fQhf/WPu
4B+ZPBXP6wUH5H4jf6Oti/jVEhHq0p0hsgJqZ38VoffuVh1H3tfINzXYl5r1GAiSLzmzmXjet3qF
PMeaokWmQfNLEhu0my806rPQNZVKJynxPis8X3TB1wlQaK9fDk1XK1+Ys/aozPA2avAA0vPD9XHd
OuuPRP6IsIddGiTWhL4CqhtqqZuDm6mofk/wLRa9z5X0EMNUbNBBbygQZMxFcBt1YyFGa9foAb26
kVM9q9Mk7EVjgrUkF6gn6Q+6BFAjmk9C3m28calCg4eo8M6ajHMlMeT7JwH7i3UCU0VgsIruBrSt
S54LIewYi57YwG1RXE1olFYj0TScgpYJ52ZKo91+TEiko0v13C/hfmuwTe7k4rPaXpkkt8NzXI6s
/t8SBVXyJDG+saAdQwyC9LcM1xnplT9K8qAChEgVD6wSeVwk06SGY+/oQkEbLjQGpLWuHkfQkzZc
1Z3yHZRwOrthF8jya8pYg8tjdPMS733UlWZf1KHnZNxPYu9kHDN23NK6J2ELsmiSlFSRdJE4QkOH
7OK1NMHU3fXXZJYPJh4FLXbWBUthdJjevyFODykxBSbiAYP8kUmiiBqqqVk69gVS2S3hgoYloOSb
iDMRYYix4FJSPIzru1KrgGDdlJGHKKy/rjdpJ3e5uuM3IW5AV7Txf8YqlmKS6S8QNVU88hqvF8we
55sdGhyK5b6s/A581taB4+ajeu5FsSVgqftMARkK6uAk+KKs+7N/AK3XM3twbN+BSWF6ANmREch5
bMNH19z6jJy0zfkCsdA4vf8T3zfckDe1Cq3Vyww8eoUtAzu8UEBLZcofW2hDHzmfmFfB1S1NZQTg
KBv71cpOVqCWOD+A0b5haZ9NE4aJiAnHzkcuPB0wbEOrujr726isyclqb1QyhkNPamQvKrbCF7A6
z+0xC4eX4QI2m9TGyq6Ce7oalOVFcEQ/U0BCYiTQixgTXOVbJJNj87CpXxIraQrdRk1tuNnPIHp5
wDO+i/NoJrwZQff0JxF/W0aL+mycmtdjLkL8ZAbEHCl8gxgTicmT8Jhw5HQt8nUYkimsxWG6FEeG
ciVhnOHnV1O6lFlFZjf/KYVU7dJ/piOq7OF100mo3c7s4vPpkryNYhHTUJCHX4Xbxd9BqNU4aH4N
JdwtT56gpBGzZ7TN5vDGE13GA/993tzqxxGcJCRlqTSy3mqzKa33+MTo+N4NVaE9bvQnffIfhZmo
1GXRJbgdmChVaThhMfU4NAPbrDW+9iGZ+GhGzNEZD87qoG+48/0KrSmnj7ta9rQSy3cOnJxi8QVk
cdHpyNh3HUoZseq8NcGD57byjVkiLO3vNdwxU9QeL2OwLQ7dvKilYL0/R/K5/BojmqK3f0d11tWp
ZNPT6curwj5PYo1yPlnPss5hqGhWFfVNN8mh2Va9PqMOz9Kz1SFdrkHC9VLBaanVZNO5XAAiSpLI
OiWaxtryhAEG8VVx0kdSpdq8RCBu5VmMVypcN8N0tYCkm/snixFTHsES9FtfI+3PSZHkNGMRMW/U
lKmYSpVVTfts/kaEMMGwRHQbhZq+vUqwjgLjLmZJXrEHmrrKwuExweYF+MO2mLYOl4NGJ16vJdMU
x4mPpKa0j6RnhWdSQxF8xph9S2KGxLF35g0YItTeRp4vCm9esWs85zgGGalXy5b1KOzKP/xbC1UA
caQKw6eeLg9BSEgoXR7Ak52xth3U+8gQ7Z0bb9MY/FVMbVAnPsOmvOe7amhLIfYgdjTQofywBz9h
CWHf1Um/p4XbPeE1Gbvhckx8zmeMEMuHOlMLymZugX5DvV5nLTTy81gg5ghnIO2/wnuHgu4ZnFcQ
6kTFh0jsV1ExT2KfQ4lrU9koSRHfgYO882vf0Gvx6pfv6xaVu7QKAb8IizDZFA02tD9A4WqkywEe
j0UhoBn3vNGLI8Mff+4BonNJnAqcdLaK8liYPFhdmZi8owjOftfQgsQO11zSMnVTyHqBA7o4bZZM
enRG6wJ7FCdcxxPVu/bTJBTTuBvnBs5hOwD2vHJAkZ8L3jO3qGpLJLNOfAJVeV5R5P+FXiaosqk9
dQ5e0PRsU6lKLbVigdg/37J1ExmZRxosIzzSXVUXB8BscFdYbAohohpHmTBBKwOEsduOy9J+iQYY
A6yT7bB2pFbPlAJhykXy6dOHkpU2hvwpXVfWsG2s9uJUyP6duqfmm3K+Dn9Q1NcFSfNq60WcuMcn
Fa22RF5FQSYwIEo1LHXGOLzmn0fm2tAONZkZHhmNZv+MfJsNHWHNDbhlKQg9+WwGENAKfzmevaMq
sgtbnbfhBTP2iqiY6hC/Gq3YyUARXMq5VhuQLpcgqXSWD6t/7ocYDV59HHn/rp6rq1MDcIKY7mb9
qZAPaoh5u28yva/G3h5yI8MPm5oWpxkPH/95G2nWoSkDBoPURvOjCjt4rSR5b7QKvVnFiO9H3kpc
ZE2J6dVPyBF1f1+eiHkpGTHsl3m4Tow6x9s/p37glxGtsFLXrCwxh9lSnP2DeRcg84iIBTqm+07Z
Bf3uhAs+m2sHmswCNLFPp8xOADN295t8Q1uw+MZ6safIZfCYjM2MKrnuApeNlqPdAhDn9f39rpVE
EBsK8swvJaFgrESRJEeplnD9ogIK00UW9YtMapnN/jqlAKJTIU0SbZ92zC1vlz9P/vHWJXxYf9+Z
N17UqGeDx0F9n55cGELM4um5xf7jYvn9hHZvFzTlUoxfjxSuhan0lPlZ4GnaLvNELTr/WrjhsUBc
FWzO3NR8HzMHFiPbtyWw48+49YdT/OGv41wpdQ00mmC9Ba18vGBWpXF6X7zLClyUpR/Dpxk/zYfP
/AmxyekvtBrPSPwdn4bvQgrlRVfpa9aKC/gupS9aM7fnKKVxdZj2J1FYwy2s8xmjm8c6/8wuFjWM
o0+F3Jplg9zUPOFgiDlCNgCODIoMrhw8hW18gifgHycPStamPnrmHw8/uU7jGMiVtfW4si3y4SLZ
xxA949C9WFMIS0wTHOpM4DAY2g5ZDs599ilSMbzjzV0APD6UReYtGqDOrqdVWIY4P0teIDBQ+/ND
EmYbuyW5oqAm6SYx15wQZEq8Y+frBo0tCQome2LN9swtAVQFrVOka42KTFMqRmLleHccqE/pwcnw
/iX9GQK12OHibnfwB7djMwr4KxFvAe2LuBPRZK0+97oWtKTcyvlLV2p70AiJE3OQ17nmbC9LvqOO
k9ngf0/HDqcae267ft5L3RhKrft2jdb2h8DWaJNbDZUcnwB7Eth8fU1SjeStXNW/V4/ZAJG1qLSF
/rDBy9OiAr3C16fymUf0wIaYx7rBhaSPonUCf6JShTzQGNRNgm6ARrXi7aPAtbRKXJKUvssFs8sg
vSC/1oTqbfNYVqtHcR9UXBcb5eLbM06y+8IehyJTOj+behPzsDL653l106JAhwGh5aEKPTi9oFQN
gJLoeohasFWLJAEzcJRjw4fgLGjF2VC46sdZHW0waQnIp1IgYpToeFkz0nVyez7QCv5aoN5y0mjb
/ZN9UmT5e0QLpPRnQkqOtoRFfNurt3LVbMQCX3LaB5EtTcvFOLAMnlTFc5iTu2CGI4dZnfyJ4RWf
gWpQ33o1iJsM6r/8ubDU46Tn7AIt6qGevBVW5O3gPAnAEciVxwLmmqycpLI2vJWx9p6Ysd/BZiad
k4yN4/i+qyDVubui9Dz0lzG9Jlm1U8MllnRnCp+aE8LRuaGQhO2zLF2WtSlIBf7v0dsIA/5sySVq
9gGuL2rDqnNmQpzljAJQy56JIxkO3ImnaCvfkCSnmbKKRgLyxLwFDvpG2mkgya/XoTo11TCoFHSL
34UWIaw+3F5RkkalT1R6S73Boi5sGPSx9EZ9IaYUXj8FAu6GtlZQnOquvfJHoZkCGZE7P0Xs/Myh
Hh2L0OKycApN9e1KPPdTVa55TCrWm0Ys83ZuJQxeuAXcoQlXbf3ZDNX2RHA02sfmEvSoaIDwpASJ
6NwC/mYWNCJ7X+tgOpmxfJoEPW91Db60jiUYLvhspv/V0fFRxWd80jN7zTT/po4T7OG1Di5Z0Ce9
+VeBzfIPhO3kX/ABYGxJLOPyRnRdXBFoRFBqNulZ6hJBXI6mfZ9LSgEKNnnzaVvA5dCpHO4sF84Z
UgJYmGNKEHaooOXbxgLYTxl0joHVmppTRxkM9FuQpJuR/eA1048qfRCF28r7ADrDSRClyeYm6PlH
ziZhSydNE6M885tgg/aBRay+UguStweg7JNAJtUUxGAFGIbf8AP0QAEFCuCfUB7egbXT6K8jhQHg
duStRPd+V9R8ZYo+OT3dfqF6IckQfK5EBZQ+dsOsoFe8TiYYnZSl7IP9MsnuP1UUzgO9DxwpeRtN
TFaT9RXK406kuvYyXOtu6UWucfNWY3Mv+7sdndzqA7O3MamWwr5S8qsaALhZmHAXTMEBVs7Bm5xP
BxLgzOl4fGfsnwGz8kpL6LXYqt/T19kEAdxJuewjUt6HyRZzSYugjDmIlaVuXJLFR65TJW9wC54r
9MSjLuo2NOE5MdUs7YPTBTbEVZ93vYqDYILZxEBCBXxi+XFM45N2rIxMyCWJ3hM8nKEATswAZCUJ
EbgRpve69DekrqUbAU18PJ6tFQx/JremEZLDhXF8K1dXPFz02ey+4metDTpOR58qbvLGUUI5QNrT
vmgxMDMkB5mCvQLTDwJxbBhcLYZJXFRFLUl4ZLPq24ZVAlLjpEItHWMb7ZNhr6dRLCPxkyTun8jc
TnvinDUSlVsBTsyTY7m4SxuPEh1H8QkQGZG/3yAFapKcr1FewBgjQurF2vxNPGRuEMDXrvmGwxX8
VTyz+PulpjYCxkxHIyjNcOBKkDWaKELparvQ7RlO02m/BIzon+1YBhDLRGwRJ7t1WAkdkdnMYpth
0oQGqZY81w3V4YeVK89XI+dK5ZOu+DWKRGBYH9+M8i28GJ2UY2gonRuFIu2/iRj+wj5VarjsN86z
Jg5IlIksAE2t16vZkhl1HbMYhYUZUNwl8rgWnptyYRjNimn55UUJTSg1tmW4vGBpMcCpGAA3z3CI
Kyh6IcVn4lilX4QQ3a3CHR4m9WKttVTcGO4lsYIw4eWp2v8HJ0FFWFvIR5PZ7OwCkzTrSufokM1g
lBf85lO58mgWJh3GnL2YUNjFMqLirf6UxtUDBbIT6HEB/t5xzdbgtmUZAhYkMqkWx1pKYFU7HMW6
l7E2s3fVPNwdNVXmg4LKJblGhTCvFs7K8UTx6OHUcdxUo11ZeE/7zYU8BLDMSUndvhxho1TrVMh+
WhLZSGKP7TvL9wZpiBW8ChZlYl3RSpoxJTGv0z1eXchT8kEmt39G+zL13OCj0IsKTwNkozEZ8Kgs
S8nou3R5Aw1zs6Gxc+O0L/80zJAnHwCsR0Xft8dp5bpERGdDu1S+UAA4MQY4mN58aRJm9Kvw1gFa
0epgkR9pAMintZserdh1Vq5rVyO3a7BDozxYAQWGID7Ba+q3Yo/CxLBR/J53Udp7m46dIdYb/U5P
VMxfUgwMmQahXa5ZBhopOcLYc0Jw4NbYdbbI7hZ1bHBwqmEuzWWgWbMomxhzo3QwqdhnyxkcqVPX
Kbj4PvJVoC1nJGbfs3QrMa/vVOgFazUe+Ep6ugTHSjFU7BgkwaVO1ltTeSjcwBLdtASVHYN17nKE
Ra5j79lfuE6vNX4tIEvPJKe8w6IbvzKc1yxkDNR+V5PqvGHfRnHGfKM40zTA6s04Md88CvmzSRZS
Q4oJ3znH3dzqym8eC3vn4ubWuRszBaZFrKqYA/hk1rZizlHsOhiNVIsLkSJ3XXMvmGPmrshouuKe
kBMwHx46wRxUmY0VepMCIAkP5OSPSmov6ksmowtMBaf/zxpqoszweDjw17w5i2obe+ytICUF/43M
Bnr9TLqt7wcsPhy9QUcWaFwMxTziA7eJig9HcIVE1og26L+0Bu1mCSaNLhefDZbM350QdyveTHSG
GM8XgmlB39P0UFP/epJFT86stORmB/slaEEp/mk5Dxw/ExcVprjAktVVzlU2Ha5F3cf6hXmm03QY
Kp2DnbPUCvdMwFYz0kasYMB0sDxhRciB/uJZ7Y+KWiRE/049TAM0hP8Z5BJ7tlfk4sWDE+37wROG
9nuRE8FizTKEb5fzxjo8gsD9Phn+nUKumuS3Xor00VJrpYlT+508nQii9950qZoFL/Sq8aCJkD1G
AKsTunVLdbfab6pB8CSz9XVedjsdoS1Gn6Jd6BB4M9PdA2vXG7oZq422QgadsvFtKK3uc+qXWZg4
T4xPes9z45PGC0bcc943QCjK8iDL4nHEtcVBa7/WBLFnFhtxzk97j3dfVKJcY/E3dbhOZJrd/uHL
BW2Nx9SGFZCG7GT2aQOle4T/S2r++YXPkRrhKgwaqwLH+sjm1t1lskqyF7tsUvSKVD1twLOOZE+8
MCNvacZK/ySUFOsOir5GUrOc5Pe9ZGyPGrbZRnBvLxWW382HSBM7SBsCYQ4ndOtWp13RQdIrWIbm
nkNTY5TrXTVsWfPHdvQ2aPnO4YLItnlwsFP4bc3PDe8PP6dyd9IhOIFXktmUf3ahv8730mJo3pHp
vh4WiHeIsvTO9JdDLarZtftUv0nJtQJsKx6aPoStN64FyUBVl29Qbxw46gx2w+DmjCsykqm94cvX
65GxttnDFHYY955aPZa/iDXFdjrJzAwZ6NuVrcmaQ4xVR2nbzPFRD2LYZz27WVXZ2JrBAFMbwIV0
b2+P2n6ugQBBi2XhmGJH7dnK//o99QdsUjSrfVpt5YAZ4/7R/QWf3C9tUwuJpgSJ/0Rl2sQxo2n3
hX5qgmc/xOUo86W9g4VLLGlqpjvv8ofi1xB8jBAJYsNjQQep7fR8MJgSVCK8ujvKLEvz3PFURJ82
q0t1PrKMIjbFZSyTAHSVOoYvvS9uJO3PTNwYUDW7n6MBuhPndZrwgUbDMw2prOCrpWK5wYB5mqbZ
14SbA9hRsts+L99XHJ778y8oTIWgsMtt4r/OlrzJJkp4ll7hOesjAE6+HsNq8Zac9qLgd1XTbZpP
ma6N10TXlCToYZvdnRKcSa/dvQbpddQ0/j8tDLM/tWafd1m8jReO4IPlkzM0yXOZZWpIqY6MbE2e
Atymd1/7v732TyV3wLY5sbIH3smEyralZjSsstmSHqZb/UYcJ5GK06wo5SUaGSMzr2plfnw/mhII
JLkkKKswFRtzadhPZFhLGZswp74KOkRH3MevyVV0r8EFnOD2OdiwnxZKR1+ryxCBUXVZCVRVlK3Q
4ny83HlQh906IFb+NVK2rAthnvHW03DFPUjDYHRVroR04OrY/JUzRP9YwVZs66aFDi89Dri8l7k9
FgtFqhSxa791W8ITQoXAHWC/tPSUO+sTwPkTdbPhFZiNrUiUeyv8WX9cBhIzY3YQngPLWr3sXdN+
uY+xWXds95G5ZeXWBG2YzFqyGuZe0IxvPOFN2NF3MiHCUfYZjdtlb0RFuLAoGnQ1DJpNP5uMZBnv
zv+75xyhKMx4XLweMyDzWL4fJBqey/1rGzuNdPfbxZOkxH1p8gstlzAdnDflCT/rqurzEN/Ia6fK
mIe8VHNNywReFLmW7Pr0lEhWanSH9iENFgpH+eH7WxQjGMgy5y3HXJDXIeDMt36/HQFawX175/75
DXO18XWzfuBUY6RizeWcun++W4toHIuMRKHUjNrNr2YhtBQ5VN693w47iv4tcN1vZQz47oZzLWqi
GXoxmAqfr43IL1BUuLdMHZy2xB3G1BjbYJSA/xQV71qkM83Zmo8+xWs/gmIvLhKmqNKO0/D+Cmyk
60Duy96cWla7C5i09IT48gdS7jNq4OuvwpzVfbWJbJlPn7IcDLncCNIVow3F5L+QMlXGuFP6wF4I
nkDfT4Bu0HbTpzSxyVNTyp+ms555dzyCvz7rhYznz11XK790feZdm5Ut/gcr8+1LUFJn8olPT2Bo
uPEOEeyW/4cui14/vSpsWrazGjVExOcGGTfkJSbU9IdrWn9HFLvdxPTRIDpidY9t6E9u7h6y0wSw
UHMkHkOo6S1usEvLGPJS5SYe20RkUEdC3GDpExL0xs7GT7zuScs2kQJfn2Vq5fjb3Oujis7FhvbO
b+Dg7mo21r5VEF+UdCqatYvZLprs5onJv/5WMBza3622IOILrULO2PvZFMnlfxwlZqOxhKc2Nos7
OL6XYNNIqcZb3uVw7otd13VAtMneS8thYkEOO5aOU4o4AUFdIwn/Qdjsse+lo9X2BmQ1lOCPPM9k
rWqCLoQ97mMW4bVZ8Di1oqfAOFqJVeAH0y/PuCIHftl140hU3SMubuUxFiaVCz3Uier0OR27/sSE
YIYcDfC7DGDB6ZVuZSmbEEG3f3YzxHfdKU1teykhtFnG2afiunNwy382hILCgcAihv1dKUdVkkkW
kmjdHCzo5mE2wFDy7XVmRaGpfKrHCIuzkj1WvhcROWz7GUSGTCYR7d1W4s+W84H5MPWMr3eWfl0p
yaLJdaGaY3eSthzFFTaMqekta26RNuwHWF/aHOwXgD8yguWjXuG0QAgiq6ArgmVnW8FxGbO3DCmw
ejEhyaH2MvrvwFR3uG7+8sno/STbYdMk5P+4BzOQZHoPv6xTloBM88u/n3f7SDOXS1/a+LNdLQar
Qy33gz/c+S559hAz54HrSN0c0HAxZSTixB9gRUM4hXbWIwURNBoqvbpZrQGRFW+2x+zZxxDJPgKA
TG0uyjgmpMZhE/E4fpHa11ZJ/k5EUn5rH//cLlKqHPMg9oLXubs0VBXEzja62ubbJy0rbwsEemBK
Tbj4FKifXZg7epDZMA4uqv0Rn58pav6hnaFB8U26Au5OfCubZHujhUgYed5o6jvP5WAhka/m43cR
BbVytEl2X7SWOKW7FudIp+IhV7icM8bjpcDfWq1tQlgjaKiEW5aM6nssHR04Mri/ktWSS6soUzdC
W6GoVEVKw3goTuARjFtjfEFMICPulsyS49bDK5DvZBDuVDlT8B8UYgW6tVzrZdhR6n4Trvq+tjfN
KDyhhAOdAqD0RegobhJ6gfXYGsIk6qnRe9CQCMFBJyN55Dc7BJWiiZR/1v7FyqsIZYZiyaQ0CMXp
RUFstkkYpnWx/M2/QwE+EZmcQl1dAwm2m59tvDPtvcKcipQOeSn0HU7eGRlajhJvX7kd/tJuJQ2Z
pgnbQPuqapqxrHsnvZSz+D6PgdiDwmF7PlrNx/ypeWQovcgzburbavNf1kczz5LE+JjFhdJHUfcR
8w2bxoNPveroq/Qz2vTtwHPy8KZkPjyLFlfk7L8tsWvcUbyYlp4j93HTPIrdmdWbxip51ur8HX+K
MHp3JHOpoIxSA6QMQsUPDd71dydO995Ltc/QGB8eGHogykPX2ixhkKgyzRrE0hqllgMea12yeWCM
EAd5jy5TnwAo0PfzBMXqUqUORcdtdKVWjNUSnibtPzfRuAsSHGDS+w3/p1skawxKEZZID6yl7bqn
KESp1vQDASrLqRU3BcAmUvyCGpiHHShhLcW0Fyh1oK9qtfUzdlUBMjL5pmKZFTA6re70I8SK3Dyc
8GM9l1KNEzpEwbyvodOmIE/dvEvEGmD8AdJ1hmkgX1SXrmrYehMfFW+Xrcy8C6730mDxD46o4dCw
QDxyA7IKrnGy4/nmExoJIZnXGAqioU//m9hv9PfKRS0UdnKM4WfqkeHdqq4kUJwcP9ArymK7RDSx
LnGrQsVrdOppMO8cUiibl2zFtarcENU8FGwu/qSKXYUBA52kve3A+tSNdEagyJbEa/scZmkb0oj6
ZKAUra3ZHes/jhQQjb6MugitaIVJzXx4cT9bRLNN6kR9oIomN8fWSYPn/jENGriHbbT8uAJCD/zZ
O8RGUGo0PQLlzB4OoSxUKahaxXRTWpPzLysxlAR/vbjNfOaBr6mLksQb+5zZnR82KXbI7Gb9X7J+
JpBU3qooPXpSYBw7h0CKloN6zXqVY9j/PIV0knjJ0yXrWd5JzZo4Bn1SVjGmXjz0OZwaanQ7HC50
0xpTYKknCVfdxaeD+6EDE6wUapInDon+vxHJm8oYxlTNIoL7f1841/9n2dvwVPDwlsQK+ZXEvz6Z
lFzkpPxC4S4mm2PaEssn9Fc8H2S2fu4pU4C6spUNmsx8Gm4iFrS4QRFCGidmKkP0jTLVKgCHFxud
+6BeQ+QZnd8iXlfp2mUWcGPYnxroA2I1mAgT/p8XShFCiSMnw60Kyb3/lVgtjN2Zh1pLsfpP0+rn
Ua7SmUCHEhjpfyftz45gF6M/qJok4EWhVc06iG5ihYdG+tKNydzq7ueiqusMtkYg03qIHQATdmDR
x6xMudgcmEK7/M7AjXRbR5LsMiS+bIA5qmUHH2VFdTYqSjhOFxATYHrgupNwn9L8O2rQW2+f+NQw
V7Pom+KjdYnWY6UmZ4+wPAA3a1W5vHSXsigdOiENRtaYXb+Kkt8q1Vf56Z74FyqtjNwtBh3rFzfe
NhysRHxWoGMCq4h1iMopd4bXZcWEZawJugjdL+hsXM6uz/QkrwK9cBniOZ0G0I79+9CwuOEEG9fF
EdVDVFXDoP/ajvVd7Gtw3gm2hHg2HGAIDzvheMxu8z5of13+g0GbXmotW741mQ+ks3CWsl3PvWE9
tM0mj2yS9Yy/A9kaK7TcTL5RCCy8cfC13tGp49uxjC+ygDcERR8SIzpfBXBwJ4VfFMmZE0FCU1JX
z8xqUSi9+uXPdwMGueLoEk1A7LZwGb1a5wgTyV/Dd504NZAQWKs0KH9YqXczRZemPOzoC0CTeH//
E5E5WdBff+FUDpm52tRnGI7ayBVoW6qeNR0zGzXhlK+VBHIwZ1CuY/VzWEpMkoF2fiFN9BYdCRBy
RUyXUKfo7PHNlg3CIxtYEN70QVilmtJ+Hy9/d4iRSGwJiMGc5CrMSruwoTFBoJYjcT9++sOerOn5
7qN5sljOeyxml2dqsAPd/S6VFV57t0BC4XHQsjnrQkSxvlz1MnVtAuwElO+AMayMmluw3pbWf6JW
yYuCKSz/0C09h35AGKCBH3cijyOJVdwqQnIogQg97n8uH96h8UsYHkhuDqwC+7u9SIs89PiEDMW2
ehDtU8Sre8kzCFuL4f6lyf0wOiv/VKzSrPwDswnN7Xq6v9IJ0XzXSuM2thncHoAwpIg8coIaFBiz
pScpT3Zco5hTgh4D11pBRLhrHgnyvHYRShsVaOBIGS/4BznrFfJNYOw6wOMj5yQVrFAorNzYcZhf
2kbk8sjxs2ymazFvIZlI35FMnFr7dM2tMBnMoxgW+0mX/mlo5WilEQZKE7Sb/TmkzIDjyShwcTLD
1fiKuizkrj5Ihg++DHyUf0ocjvI/nuupTaRyPT3KD0HyJz1hywBKoZBzrZuWbSV2jCHGC6CnoSPm
lWYcWPW4VNhYwyKiO0FBN0IQEfHgrGYoAHNjF+xo6O+GuVUwK8npqh23siviMZnMwpbiUq0l4UEy
Az+Rkaji/KzSi7n7xRj1XiX7GWapvJDE9if5zIjENLVUPPVe8CX51A0nPSpwNZQkN59d7tyfEDug
Kr9ckDcD+pTP3UwV2nSGWo69JzSSwvPLWQbwYJA9KF7swwVjXNWuM+rOmftRC6aO4IaP6CPC9tJT
KTkP3oSiLVRrEfDMLqLwqyd/8B+aCxc03iZnkOrMBIvBPFiDbHNig5RnZyurQphU/b7OCI/7oBjq
8LGtsYmJ/FCFZ+5y2zPAD/KjLHPKZZXKL5M58d+B6gBXiP3ui+KevtTc7N5Z0WbLA7+gc9EhwfGR
VQ5BHUIFockGTqPU0+Lw6zF+z55hnBExklQstz8fetFK6K35DXBq+187Ar/NeeZuyJtqJEqFDIXK
/aGHnNugUKICPy9eJRGSTwnQODpYhe9KB3ZJhQdKZ+Q4K8YT9PE1T34IJ8L+kNz4Lh3nA4WVgQug
1iQL/4FQ69/dT3EGESyulUMURiDARrO5mHVbKbPeogmF+DWN3pmRgL1FZJJo1IzMqSyMnKVHSGix
sGpovGMVvxevtfBHfxqTsrzRlbIZip2g0rrlWWS9hQRy1i9tAltSZ9rhrBrU92X3khDgTsmMtpWF
dDuCE6dvIxCStW6Z3oMkeATTVL2zhJ8yb0bfz1/NgX1sIKi0VjLLxSMTBQQkxfcWzq3hW+xFwKKe
Vi+HrElh8OgrxuD7XN7yLbV7EAi2zzzAH87pdND6EWTkUwyFHBIynpjXanT6PBtJF+CqB61KNv17
swXAu1Ez8e+ZHhnQIEBLzel3NNwlTWo4C4u7XyD5BsSZDW88OSj5gf0lnnOORYfWlE4TtP8DAtQc
TrHzL8nB1xyrvywFsw39Rxe+P/TTFgvA66cicj1KeH66l/KhWhxhW7QfORchEaq5WG4S0rcYWH04
xBpo9uXElJZQGKWV3+RKPgFC0PI/xSKRSkcMMwI/Ax5NYqtQ2AUaITkOAdorevXOl9dm/+GUEiY7
1xOuC4kZwJ4d1WMIEIHUmAbwuQlePXG9tY06Kg+/U59cU/ZtSV5g3MRLn7E2iLGUXH0TXtrUKnuP
Lq2BOvUmI5QrOGK+pnJ9ptbNZvVzwpc14qAX+Htz+8ntWCREgCs177Jx/BBA8muKJe6XfEPW/3kU
iaKsUBUBRbjrobSDl5TygcbhT++FULGBK22NYazNGvueFDE+hTjpGGfA3Hrnq49lxexz19x6W6/a
GQ+59FOLZR+LF7Q8BXmwqS7IICTHMTVsyQuWBGYbA8Fm09z7nvQXRRszrwYZcH+lEQeEYQkpI4Dh
7GIf3yYHuFg614zKPYgYV76K1Ve5Olz8hUiQ1+jPFs1siBKFjwDDdmPzO7QNRmqOqNPjOTpLxf5o
Wqs0dhUNBaip8qXtII1xa24MFgmhb84mFr8EV0hXAnPqc37q8DLnMFzMTNqwW8g/edEZDujGnIHU
gGDw/QX6SNWh3EWSoh8bha/qr7bryIzApm1irX5JKO3wC8UGd1BaTlc4NbqXpmAkI9/rVRg+WKbK
pMju3GkoPdWJWkVzTvsPw8GwKklmYhJ2RpJrXXTVBpd6n9y0ExfyS8xmxxAzpKwz03rd3h6aXnxA
3vZ/Qhe2SdoZp0xpJbMSJfXENop0e+9R8ras6R5Wvc0DjsA93OF2HBUgtwOFLsuO/8hp0lF+HvQY
ywO5FoMACuM+fm9o10TYVuB8sFz0dQJwKg+g/j/zatiASHqiaYpWG3BCBSrwXpp4evB4NA2M548H
G4ePrM2+xca3DyKEn2II3jICiZBRsYe/qlfG6yAsIJ3v9xIaAQ7uHvgLL6enYIh2yQCg3W8RLvVA
VJZTX29wbT8mu8JBdl4uZVnCb5CteopMKMwr3AxvpJ/GfbOEzElvULsM9rx3iKInqkX89uvhrAoz
XaPAv+QP8LEy0sEOCEVczAWHBTCeiWjH2PjxixXG6kJ+0+cGPOXRiHdHPBis5nQ7CjEodJiXdXbS
Uqp4dRUlT/JmIQ0AMb9fH5mAMmD0MKIcfeVShrkOAlARD5BoFOsq319enOOm/1/KHKsLoP08JcrW
Y1FvIEhRMc0MITYkTyKbiNRUVdWQL4e6R7MrXljFEyRYbs4+PruB4GG0tPPE/3OcAzdvV+aMZjYW
+wesK/Q+s3jdLEly/r76fs4DcHgkG4O9bdYIZlWO76MCPwaPZmONPvp1Vpw8TYNvR0NJdiCPZWZq
S11EfyWvoYh1C0/gid0OJdrJaDMLI5JwOl6i8e2AdjeXlpAsIADxnWoq/3XAoVCuP+kH8MyOZ6ho
SphUIfoPmuS2++I+YyjHTt9HyebxzdZRUP41to5Ss1XDNtd42i/I7gtxEQBx9bHxhJctdPWw3jat
95cO8HicqfYj8dX/1VFbX1mtFEJhu+Qpr/o9RLSa+pVTciNDdlLYzixttz2Z6WXJvviiVGFPCEFN
IZPkRi+GyNNIEkhrWjWUct+nmQ9JB4jVRr89ac3KvsVeuOYZAvAxSnP0jEHpOCrrNcNrkZ/qd8tm
xLJNrzwZV4RO1qnOpNa8ITbCDXLQQ82i71AZnTxMgyT7Xo+5xaaCFTRjvFkApfH46syRYJq57jL3
lLzGOsLGPze4JvikN5lh8hd9BVkWliGGhZ4bjZ6JRrnwPUOlhemzQOrvuVYPq5B9bxENGVQGScM1
g18b/5eCW+cTBZoxhlJ9pss8n9fTDl+YuzGle7NSOghZ5/sokQsvipdHi/bLCGGtVtfI93XFoXgX
BumQA6xjz+7nD/iXsLsVPoLh/MC5ZZN9HFiFGpAtexnxaJByUbFbyk2XDlpByjdqbUfKZBTod7UE
5/81mZCxSUbqRp2y/RGOylPt5ChrmagApzSvYa4RRbSQ++YoLcOcPaJXGZY4BSBedkSgf4j5SqJJ
hufJ3/2hf6fuPn8TrxY0XisRVjSsGwRulCVxL/8/jkgoUeiN7tQmUvVxQuT6+pa1t2/kFHcz1KTU
IQM/rzUS47HTVRE18Wct0iRy+rD2HOc5cg1BWk3VSEFD2fNqEb811RZLciqDRIBJRv7BM2DTdccd
crx7qAiLH7OGCTTIMFR7l3EzBnSpCj11BJEj5QiKI7SD/AKyIX+QWgDszlYYhVG/yjq/x0qtbHZU
QCveN70cR/uPwjlIJHhGsDqK4FJ+jgA0KbhVlOb1FLr4L5V4g0j2xTxzM4bG3ScLTi4GiIZdpel+
XqptAW+HXxTAZos2PZAbTRClF+xSt9rVG0TvxkxzV5Pmar/pljvEZsnE338ePCgOXnmGEkTrqkay
/BfDLlUl6wMAMCRVj44ZhPxyAR8pMS0wHIHZJne+XpltQvSEJOPHKSqgH3b5Bo0baMozdiJVeazH
b/T5TtEdTVvBu4YZMfvFEZzXdklJA3gJ1mlfSEzHOO533fmY+abcWzZiZ2V4Y3LYJS58ZRcMfnea
67FPWwD9HUSS47c+A8TGYJYbZgXm85WJOpTfi5APzMONX4d1p7t0OyVOimvqP03Zvxp9sdp6ZUWl
WhWMxlkmAAFRXNupMfUF6Sc+qgc3lPpYexiVv1Wzlhguxsw5z+zikbj/wZHtvfAs5EAFv/aRds/W
NtYrFOHEEeAl6sI6sOCm5WjtRRXpCrr5Kf9bnn35YtOAmJayrcp5H+nYR969vC9zdKq7Ob5a4HHC
lEcydWyFSUvtRV43pVN9E9alWWsmObcDmAjLIHesO2YAe8acB82eqmc3xd0i57CdMt1FLWFo3XXH
M0LnQGSxhSJonPD/XD258TnjmCnNU47m2ynMx+MgHChFjXXWzETsnCnfgGt/L9fyEylM/7Wl0ou4
ZyPyziniTHkDfXPwJCO70jOyVJr8RSrJszXotCy6SgdzZtDGeI+UrHrJAXfgvPL9oTGqMYtYZ4fE
ntU1/W3oApYPqsG/l3YwMhtkEsOEWzyKEPtdeBCg/B25qoZnA0LU88EG/hv1kthORqIEARfWoSZ2
supFG3ReSAA1QIV6CdzCjjjPvKNi7foou70DuBSzSrEUzhIBU6vX9gwqZkNlHF+AYkewjDWJ8BtA
IxVMNg1hM9wbRP7IWyvFLfQgwn3kQZlh5x9JfPLSgfM9zxYZL6BNcK3F3C7C2LUKxkM+tq24sMPv
1n20cSpUH0SElgEwF+UNXsYoSLlOzQxUvhE2PG/qGm+SYJFsSU1S0NBhiOcF8It6cSP9PuiaFMZa
rlzEooYATM+Ys+f2es1O9HTjiL8E9qICAxANQcqLv/kVpbWiDwUc5Lgsi/KqW/Dzglx2lbw57VCA
EkZvGZhKEwL6QbGJl8ZTE+yL1Y4nJTLJWnXOUDuiy8pO41wC71tsDibsBjskSvgqUp2b1XTJjK4y
w4zaa5E6MtXo07mPWWbcTiiNb1SMiTcNcm8sYuRPz7s24jzDJ6gVdzRWojIiw9okqKFN5UQcPVKi
Rh8+La1m/Rqv3DCef4xlZAxHyLEWeJWJCsyFqr1LDbSBzkbNRp5hNgUcLAZbsGgIxIb2d7XIwcbR
aKJ+262hSA1tXDipZokqMJc3n74cKAyTWlne8k7hFw6K622b2SH5SuAseuRXmYjCH0lGqA3MChvR
Eg8NzOrgtDXfyVhbXJuRCaT11bIYApOAfK/QOdWlakC4VFnNfMidcY/Gqugah/RlgW1mqW6WOjGD
eqX+TldYsuDtUgMEKX0xL69D9a2n9sSlgEbq/FtqjkZZDNgzhLOyuRgckOAcHtuKJLO7irHeVk++
kyZkL1a3yzAhC352uZnMrQfRXLxwAbDrkfuetDT8RjQ1BB+Qa9gCCGkzNZ02m0OGlYyXKeAUD4Lq
2BERybE0R8BGi6CLO2+50LbOtUrbe+i8Rc7ROXcQRYtEyLC1KAnVZRyzkYOrCgULJXAjyg2SZue2
rIqqAG0AjHFa2HeCxeFT+CllMOV3gQEI+v6wrjL4FADRjCIm13qsHiXdAwPbQoS30zH2hhRdJ6Mm
kQ6pK6Rmy4u4g/OWVn5T9UMsDgN+aOqTCbSDX5pHUan7aYDnbxGvxGccbxXTfiHvVWeck+93h1yI
yTvCfCbSjHHxsEdifkxz+VC0vjRKXCmY/kKcBuudejDJ5yLwtpY5BZE8YymBzr6GwWU/kal0nDP5
n271TStTcDUq4qDdtDPt+v/Nc5C8z9mks87zojpWgmpyUyZPVuZcKwyINbxMi0Cr7/45WHluo5F7
t2SaAocif+AaLmYv0sIum2gHOlo6FJWomkgSkOcpgw3xXa7Mlejpq7mIqQzwKOtsasPUWtL4W2UL
AtDi7uxbQ3fIv/5Q+pn3oz9Do+lCu56VVxEm1GmFT9Lt2P2dHPh94Kh/yXPJ9AVrPlsf8AByFiHi
Zd1zrQ2JEt45xj9KceGO6fkWzsbYPU3ctUxGjR8Lpyv8UJGxeB+rAkBi4cD8qaK+bnycGPMmVbn9
UXC4O1ZMHOpNgWe4Kr8dbQSDrydK1ZnZhoCop+b5cKHu8jmZk2l+A+kr9dpEYT4OJlO1ATG7T+Io
ZftCgktMLgT/J+1QCJLXONPBMISM2M6cZjUkSXyPcB6tQnJUYnfJYFvXXpl2cZXk2eZGAxw4bhzq
xTuO2j/1laPt+0A6Xfi9SLXbvIOATyY7wMsaurkgG7Wj1k0J+n2j4HHOKh6FSaTgDMXqo7m6X+Qe
v4ln8M5em7zax8SwmmcTTnjIDLL39wk/aXnfFh0AO24J2bpI8K2tzEmsYSi15xdsAQTemyEgy3lk
zAuHEqlLbxRx6erYdDZpOq7+1TS/GhcNCTPcC3YeR1LLSDVLT1K9DMCpGV7D336ru70JRxdnR/Ua
OdOPvaTN5Fo1LFp0PzRu2rCKFGoLRrVHHgS50i5iJWoN/HxRI2p45WEaXh5V0Xz0EBOK9r6Y6AB2
QVRnvaFT/H2bpstFAv4g/r6mAbW9tL5+r3Za74gCnmdIRV7iUOdkvB5FT4zWxutc0tg3KAe1ewMa
utEMl7haGYswC089LbzyHcBPpJFfDO2bUJuyPavu1tzf6Tg4ifxmdlokPfZvSdjOMdy2y0fxj3hK
lTyLUYlvrj5NQXPdtrGcov/lFVCBKnWprkAWeq5qZcrfWYmZ3AEglBlDmLLLz+Fxk+8BzFXp2wTL
UzVVC02UuXI7p2tdjjgFGPIi8y5BWQWK3GDWrtGLUJDlmgJjTKssjos2Yq+9LT4AhHfhGC27+e4+
1Ixi+Kvjl71ULgdwCLkAxozhE1k9hNlR0WGI43K7134rrSMaKQiruh2KG7YFij7ZvqY/Ih/L3Mfk
D5MKvayf5BhQzBeai2pWqPjvehzOhDpzniLvk+ct7tCGCmfndFO0zU0vy55z3qfxBrtrSvPYoWHy
d5RNPkxibUGArhB1YlQkEGvBV54FVp2sg6gWXKIqodfpjpUxluRncsU7hRMq/sCE3yXmyUlZqJzV
UqXj4m0dkidiaqPUwtANiesuPc+8iwa367XzQKK0kcBWsHToVK2r2wJXmzimddApGFZum3mWMP6d
UezlECH2vPGZ5kErnbZZso47tOI1TpeSTIHrP+AmXP823odZ9hJGhyK1g9N9Igx7FlgjDl4EAwsl
MIWUW94VRJaYtUstvWDZzHZtwK9BKYctlDAGGWNg+1Dz4elx8BDWjOnuXGZiMV3ZksL+I213A/hZ
WSIznwJaqDMEX2Xlmj60S3KSudO824Gqq7gDOlQ8TmZR68ic62RUtNV6YHAi7p4IWvTb9HeZbDX+
OKqotWGV+iNrlK8OT65c2HG5uD9YIC/iqTSHemVdYqbHGoRsyTJFfvX9cTIbie1vSLQdR0nxif/R
5E0izkYTFuxyWKhrNzVbAZLVKzRfKxVquwkI0XmfKZaG4ok5H9JQpAhD2Rpj4slxSleyal/wQWa6
c54y9PYu01k1BaHXNIybkBnZlzV6PzI9PZAWHu57csQzKYwG0PLMYJUbUuxW3OAEHdosgBWnh7ZZ
x3E7j43B0hh1uA/zaSSxNw/Mnixj0EK4TA/5NFEMRdi4DQQypZLFbUnSvvrhJ+0lRe0ZoMmayFF0
dZJBGoR9NTpbg0emmcdzl+VavMNX3pcnA4OM8XctoNsDz3Dqm+x9fM1TiEL4DFFmfS7XILVjKHIS
4+YpNhda3CrgZCqwJW7sLYIkXxdGudJCC/b1SNTtGSMFbGNYj550lSxJAopLWULk6xR4grUjQWCK
6mgjCx90H5+lAcCGH9iY0RxtBueCD03PchcaRI87PyctcBo/Zye3djmWLDV1vKtnbxXZKcnCyUKL
2q74swJWbvlXuqV2DZ21mlAQboLyPbOk9nV2MeGFXMwxJaVIr/8WsqMC4cF/Kq/rUH/5eqVOD9gb
uu+Z5esILCb5cayatVB6bJQlH1KC5OwY6ztwh1dx2xgSGYstDSTpq/hsurFORyeBTaBF4u1E0/hY
VhKVsBkntP0pKQTEF0vlUr+8M1QZkudLOCqNG3iEzAMJREwIr2/HgMyn5SoqzNb9ob8WKcRUoPwM
ALZa8xSM4hkieh+lm4PozOmMTkiTGER2/qAkJQ8Lkhhb7FpZ5s+9OOQsKP8GBgEj2Vj73xSdH+jC
ZSfdZJQ+M+RXTtZB81bNYpn2J6dn5VWy28c0ahWl8qWiMpD5ItP9CaKd5wEnCpV4wgsT1+5GCgL3
4Srm63dScsUP83s3orNBxexRan0G0lNTckdqZY1SrdEND/BR/B7g6YuZ7q1X3ochx37gcTDl3OYR
R5AfFW8GPSYPRlRyAy56Z2Hu1G0+zNnBDwTSS6BIYVQstqKzVteaofOO1hMIl/oZlToM8noAiI/Z
yDgWeWEdt8Xe4KCEdBvVEHCHA6FMJxPt6mhIbbUFcq5WTpRpr8E4SKb/0YyblPwYXXUxOBBftYBt
rZAlLMuH/MYDC0nsljfeDf2FL8TpJPNgsXm3XcnOVhciEPhp+4enB5TEKnwa8LCyYMdD37PXF1Id
aZTXHegC1KtOFfWYY2MPq6tsQPiUyVP6rD0YHc9Yyv7eazraIMP9MCos2LJSl7SDLNA2LOpekPZl
r7u7bliA7BQpyPSRAYRDKHvMvaWxgW8OdtGvqZEH+HC07raK9m47t7qN4VKWAIZLBK31PCXBkqXI
oHuoCb7qFXtWTOtm7UfDM0/ScR/tXDYOKS3hBcEKGJWJLd1WX1T9V63VcvkZOZv2/Zoodwlt7me5
bl9kgMxbffyF8UblTc0IxKhyO+/ScGP9gNbIwPoRmPwzi/OKLBnW2Qj1+9HRf+0Rh5AhcEnxCKdl
09mOPxeRmaMRLAvGtNxZpLGfzs+k4x7nEejKdavoycgVxR0GEiqTs4qw6qlv7ho9LvFgBZnzkW9M
I24cnZbN7pKwEXzF01oGSBU98Qwg/FPe8MGqTl1DV4/z6ZObeRGHgGNQ+wQkfK78IivKMRMdItwV
RTjZSQLaNe8q0K+85Z1ga+unmdSfauJEC8DdfxtWnUJunywNmLjGesRFfkxaFWEHsnoZSjtXcM6d
MnvIkpgfFBPEMY2i+6U/gz+aTXJVLMcyP1OJ/8Quv05K66S6pZ2v45Qx9qC6VtQCLepOukT2FNi8
8X/oNvghWOqWP2CYQp5jcgPVhz3qZXwetAaTqdjRacFz6ErKqlwGVTZahrAT5J9UEymjV5YUxhrE
hPB56GNQIX9AiQsX454UX7nVVvceg0/Jv0EcxxUL0yzZ93rCr7HZvi88bQ46J+B5bUjTXGvlIBVk
WVmaGSH9rjzE3LxnORSaL00M/6l2xh4+l3tXPbFmeIN3D2vzIoJXrqgTv4HrxAC6JncGaSkRE2hh
ysnIkB3b2Px0F5ZHpE2fjs5caE0jc/61E8BEciUkiuC01ome2tUrLTG7QGp9OWX+KDWxxINZWkIo
80oebcPgiQz6Qj7MQO2xM5ca04k0yAmGFbHubGaEPHSHi+WS0+Gs6TeRCK7gpluPygvn+wn6VsWn
FWmE2/cxVkrHzC529SBuBWeWKyktOG07C+bqlGyBIwC3emUv0AZc0sdsxOxvHRtKkbVbMdfOB8Zf
xv1BERB1928kcKt7mAR7tCCu7FWQ65OE2Kp+Ud2NIt9PYQBY2x8/4r7oTKIsI3KcLK0A6TOPDLHm
hE8JaUr3IL4+tzwkCX4ITow4kWuPtc6dpx1d92N7VTz0oFQpgHn5IahN2iDc6ZUobzFB5wfCichi
56bqQLaKAt5rSBRZFf79ubU3pVp8MOKRum6eGONbdvPxR3fQ8FeG5lgwFXwmVNtW0BXVqgkF28v+
q1hFsMtCTn5GRLf9GJYzAT0sF/oIetg4q6ycMti6OS2Qq4GWSj1cNb6GIfmvguwvfLFvE0va7Dhh
fHFdt4oJycsrdpbdT/qGlCt3avcFHfqYH3ezLsFAIoHdjqPO/v9+wMPy1fkB7l8GsS+8GEBBd02A
sqAtwUbu594YmMw9A2WXOR+7WxnlLOsp2Kd2Kc4x5L6s4dvlfHRtxsYikh4T0Iz0ni0j1NjDNMyH
cdnnHEQyn/sva8pYmiCnCVLRhHmdYwj/7CU4dk8HfXC++y4kcH7t6t1iTlelE291WLyB7fUtmdVA
cYLH+gZLcA8+2ZBIjTTZMeRJRf/XAA1JfSVvbdHDikDvTkoul8JbewRV24AwWi8Io0sHcDllppa+
+eYU1OuVW38VfkdMidAV5+dIlOWppY3mVpbGcFKCbi+3PwDEZIObX/Sc5jwd0Y4Vd8KzBYjEKmBV
V92la7BOZdUm3r325XC0N3HbYG8cvNfuJrkx0TRo7aoec9ZtwRD44HHTSj2368OaFUpFF/Qv01Mz
AOx51SfBgHeyCKQ30Wrn6/GUWqr1tGTrvapxEUhJOFTP0oiga6xV13zIPX7Nx7JFIk2CkvtJpeVR
5tRh323+KY5ZpEaM0By+SzoOccezYoTVF+0snaYwv/Ppt1c62o9PWvkWlE0ZYvSaRDbFuG06IxfP
/OvrxUPo9s3GUJ3CyuKx1kHt6hsKI/z0LfDGUzVQuuhUKVqfPRdFgHbPPbPZv45XPHc4vH7tH010
oM7x+NwmEVX1QAE3leRQxGqH8719go2NELs1hpEGObLylyUukbW5HBg6pXXaSp2r4ezQ7YVemWZ4
55LrhwhinkqGQyaE9cBXZriK9GZw1h5/1F/F7u4IIITYIDfI2dX5UBfkIyyzziXNuYUvqJUh1wyb
uAQBGHxatOwDlzz+KOkr88RzKq3VLKHcmtiz6jpAmYepB+vp5+xVysrYKmVvLBtvVyCZZpnKta8h
solvioLu8oXix+APXIt/0lGJp2ZFZGK6tFcqzHlAKLA/zFQb0i7FluZpIgWq7EN+scykllGWU/gL
+xAaXvMq3EZqXpCrN5iR97xHaJvecwi1wq6k8TFHW+DudXjVCqO1ZJchLK7HiYl5sDsk7Pe1l2r+
XJsueb9ZUo6ECT5ISGOMuQDewa9LlFtmM9dZr2/2QiDl5+Z/1j/uUGaEv5dMgDioDoMzNAfqr3VA
4ZdTzHBZ8Pi+tKhP265uoUaqMzjXLaOlPVqTTOXknUnwLxhleOwHszK2dTJ2wLQjE8RaOq9MewlH
jdSZ6e8YOqCtBKZ6+JKkGtXZbGT3/hhZqO4/ZNuGP/cWIEGEZ6948h5d1b+WXNzRcvMeSLC2t7og
3K9VDZ3djNfxW41CY4Y6/KbfRh7HDcO2xg94X/vCEg/yXsMWrHi/Jc5Affn0eRhm7Svrd1NGuEai
17rWQHlSenlLsxdZxwEvXV7tWgFevduJCXNGkvDhlqBMM0UZof7QcLynqvkWAXH1+AgEhXBQMYDD
06fYCvouM0dBUxzP7/vJygRwtAxdjOUqdtktt72qHomIC3Jixlkaw69yUvGv6nCkcr6R2nQD/t7F
0yaDuZ+lJys9AIqK+cZjioSPOCJuHPPpu55pU4mllIFalWuDggJZhqV12WTfGZFhpAN2GPIL3M/K
Kv3yH1q68S9JJJxuMnrDhK2dPj9fG6YM7LYExuTMGm7xiIdOPRYb6XptBjZ+KMLCau+QWA5y8RUr
HpG4b1jVKnJJyyPDJOwwG1wQMNT5fAk2jD7m81pAA/u8hOPt+L5yft0I9rNQdA4JAxyVND4/fvji
cgm6wpn77iTXsQvqVftpnX4/Oj3UB2yHuzO4zPEv3EB8tfbySjV6nwy6gn9P/5a7KSGGxossiuIP
+B5rSCyIxrPx1D6FfML0Xd5s9Df7iBR93Nw7mAi1umIRNxEOmHCqZ6ATHS5kkfpXSAfHcufThCT6
KqCn3132h237t1/0kj4Yp1vi+BdEqCSYPkgi0icGKoe34VzI/LaUDBekd0ieGOhe2X6piAHd9kuu
tOWPzEUN24MM1MDS+jvlIhL+2ooPInBzoEGzXuW5bDuAFN923X6rAgMKQ0kbusJcXRN7ZWMA2XFx
8fxMv/YgvFZBabWMq5n+XijYRU7Cw+XOh39bv04nCmSipp7spe6ec6MObxTCqHxr6SCqW8ulFNMk
0niWfp++3goNPjzRQdOxCvDPb9aM3CiAA8+vK5vs6aLAQTXCFr1nQlPoXDQIR1oH+thTKinbJauX
Qj6mA4+iIFAqWCWjLV2qvLjmj2SwNewRejtI5aLa/PFpWuO4BxIKGNFWPNMXSPthz6K1dK0KOHST
143/nk6G4/b/MlutDmmezOmOByktJFm1/8Otlj39WUXvg3IvgYvECpNnvJJeMtpHIE5TLIYPuTb2
v/jyeOHO9KDks8/yg2fmtIP+aPTgl6Q56nVXZ9W8ST4ugDYfxDlecv560nS1BDo/xyPNiErZUDiO
cgx46Mcyb2FLAiqx3mU8zsZYFs1Z4kBPyrbr+w/sOoz3ycDfZxMQHjYYjZYf8v3mgOYURdJeZY0U
PuOUMexaNmQD93ptxHHqTLFQh7bFoLBxAOew7ILVZOdZfORGF2HfPT2YXoUaz3P5R+M4N09tNMnf
46tTa3RjPsG5VC51a+GSmJHLzLyehZqAB1TfTwy5Ua+HL/x1tp/n9vV2Qru4GD83aZQMLEUe6Scq
fT9x1KixyfRk7iFs6rOyVSkZ1mW/igBESM9d5+PfV8Ed+/WWmUVQXxCKzK58VYaVc5D4LJkfboU3
SbHP2ytifM8osq7LCXmOPr9Txt5zd5J2DnMw866+JWmEjvWCZsZNOOn4x4rCg+MyaLjDaapfaC2y
AqKkKlXlUCxIPUgEqqJEM7yVfxDOih62e5EDDI+bSBMGcOulO1sKBNoZvKmpe/XycV7XCCkyy2Xz
3HCseCqhLWqB/f2hSrbQqR9BWrkiEayvgbdiwEjFC4+LbViQyQyFUSFoUYiIdvE5xTXT1qvvIo3+
hkQag51WAf3ZEpbaI1hJeNllX7BYuVA8+m6NzCBb+ZruhloAIwFgW2nx53IiVwEpYeolI4S5mFsE
O9w72zyAlBWc2LwDjhGLVQAx/r7FgO9DFzw7QtgPw9T1vvSSvpXX9wEPvGZ5BuUHguFUnJtoDgdm
afS5qiY5DQxWbi4PK+hFIYU90TPaW5LOkzwTUEqVGsH21FnJRapVaZRZMLF3q/kFGk+1nN5YkZY7
vFL/x2eqH/n676y0CWRbmSqisbePTgsfVKkZh0JhWgeFFYZZkLaDn9//l14wX8GEoOxdqqcrD4Qi
0Ky1J/2Mcfozx1tDbmRd0xU5TBzKa5D1xSjKnhJgpgQ0bsI5UIThWhshJaZMpAP9RyFhlL/JstuN
ZM8Z1/afRAwIUhbYWE6n3spM7kba8OpaeMHQxvicfBRnfyr7fLPKXT3fJ4HgRDpRknjA/g3GRtip
qtGzAS4NNh1OicYm8f6CKclRkyJDebbqXjh2tcobQQdEwWG0vDcUHzglEfMw1Cdht3mEt8wVz+yB
9375iPmdLpacWBFj0IeFeKsCKUYQDb2P1MkPQCoDcLbeiD0OpmGRJgznurMiBvU8OL/ZUsYrEDoa
vJlXMIjWJ4/vyc89RXTz8/LvDr0fmttTlnVp9KDNb9TjC9301f+h7xlLdkSCajKd1cdQ5CWf8Vog
nBajqwJ2HauAsyMhacV/IjFNyyZlx15ynVZAoxr55XJVzQn+MhR4f32PEU9BXy3Aoqg/P4hRune8
cCnpdAX+Abwcy65bTLk8kCH/dPIlCqOW/eFa+x1R3HO6W5Ka+44u18b4Fxv4n7EFdSWav+yAP3b0
F9Vum9dBkpMU/GBofelxRkCInjyNwj9SqIqo1J/+WOGY+lElCmNpfcaBC/Tg4kRAlRzApSmChow6
2wZrl2tXzm+9Spih4M36hvSDAVDB1mQVIwT6BnwGiEThPMwq5UUuKnp9ICBp/Ty2nvN8JGj1dEg/
Np6OR3NTGEOBTuO2e59adRjFCQTBghTcbq6s3d/wecXloSv1TzV1NH18gE5TES6Z+M7s7l6VSzXM
CjdPUSwlrJWZzjZrE3Fq20ZxrTRjpGs+yWXSxqc5LyKJZ+NWBPAzrUKYtuEg98JXI8opCE5Deypn
r/op2PlwPJeJkxDvwMotmiSDCtF11NuEvGYoaXkA85WPstbAgp+0PEdc9h31hS7dBL/9+raL96m5
dye4EnQRhKR6lLghJ/EqLdRZjz2GkvJ51NdjPJjECkyj0xLdXCn4ff3Ebj1AaFvx5aJPwCaKN4v5
ym7s5qzJGvk1ayTx+8jftEVg6cw1FLCQv6KqMbAUAjaZ8JaZwCXS99LGBhJ1pwypGRtSAsFQ7vB2
FXW7v34cd+DJCDLIKvawfUlNEt1Zm4OFPTN2A9J1s/NiN50ZV7JiLe2e+hNHHmeTmwncbC+O7IRQ
GkcG4Fmq77Bk/agA7X/gMTfl5jFixQtP/o0UKT6F8bolpYqwuDyTZZstapnERkjrWv3RsmI7zPq8
1MTrgHELCwaaraU09MkiaBvrwKHYtYNgv2X7cI8h+dyKEtQppj1j8YBCfLWknmaaEXMkudBe7+Xj
u+CZMwq63fBnFA==
%%% protect end_protected
