%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
J6nPmi3a0wyuPUjS9soUEzo/IcT1O93gtaESL6B9QWvetkHHPV2R4+EumscU7SQ8MlBQ2lXjkpDQ
ZqwpD5ZldTlZN9CqxGFxq+yesx1lYWCalcr0Qe5oTPbZCSnsu/keGHkh18xzmIPhlWkX6SuzJo+r
MbKNy5D6L601z2TXWmeKlY2GsBSBCnaogPgqNlYINGA4q2UNPuR7uQZxMsowC9laCvK0KbhZiOD1
ywv3aEy2JWpvLnzmjiyMd5LSoJQJwE2qplq9bhqO2CNBChWJggjkVc6yCZO0IvVMciudDtCs0ErU
ju27A01miOhSHYAVTsGcuNWzpdAzv93pwl3Sgg==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
vB4EcpCBKoeCFYmiZ+oMuEj6dZmoGdnSB5hsJ1pi0Ob2zFx5sULPZJzV6ExQMhbBZano8JGnhD4j
3OafkXcmZITUe6+pOsW10GlyDSEC5Ag2SORk4mNEgnTsfDNrZTsuxO/YPmEMd1a8jyuJ4Kl9AzC9
n+OaXWWdPK1JAMJ2U6e8ZsHVVKjbv8RFl7WA7lctQ3XsWTsWNcIpI/Qt2dKO43aVesO4dzQ2BUdc
jwp+CqmOxJrklm0PBIUIMNNSEHmEgJTpJsMqlwjEsP7/KzGbOraQBzetXgG9cPi16+3dSepf1PW4
emgsKbRjUO666Qt2d7nuITasGeUZv6dYXqyRFhNZ+7K4HHfe+OPrcrTQs52hRJ64o2KQsk77hxpQ
BEOKIsg9m/InhRJ1viQZV9g32ihIIKEVg4+4syVu2KxuCbtS2XZLfdMBk31hv/VuSzoFqCFmEUQu
tf3Dq+ci92EhtUya8INOlBOCVWh+qkeOAE6SCJy7OM2hAKLjfD66IERCtxi9CfyC4qFircladBxO
5vi0W2AZ0/BPxFoHmL45H/27GT1ZYaJUK64P6hDrBF12URxDuipi8ARmcfbRBnqkEslUcrBqD++x
MAZlM/NSOL/PaX4XLnrm0KkQWmrpbA8XIsB6/onRE0fuJQTAlyGUGoWtWEgsT8/2Di2rbtcvtbMm
oT8C747nzkXZ5DGejeDo0W4z9XKw1M3OHSHZNFG5Qwg7rG8QIZGscHfgQ0aFNxiKdmsIj0jaHxlr
c7bR1ZCXeyO7wfSUUDQKSFP5zGkOBv7YhQsY+UOPd4+/79URPWTI8Du+UdUpo9uqC1uoVq1t5qRy
freZGGSJ4hQ4aPMVvr2YJX44Biur25gnhKe0JVxlC1ktS8wYu2RPf8cs5usYJaL2LXLzP+dKkEbC
Tw/qmFnF4TfIHjWl2KZ2TKcuhRWj25Q71wsuZjLLsUVDJJm8a8/DLpuU/78LBqutLuKHgcs9g4/u
Fiu1wYxNVWPUr5A18NIjlBi7zyLQKzfgKTX6tGmP9gij1RgGWIOnyNxeWf+QUvetFF3q2x6lp3Ig
XJZz3S4Dv3AKW9EMBSrT3Lpl6mrb9+C067zuLuybiOGvCGk2kU4tykghB7lvIbGr83U1ntKH2BUN
cI23y0CjGf6SY02DwhSFzDC/+/Ae5Z9jeF3HzSHV3zzyxJnQlk+nQrxQWDFUjEeND4udBheNR+qV
lOmLbmWIBIEGA7GFUJzSHOGO0gInkZocqMFNlgfqVgIT+b9CZqsoaEU7IzGBl2Cjw7n6ZSshdS2N
fWdMic4wHL14lZ5kWUh3eiT7w2VN+PTE6k6vKzZJWMoWTAsrB9TJwqGxMIVc9sMxY7nM/Xsj0QMw
iLQLiH4AzHwFFJcV/Z1SpHKBfGD/6uHNVv1ZJ4UIeL7UJa1XGjZIUFQ6bsL9nEqIgoAu9Tl4iVMz
3Zb3ct6nZtcaAh19RDjmxsWo0ssF9wRgSMJ0YiRRcyES/ERKQ1pdUs0DRZci1kENyfmeQyi28mAb
WFpRA61YOyvZHw/CUobT6c71vtP8B7/y0eI1Z3y2tQMYIF7hAaL8+VS/mAt4TNwOwXGS+2pMz+J7
NfW/UTquT4WDtsLl/jsYdtMcN6fB7yXSk98IRSfAmsolP6Sb9kQCC5u/BiN/JCezWP9niNApDg8a
M1fF5QOlkPwKqZR42zDFMQ6t4lZLMXP1JLBKAD23C64yjgbwwfvJk3/wk7cgvLWbjkEJXRslN/BQ
QKl9HFDFcE2EqBF8YZ0v/jheZMQrNDji+UxGRo6M0IuoXLcJBPHdI/e++YH/1drvWdlQrCciXeRm
u8xZqLhAjk9+MwUt3JkjMruubxFtPmOkije+ZNQu36fH3MYJ2w+dpymtIAq10rh2QqpAEJ6or4lR
IoSGeLeBfET8nVK4dZLtbQaUnrVahR8CWiFYBzytU+S6Zb21boa6jMrl2OVCCMVnJfwdZ80W2OWF
Si3q8fEh2e2p6WFJmVFTc/XhR0r1e2ezXzJ3CVlvroUbSJrc8l++vOIF5jrn/+PF7M9QEXS6zOv5
GxPcgZYZygPnpxUZBFG1gJpeiGAb6npAyyxM/p8VW+ItXaOlamXB7EH6+pexX05f1uev6FpOD5Fs
7kilAVL5iADlarZyaqswb28efSng+662IfRvpddnnm/hgVHp2zDPrX5tHNFlYGiS+OgDstQ7x54v
FRcynNiPsL4pBCkhyTBtyVUci1pfjAR0cLWAY4Tmq3QfFo5zYwlA61kMis3jQZu3X3yocb1xCJr6
eGlPR1JLSIuFcWHCFK8R6H7ML9qxXCXwrUF/8To79/FKzLnTcsIVqsssStrFpdawsp+9xNGRj3EW
iVDg8+pRKaNEQOrW6g0DFZXKvsv3qa+HPsidAqPT+p6o5QKKHIaseZKDQse2dBknyB2UNcwgWFKb
qKxhMr7/TVhD8gqs6yTP8dEWK3PPO/tnGPzoDFvZUSUCmH1Ozgvfazdl9jqwzA511zjiPyy2HdVG
7vtqIuihxw7WEijuk955mMqOKJ4KIg02TU27tLoAwfpSOAfaLS3a1xij7xbGS7eUz3l7Klpyj9Fj
o5Z2T8ElVHbstIYLbPnJEWEDHW+ZE7zoDEA7NEeuRz9cZAVxSynS+d+jqNwl8cTyPKNEZfyIgGlB
l2Rwlh4Lrk3G2OvV3wKR3DBMSbh+3LAXC9gly6o0mqiUidYAXKNGkOuBjTs2W8GMErQOp+HtYKrB
Q+1HeHnmpk/JSVyxHjjoIvva5Wo0BZcaQg5ZroWVtYnXwFRg+E0VU+fgUnQn5LsbwJZobgFpRrkM
Qqm296Vj4xUF9Ht3yYeb/JKQl4pt3JoBwQ/nhcFz+wYrFPC4YN66mC4fhjt+xIA036O2P1ziByn1
0rMOA0QS4HekbldbjZzmID7698aFjI8oCz+PnEU4C81HZWFyrgdYYhkNgNc4sytnL4yAgHy7V2AI
jY21+Fy99KIVxaLz8QfKed8RNO7dH+P3Il9WYvt3MbdB07ZrJ6S3y1iYo4Sr+KqsoegghhGXJk9e
Dx0SZFnJ5d8QGAS9MSchKe83GvxnqMZvBUJdxRIMgS31+W3mrF/sxMA9vL380E++GVjC4lYlS5DF
s5cWeUp6XdNU/5uYY6c4jKujqbEQPW+eFg5DCI3EtDB3xH7iI9k9lm49/Yyk3n8p5YnFMmO3wyLI
xFHjO66PgypL9nDkv/v4kreeP7Uk+aONQ0fihLGAseBa/PeYJVyt/2SR7z8zrZr12v+XM9TKh+mZ
84Zw9IexQm0tl2cPJL97PdMcbvGX+9prGmK+LJUASe/2+Q2ZDb8VhKnYHmsUGXhSh4Lw59MpWLME
GRSEr2lQxKCfp9sYHT+EhOzG77lVlf7Pf/MUUszo7MVqGz2VCY8eY/ghi87Ksgrlq6f3mxXcUVAN
V4dF6lAOY32Sd8SBY6kzsJ6gwseXkhy4Y1Tk/MJ/O6LAlfXDAnNuXWZW2FB0Diw42wscibooU6Oi
eybXjx1ihu34EkDZmV5s+THcoYWl9qYRpdVbzad1IMw26P6f11fICqas6j7U4DPBaorOK5SVDkp/
xLiRgxSqN8Hu92bQ5Gznl0l9mXH8LS6GoH6htyUA5um1el+f1rLeSdekXu9RmOb0A10/2ZZPDYiM
4TJ3tRvYr5q//2UwoYMf2cUJWdjGcPl6BlkI/Y6cTY1wJLddjcHXCRCQWb7Ltt8Ds9Vjf1XmHukq
O0Hghf/RSwAW1/tk/0u3KfGUYDIIxHx+AYZO8BDoacd+rngNl8f983QdbDhJV+dmWUxcLmwmmMC7
Iz2xV2IlO55XTVd6jsz804teJS5h9SxZvnsLGCQlEHUDCY7jn8+0wGN6nyjEXofTnO7Nm4cKus3P
pYOQoBBDpWmpS8fgraCnshWqLR7HxS8dF6zEfxp2aVS6nwt0cfTpVdtt5YID0eppuQFKrr7GW1iy
gkvVE+BPON87oKsXD1ASme+G4P5JQYNsfmMnhrpDR6sPCz8Oski/hbNcz6+1vdK3Gav4TBn7NZZz
UUvLfK39EojuhXAS7S1pESCZGm/DVFgAxq7iEq4lYLldYFLtQg9NVQg5UR6RHZVxgq2FJDBu23RY
Pmf3Y9bkRdn6082YW69+uprsURCZ2fCSWCsG8UjQFBY67poUvzXDaJOmPo1aP7/VpqUYe5Z3eBUj
SXalRnqLdKQE5a3COp8PTjly1q52TAxyqtAqBN1fwaLSRMoNLlBs1ODX5/t1yQMl3rohLIL1YNgy
qphJTLGTwnaROFMzGpA1gESPdsXP2n1xvJb/wsZXmM9UDCB2/wzsZdZ0Iuzl+nwMEWd2MuSTGTki
/MzrAiHa88jCrvuEd2R3ibO0r/PkxUmcWnAJphEs+bps5XRVFMbGYIXGA30zLSlxADsY9ee3H6wA
PD9MgVqpS2fKhfiovzCks6IVN1VDIt9M1V0x/6YtKFEDyhzjtYBQ2DVdLA0EHoDB0I2ro7EpWn5d
T0gQBWxRetoGsaPJiQNg9s7c+XKhzFLlsxkTkXyLS2VO41CgQ3+Dyl+WuOCBVueL7KteWF8Z9aJa
g6hpO7Fz/fUqhv3hFSxDE4AHxgGT66saVas5URtE5oQrf2zCh7oTKVe/ZHZsgn/TKwOJP9zwYGz9
bgFp36/POYELPg5iW4kuYlRSs1y/vlkvmOblN8vkAg/DrU2PfYlfyJR7MRRwCVaGU023AX6T+VXM
s8aVS+VBgb8v87vONxX84L+iO5OUJPNUxwdzG4or3dNFl0WHbarvsP3Lgae3MR/g2ZpT2LeJnbil
kELxBOcsqYQMgOnDCO80woqPl9/Rf6sc3lWwpcOfjIHZ65FNCdTwxj/eRUdwnU+RepckEgViSgDh
ZoVqxDS0p4dLCnl2sfl3jSw1iTY5lVnFn/dEMuCU1vzK0GOMN1k/HPmIia1lmIcH7K6Eb+v2B7kS
ewE/vPONT/BavEsF4bAFOnJlO7M+V0UAfXGiqq/uNumSoaCCkNDhcoj8jvxn2r5ZQB3csm6qVEky
jborD9mNPBQ7+RUsYU2IPKSW7FJ/VUvd97A8KD8zWcTm4WU7qZNOf0k9QmqkPthd/BIbc8K2Pj+n
EJPG4EqK3Us09efNRyltG2uDF1tAbrVcJaQYnQFRw7RJgKvuSQsVELxICyshwNoFYwSku4dAIG2h
5V8ePPXM1B+oPuP3PVNTD123Ui89lI5YEekyiv3nxLMhvSsg/GDwHmaOABexlmRn4zaaz1jb1E1Z
Fkm9tcT7sjRWGnOLT6YSv7rhY6vR5JjxOGAGyF5zeA2+8tE5y8CHbtIXtftSRLYDFLkcBpW7ShvF
X07ejzCrma/d9j++gE5LZBs1Mn3c1UESi1Y9MzFCn5wQUdYV03tZBlThXkaqZe+I6f3C8KdjEdX6
zs3k9CkGGkVCE/TxVB9JgBAafmT7qF89QaZEvmmVTbOhIWk48dyhaiTJMuNzI6/qHGiy7HJcENMa
ENPIxWXPa5aDJ5liqjxJvKYuuoc8gXqQCy0zGlIse0OgYmY/2K4pK7KRKkcRgOvGhSdkhtOJNb43
Ia7dsj7bwaWKL2EauFgXjrud614+oJBy+GhJXcwPcJuwPX2ep6+bwLV3D01wqYqM3GYMeSmpqMU9
eM5DfBuu6zKztqU0k6HoDkJYaSPv5yRDp+0Wc2IyYoqFF8TMXpmGsng3HPDqcZtwMAc+xTHANID/
nNAgNwPBSI0LMzYIO0ng8zYaf1BZ1L5/eWlyM0g5C8fUBTH1qNTdSQKwhEIIrOirjDCnYbsWQgz2
iPwoFrzGd30mZ1USrdWrImKIrmQXOPzJb8W8gyVr+ShsXOFyZmFlJBOTa9e3/DjWeil6sIZc1/OP
ICSKTyQdEeHwVf0eTcUFY3lmORG0m58VNKYEVHUHMhnVBJa7K9NX4xLJIZ65lHTn5U5PqYti2AB8
LYcX4ZK3tGJqUGHMBESKJVeQM/1BjlUtVYXQtNSyckBBW2uEGHgGm4ltqzXIpjNnmmcKzdQIVU8q
ZjqURlovLrvC69RKOFmEoXPuP8ouOXsbAS+STFEOot4bEmT+NKUu75ALFtSHWVharV6SaNvZqPEN
L7a/pm1/JceHUeXUYcFx85hzTskrdSqdMue2Jul+RCvWNcL7VCeJ3hZQGveQXOURoQk3aYCCLSim
m1j8x1FOuBMVraddOqybOj2hdOzm8iLlMqggEeAUJWAaB+FGf0JgCWnOnbGawJD6T1Mki4ACGDZz
Fbk8Nz+d2S6jjbyIruT+hjD1TtmrIOTVAXuL1iKsS49IHlfI9CLWifugdnxCDYJw5qRI0FqaRN4e
oqyOpHXJRPcX2k1lsZQe8tClXMnKMQzTpN2JeVbX2IhjOSiM1oiDSL0V6zf9ed+jZFFA6a0KRnNH
6FLjsPgLpf9wuVrpjGxSug4QZ/6qfjkhevsgTYlTU+50dI9DAfieiP7o39hb0yiojTY0OZmlVXeX
yKKY4QV+reUYLhJKODnWSpZDBRGX5uzh/btoVbTsm9LbCNQQlcOo2EcQbVgeKEH6L4ggQoVmKmjV
sQ48Kp2X4noKfyO3IjdZy8IKHiel6w2XVnp/nC40phcAb3SVe2UjqhEYjzlU1G9CljBRloEbN0aV
B+/VQkRG+K5gWT5CGLikXd7Ksh7ddueB88/bn3EGY3NbtrUFMOtQz8lruPfyHDt6c8hL/6dmtJrc
4ij1juOEpu2XI5woIVU284OrtG+KK4FhdsXVLYUwPbaqmXm6g2eti4IdOlC6Qrm/QaidpGQBT9S+
ve53BiTYjsTPxnuD0+cT78uc3/qUN81mASL5+JcSao5xCMUEUcvAxfz6ZuL9PA3MySO/YDDYsWGB
FQ03JRQr7cmAF3dFs732kiiDhUXvx8H7Rh0C+spFtj9gUA4K+YbfuJd7LWuFfzC8hrNPGC1AQDVy
0o1wtIW40dW2gLu1mqv3Y3/fPfgzj6asvOTui4aHxPpVXrWXhLQRD5XlpWmPRbupEXOBVhoSoyrL
nH4InwhrCh9wjcj1WmqfNwmraKO4QnlHptM/JiMU9kdns2jcf4hI8iBDynrGvh3VXPYeEnpEwQQs
U3PEcAbeRHpXxpAL7IGXBN4BFcSgvvbSDll398ekH+viAwg0gM0RuogDAeYqAWqYlQVFd5GnbD2K
KRFGyizA4K51M4b02vSv4Jb8BseGSiBqZh9j3YOvmM9mIYGgePMt8ZmkV1zzo+lUgSNHrbZBYt0W
yCoHZ6IwWtwYcs7E/wHaUAMZFd0W8iIGNryY+0H8+BbLP9ip3ODSw7KWbmWbLTQrq6tYTCFCt/CK
qfRQelrluSSTaISV27/XmzEMv3dlA8DaWD9FM67XqHLDTSkK87nRu4DngO+LcyfPNTTEQOSGWLTN
3dA864vlMywSIw1hrdpqIPtSiRi+gGROwuKm6NrjZ7b4RWFPh7vm2tDM54o2BkcZzhD8GdKAwt5N
oo3X8kdrRayz8CNPUjUokkmq8JvHiYBtn5ERH/ziTemgiRB+DW3vEsGCRzjN04H55ahRlpyJlX8S
YziVCsaJlyRuoomXWHmr6Dv0uSn38mkyYqv6u/ysQR1vXttlhgxAzHqYbfJ54vfux3sfMmPU+3M/
//3mZPATRd0B9kMd9C9xKw6YH9vrl2GEmQHBgy4uSUFD7+ZpSUvuhPlR/bPyFwBB4c2aVbcHHxSb
wfO7AHXDYpkk9QBLWTdqY0G5aITJAz1NcO/k2RR1toVKAGZCPbSRmrSTUVv6ABttnZcjSwTwSU85
U7/IbXrGDv/in6noOi/6gSbMo6zX4W6atyvsOooDvl47FDchPD3UBe04Sx9uJdPmhNYhP9Gh9gNm
BAOREUcKBp6jnFVxmQ4T2QwXb+aP3+YtR/vR66V4EpVQJ2LOV9CuapjrWNip+8nEnSB/dfcHgSmp
9d404033J4EyQxKaL/u6OfSdOqg1787viLCNg28wfyuTiIhevjRgkA8v/o1nnwVuULbKGJ6GzVL9
TUk7Rj9TlDwcSV3cvmznvMEi6KPsruFhs7qv/mpBnC5GqD9UZYZaZ+68lQKK+6bkrHDkciLj0SrY
9o2TZOvXYV0qV3O/Kf8w0xiY1KQ58X3EE23S1ce9DaCMU+PS47VjST5rhH9sQltajEil1xrq6MDp
Y2KYpqUM8LMZlFPKDzvZWQKdIf3OJ/9uZsB5mJJSW5R1VmulpFoTuQ4Xuobyhkx0vnc7aV33CChI
x06XcXI8jwNCoItjev0JJBhUfftZlHbeC2ENGbPwNPOgkDsYWov6Sx/rm3/AMM5S2PzK7pCcklTd
dNVXVEerSrj8w0rup3g7jtc02epeSG/su9II1PU8DyO6OIcPGNsOCJ0q/tJd8nFGfmjSJN5or6xW
Qsuyslcia1wiwk/Imvf8Fuu1Ej09f1zgoDBQ7Pte225GMK6l+VfXqKy251uxAZIJ9vuUUiZTg1vN
FKt2eFcYVcHnPd8LKFl4agV56aci+oHxDMvzgsmKXKa7q2ee107bPyDcNFc0ToobUzhcNZdc8H5l
ufAPMjWOUhm+mi4kpWKrFfBwEZAMVSS4++JC8RKBh37DC1pihD+vmSEMj33x8Hb5hE58V4yBcidj
x7T968G6VG5YmiVofseJo2gsnSYTwwxK2qzPiwvA0rco4/UphM4m+qpVqu4YTwMtCjcBsNT5MLGA
b4M8U8rFVz2H7VuEmG+fjdM1A+5cna/sU6ueVl2jhWHpXGWuIpJe0YqIFI34xm0PZ6O+CLwH7Zj5
6UlKQ1U8IN9lZ3OLDM5KKoQ64Vfyo80aXT9gEsVnBgG02KD6PwXuuru2c4Ty2DN+OnLhcfv0wQ8J
ErSsKEnsZt7UFzhlnv/srh6hgcXbgEqjpUJtRkSck2QvzfyftJNlg0yulJsr2Nun4k90Ff/aX0eE
lkmSQz/wQtuv0pMrJ3QIeaZOT/K7qb2CwLnAsKuJxW8tVnrNhwODFoZVGPi0RU+hTtSqnqJtFyn7
d1JCDruub4S3Te/1iTJ0WbcU2gcMV2HUfuISfzD4i4Td6hRaQBg9dO+DUAbGC2x5ogwRP4h/rkI9
0m/eWygpYwEyqu6g3iPo4UuvnotRujDON4biNfERhDyBpNtNB9B8ZqGX8jiW6MOSi0ANt+VleVq8
J8CTrF1/rvqyKtge108F+tjKgt8kSSccQGsN+st5PI+uKhk4+YAraMYT7TaBZg576+jzwMFU8OHa
oGc0xhTOB22U88secDkw3pjGGrTwLBFbxG4TQ7TQfw5x2k0PMqq+Ktlacmb7ffnWku5RRjqDArtf
H09SkaqjPSt36iAJNBVEJIBUUx529wZ+/0rM5vsz+mDdYmHR7B16O0QhDUFdD8YpHO1C6H92JgM4
YnTSlmFo0s3b0r1WSl+V6m7O64kuXpOpEYfENt8rPLdDBE5oo42VoHbfhf70Gy/5Px6pjQfW8FEE
wYO57B+tmH5Ud1E0vJrgM7ZIBiS6jaAQ0NJiXlypTT+hJExa7qNtdoy5TH6bhR/DzdC0JfFNNhat
SdUX4EwaxHybIdV5/IV6EMBpPka384EXPXvMF3JYeIplFMPD2SIS0GIYYBGhCF1pQ/owtHvOXhXb
jF1CXkaZcMV8o1O+X7PkL4RjJUosihD829lO9RgPgHlB/zyQvFgRdiJPHZvhNaigA+MBHOCc2GDT
hudz8XLWrSNr4QLs/IaIaaVmB5LeIDLfm9bxYdea/16kC5OBM2uejvWIWK0h+aDXMPOmesO36d24
IJnmPspVZ23gZGNANqv/XieCKXf691BAJ1vfVLlnTAWRTkJrheHPyv39kUMxHYD4IAvfKZrpWIEr
2l9gOPkImXl92fJSQ3uWG8bb7U58DSjGyDietUk5aIsE6zEX2njR1RYdbuMah3NzccwSYoCGvhZT
NIbdw6PUo66sybuTdl/AQHoZFoZntEUjoT1os9vpxLUthEu5iZKAwh9oQwmQm8Al8UFitqT8yTcW
mzVzmyWlrC/nKvG6PPrMRILF4smgbQ6Ov9jMHaCMnIdIrBHr0SgcxaQ0DCsCoVnmhpfZIlqLARh7
KYJmFBuw2K7ljC26+3eJwUHu1/BfmHZuUkn6vwmC6f5IPAOFCxFiELZ04cSNaTRiDokuQYnl+7hF
R+Ky8GldHNbYPnVSjvPNVzKGBuWNMJvfFALJ+O/tnXz768vegQMpRHqp3rE4mUEHo9q4zfuU+1tv
oszatkFYu8GB2Vu/cwcGYKR9MkuuxEwTK0bwMVbQyx/MinFFb6n9EcFgV3lAgoD/6UOuAYx/fX5K
ofVgZWI5qVizt8fj97WbPHy3IXjY3k9lfTxDrI9nlRST78LRN4pjK0Rd3u9SSSo6MeSQn9ElfRwn
bniyQQ1eOOF+yMJu0Hem5P2Yz7VKrDlIaUl7OyteHTzyzA6enlwztwpvf7upNJ3IZ0Jmvj1M/JT4
roDIE5qSr2NFXKzwpw2gFNS9iCBPDNFZ+cEPu0NfqUsp7i9GUTG3qJIm1hhEkbk9d0XcmKa5i937
sWovSSU1tIebqalfWfmPD0mYmnCR7SUhCELjS1m6Q77d+AfhA0tlkq0Ew4x79dkcT5OoliQa53wr
68po7zzy3C9MFumxD/3DGfXOF7uSIywZLJ2x0r64Sr40AgPxSKMtcPt7S6dvyMjoLgGwUSGQFSwz
fgBUCijZkfkOOdwO5W6p62NS+GpnHSoPRBo4uMgPUi8u5Ln1EjYzZJo/1hTyWbeo9qr3E8O3sEn3
5l0vy+ZlDaa1nei2vf7DMmBPmZmXqKecBlHe0a/zij/+7yo2KOKS0Z02ebjzSguo0Q7BkszKfROE
GQzEFvXmOzqYw9U4QO3+BKYTh3iaTNbP2sLvd3s5/2tt1y92D7jApxBM9naIPc4BJ1knKmdDq3aZ
s3CMfH6+e3V/ao/a4pInCTW1gDPMtTKMjLjTnqY6flDKCDu9ZD12JpTqwXzvc8m1t36I21IvyvUP
NQS5sFEaFcFLqkO4gvqgvMxyZhFwG47WL1U5UiGJOTmrxhFgNzLshSftHkd9kW4ZeM16VngHnlmj
VgjbPuLlfzN+kkc5r/LNjbNfzfci0M4nFYeGSXlfLyKt0FdtqiE3F0fM/aYdpHc66cd1BLmqqPlY
zqmFOuSviI4RJwg9k7YJV0oTVbFFuhGRdsuML53IwHyPMXEwXK4oPaVsgNQJO8+e+mTRWvvgcB/0
CZz/yCifDOaAWwVyK4/hvDJOfu2mEGV9E3GbhkXAFHdFN9l/xm82xGk5xW6oEtsmQ90vmh8R8JC2
oFlacgy0lhlFqpnGTkaIPYO7TV8eMYM5O8YsRVD/0lefERQbKd/e5WF5taAORux8s6/LAAhKoZr3
xnKmqNyASvy1VLrnxv2NFgx1c8Szo+jW3yvvcoQuOee6yWfImhBm5wT5jWikdkjaaDm3OlKoFFW7
gk1acwn0IhdJHmnFqLPRP6GVCbWE0FL2+adzDONsw7wHlTKXsUb7QobUWWAmcCKIAWlIokpGd/ir
HnneRmr7LqwLfxyo+O80KuYZLjhRcS8N0iFOxjJiA9dDyqoGJtE/CfgWTc+WDO/cyDdjRfPkRp1X
mBoBeWLhV44q7d/Edblei+V6IND6k3FD0LWAaNDxCpTwU9yKQIdbNS77n/rVRDeOOE8kFhMDBCCl
X11DVjIbPQTJHqWD7+ffkFl7ZOzK824uDpart3ppUn7Q8ViUhVq3iFkoiUsIJgSsQ26ssQ2hejZw
se7tBX/vdfRZRubEC1VGmVRp1T5z0LK3FmB4EtlQD01ta5GuJgOJk/bWvwKHsDJGKw3ikR65yoaw
ul0qZCQIvX6dc910mivnBq0PmvT9dsR1X4QTsZ0+pMQE52vTQAkI8GMX+IezYSKMJvNn532SLT4H
IV/wnYkhosGo/VH+lCJ6/MGXVSn9OknPKP1yIp1KSqjPUREb2ZPhhv/k+tJQE3RY26oI+fFjkDlt
kMx+QRg3fVG+AfgvBv3lQv6H2nGHdbvreNNfklM54uHc0rTPcTDEy9q7dcENrcISSJXudevgb9v5
S58dfJG8LC1qBdtcfaMdOhk9VBIFFCfGvH815Esa5O0l0TS5uiHCksMvR7rbEcZFfUMhXStNL6Xn
vPN0I3eklhUR7mLRC6PttAFTecHIUOrKAuNyKvC6FbTC3YwIUxmBC3F7p0PTokEZIUBZFbhuOzqL
+MhbkcC0AoUfK8KvJnaBKLdtHQPrjCQxpYJlrOGH+i/MKKPhlEOBGz3FqNY1eEo3n1vVunn/BA30
1rLQzRQNvACVLbU9yUTezgV03XRGzQBy3HYkbGQ0842hvdQo8rHfLLkNsLvF0eAMEAgdnezMdwEc
vjVL+IsxoVfK2zzU6x7biiguFqtBPC6ddgFPsGZyJfXuKgk5meFuh/NRdtbqkT9IGrZxai6TiNlD
lzxHNSlOvi2W30mqYhOxlyMULiHOVh8BVubP8o3SH3ygiQlXc/UOP/e5K1soNXX1ebWJ7mpjRAi5
WbqaJJWkcSVyF+Q+QvYr2J8nwO1KDJpTp1auZk5Z9H/U2I/eFcfH2JzBx+Gv3u6UXQKeZCub8NBY
7KR2V9IOBZWPlTPDpzQjeUVgao3RHNobT+bJ7cboTO9nhu3vAuOeIEqSsaDNUZhSUA5J3YGSmOLD
KrdNYXUHm0rk0ZO0qLFIiqTaYFkS/BYlfm1fsi1mxLdDbVl3XZBtgeDxIkzrK0cqOBivwq1RBAHh
nKmTzNdkDkrY6E+L3FZWVyFnMIyYgnl8kV6Xc8Dy2oxWiFNnKhyBt1FrtnWAEvBjtkzYiWz4DFDI
XUbAoOhsaHbSAlPwZy24lg3aWFAtBC/josYL9ccgmyHIltxQSFaoQVxu7dU+ITInYqaA6OxU/0xi
Mgig0I1V38dhBmItgWCoKqHh07zzQ9apLk1tc+WWgND5ne9o8Rw94/qgPDxMemKpccbAXEg1hF3j
FWQsfEK65RA0RYIpx4ZQ2S9fWaJnJH/FNjNRJtvGKHLyV3mT3oFcirN7pIeFUBIUOas1N6HqbqaI
skUd3udnrtG01OqPEu3uq5zK94RwOL9oNr47LBkn5AF1+P0nMCzDHty7JXImGoyYzCuVw99ajbZo
DuzpsLuR4tz88Ki1gqpjLVzH7SPk363PWZBEDPo/qWXPkQdQxDO4m0dnED+vHTzuUvSxGIHPctH8
RTx4I9aCLl+XLkj/W6z6BVLMjcnRvpr61PFgVOFAWqozSd1c0q6b+/KRzQVUDWMmGbBxFvCgr3Tg
4CyvePj1wYTYFbpL+L2tyUxoi7sxBoL6OYz1khQnzZiBUqQPC0XlXmOZv6S+TOy558dGxkdo59F6
f7QeT15Li46nhR7SV2/RiHuT8mXXloxPqu343ezyUZeRwJ/B7Te/yjp4H7gqa3RF2p8/JSg6KArF
sGNddg1OoGzYvptFsQ0gAf7jzCgvXPkmPtAw+ohaFm/Vl+VTbRtcpNYLCUYJSbhriTKIKom98FLI
DGrReT0BKdoLk/ECFO4lEiaPfnp/t2/byGErhDb/HNTaYFuoJKcmGZdWr6902mYfne0IplW0zfv3
hMivkCe1D7uDQIik8MfwKre2+Ur4+eFvxrpEzEJTl/4B0ZgZKIp/yLb3aBxLtPUVJvkXbkCiHP3p
BlvpBuV0wmT4iCpm+03Nm2N0Qp/KDbtj06MDBEzYFmwtP/d11m5blafFACCMy6qemEvuT98qqRf0
ZyYz0YB+M9V6v99VB2GDhTvWS4jVRLQPWP7lKtWTKrnfEcsN7ZTlX0q7Xlv0Sk2gNtUH2EBHfjnG
JsZTp2kH+sXW/yXaGZc1WRN96SqQVxv6fsfaD8+OgVdCHhPRnG+2cw6+lEXyGK73LDYyPoNO9kYA
x6egYQ+kHQE+LTIWXhtRLoRDjFjJ2gF/yZ5LK162JpyrgMkNIQjVsS9YXDv1MuxLs5v/c7eSn39P
gIXCWHpwhUxzt0iXfAlmcoZJZk/btMUgutFJ5RuJ2Mv7Q9uY/UDjkQk1v9VXyVbFKJ6pvIrLJ1lq
1ox7i260wye2wWDyX7CvturIsAEpTnWNgy07LigswqjbqsONrkyExx0wCV2NqF7qYAWLqGoFMY/e
Gl2SEtkMSLSLg6MqYZEGEtoy2sZkwM6q3/aAH45gXMX6Zyw8LVNBBacyjfPMKeW00VtR4uF/cSZj
yrlGzSO1CqDukHZd3M0o7d+WzwzcJq9VQr9IXKBdu7XlJMPl7BWooz5kbhGxxzSlyYM+WEEvHctH
TzpChw/8r1iAMg6X7C/obT3fvumsbJKIGksbHWGTkyJMxbkXonFofXfHFrvWUNeS7lQwuLt7GAO4
gdXYKyrzxIzUFD4d0RQpXHgKv0QAyMVnwiVLDB0abeSyD7MlMW32C29Tqh+be7M+eDinxllv+3dV
8SWzFKwiynOEIKb+kaKr8LycOaxPoQAZNHSbdgu5QAgGzLcNM1Dyjga8Moi59XytC4VAdmlFhNre
kuWRZnp4QeO0YVdF7dULvwzAR+9GMC1jk9jAtSG3s6t1kHCp/xqOEP6bEovfXJpfdhiylwwufnyQ
WHA1FWKgyeWJJ0VznjPFWdRjde2Kh8Z68mQosliuez3Lp+o2caPCWi2Kf9DpdNLr+xEJBGMUkcwf
7lE+E4vguaJ6KIqPWptRc9/f8zUdN6E/jyXgNOMZziqRYCpA4EZW468y+jKP8SLAHeGLue4+TZ4T
3/z3AP7gzohocyyuVZpb9hvJQg4w2G3q8fQuTXFqCuDbB49LtEcTpodnl77PP/f5H0QT7/0kpyy+
xnzMb+dMBrE7A4T+oRnFMSUIit1ki01WfxFwwmAVrHiLPTEmvqiUNG9ort+dFAKYvaKVKqdEkFN6
3ljlxJxhjRx9TGlvZh6REAcr/e0WYoqz31oqp+JRcmcE3Rj2HnmvpqUz4tmNfLV/PMd5vcfOqToV
gTy+ymwPwyHqk79aLcFqOFHapmNsrdHoKwqhcHYKqflBOKPgveeAy2JjmShh+jAKzGK/tJpQEeRz
fa/XDVMwKM/GO5jkeFUGlORb0yJgZFuP/KEtmxizLNRhucOtGO/8zPln6WWBS+zI9yUYnjkXNTcc
up8g9qTjdFLnxzqGPLZKefKCIa5WfP8zoO0Ma96kj+BdMX3fFPtm7SidDHSwHejqNpZC8Q6m6M2W
h4YXgBxQDv5oHd9xlp9lTJkd/vc/sKoRJf8w50Zil15EoQcdavRk10wVahQvGmQLqfqNnNkoH89y
7GGLmu3u9aZNaYFxZ1TiaqQHL1IAKEuUgv4tMQvekwgTdI+atW4REAcffaNCc2tCpDLiD8rWnMHc
i7llF9rYSnIDhk/hR+rTGsUBhijCzAGV/h5PNmFiMQjf2pgJMeV7BmUs/XPEELIbrc6Gmtkxxn0N
3mtXOqEUrq2VwU3+F+wA1lsxje0FYOsoYogn2Tx/PShPuybtb2fk9tSdX4W/57b9UjjBRqfZKEhZ
hblWG/qdrxCc+w7K5U5VN9G+pGUA3UtHy+U9Ezy+nPqavRwlsp7x2d4Y+H4rAwW9ECSVDW3a+kid
4MbOoPY+HSH5iNRG+iAc78enHxEd9t8rTPYvXgaDZT+tO/9sESvqDKsQPqe8i3UbNU9HWYbDD57K
4wNAJX2pFPPZ0xtd8/tKPcXA0bNLoXwE6+FFEe5YXwn4mD5JkLW/mmzrJzs8AVyrdVunX/d9Effo
IL3J8c/FrejH+2sBtKx5OsPaeFx5i1V07407cRAGg6cJLIwgFjh4ERFfgL0VH/Z650XF/a9cnX5T
QoKuNXQsx3JknTeuUiY6048bF/KTkW6j3Zuxg2FPKzr0u+D5VejWaaudky2JLC1qDC1ftqhb2LdU
XmN4jj4zPUmCWaD7/dLVT2+Jm4g4zDIQC5Jijiu8mgi19BOxEHgTLEiI0JjtF0DpHIwSfhdUYWEx
R7ZBTuCJNaU/EnM6qPfqgCQ7rEQXB8z8pslThsTzh/Z0duXZEPO79BqYihzRDRpfvj/Ftutzi+Om
zyoATLhHxQA8EqvWWVVxvAIwo0HnRnKgJEG2b/iv1r+yNAUyPvWYhha6gQVY/8ZsvwibnCMd276i
2B4ow2RwtQomxxmccTWWB8hR7K1fkuLW4kgXVzZFUvjX3JX73cuNwzT/NTSNO7kwJL7PM2F/8anM
7dzza3lqN1nz9nzCZHMqbvXG/DH9L/ZVDh+92VhFnfwg2IvgGom/zxRb/0PrUP80m1ccfkUzzxoG
yh5xs792ZRoZc9yhm0LgeqIGMiF3XYc1h8+RxVD0hbiYEOOiTk1ucQc20haGZeZp59vLeuObIC9K
Kr2obBg3krIOoRgFNl0wKZPEa/SC4qBYp/rDj6MytvYdYS6NNjOYr2Qq0+RVEmWEYsogE/8tNlnS
TKp90PQnNEfTSYYGJZsJz/nP86uS/sIszGSDswariNbSLmkJ70Di7OGSGtOVCVz3iL3c6d2Ix8M4
m7yVegCQkRhS31ag8+TagArlZVDEQMd6ZW02NZ1sWiZJo9zePfIceqHCobi3gAkN+4aj9SFeej7e
SHL2gL4i+t2hwwDW+pPZiYq4Rlw/ZH8powy6TOeXILpC1hxy3gTDVzx5Mdm7pewOiRH0v3VrkAN4
ulENiWr+1XulhkhhKjpJj1JArBVYl3hi3mW03rU0rv6i9IKcbDCdfU8bK45bYcLYSV+CThEqM/vf
di4/u23/TnorZhIi4N/R1Vlq79cQLdnio/f4oDv+FO7mfEgtPayirJQL5B8GCoJ7EmRx69BmZpIz
pWwIPk8V7U0j8XP/uTmdVn1FlJB8P76oSyBB1QXalib7cszy7H/k+dtUA8DfRuYn+AX7Qv9W2yqs
vWLERW75zs47eHqA56OuaJ3UDhb+9BOkA6f1pKHrWcdh2i+xZ92B6dlwdL2rWyfwV/9jsSAzL70c
qYXY1NlTmT2ZGgYyKefhjKUrmUZ7J8AO7Em1Y8qnxnakIEpNYndQ9M+tRf45ZcLUruKHym/EOSBQ
PYsW+sH0zGaIEES8GOVFRt47julCA1O17gczjgR7BZXSJ77+xS1VjJ7e+R5VhxTiHsUY1tkdFhvH
MFhFgGUatttdT2Jsr2stUgDQL/7CKycQNRWvZhUL78GKzZZlJu+3UJLyS9X6E/fMCPQADINvuk/4
nDgSsqdG6HVGyaxl/SxznZKvPy9lJ0ieMUJiIqrCwAc256yYJpdqI3RXgYXNQrOAEgcBuA7vvifU
v/GrIeUavUi+5pvyBdBVb1JZ7h/PK9dhpPWnQLnQqcJ/HH9OsLtR1yurjwejZUnd0DBeVq+rPDpl
J22PBPnKs2LiSmyOxuyD5QgqimFmgkineHZxdMu2RY3tP6QdtId5tAFnKekVgu0TTn3lb2dOs2nr
G/HXZRH5K548LC9Nsn72U1gbyMA5+MDk3puRcTVpwIoDhjmdtnbEfcbULMLpNF28I7vzSKWriYKK
W1ucB7KQho59lTnFvvJjL4Dok/Btb/gU7LrHbAUZ6dkE+Rst9TyEtjMHTTccpuNAC8KQa1cNxeb3
EnX0yrd0xvOx1Si6SnP7owfuM5h1309xzscm5ftvSIJ1cC+B/C/5mAg/TjFgSmw39XlCc9cjsbRv
EDjskVW8vto29Ec67ThPZ3pwGtdz/PJ6/9yVF+iwhysIaj3suBxgpGgWTrX4JJUCLy4YpnjesHIV
b7aJv3N6glpzBBo8G5sGidOCRAgw2pRWpwowSex3BYzZMYu+DDs3a+viBH8+L0ZH/rINqLCxH8Br
CTSPhqp4N81cTL6RBcecOFlzw86psyb50onLePBRfLdUOMhRcoVWNSy5KppdJwA9SiPWmiKdFKvi
x4WlckWflehft0idYilO1pcbKLmzLvQAR8v26sH77/CUXHGdtzNqJJehUfa325geAX52jPmRpaME
jADE0ikMCOxJuqxIHqldOwntqkjMdl6fo7DyVlnn27rmL4t29syl92xwmRMfZdGpGacxVicZpCF5
t5zocwOJVaoUTtDI3DrpayfcUapoVgPlHEIb4Z2hLsklEk6y/3KKMCcvEyaoQyNkEfBcUYMJPF4D
bq8X/8kN++Fx+f+czkYtG0hr/XWK2x3OGPkUNJQ9h/nECbU0RrqR+xiUSe7tctjxD7jeF0IveJ40
sYgHI1XdeLrSu3vl4VeoRg7+x6UlwvOLsDSQ2lSR0lYPBtnETiXgxS0WLQC4qM/LEFAzk43YPd8K
ZOloTFHoPivUC+yjsdDPus9wQcKIPqid0A9/RR0iMq9lMYqiCOQqcqoscueDrZEBj4DcYAnhQtux
W4vV7ggNrAX9rsEbeecfNPRWf7rw/eq6by0oBBEWPCp6mra44Kk8tI0Ii9uNw/yVcUZPBF6yPfjo
Amv0m8EpdpqnbKdcvp05fr+URNaG/PYLkpo+k0lak2FpM2NjzH3LKAhyWJnJqmgfJli8jmyaq2QJ
UlBjFpI3rCc+VRo/1Vowi3wF3hkvyTdTtT0Lf+XIgeAaTUq67tQQYBc9/m9tn5D3jM+kEhTkS86r
Z9qJ2DaI+6ChYLnEqLTxPH37bLZb9Np2RodNOOgJxgcEjeenLURYquOJoAqqb49d9n1ck9kI39xE
F6EhpVopD65im0I8GGLDlBTIogjiQ+J82K1dir5AOpAyIeQcrRbmkETMv20Gv7nzRzJ+nOtwT/U/
0+uNtp49sCxlsbjnmc52PT+2x3jubP4pL1Kn4oFBeeWIxuixqPBqumNGGPaMlqw2220xZrLVKcGr
6aKhJd0MKDWx4qr0J0NVOYmQIt1ZdHwuLCvGIc+107pxMJXkIpyFduKu1XFua22zxxm/NUE8pP6a
KoIvKMf6HUMcDPOpumYptn7YENI9etQtgoRWl+8PKjtyvuBgeNIiOqMmwt1cPVRrm0SWmf7+Sezw
FxT5ijjSuxSZUkcoKb3xObFZ8RbyJ1XXFfu6gKLLkxaZQRPErplR+yHUUOJoMuXNBlXc9rQfcemJ
ZjD7q2jdR1/GdYKiA8PNOeu52xSnv7GoKCiZMHA1BMQ8GCPYMhMSathQenGZaCGTdZ0/vQIaA73x
0Vo7jAJUgKeIRhYT4iavPsw0yF/ed2kbjG640Htm9ZglsTN9kklXiSCljKbNjsJCXNScVGF0UBjg
+ng3ZFk6N0M/uJFu2Uv/4TH0ND7yciCVPA2NskbuZKSYp9IFXgmqA71KKy80l53Xcq9KkWJnafY1
Q6A9LmEKQM8YfE+bsQ1kBHfU0LahNj07kjEFQ5q+M9WVqXYcIweuZDyTfKx+kn8URK9GzPhLwC0+
wlmUXlsYT5WNT0LthgTsJnIFycyzMLq8PTSrqz2+J3T2Muks4UdAiSTTpXUxF9xuDJKErOQmvUqQ
hdrWat06J1F/m+SPyobiNKDy3db5TF/bWx40XJqNNMYfVe79kqjsgIaodP1DBTwsRbDZqvtU8CB+
jaNek/i5hJuWblIHEeeyENYnK9jG6pLtV5+8RysrSEYyG7dqGd8e9ERc41n/0kyfEq/QhBRGhCnr
21+AAk5Euynb9w/vmT7xdFCXebfaT2SNvbLI1HhYUwmay9FgZdZ7Vclksjj1gDK46aNVL7uPRcNt
IVPdHL0E6Z8zvLRFZsVBi72V0OcpH0MtTv4y526TM85FyfzCgF+cC5sgKQbTAMU3PyZGh/jq41b3
f+U9C7XSpD20XpqFy7E6DfRPp/Mzr1Uh33f3YwAnA4KxBjQ69ivltwKX+Mr1SAzbnPiSSyj4Nvi2
v3mnEOPkvZWX7X6nvfB4hKCpwHTn3NhNDYSEyOqt+msUVj1aTzStf10xKGCm/iCWXBjlrbyKOxEO
cu7Ih1lldtVdI1BpEhgQ18CeQpTI5Jrnl+/jiD7IIrhLHA3ntaBqrqxRAktCceRoHhEFP1dKlgbj
bJxmU8Y6jR9YyW4IaJGzn7Qw5EiRDwPGGRpmRUtzQMEIyR8aIqm4q8Ji4K+MH95OBPCdH6Q1X84E
1gRi8zyVEVzh4chr1PKqVS263Kl99erheNkpjxuLGFvBfq7AWgY/JqTuQC+ymL0CcDdcmFnNl4Ul
U6/cPrmI51hXoc7ouUYJPJZEH/KliIp0CR3uMOT6NrRmZYNGQyJhn/oWa5Dn3aIBI68gzTij3JiQ
lhduGnzfW1aCUr3BZ3wuy9rFUYdApU1RTVNmVHY5yjLiGsAxitldlw/VFExD2B5oocY4z1brMKQm
h33hidD/plnaTHbWrOj/YGfgfo94naHz5yjha5H7o/WoyPEh7ue/GcW2QWZp/zwqyAdqx4IlfHyC
MYjnBG7wt2IV8j1l+gBdVx8qcX0+bll7SRWQ2/jF5xdIKahLc1i9wWET3YwSh4Q0zBM+N+owkguH
Y2AGDFmrNSFELtSkV2J0mnQP70EO3J/w+SVqaqQgo2cbhX0maC6Pe3bfZnd76rkvTuVH4Q5s8vur
8iwyAyb1jDBy4hDY8oXloBofa9EZ2+jaVvxX9PYaPegu2Qb3Ro+GPsdRaosAd8EwwLahT7P4USqJ
LBHnq7s2ziPp2J0OWtK14sqIiLk9z1eci0cJ18+09FjCSCB2LVsk2qUqx7QXoL+X8GssCz26LhCB
OQf5STpVn1VwYqP3qI2Gtq/OMBYqsvbtJP4NPpQdj22O5sj8COkF7AJ2VAtyyBu1IwoX4pUajI1m
H2Q1sEV6WJtoto3LiEKlmNRVxfg0jMFFMAp2zkCNgwgWqdx9aGQWIeOFlsl/7gybAgx1/rl9lR1p
qFgGqv69pc9t9mC/NW4jZEDZnirrRRKmSACthk8tcw9ZNjIR1Xr+rMLNokhFi0GSapuwtZKzy4G8
uEwjX/eX9ULr7Uw5BXHki3PFuZpLV7+SvePWpjzSnnUXgWH2r2zzQKUJ4fYiTdutqUK7ZWG909oe
U5exoPUXZ+ygBQfFMYwQqI1xk+/StYyX6Wp1ilQrwJbdhdCG1KBgwRFQNKfL7/o12FbJiHrkT35+
EMqYZS8BvtWA/6ElOCithUQzdBucgQ0chkJya+/e1LzrxAEkxdkefT5oRfe1qjL64jHq/V14Ovt5
ZFuBLI0unNc3Q82/YQVFqC0f2vME3/DQj0W4TqIjYU7gBWPzfox6Jd2Fzf7c3vgwTPjlSvojCaMv
6oWGUb82GaGldDmVipHdkx/qouVAwA/IIG6H+QbQzWpYU9+X3zHWnIAynoFMvHr4tWufNb5yiVHO
tKgkyTt6nQx4gpHBC9I+sMoEBkVnuA0EZ24+dXnQN5fJBt6go3je8QlxewcaT5HuWZtSK6wjr/1T
9HwcvAi/ITkfKFaaRSnZBXB9NfpYqbiPZrdWob5Y51ItQ6kutqYx/ImEUCOkE8LNQotFFPmH0X0l
ICypZ3O4qCK5j3rIwKP5a37IAjGeDr+H22waMeVlOAvXI2MJcD2DjvNsgrKH+IoxRq5RDJAmfcme
7kdOcI0AnI34lf7E+9/5rMsApzmqPxBtvwlS3FHl1EeqjjzsLaqSgHYr6ifV2B9epEZcHhkjT0nV
RKx+RSIx6jvK4QSWCgiQVNpfFx4o7tH2kIXNBxmicoWl8HgenzCVECuRH1zSrLPl8LLgHNHIOQBa
HWJyUSUwWtALtzh2UisGoO7Evr2hYB3I5BZFoTWutwVKfP2CuHZrMi6Gjk+qkgdsmwIZiGQZoPE4
ag9eEHnJsNm3ftb0VMG+6E4jOcx1L6Q0dnOZLWl6bm/nGnxCXo91JEy5Us6dPyNN8IKOdKQb/fxO
j3fC+PEoVq4aZjPqMJHjbjI3vWnRNy34EJAq/1dXple5FGWLFLNyrwSMJe81+Atokw8KaCOhgMCf
DyHodZ9A51VAPth3W3sqGzQI6FEA+OkouHxn8IyvK6GdEQa1EUc+yhHANvS8A5vr07DGwqXMvVLu
pV1JBhManRk7LMcn/vJkPBXzz9E0nvsDpxgGxYF4Ce0ZXdIjC7qJwhCsUkOGAakbl7LXJlssijFz
Uaqbp/NmwWoO83S4WW+LFlO3xskYfJ3TaakbjKzGlpteglrfOHZh+GL8j/lrme112960y80bkHif
e2CaiWFe1O5eXjujluI2R+kba5GEMQEjRb235nbZA0XNDEk5IIh85T5NwtPBg5CvBtuZD4eDQ/Uk
bnrR1kyIz9XXNXJz4DubjJOYgfJ3TSzwKTPZpKUYvrdxwXnZfcoZYYRJMbTUpYXILyWpdVZqjlJT
h40GY56KHm50Tj0T3nZWEdOVMH+W9sLg4n+FvMjzQwQ92Qon3rlyWu1j1J8bVCtHC/fLd8a9QAmL
3xSgzyX+n6HmS/D1acDDhSTh+gd+SYfvD/pL1Y31oXPlHZUqk6KDNV6u+ENMfR2U8zL4uft6ISKR
Zwm53obGJSaCJjCG6UV5aMs3yD9dN39jn9+MiQ5PfyDjEPyoLnSkMoqRLXHu/eGa2/umaYbjpF3S
93DUkggKE4tBAauFTUAZYo2EnaqUdaxw2taLFZ1NFL5yCN++btY8RxQGGDUNrrKGXzGb5qDqo5GW
uZtERxBrJ/Q6C6Xl+NuLYX18JuJ21crI++wW9wcyfTn6UifvRVIL3hzYdgBIDikXDCV0brrkGwje
Az5Iuo9IZ2hDgRQJuUW5gELSe2bwhd3tfznX6zMNMQnMXafaKi05lh8OMWypZGVGEElfXPHPHtVK
LnitgwK1tTkUMJry8hLjq6wB379+nzTV0iR/x3k66VlXiCcOL/zzB+TzQUIMYSeFpw22wGFmUm+L
jsMRiAKeEWh5mtNcBhHAVtvS5rlazhMzcQec4+EzYTkaILXsnHxhouqUOKky2qHCZoBzxdnBiUMA
wUKRzmZx3IysYDhm1WE1R9tBRGsLTS01Y/c6gH0UNHbM7m1PnXjaTfCUrXCWbJDE5kelEMpyTZUQ
qihP+TXM2etTZnZhwzz38vgQkYWu5YdNsXXUt+H+3vXlCqtgrXrwuOoM4qRHKAqPmgzPv4sOn6yy
3Mxc123GLf8bV5IR2HpVBKGDQdTvQiZrjbTvu2+wflNBgIoJCuLmE1cZ3ZV8LVfdwzy6rcqhSvHl
qY6hTviMkopU6+/HZqLb+AonCDDrgHJwIoySGUTHxyvjQhCi855x2wvhrdMN+s9u9zPWEpFt2M2O
kQGVCXTt35/v+fLPy2y+BSZeHN0mJpYpCFA8kkQ1+CCuG/lTPfznfm0sH3AzX5DFhFhgxVD/Gx6j
XD5A8+KAmb9kigYngL5GyIiI6Jwu7/7Vk+UZjwuRouUVNRXuE6sHeNLuLKjqHhAYuybwXV+8sCcm
RVxzzqUTsk0y2MbdQzrMz7UZ5a0zaJEicWfKc3E13C20wotVHCnTwn7I1vbU4VRPIO6kjXMceZqe
CNbsNCwc7kEAlzOKAUipovfkejYrmyM4ai7wwNphb4H12yx2LwBcG3F9WFBAfQ8k6n1HT6X/gqMZ
QP3e2Ky/PR/vwwN3nQmsBUyO6vrsuhqhXJkyVkouKMRhHx5hWJAS2eOq8jB9SteBY3Y1bKfYs65k
baX888KGt0ru2ZcDwSP1RN3vMtfw1upaZp0Vz4qXs7PuT+LV6Qki3wfLPeS9o+GvATSzteSFcLP8
m/z/7oUPxY16neniGnN8Z0pLWXKZVmkqcgww6hAVSR9aJ26HGMorJZGVHUhCR/w00qIrZIP45ZNg
Ua9AW+ElSrzXIPiVPa1chtjnWfWD/SunYQFRDbX0rjBvkESeb0vEAvmbZY0QfG54JLgpubWpVeEJ
8dkqpld2aI64y1osFUK2+qw6fHKkO48vr1k5sa0+o3Ih9QbLDTJ8SFvJUD8evRX6+zZQqoDzYt0c
UZqmegU9ySVkzJuI4/IOvNxJF8MOKMPnSIVjb5VmBQ0CLhnflJpSYLizZ4LlhbRGOuB5w5RaGlqR
zq2QTTUzYBnYBljfK+QhtCQN2VTRPDYfTl6ZJs6K4x2XrJCRDd8Re6d3zy27O9wWT3n67aVVVuvq
9m+rDYv7DB8rtYzNCDV/3Lt6fl+hzIf94Y9H08PGLHm1TJfPewK9Wk4evYcjduMfBNuBBeUg/pwg
69hAC+sWkpg0Xr5FkJ1IbVslROXWlEc6Ffyo5FYldBUV8BwCXeND2yASnX0TH4ytKdPb+DY08eiX
HjKOHj7bnrkm7/Pc30l1iPuwo1MLUAuGoStHK/AW/01UlzXyBLgq4wgYDME9ugpZ4OchYQVPU9DZ
xqs11wM02NkNax6U8LFx6t32FE2pmTiD+/xPtJzaSf5SF0iZT4o126jwHcvgYjFC/lOnHSBpkjjJ
IFHQjAa9m8CBMVXOySuxtLaZr9e1RYhXfFSGeHx9BTF2z1eQMDZLqweOxVPjJGtJhaHO5TI4F8pP
+V3ZUb0I/T3ccTdm0M28xHvwBmlry5i90GFCk2fG9Mdt7OwT3kZA0D/5jlZb0Y8tzcBkNgBeUUqC
b2Tk323cDeF5j2vatPjYkK39Z0dFc8R2UeYnHyqZ7GoyoUuPEL3wBkOM7lhdbVJP4REdVvS52VE6
Nsd4K3GdPuN8xXhIPc1+8AkghXefa7ItF5MyHUUsy0kdnxQc5gXe+ZT1DoMUhqsO+pn0uEWhosak
7oGhyTmSS8F3q/QqgKWAiRAclJi5bPlHdS+CmEcj4d/8gKna34ZcLAykrlqnCjdFVM8oAXu1QEiW
0HIBzhcaZM2v/Nbc/cIJFCBaPCoomLsSdoxPdOR0GCmfA+5UIfNB/iwgsdRCdJvXvGUqm+/Gx4oR
LkaCMIyZWRjc+J9OVf1pj+cqSOFugzuVdGMUjLUVtGgKoJ2SarPEH0DzaJerjyakhp7dL2AEafol
JR/8sKY+gDzKJuphLn3wZLfT+0zBYIklbdiSD6bQStrOPi18c48smTDcU6a3WqiZmqJj4/e/Y+2P
5hHZ3cvp8SLga/+P/2eQiSUZu2zNLZFtEcyREZf4UrmxK+6KOfhaxOFF3O8vC/dAKWZujzUsTPx/
ONTZUQeJKrPYcKWWdh1abkzZq1QhkEZ+/NvVVfYh7AsiS+HkKrwlMfe/v2e9MeKu2JVIPqJ8irSw
9OL/fnLoko+mY45bt4Z/QArIOFlmkRtEBZ39k03fCq1fWaNfm6j6a/jJGmgh1dncBWo+fpIvoyRU
BmzJSAxOVtIXfzpyYZ68RJaxg+q0UneEzIevAXxUOrXAK6Tgqx1B1y8F0Y55lOm7RcZqdXu9EYea
X5yt05SWdjP682EYM0+0A+NO6mdRKAbRKE73NCHgMmr/CsWyfoQwvsrZ9rRWxGb9cj+yXkIW5CTd
dYrn0gr2NRb0j5kk/GL3mlshvEkZms32Gz6dbJRI4yexTifzgSUhVnFVZx0fCC8cPy9+paYfo5lv
QIGC8h037YdOXfYs5Ohnifyczgp45LFIMg6vmb5T7COdhkV/NpGO3G2z3Q9d6uzHKzBit/wREJ+1
FRE9pXQFKS3koK9v779V6LrUkYY5eoZHJUnbtkt1CTot14i1uVtUW8TRk73C7WJM6AgRaOq2Yg3v
pOOf8iw+QeF4Ww4jIqM/rnfdBpEYusWW9uHG6BWvL3MwdA9Kws+eS9FKyF3uOP3LpHUbRcsKHAS6
1T28P2sHm+5Iu60Y+3NRAzM9ak2hlwrjKQhuryrp4Kk91ALOuE16HRZ8bo7dtTwkbl0HZxbf7Vcu
mghyJs/IN9p7M1mPAufMsBlwnUlvKktrE43qDtKZ2k3SmfCZ+5jkRZ3+qsd4F8UM7b9XG3fh/vNF
hLSc/MKuPV2qIV+lr8tB1hxblah6OJLrTmZnF0v4wDYsTdpwmlRyB0Ti6Zu2rtl7tKL6jYe0hgc7
LAEDSH0LGQG4nWBIXepJuzhk/N3FH/GQ5o8wA3kr+XiXcl9mQOuTeDwXgoXfU0vclmQnUf/okMMF
U1DMdwMLoMhV9WFpH8A1X0dOdt9rke3HtsFP3ehhGgvqgYhZtnTTXO0Kqt6hyOE6ishcxNrc/3B7
jFlIP1yHZUQt3hNVYEf7yLIqnNO2f60gu7GU0lmh6PnPtcYzRbrRXgGmXW5y/RUAr/hsf7EUUyEk
8UqgrTT0ZeavIO/f0yd/mkI0Df91Xb5yy5wnERVZfhxd8GC167NReRifw567nq+HYXhjnPZ7ckOl
wXza98V9Gedn2Z98PNKql6xRzhR5E+9zcac/msLwt92Eh/w+GWvQmjWr5yZ8+mGHoUYhzxBeqmSK
fuwaFfnYCuWLvimhRkzr+6or+9w+SQteT3vPigP0ud3DTSz9PJcz4caiWnb/UPrkAMadv5+Ge1vY
K6lbX+KjNaqWHqBr5SlJPoIzGoyghfnRbT20iqS0WXCYYcDly8F+JqXfGHRrICtxjSDsD6lb0NpV
rwu0xXONCzwSzz1BsFIh/QDNybhga/Jd+FyA/Xh+ENUGakYY/cQkdQWRBlv6F3TzAXFJOkSrnTD1
ADyb3J3rwa1ba+XmVPEB3iqPjhSX8ddR4/V3ZNbEMjhQndbzpa0d/9Cb5JTxe3RDOPW1dZFVy5EK
002LwfTpZAbRiIFqpaKhaTo2NMrG1uT+I1mVVWaCTneQfhluXMUipz8fMbCEsg1w4LGmV+CMEJ0P
knna1ewosYih6zLRYBKk6QOGIDtWNZ0YnF7/WBg6jPWF60rU3FInj/2TFK3vs6zYqEH22mGbRUj1
gNSJIfR8+S+Qcb+bkWqO4WS67AHrDfv0kd4y74DxqckALLz+lLTyGhg+VeLY/7pyTNrv6NdQrwOd
guQqqR1+z0BW+SPxejGEBe7tonTswctc4aEkE+4kRidsGPdxCvzynsJDtt7CcNcsXoRDeoIl/duY
2atKehmWEpXMl47tn7o7rT/Tm/m5wiof2qD6L42GwBsfMyefwOdjaKHZrvkMWK19nl/Hl37juqDE
HQ7kjTH3/zPNlfcs09+AuRuywBPpGjfGOkb20kTujBXlX6vShh/6QY85xCqi6U/IMWT36ZY/aw4/
N3a3gaPuHuUYqC70oRD0MqOjhqag05vWVC84Ft9BFT2d+fonaPrzMMczOqffjPjsjA3/sF7qOMg5
+t3itKZQN/29rs1YexDJGNIyLNn9PbOQVk9lgWOjLI3nOGSgsmKOXBFK7HVpVZvGauxZKu8+eSIK
DtdpuR63dx3L7Ph9+qOQtafBr95dxkzqjRZiklJZhZx0uv8znezVDerkU/kUR1IlwHjYfIuIZsFZ
NiaWiD47kttisOZlgluY3U24GWdFeYVN6jyBdCosInGP+E6M48aAzf/+Cf8TEw94xFZegzXxktFj
JbxyzZtBlvAZ5KS6jUKLLs2/ymtHhNg0e5HG3YQWsAyboZXM/ALc/IjQUdemikd2nCZHUIxcoO3W
66XvzgyE2/0rneftfd1xMsqtY2gOekcDbulLg7WHxW1PzUkPmAygrgrFUfcBH/eh7hUKWcuU8hVd
sq9637TGZCppxX31K9wm76MX0Elkf/6t07gC6taAWZrkIMP4ETWO12s46vh9pYIACnYGNpvYGpFl
eC6XHDApaWkIdSj0HCjZkHtBlUgbjYNDeVI3bSB4vRX0y325+/BTFxu8skIFdcxGF2xc43lJpeHT
MD8ekaYgRe8eZcTHeL+mJ0lT7h6W/tG0t+L7lGiPakBrekSukB16kwZrxKT052Px32v1tUfdVTcz
Pb4S++mIieo01nckmgPFV4JfjWF1cPv9A96lyxGk3X5JvCgUT9sFOn82AyelN2Wb0QgE71R1VuLn
GxjSdiz4mJtOQHjx5Ok2wTtBvh6RORk2AmbfzpNqhyAbbplxx3dZquQwicvrV5l9EyiYKYpkrzMm
lLzwkxRnEx0G7GcD6u4Tk+tgT72yJyj3hUOrWA7wdQniPeW1yjcQ9VwglK/BD5XfsKkLHzBMGfn2
XBWNMnzsQaOXqCdwZkG8+WFqhdquFhshnDZcPZ5Mh40uDwD97oGJJgSTBvJrvgr4v5RG/7sT98R8
7Cg9XNQl3tGD57C5gEpWxG/HXZreQddhPUxjsyFMZJxvliNp8avhtaxT8FCrgB0K6cS4gVam/AyY
dQaqOeBx8mNVGXotGMAtGS6qAgDU/TEnagBXZioHaCjhL5OzXtbsSQMn8JlYxY+hrcq7Bst2sB7E
8C7t7wm1n+zXxvTZ7q8liilwiS41ciKQAMSaCN8LB8HDxcgR2lbOCysMlBMLeYMlIv4ezzzXdW+5
0+th5uQ7r+qVPI/nrBlfiTvZr9iyZkPi+ieA+mjoZPoMmFvH3ashvhABjLyTLJvGH0xWIrYnOx9b
8paTEjOzXCc7uVZklSRoJyM40mCRqj6J+JtaFH9nZES0lD+T4/jnJaXYv0so32jX57yd7KJNxArX
CFfyMl0J7icuYRy9pjUTHgB6XfWsq4fqkCJN1G0/S3XTun/k/F7meNZQNhfKULd8BTWn4UftxqZG
7QlJl4QMXOBIabITHkOr6v5SP4sb4F+Y4g8KVAGHYwEHCP0Vf8VqLI0KFmu993KxMglnm2KncoYo
pLogCmacDcbI7DIssa1jyv6Bp5HvpuYZJ2fQ0ZlRFagQawpJILNguhPzfqbTk1nhckDLY2qBlCaf
HlpcxRNIJqcnBJKcvvxVBGXqiWV/CaU8FrOAC7BwS72kTagIpIrt2WxgnOy1irAMfJT+G3SpKHM+
4UTmGiTPH96ofRCV7dpsItgegfxk8mXsWUMHRVMdP0l49rZvwXMZKHIAm8FvPIjdNhBKhdkGkHQY
IEtwEXvo4vHw9YzKEhgtdA0/GY7gTTfQ4FLpkezH6m4zmBOtG83x56Kutn7/sJrXdgm0uq29o0l/
KR1nYVIxgxpd/XB742WqbFdogOpqC0VqmmICZqcwIY9vZnF6ZuIelABuifU1FD0lcsSHQgqKoB4X
D5AhVrj/HdUfo1vV9xHZtC5XJpplK/SVwhayfmaWgfnPnXyDNN7zpwBv0ukz88+rEr4KBlkjmnUX
Pm3nZx4Nv+B5SBJOyWnh+rLiIxk2DrVj0GlAdJKc18QQU0upLNk8Loex6+x2FTWVwFd85E+eIoDv
VETjy8FXG2iE5xiI6Tw2vc0RQjQSv5P6HMAJP0ALRg4xFKsZ85DsBi+oJQysQY+Y5slXpLprHQ7c
TPT/mmGSecoj8SmRsKKQVXVcA4o6Si4VfIDbjoI34BljT5Z/SqgIT81uauPFM8jGD37Mh8OJ9WB9
XTlE69iLXT9JPv1s7Lg3bGEpHQtYSNlNi9AyZpzsuLYXvGWz5ItyGIwApvJUw4wX+wF3posYGuPO
vUMLyNkoDnZhZPLHfg9Jj7t08FVVV2iOdvSl84zZVBPEL+AeTUfcXkJbja41/02BK/HMBIR1kv2I
n9Qx+94GWU0y8q09oq5V8DfrpQ6xsq4Rsv5bof7UA2CfPrC7kqRjRindfjvXM9h/yo8my5GFqwA0
xq7rOGqcoi/7p4DSnWDJu47/DUO2YlRA3Gpf6NGqRqv4E/fdrwKzTIof0UuiSEL7b5xxq82oku86
+20HbopAD6Al8X7JGdltElIGPTsUhW+9KrMU7p5YabC7IHwpVzV52X5OvrpF8/X21iMfLI8ifGcS
lyEi/9EL6U/MhkHRyX2LcneQxn2f3465QdWv8YTVOy3kIibTp6enDbUGMxqzqbSxxpfrvK+hMQW4
mNxSWpqP1B5lWE6JgUwyq4b1cmfDvACavwt2xgDEph9fT5ON77Ff2aeE3OccBk2SIsqG+fVpB7/S
NgpOnniHlQ/zQV49BdzTwMbexR7DWPYJIObJVb9winXPKtJhQC00jVmZrghMSK9ynOaCJUE05GTl
e1a9WauPzcROjKqmzkJXYW4iKelZxV6Nnj9d3kVfSBtGPKz4bteoOeK3cp2PDaZXuxCWcwFyhL+n
ZuiNXkV1UAaigy0ooEe1HtKSMCMJwX+FM+0IT2eEdXBAAEBCXqMatw+32HCCX9Pwvyf65TibXiYv
38oTKHvOFeNf8Z3kchFtYyLngagmI3PWjmcRBh70jUUW9X1t8y/1F8lyUou9yHBtXshFHQk5sIUK
GEFi26IdcmxTqRdKQB4WZOi61Yp1MQzExnXMZD3azsdNdQ81/w49Xs7+Dz1+qM8IiDS00Muk77ur
5UzCX89A6ZmD2mqm4emb4L2En2CNnuIjg7xXLdIUGc8fd3cQYC2lY19mjTFen/jgQeWjtDgK2TzQ
OXlUJ065UuQ5DOdEzhkEqecWmECbp2EA8meecQ3YoGDBX/vdv6dHtoxeHmpfX6p0f/B9fmmfooAV
1msTM6xz++/A+OtFAYs5r3bTOL8nB15wOGRgvCJvOO4Jlgd1bxRbpSt0Xt6xdgE3nhXI66Ct9vlk
akiUQU8VFbgBUuDB5YteeEh8UYJMyk/oop0NIYaDJkDB/oemCNMlEly4ek5VZQaA2PTzygPIoSBh
i/kedBECbAUd+poBugigYGkCZ2uPLuSLQtCUCi1azigwze6ng+/YWZpAaJMc63kmwnPpY1WQjreh
+TwbBlS08H3Px4JgyrikY/0BAYesb8njUp/PdujVW5ceK4IOVL/Gq/cAp7ZqJVkyKuutofrbOjPw
xO6XJoGJ1ozMg1SZerEceB8twcZWkXAdSidAhlaMJU1UlSxGxtON0CEg9Slo17m0jXCoOgcLVnTk
omKMWaVrdidL07jizfSDCcV6fIHLyxo3ksMh69Ckh6jwKm8NgRNARYinlyb5FUO5UpZR25Ld87le
+ptGDpPlL+KymR0yhrl37DEOaP9GuyQnQJakWWA80AsUn85PCABtLAhG7k3OTFJ42x08e6ghFQET
acOAjyhrBzMtaTGQW2rKs0fQ64Cdhk8cKlQb5VFjrPIcHKTYBwNx+arzqyBcykFo9pHUg3OmpUpi
l9ikpApEDksIFcfW4vDIxAzrktIkI5sP0fZLYb7gqEzWZP3EpeV1X6BAv6mivrGp5gyWqRopKiFH
gprZKNnjlW/0tU9YELWyw19QnedDdhXtaCv4ePZVfQXqfHtiK08SAYqg3vUp2qdMXHsqKkx7Fxki
TzcnNea6HnobfGjrHsNbEM8nHHRECzIbVfITlA3iNUCLgO2CRiWaEZUHqvIZfX7/PwfzkVrUN/S0
jKUXEZK33wjBecYoRpYQe0HjogMkVmln6ByCkEAaDTibfIJ03INmmBfYcXWaPBPDc5Xas0epN6ws
rJ7gIc/r6y8MqjA+eHPVXDJTPzQ3yMop2fHsJUG0ifngZ3fzNqnjx0a8I7BHBQjo+XrvnnBttGyu
Si/p+cg+Ar9sTCvDGB3As3GE0SrGrTqgRD/MkGZUk0ij88/C3H0h+aSxdQa/HNhlfml8JHD3LNGd
BGjY1bxXNNMSl872eMVP8gK3juJZgoPkoTUEiQkgn/yoMu7fPJDRE1BHJcVUyjfXvKd5oDPd1kHh
XCArWrUQ16UWkPSqTilBhnoIGqfW8/6i5bxr+sosHPJ0eK2PlpBEW7mrMGg6U/sNaogqcvzClp+7
sxBO7ii0IqCqsWE7o73SmkM2fNg4xy8/m2EzZIHeChfjKu/TGGe3tpxo6VTxFb0O0xmPoaynzcsb
pKMlrCHp0/mifFxIgi8+1BYdTPtu3S8Skn0rODLC4rRvo/p3rTkbLqeJl/0vNWxrjLiuiEDF8Iz5
FaJiQ1UYJy9OK5E6lZLEOIYKbciUSgevgOu9GUCDM4sh25HiD25yB9bXK8U5P+3AQEtiUaGsBIud
z+Mdn8Ebwyi5HAgSP4byPP7sr9hGLpkPUDo7Y6vBDO84OtSHio3IGlKO1UpcC6yBLFnM7DLezSFN
ICe58r3ucyUmn3Zm5GNj1KYkd71wpV3ocTQ7CqlKirElrBGHPEn/2D/3KvU66D8WarI+vgFhv4VZ
aaW8qXB5hkXCsy+WxC9+A+B6hXUZJXicu3bsBtCP0BhCGbAhqv/UvMA3Zyf24Aovc/lvzi+XHMns
x8eD2L6tiGunCdPEBEPjNS4AL+QiHXTKhehN+nyRgs0g2CSTBcRmgp2Uoj2rrQkCeK6x7gJfooqL
y1olizt6DtphWpXeGkP5KgxEZX5SYJ6fiqlYOZbfOeWWZ8QQHjlT99WsBi0wX0fsoRLEDTQAFcS2
CT5Gk4afNoJUv8TUC1zaEOZLYioMcAzg6XVklXEATi6OUQBMiiMNPWe9Fd6LDsKpgxYvUVt10jI7
HFNPxPstF4HK9x5kTAxWoOfO2uuZqimSiMyPHbaOFQ6egT2jgtR94RzsTxL/fW7q6GD7eh0gTiWG
dvnKscp0MMpCeI5LkDj/mp/lMZHPiWh3Iy8f2ID5qHSk1mtM7RYX0IonjyDLlqV+bQrRwYem0hGD
8yMCrgG+5EMx3bUBM3W3sABwcGDe7nlFyuSzhrY2Ug3WrbySkg+RhKOtjh6QD1edBPx0g40X+Y+G
GbfBMpd40l9jY1IZXSMBZ+pSIWy7/nPv22UQaApk5iSjT9EoB6akn+gytqDycCtcvMuJBVVxf1qM
U4RIeS/8GOM85SeF+MntvoUzBfdTzmDC2u/4ELCytFhgNeRKow8o6WFmeK2e3pHrMC+AC3pDYQ9D
5HLznDEN+7798x8yKhJ2GcBkwy0dx1Y0z2XgupoqdGnBmbbzcQc7IWsZfFMNHXmH/zhz73uropO9
1XonyO5/PpR177/Z2m2CD0cK8JvQxI2uejrZJ7RQGyfOQiGYsxsb7p7zqnTSW4gwmnKp7zKoM84I
ZToEG42e/kFHV9irfv1EBC9ec3tJ6eWha0pOZaLNF4AaNG/EgAdZYX0VuyvM2L2V4kpMBkNDtuAK
83SvZzBY9MtMeDyr2wD4mNkERPV8QWQ9xZyHbr9rC40Nxu+aMIoF36R+TES75cRzkDhWUrbKejLL
p78YbQX6qmTn0SdLkqMZzm2zKrEk5Ih4/6LOWFGg/nrCZDilU51VrwNnEBumZbsTOPfMUEd/Su5g
re6pGBQU3AnBANWaAixcyPjbKPLmLrWNXH75KGY9WAlsggNl1mZP+RlX7o3rzpDfjqH+XDMrS76F
O+N447wDXbouQTzJDOkEOptwnUYjsSqnbdyKZBOW529yktN1coehqbUNDi8y77x++jt+ru6HoU33
yNy5QoEnDBvdD6KDcGVPZRSvvk7bpdQWZvJfBtio0EfbbE6G70kibe/P9lK1PD+UFhdvXlMRKlmo
G7DFbebbG1hZhQ0KpD9ZiYyfaZ6vF9fxObPaPtiR16wxpMoAbl8RGWTT3TBlDsQyI1+PtjKbq0OR
19QIkeHbYTbs1nAns6hwezyhmHsfwEnJHAGLNwcvfdjQKdlJJKfrhpxYhGfYVdzh5TJ5XE40/m6U
aBHbRa400kAI6p3cVfOU05gfxhsFQc0+NfVtNDdQSdp8K53CViSEd8vNlNwP00RTkehrVlGv+vaf
c4MnAiLEE66ziKls+9tBLQCNCcV/gVeXZRydTPLP1pJDBrJJAwC6F9MiTDhKzdyyxUfWShbwvoTk
x/bqUrsY02d0XJtDwBZ42Zk6HhJnfUt24shzah0zkqlumUvBQVGtcd1qKpV0IVf5uxyDXh3forj1
H+uho4GcmX8dfzxeScl/lbAKLokTgtzswUF2lvN2k6OouYtCSfagXz7uemtK1M5IX2ppD/9AZW45
lGuJqRcvLj0sxGEj8cuq3RAVM7Xoa5guQtuL8egKJtvSNEAotDrL/mGcqrhYm8ORRMn7Obzr5Rpn
FzOeS72KU5sOeTdICwiG6RqjneV2hZXrTok3BUJN0cOcipkyQC4x8WTSz1wVXxoY7HtwbmtDXQ08
vKJny2tO9UXJrvudZEqe1l4tIZt3rRjvDJXy/S5xzUrdW5fRd1IQeCz2u7DYXLh6N4HG7KNSkWvv
A+aU6bEKxctXynrDaKqmanRWplq5gx2TP/wuaW9V5ySmAUNksLkW9HWp02fo5kewNdYW3eS7g0xL
/KDnkorkyNRX8QF489b3lKDcwdLDbxvtk2Fj/QBqaZmleXjsJNN0tKMraQkAlF156r11RQo8Qa91
cdW5lpc8L7gC1Hzsc5Rrzune+23AyVlkvV+4dM2iQf+zmRD2VEOxRMyx1VB8KScH2DZgk1QCJh4J
BIO5SM3dcy8fhFJla5157yAW4QKtpvC8bQxniwNWv3JO6EebOP6yOOSArVIpj7Wi0CTnJVhRDe53
FHP6Dl1ziVRtb2eJASmeQK/PfeS4Oo027c18PQYvcmXuuLFoQf6RT7RMpqycxFTtfSFGvtT8YWy2
n/E6nM/3RKiNiLKTT0+ngNj7lyrGWhnQixB8F1g71GyVitMn1mI956MDcQTanT5zJrsCcGVaHTjJ
3jXc9OdfEoI5I483NS6t4olTgcD5EdC7R/4feO0YbJP85BxFLxj5IqbAYgGx/R6AxXzp6Yq/RgDb
kcYF49WmWhixKu1Qh/zu3jMObsGwqoIzCwDNK6klaKsQzlcdEIoGSTGRRUhnGSHb9iTJpHmdNo4K
wW/5cgpMHe0XnzxCTIkehjqwhZ8XSIJKUNPcEtN97KeusvMKyk8tXGQ4yro92ZhaQGd2SRDXIOTv
gjyR+lkRouQV2NMSsNDijyzkQzz4YHqlQM+9VIhHiIt+PbZxXGmmnabFAQZp3jvLerkCYOkh5cHg
Z48H8VtCUOOu0sDKbYtjrBhwwGAI05cXfdX4t5tzyqHYpoR+jLw11xgRH6w1+BcW2rq3JQzUO8bE
s/29vBvX1ir0tRx8ssgKzi1tS7nlBwkhYno7vsoLUNr889Pt2QRiAKm6q08OxgjHyQn+iw3DTNEO
sQrycnQ6fYzEjpCYduO3yXRKv36kxKLu9StX1KFJjUjDxaLfjVk0v40L1gRrx1fATJYe9DRXyOBe
DLUuossSqVIuI1PMrjwM2ciJkvDCMja9Ss2w+PCrqEcbCPHv2H4fd5zWH6VbZjUlfqTkv/ytHV4y
Bgi1E3DS6BhnQ/VjsA5ozOxxLPoAzbnScTqg95Hh//ZC6CqYgUYsI0AMTUO86RbnCYNazto9Og2C
Mh9exrxQ1sF86wpY1O4rr1YL65xm5HUmmqwAsfSObwVXaAig6Cutq+ndssvLh3IRKL93PJ2fruBP
UvG1JRHtI6ayflkq2UPqUlf28tB2kSW4h2ScS1gdWAxwToYVteooVIJYr60/1KXq86Nsp5YoTg7D
kXXXJMPUWTCoRhlzNJMWmRsyOWmcO+KLX/nEM4Xmj7h+hGZ8caRFGzFIQcqPkKE1iYH1yGKKDM4b
myvr0FuJo6v9Ue/4HDTgInFb+FwFUDkr/DfnmpqgBnjIh7f4xOsB51Tk8xToNk2awepbDmItM6Z6
d88vLsKIOIcW5lsY2ATqNx7LLRFJqEZPkRaqb5cDnQrO2jsMAJLw57q/uWZvTK4K/xkEp3ulZHH6
/3U6dJdXuEZx+pBuBDxuSMA+XukZT4+7b+pA6Z+0p97Pk1IHUHWUKd3AxbAtTFm5Uloe7og962z8
80Jr+kJX5j1Abf6IHywvhC8RY38Q9CBTel4evEBSYVIpgfpEILCj2MKf9A3MAKipVd+oT5sDTjkw
mcIDi3mi+rSuBLOFi4vz6YSOsTcCyEWuVoQTzR0OLi7Y1gMI9bmgPdPOWvJtK0MafpZoOiuyBkiJ
ShAd2rJ1jyeNFaDhUak67y16yBEmL5XRiIuREp3ocxaZGa1GU+zDD07WZklWOp+41blOV0hPG/6Y
S0uzIqJBKfHf9oazdzL1NrMrsP1+UwcX1v83rigL0Wug+cIWTDBrUmIoyck/kmD8f2Y9TroCPH/P
vLR/LjKqVmbL1CsClq6uc1xOO4vi7NhoM3MnWxdMRUR7ofYg0hrvG1ea0f+4hmKOOogspd1NpbR9
S6SlOD3+JR6M0ZgZJeEKNhETmgFZwOAwyxGnvbuHtatZro2aB7Y8QJ5tASWdBVKYw9aBWI/5LPlw
fjPQ6fe3cAS8LiNToZ6yBvr/+YwLneApWKGAQDAT1ZrjIljio3yDxSBhpZNGjUK/WlkCCE1vkTY7
v1RYMINZAmfmH/nAgPJ1q/v9LydlWLszXtRtzGR1gF6a275/9KZTb/foonHCxWfgN4adAK0b0Q/J
iFvCII1mYKc9yYZZVf8pBwE92WV2ZOsiUNBEZp7oC9eeBj3ov3lA/2O9BzQqKNzSltEN5c+amz9m
8P30SH2vRXNqysP0EEmQV6+DBCb2vgwQ/36G2HkYRfZtoPzDXAmkiuBHB4jVkksCEJUNzkhiet3V
rmcJFOP9b78bW41I3N08tEAKLEvnAhmsBoY7eWbxXElXkhbprQkzKGOs85+t2Awgl8NvpLkD5tW5
5otz2rUlJzpMZxkBlKGsj5b98FnTCP3owonpyIWSQD+uWwrK1c5TG2VpDxn1Inq7uUhhHgDJRErA
jxc46w+AqPsFQrWwJXD8++y6/pLfg419MMNoI1TNhHXTYLx9aU12tmom3sgBbRMdt4CuiI3LxGDF
t7EwTTTwWdPKpuBS0+cRn+QkGaLs5TTFZFgpCKCUzd9H+g9JYbKqb0k4w3r3Idj7WjoxHRSDtQek
Whthpgufb9aBgKT7GTMmDUWRXIYYJVwtdK8+FwQ5HvJrvKivlgKOq2gmZMsXF4Y8IQWVh0Ae26y1
YoQ5TVQYZBtektF3iT2EsgbDDasJBAdk2rBLp8IJovtR4YcVqtkgzKH7EGNunNcDNfc7cD3ngcHW
vAr69uR5F1Hg+T3xOVN0Ad4rGG5K+GsRCTehR09rtyc1KeJQ/6klJDIrnEVtukIC8ZZ1ix7/jZ5Q
3qzYjLEKEH9KXDTDIjmTzKxumhyfcU/DiwH0Mr+j4pH/RpLErTAcYDAWajO+hekojFqCL0954qtR
ZkIcf5UuHoGzq4f8jQRk+MKe+hOVOX17n3R9XECQ0Ih7a79Il/gg/cXhw2uJya9XIgOqWrsEgo+o
Ogzf7msl3C+Jj10WW4IU4lcokGjpFCL1o9GmGsEQzQsc66ICebt46mROBmld0RYL6sm9CL9AGOzv
LyZhtBsbNM7l3/Isuu1u7Kql+dumI6370kfICCZpT9p/Oi2k2aBojH99AS5xqsm4BhghdrGPQ9FU
L9OlsemPDZZ8wjekjz32UEAIPi0VeK6mq/xVAs9idx0B9f82gbLH25JAiwo7W4KwHqYg0dP2shQz
AJyUVS+oDrbj1KiveCBGCXtHik9d/ajINRuN4ORNtes4noyumbNv2XaA9Yc5FvUCY5XpN4z7ZdRD
4DJH2UrpgmNjFWgnnS9wsJNNPpipVYwKLyTUoPgTN8Bqk+cVfUgdI+IMi0Sn6Bj0kOuVfDpVghUs
/Guq/ZgAbZkeBBrglWVLXCJlnJFDUVL/83QlYa4D2NqMV+Ub+E6z64JKhNCCaqav8gmljo8Lu8hD
SdhD6RWXWLeLiZSCji+iHSqvp+da9w77rjA5Ics+zfg68yaibHkHIK3aRow3M1XJJlr1IEbPRWVj
K173s0wyNIFNKdDdN1Ymrb5ohscwTSdCwOkbq2Ep9vuwRSNhqP7IxG4a2SHZ0utRxIY3NxRlB4PY
OD+kpHKYhcQeIw2xQg1ta8NVO5MYu/YASoUWMl0Vg0AZQ+DN2PQ+z2feSUrA1HavPxGM+y65zVZI
TRWMEjsKV4qr9/U2xT8crGYtpV/YaKF0BMy1bFgH4MFoW+/vj15nX03cKEfjZP1XwJGtzE9q8vw1
xJR8iTqBLRaSzbtv1q6d3GowsptJZeYeechb5g0KIjU4+5GobYho0ERrOPUnO6mtng9rJRMNmQv1
2Ua1sKDN5kbchuMlkrQ8lNoo5zyAY44ubGY8BSbDiRrWmFSq/qjlLcqORgfFCCBZJ1MKi8wYQkAg
hWWhM9TDDYqH9alzGYHtj8sbCsD6ikQizj2+vLtpksKRzu1N/KG9n7nd/tP8k8VX97jrPM0o+Cdu
Dqa6LuSbQ8IdOqXznkkYsPQHrVmNg/P8fTpRadCXTJBNog55rjNqtPqwBDjkYZ+x9g0tyCQABF6I
fzomjQbnFKi6iwdFcCeGOldjYp4nEgQlqfUfgdzXnOBnzeh/Zqn7Y3D8cGsbOLz64X7nqO7rYs6J
COCYJ8LfTKSoO+hz9xAFWV0P/WDn13MnpP/OEutD7Gp7ZHzDi7CSY9YAg5KdXKrnAtIKgkiJI8nz
SSBcpVqumKBEOc9EJb8BRKm8tUdskVScsh/mwgK5yiIgfdItCpMHubdx2Ug7EMvldJI/JYwh38dy
a2OVAVC0XrMiV7xGRpzmV36VBTnowtTz53ZsED2SSRdzouqT5UpaSzJt5BPi8Rw+5bS1T2et4AoH
hVixqf4AkCApJ7+yrgFltTHutfxRinRr+A8uUVUPGlPdS/BSLfgqgueBj6zZFuaARtgGXTz20Msn
zUu83KUh/JiaXIpTy4HbB705XJjNGmYnLIREJ5p/acZTOu3bEJ70YZ3dlgq/idf5rvRSww+0ZK9X
IOtixAEUBx+jJ0ZX8U0nbv1PwWdOB7I4Gv5sLaW/GbkwXH4Yp8R2w0UcQ/Ma+mWn2QYAwVfeDWCo
HM3+jgJiEjXBjT/ufyVR1CIf01E7Yc85oLzcZYzuU65SxeFPVO2KQjBe0V6J/uGG1bIjklTz+DaY
f/1t5bub1wwublo6/fJBFyDeAg8T0Zq2B2uv+Iuy6Rsx3iP6/pHMvrPueRCk/08W9zFXuqBRo1Tv
zLxlIL1Yij2Zj2Ug1yeQuRZs2rM3Y3WX7J4M19izsDyBmlEmKSr5+3CXhDfMA5Ut3syc85DBIZlU
zrjVf8fqWd0TzpC94X8+H/YgHrFobODkTAMYvHKppeRIwI2KlnLpJ6G+PomAVodVCgmAKc6edM9X
Z5OXNYMIuwOliRH9gLAJvVol3A+vIz5McVBHTtwSlARcZQfkVMKSlbjISHcHBbbvmMdcA+GQ2IyF
60wAlF3SFpRVFlvrqZ69OxfSPYEMCdAC6gEOAFlWbz0yI+aZb8D6G10wq+q1UHjK2PEDeWl0MUMf
3/i+gV3lKrGzLVRhpCMakGQfj4tG95OehrYW+n6R57J4vah36e3JvD0XX7cmnIuIpY+HPP8AO9HP
+2guw2RxUK3rbEjVTiC3y/zNuZfqbfkrvHd3H5OSe+A39RIV98qZcO5WCdOw+pYjDcHQSFkSr4cl
QqRFMtp6bXzX9wP6m9s3KNgNcckwxm1VhWYohA/HIlaJoRYo9WqmE/hItqPb9JHMgk5niZH6eMy5
+caDY6bCTfR9hcI6/UYGw2ihyu5LGW8ozzwfVLsEgzUNO5oWGHUIN1C7EBAkWr5C8dOM0o8QlJlc
OGvLFj5WMzSO58pjWpRvi5kt1e8E+nY9IEO9JMRFGr8oUUvj8FXxUM5lS3GIKS2ImpWUx+LdyxZO
aeRhZDiU8O3sr9ciFaGakmesC5KswoPN/6+oqoiZb7nx7Ore9XBVGRLZrPT9m/t9B+EcjyV/YBvA
RgJrDPQ9ipn+Waz03frpejj75Kf0f9GWUUlgGaYTWKpP7s+28AwIaAW7p4tUjTlVKOPY8LsQz0fS
7fmyk96cRY2EGe4NwMTV7SPsaKuENbM3eSmJsjJ9qqFj7LuInKl9XlJWBL4+cK8aG+9dohW7ZRFt
paTjWvc1pZVKXs50L7RYUIpsYFx5qFICx8gCeeTIG82J67ly5O/vxHS/pc9zlAfAzWD2h0Gy2ffh
s7dYKDbj5rTsBs20wbL3a5ItH64xniyLQ+IMeNiE9fa3qpbvWiO+6ta71CKvqFPbmcGqnuBsOsqx
9/ELtR40JWejaYrQ/W/OF2E+5Od9ZCQZtwsQkFshnQejpIHbl7dMIuc4ltNzIJwFVDYLkAZtykfL
QRW0f8TFwvCHtTIQ606lx4BVo0OH/zCdrbbK1Jp+R+9QFg5pOyIz++xqvHLh+xeyokuYkMX6EQx0
bhnbFa41EFNYlq6aRx8GjuZQaTyq3hqI+ydLqS+ktm9H4i4Wg09J59gOiOOBpFZ6/CYzs8dwDfR7
IKpYqu0gFCp2pLIoJiyQHKaThUoFwImVRPCW4V6ii57Ztn/Sy8TL6AA5jOnSs3ovmYRuU7yJpLh8
GCE1sehtOkf2tbdLV5CG1o6W28VyzDEVCFRwX4sWrHyTFLV1atb2umWn5K9t3TtzvOlv7PMzh6UD
6IT2esNGRyijgzXPU3xL9wiBoeFbDs/9xUfc5Fp2muXsPa5W5IuyMdRamZZYGRixkEJfakR0uF0B
vstNUGcJhyCK/B49+iyphSMVZKTH82IQWPECrNK3d9Ui68EYoN1utdZtqjTnjEajgfNDTh5NMzQN
eBR35No7TGxBtMYVyisl/EMcOaf4BsB420IQ6DY2OMhbXOi0DD18WzedM9X06vDZvxQbFUJqoO7j
kwkTF/ZwUoZGxhXURLLa5Dn7lUErV5zPWTF/d4+jmNmH8NLNw262R7yYCgXkfU+7V3KJVoO+9+US
AnTK1ac01pjuDIz4hncizhNfC8wnThDVmYjWrETPLcltx1yi5OYz4Km4Dngv60XewMt0l94JQyNh
uPyTllKHYGMqonv7+rjtgLJkd5iKgZTzldBhRULAxDLhVt92XT5husHFeEmz7lNHx9jVp9xNTzKk
VA18VO7nX12HVeYymtNDQ3AfzNZN6M0FeYpMOm2eNH1fhlTyZxVf+l4Zah+i2RkFyeZc7aCb6Z9l
30l/u6LcK8ZBG25/5GHRLTRjhS+8Orn0tz3fMixbh8P5bxY8Mkkm5UkeViA/K7VEff8rXZ2Ldvcl
QjO+4MoiPhY8MDZolyUEykR8OihCp4UsMKzuvNR1s+r9UFWzTBG+0Cn5Ztz/qz2JU10MYnmUIXzY
JpAMoLtbnYeCxZNGjQaFeJqa8M/8VcxbcFEh8O9FcjjQf5rGSyedfSI4TJoTQzsrqG/kTL+p+3KA
wQH8s9VzoBELQdiVbT0RqfWZOUpriuqma4s5hhMY1TUF7EUjoFnNAu5sC74zL4voJsyEMvRkHYKd
eCWYKlrzjtRlIKbVk/rbWgi9/65/yhsPZ5tE0HCflHA9eOyQ4OJlw1+w0EC8PjT4seT/FTxN4USn
GGoo9gYuH4WjvuaLLbrtDYokw9ILLHTF+focAwhLn/X9/+nzqgioh0UNmcx7vdvr4/A+o1DzgJGX
sGZqqoLfGEoNshQfHojAMljKqAU5o9ElYuiP4yc+CQlg4B0EVLkuKwpcEuEkIlfd4alhtemquFnk
F65wBz/54Eh04YN3EXlTKuy/REnPHhvd26B2g079trHFN38PfSn7tvVLOMbVaJVpfmJ/7OGRpN63
TgpK7xdbpl1dvIkb7IcvyEQnraZacA5SIns8DM+glQA/Jkx8d6eNLgU8Ia6XpvpMUGxx0vpGl2gj
oz+V3pqMD4rnxhPE15Y74oOyb6Tfhr4YgnlJ0wC1xYBNJOJKgRmf2wo7tFBcwBsbqudoAapWv6og
tIYjYFEQKcKtLicjxxjgpQJKFtv3tRf+ceCUFFcYaEJfHHDhRikCSepzIhLFQbmz7pUXpcNa5NT5
C6AQ5t9zxGEqhpr14wdpcBi073VosTPCsKuXbX8KAP/Ph/tgdGqFneF/dOjZwnRQnqWq9RVLciGE
BBvUti8tcED1ehBuT/FQ6CP+53k0qPcAR/eeiOlmzMyZAh0VkSLAvoa3F8DKnqtr1ZzUS0rdYkmD
KZmZmdlwNl46xVlMEskWT66ZJmVxA0Mt5ua5KMhL9++rnLGuL+Ar2Vg7PiSqnhGbJvfnuhztBbbk
QBgiRWqc1YGuPWdMhclHx84na5OxOGr4IvEfubvyOFlNLme321uNSCYiudOTk4Xo9rbMVkOxoGJs
bMKAYrttXY4o8emc0++w1HXgpPufXs+R3Cm5q9gK9tjjG8WZ/egJH7iZye0l2aAjrAnV1ZBibt+f
r64+c3aSaimC1NsO5lqZaqim3HjPSCwd4l9t6zaxrFLSdtKOCbrx6fPtpmoIo4+IzEz8/Y9/K16u
OoOnLX6NMcLdV6muLlvXC8Ju/9gsB0KtHXFKIn8H1yQe67rE8+mQeSmwMZhgGIDUDp3bj6VKr5SS
Lts6WoHaV/msWdtCW2HEEyvOiXkyI3Db8UKdpPZ3qncNpGGVClgfhhsuMsIF6J30ncBIoPnNhOAa
HgeD4dXBk6Ci1lbUuYP4STmxSzeYWVXjmzJ3kbzdqgDJuY/Hazjz7HOeqJ5jyDdQpzwtQJDHFJet
PrDWUO+eFa+8lIFm2o4w3VOhqnZF7XjBEYyQ/UKxByckdu02rFLGObIacKjl+MCu4p+5KV6K+Inm
ex5CrFJNApP/VP2y3hpZyPqAP44ryhBvIalBuGtS5MORqquNRFyukMjbeTmWZAQbLWuNrNrDMDOe
CZqlyXjl5mb33Pxksa9JavQAVdiHCbdyJexpf/hV6UWRS4IBKqH8GRuQZ7jOlVULilSRUib8nq+3
80kjLKQh6j7hwqycaIQXC3AIytNT+g0JVCWgikc2oi+tV+JzZLXttuyHsgdQ5wnTqoSsK9rKBLGY
7yb0cuIUx3d6P9jI5ziAgWm15LGlhQ6LgOAXrrTQApkb5imqr+DqCFEYOvlYZhHvXo1HDW4xmOGz
H+asD1Umzt3N5PLwD1TomIZOAzDoU0a0HcGCesNKR/JNcOnZli7fPdqNrX3bs4gXyicomJIOm0NY
Bceyd8Ho5O7co7sayHMVuT+6YDEhr84qWypP3qAoPb9pBdyHryaAyjikepx0l0Tdu87FuN/CVfF+
FxPf+sZd9ko5D5egzD6hQCPRQ1cwCW4dtbbf0+MVdsQJG7R5xZIybbavSArh78+AHeWHz5htraD9
MXr/pYx8mxU2JSIRLAtHG2CWjbk5eOxJWRmUbxWRVlAKo6fZ3TiD9huJBn3Rd8GgPzngjjBh/IiZ
QL/PE4Jv6PYMI4cTEhCD2BfDB/z2xa6FAynlX4eB8SxH3Az+ERbJzdWsX7A2YSrI++36GgMAJEFh
RsYu/AItJWvfcRVjnhsUAYLnNjxWeOcvVmvpPbZ/xQAzS8ncry8GCeER/a9onLgDo/7p7F8HVjyf
2U4MI42BRJSArn0PKwdpoBfCNVPpJ/7g4+uvAAd5lXyXtFwu9SHyOM8ED+DHDwp+74dlkr1DeK3S
xkv1bBsx+49zzdfy7HiPaOrl/o8lUpCXtCfVOybojKpH7wFDk7fTIw7Wfe8v7OaVjbukKshJLETj
U+T8uShsb/I82oDIFsO0vmtGzsXTV2GR+6FvR2g0OMkwM2J5gEj5sHYJlJuF/nHfu2zN8hlX5SUJ
T7q2E/PcAPi9pBQh9fNVMhVmjnMnDtA4rdvyXTSFNOv33Zp7mTJyJowVjtRSAW21EMCtZvCrKO79
yzY0Zio4gXR+608FaraZ5iH/8sbBj3dkYlsUFvGw3r7TQ5s63CjecrCvDCbN0WqinU1Q3EcLLnfv
GDfIT4FrtzlfUzxIMZdSUKT6f1ixlvUSvepZFeWQJV63w1Jz7OqZiu14hzoV2ogn4/asgfTZ6DIk
I4T0qn2vonk7xM5C65vZ6wcKzsMw5p3InwkAprXfCipqRD0oUgW7/wY3wIbpoSkg4DHkfQfXMK4+
BZsrGCDLgMe9UHOLxWnlwxdOENFZ5hZMOOiVzj5XDWo6fnby+Vkkl0+t4sqxQvUaKy8lV7HBxkUL
wYuDNhdcoWg39ok3DHYnRjNOafBSUawhluYODCXOHcygtDF0YRNmYWg8bZQ9KBR+VgQzzcn4ltKa
LunFev9iNZ3z/SkJR7Q42uvQju6FxfBWH8twnjl/JEfI0+fJqRnz9jjLE2QT61TQtW5027NZ08Hc
xgg35lFVdGXCpK9qc3hJHyIURjrjRlrSShFMlXsuvzV6ELovxOk+qlBok3ViDJdCYV5FcxcEmcjL
iktggivIfUOGCk0VjWVGsgrOy3ih328yYgm/1G8MeTMw81ncRXU2lSdt4MvuzyyohVWEQVcBLD4t
1CJ7ChLjD+9VjSNB/6Noekza2t3hgeLxvFkGpjoKYc/Zq70hI21170ZcQM2R/FrJiv6NcI9Rfd6S
dwc/4BAjWjDj/SwfzDi0Qtb/MNN1ZKpS7Mn65OHeUljUnPxgAKl3gfVJSUxiAT1B0pYBDuG3egtz
TOtrh3F4GVwO0MKtKDdAgsiOYrYrura85/XyJALrc94yWJzNqYmdSD6Kw+eYL0NIq8hoCI1p7jfy
3KxcupHjkb+5m/tacxjGJ5MIsPlY7KSb+OUfqqN1MxxtlCrC/XINbEC5LD6G9pt6ScZ9bLDVl5Xc
khs1/hlYLiacX0EjkwYEsYOG8XadzUsZF8GKdMoKIWDwHnrIyZxp1J5OglMFSH8Q+gvmPVcxB1Hn
VMYGwvvImRDMbvQSwFWFiGCwhctiwShsRNskLnGDtCTPQQv/e3cqdk8mPtB0ro67zILW6IDu0Yos
2ht4Z7y8awiRL7IOOOivOJM9eGc9XghMRqJvf9Tdqib+mv8dSHWgJKbGS62vHOo3idZyXx+tOBM4
hFMMOkl/+cNkeEl/1YWHuJ+g2HQTYdlO5SW4EPohJAPkx3wl0GmDA9RXXRh30FMZZr5ElUIttCCm
vLaCGJRhTEho+XCBpG0CZNRykJL23sL8hiLZns8Wn7aEMaPfsYQqLRln9re9bw8KmIXhF8zFQWR2
uAGN22duwbUVsIhBelY6h/pmDgXtbHTFZR65NTyyyMGO9fy74I4MjUIhCWkUA0SNTfJrRWh1LK/P
ltwTNxgYbvt2VQw6JwHOi44SkwOBboE2TVaELPay05DHSBKm8i04T1xWDiSPi96gSN8fCR2iZxTd
gWOY22N8u3tkoKqMlgTPfOzosmdapQwBAFg2pZ1cX38riD/N+TYP6gZgH0Fd+ajkiroVgk+HsAw6
p8VWzyVeC/wo1n+fa2pho9aXI+m+NaCxVNVtWgm/7Tc0oFxkio9qfJpmrFNorry4aiLjngnd5Ceu
afBferuAaBh+dTArfEW55qdB/JTjKkJBrUIwcbgHoxW8Km+lcurxvYNy2to+lT8C5+vHNvQpVk1k
9KQt+a4oFIqcFyuOj641IQzHxq1ghEGysA47bTOxbwvSjwawYgGp8utgAlZMKGF+aDjHVCBnfmvw
a3z3OHj0e1VvW5+Tb0uIWlyPCb+S800RlddH2Fr1sRYceJtfrYyEGmtpGYCMY3ZYiyMo5qHjQn3z
/ckpm9cFhPj7RpA/9SMCzy/jb4cee0cZ38FPU5hPLukf+djwyOTpaK9fnxJ25PoplN4TQuUGjSOx
+y+Arm3+396v0/CsldXyins1GbEbIyWBQ1Y7Qb/m59qJ0k+0Q7mH/LWqwrCf5z0eNQmJonDryqIv
OuGtHyk3W1vzPT6kwwckpqMuJDuERCtA7nHVdRQH4MEBkYAXKJpeUFn8awPfiws1DE+Pa3KBgLPx
8KUHL15CWilTnJP/NW8p2YJeiWSUUyZoVzd5hLr4iQYHP7t/fABR/rnFmFeupU7Yg8IV0pi0zdT+
CLHhC/59Ut0O9UaAcv8TilcIOG7zn0jEMfs/U8gBa5jGu7y+WE7sP8liTbY8/spcYKnEw1BUEv3K
QPLsUDYSxxuWZc4J8m86AvPZLJJAGlBAXldtF/TvZsCJB9ta4/DFWZ/CSI8YStfUErPFDKQWSI5e
pqP3OXwHNIOcXc3jlC+OuwSGdJz9wGzP7KQONXfeN0meYGvQ/8Z1IpbNtyGzOpmSzL1j3nb8pIyb
NAHzrwXx4YUYH79PsuLxgQZ0Is5OuAZdRULv32g9JFlGkdRucc4KSXfXjb8cyhk/VuZCyewpkrqF
GrEo4GSmDEamxIyL982K4RG0OnT/IRXP0FX18nhcejDgvFkBNOaXW0L7ETYIta0UoJ/9wiPzj70o
Vn6BxBzsl4wAoQrYRIPkxHDwBBDFqCF3DTaITEFN3/JnCIzfXgaoDj12Rv67Lsp8UK4gxaddmHd4
JAkz1LRhqmk3E/nCIw9sYFUE1q7S/5HleB7k1EV5/zeJOfrNKKtrPFXOqzH0polgcHe3S/F5n5jm
lST3NRpeqexlQkp412jCc0a3b5quG5mdShYpcW3dFVLuui4clqJJw+GHE2m3LfPSZdAzs+vbz9oh
JTLakg0JsgYTKqMaGdAQFX9HElxlVFI0b5L647ko7TAY7M2uTix3ebNJoyJK8cwTBL1nUk0QRwjN
CCV3ivhlDAxOBfQnH+91BaC8ZHlUMdr5ig60Gi8+s1HsBjUlm1uGRIkgqvxLaUuL4SoVHU1ZvOja
gj/17g9fKyRXVJujXAm4IJjrCglsJAPz0UD8EfO5D0vMBxnOklcqE09Yk4svNeroAr3j9HhYpcI3
hVC4LRh7qX/dlaNsJ4/HXUUJH9yiGfLlUBh+dIMpI7lzavsjKT5Io1CBaYWTy12eiBUxd4Jp02oq
ompCGz30ocw2hu68Uu0NDX0Ewt15uO+YSzEpQohsgO72MjfsrZ7/H+Nv9o9walUS4H8GYkS2zJ0y
b056funyHwiNn3VncrZcQi/XQ34NSKUw9G4GcXMm0QrUPpbatsnJvnzCGodwCfWqALJC1qVKH8YU
7jlhKXKo8u8pBFrUbFhWp7VdMctpLLh+AtkOgne4aixaWe+NFTUO2DxWxyy0+sScN54IRTFxpRd3
71n5fb5P2Mh2oWmEGLHqvZpGmHzoDC9kSRA10xNwCiLHyldcxfp5ERw4h24zWT0gYrf7IFH9IOy/
fH6M+2u21Hj/jDZHKTnXPXZM5pUocStdTT9Mg4zvUjOTyicOWLvDTs7RAfzNrDF6XPzWpGuWSA7a
CZ++cYOnVBA5BLDwgdCryLTZM358vGVJ27wo/4rmwBz5q9e6O0U3dtgm+YwlW9b6QKVnwZWVlbMP
4sYIku/vFVptNrvGDta6eEMMOZU+kIUZ6runAzE2JbNyFWnJou9jueUBc56JdIBSE7ZfgbKgeMxD
Nqi9AY/3wdRANyZlkZNvdGNen8ky766ksug9YcYYn+IQASJw8Ng1XAOJ1cBAphyly1ozNHEJRsOz
rR2z6v2icJad6pZwbzwxeufai9+WPn9Cya4E5KMiLBnKUvPiQiWc7fIvZntyVsFkisCDYScFCV9W
pm75szjFQGeMCi1y4NSIM1VegCQM2G+9AuvgOWTVGEeTYidm7gShIC3ZcSpBh2Ly3gt6xF1pflaD
Ltr1R2Dv3YIaWHF+rV8xZnpco8Sqf1UEpwmBswgWJQfTMgC4bokLAgMZE5Hw6/+Jy2Q9YBrRfsIX
5phDT2khuDaj08NTxBzx2ckE2pOZCNaLpKmOy9F3d3s34qbKM+wpLKdk7B0nGqPI5nRe8+stC1CO
IeU30bAdrQ+FY4BPe2eC38QCysx54xtIx8ehOyQytM705cy3vRMjYnQiZrfuFfAKCHn79OpYedLP
MhzsjVVlV1CHzmceWTwMQNJ0TDQAqL3FXgCQPmePcQfo35EFl1dInk9RVTgfbC1WPYLL383gQWDP
AKIQhAwU9ZmNMPyw5HschoYV8O7/hQd39CyS75BzoI7+MHaGCDl4ULfe4HKbLrAkHnb3JDy630eI
srfu9Qjvx92piXEIm882c3MpgGAAgGg3IEr2sg2lAfFFTSH3PO9B0ef6/VxwuY3IGGVSVvAR1HGr
UHy92Rut5dH7MnDOORUZ+fCiIx3RPCDKP1IeXRiXf3+4fdVm/UduWAWieeojscJe8+qBhQNmrypy
j9G+Lqi3M7ttQUFzuyT0S+lI5IlWbCzs/FScwZxmE99MAThvsLt8wVbtNawMCSut9UgEwiqvXZXS
3jDLE0WHK8JouZ7B7ddnL0YBDZTUk7sVbDTZhGcUZsTOqfOFy/qpCyBY5HN/LdD/1WRaIIm6vml1
8Wm7BDwu1sDPcFPRRLWOiszkePS48dMOec4C01xAZOZ0dkZfmQDprFzjM42b7yQmXfNjsEYNS263
Bawi6nCEEhBKQhg9XJGzY/BjAD+ephhB+7tPlT3gGmWl4xVBjTJOoHtwEtRXd0jPG7l8AKKIkVsZ
Wm1n7K6dTQETY5U6u9LlfikDG+UVahEns9+qkManjmMPuGygI/UHznLufHfb+Om3OmcrNlvU7Tj9
X90YHuOw9sVS4F7+6TZ4ZJyjy9w7bgtx+AcWR2pArcT7HfU8EigHqP8d1L7nSrfNU9L9rXMj28FN
bZieql/XsoT4hFw7ZpwOuWqj/sQx1mT9WYZ1dZCz41yvZmVsQ1h81rc/9xArnfnIam1q4JPP5Mgz
j9mlPQBsBxYCjcNqQE6xbY05fzZC7OpmHBQE+vsSp8aExGFLJxvmCEnfLR3XkOEErIBZEXIez9Iu
md41yPpYmczB+1P9LOxUAsPYiXyLVXgIuTWWUqYqJmJ8OkgAAlSOwXapwujl07F6DTv8Mnbt8rMA
fqpHyt1qxpukfb+Uxj7TuWWgq7sJWsbVS4jQ5vXSKvccXRNATrvQVQsX6OZkP6XLEoC9esQA64nz
DJ3DAXec0J8odOdrzwyKjiExIvxouLGy9NmmEOWk7cczPEWbZvFI6djZdkgGHjVGxzIkUpH0PV78
h7UOfmhKECB25Iz+YwL2XCQ9IoIlkN/YanJubTvKZWvQsSFTCDXsn+yJ+/ca9m+/wubXaaI5j7Pe
2tKCdnggxbHDCMu/CIo26lldnsgaOs+vLNwfdSlF63HI7buDxAubTDLh+nFUsDu7Czik0ly2dgzD
X/Mq9V7VgvAWT5Y/KZwOHQnMLwfnXRP8luF+OFzG+gzDrjon5LnBcf4XYpW8pSX8FIJGIrnJYMUj
I388Mjuy4YYFIfcigWvgCNBQbN9F/1sCfTJ+VNKhbJ0KowvO34U8Hspp8jp42l5MCbhOGldqoaPu
BwUKBpxV3LJPQepfo8TzlCitDMNiIdN9LE82IZJg43An8HH1WgBZoVNVp+qMlJIarh6wjznbnraY
n7QybJMksfIAApmuKc8rQ/c7o5sfZou2mX0SuKW2pVu5h89pHqMNu/r+P1iDQM0daOJNFZOtBXnL
yw5xUXcznXXV9jObNfnAQrQ9HOZPZYulZAN89KV5YvPmexAmOCRw/8UISKDmRlSH3fU3YIc3p2sF
2C5wjRZTdBbWBgMyTvKCOIaUpBTVtdavGPSeXx0lNoEHBpRbZSaWL+mogjxOp9ZzP0A4ZCk8S0aF
QkTswULYOaQ3ELIOwuJNWstXFjqNOdtnHjvDaT7ixEeJSLhOxeGsVwCPaeveE7QiFcHl50pgU1c6
Mr0e9mih1cNnGqzq/sdJm/0B3oMbeFHD5AHGf84ZWbGlxWaPi0FOdJ2tFdQ21aVkAOb9u256t8Wr
cUtWNADKmrCiQcCk04SK5TJhMLhdHaAj6Ani34MRVEWJcQO7dwpj9mSTphVWa4DK4TrKbQ6TZSvN
kRMvMyvH3Jgby/SbIg8sjTwzw9ft4p7FZpAi2qZEyGn1JiveAcBEXIZtf41MIK3ttEFV9b3mlcoP
6dhRybQJBQQPt30y5sAPGgoQbM2QjtwdQUUfPCq+qlw5D/AnMzaiUK1AEYLwhOMa6YmehwFbYqBm
Zighrd04WPFkaKkL3JW1ImD/+yQhhGqlqia28et8nq01Vzudk58Ix9O4Bd52YavyhDLsxFahTppT
0lR3FfNgYR79Bj7HIPMnTW3YtGtf4xU7ezjA7thZO4VwgyEP9+IxTFvuVUDT8u1bPsiD25EJidz0
pcNsGI3apr7zPB264L2bbWCiOk8gjkhV/ccNCmwnqvBHSQk5/7uuvN90TZS7JMAl/eB9oQhAxyN0
6AXWMtOuY90ZTgD6i+YDJITIeP1hxpEijg5M+/uek1BN+y2epyx7IjVnqnYbeE4WeXF+3eNWk4II
XsOEStJ9cFQebL31EWRBj19XEcvY0yfwcUygq3L9s6mLL2aR4J76R8gyxHbtyyXk2DKCJqiKhTHj
SrwMZoax9YOSXNOMFzdILM35udQMG2iPoKLjI7DzBgsW3eLSgHkKO03cEANdi+sDGLvVMXD+Y1pP
sg8qfEKsSv+it3YucuOz0CRdAKnDl6UP+O2fIZ0y4TJEgdZ/xTycaNrVmSK74wq5yegwCC0LJM6e
OnN+7zNWFDBLN4vKBYWZo74YPzqb3QXSMFm1OR9J2Z+jQkWZwdylRLz1fN+5i9807hoUxsD+3OXg
IKaKyJXP2CzZTHEPInI+MM7cP2pHzPZi/7lvWVV+EyAft1O/vB2loK860SGW1Ku63WidZ63RrUm4
URWO9C7Lf0cHrAXwdDb5fGJkTYnD0M88KBRGnBKgBqZuizXe3C50llftjh0hbyiD/+KisyGtmanb
DQaBOzKZR8t6hKcTU5qtfUOa6T3i7vbnRFB5DPEJCylvvK4+qI6LI9g9vjQZjgTA2zY7k9Sa8rik
lC1W/mbLNTRSo/5GA2n0ciACGy4ATVGadgGvb7aXmVZ3GbFkGE/Gu9woR05PuudAxp5Z5h8/COKv
CQgYfjJET4gerIHVEVHj/WrI52s7gGAIYh2MMkwBvvGcUUQefVu3zRajS59W01NlI51VScmllZpY
ZShJZ7AoBPccUfTn4XYq43F7VdE1ozQLkHdDLC1T2/AreJEDgvJ05AETQhp1k4HrAkUeNxHgF7od
T8jKcV+uTU6bhI3etmyJEK9fzl+h7Ip5lOYJwd5PQvEWuxTh0PwpaL/ewshoKhVh6aAzM+ZZFIjb
1mk3CtE47sq/RHYOUoo3c4v+vM7DcNXMl6uUXy6ZUsonqFh8A38510WVBO28cPijL7r64g9MuTfk
mlU61Y7zrA9fXhB3MsLf+QYBPADJVd8h6zF7TAX8S0galvzX2eL0Hn/GT/IU6Xy2DWgqt4lsjHAF
kMNwk5OZ5qCZuiMSLhx+++1yVzQS3Qn1MfBtUsaY1e1LY2/u2ekcBAijalfKqRT9ipf/oVg4yLnW
u+hT34lQpmrKlP5Y/d2OzyCNEkcXmW6gqXN3y5pHhSDmOqrZ6LXt5z5U8URReGlHTl99YTuNLU+q
H21s53llgTbQHuMbSfhdH1zzLgW4wGZTlwiqco6UpnXkuT0J5pgkAF9PAJjCpOtOnVI5oGfVCBlI
MAjntG59YEniBSiLgCVvGRePqaFzhb/eNItr2x9hafDNO0SOQbLdmwHzqKEz6LHPYMcJwCR4GHp+
UWHUQiAnNKluVLsECGDKqEybiTSUro5w2yAy2X7wjZBk7PJ569CsYMo4yv4H4/fzCr0YBhYk24XB
wnwMZhB0VOJtFCemyXlPsvZSxMZof+ktm/qB98C8LwLQabmjXNJNqInZ1fkCcG8phow2feiHKD3W
HIfuuOBtSUg9QyCbDtFBpuTttgirTX8r639LEt3tU3CHy7GvtXC2JPaslSR31l1dFz2tV9oJXPMf
gR/Fu9XzqLSFxIP9ayTayujUkaQhiZZo7CuIWc8RmiJcdY74o57JuE6EInTSq7qyyj2Lx3tNBQxe
hyfEO5ZupocZyBzsvjhiEW/Vg7zP0ivJyuxpsuFc8EkwhwYklw7kjPpBNJ8TKcSrfw2zKAyMOpZV
0ji3mV/DUKsGBizKXMzoONE5MIppWkgIAfOGRLkhwPuo350nc0oSvt9CVzyaU6W/w6leMyTPz1ha
hCIifjLtbpI71Jqo3MrvQ4az+lGrSy4IkQh6rzRbKA0AxWbvUuqI2pu2U5oqZdSbJRQXZB9kqXb0
rSJrDuCcBpVva/RYhqJGfxwj5UmzvCwK4PfuRhMxGqljvju+N9YNHO7EXCutZPEs6LP/3F92gvzT
xLyXktF9ReVO/ATKeWzN0Lr385862bIfpEBWFLpSYG/497ePVuemg61Qky2t3tJl9aMbqESJUSnl
V3oHpzoYpFRcC+DNrt0XN3R8pyMPMprQEBHVXYNakilSQw3tX+PEQ7jHJUXEdVpLPBeXTGEXAo0M
PLa96uVYJ4KIV4t5RwUcSvKhXLiAnNTW5ytaHReZPu8vZ07oIJf1dX+mw3n0ig4okBW2aykQ+TBU
1EsDiZ9LpRWHpxyWaY9eTgSASujoMJHQ8hA0pdfe25CShZnvDWq32dfw1bkDqes+U+lBBb2UgpP1
u3eXFBuzxeec+uInQPzUUazRj4yCJmdcqeEwgX4j1u7KcszcXH5UTar0lvrWWDQc4EtGlkkSbr2y
2FRYWJAkrJ1SIlOGGBsEzM1QQEEUzTN/1b9Nxq9Wnr5tYhimD1xINCYdxFej03tJgVDUcz2EDhoN
0Bo0UAoDk5U6J4YKpmiywVUzonBhwpKKlQ5BOL22sIF38yzL4DTIH1fv6Qbch70J3AvEHqNXES94
WVDBh2gzjgXIHlCY/laN3x2UmA/Z4ITlyJQRR/NsBy1YmoZt5sVEbYKNV6Mr9CkMtnsLMKnOzeNT
yebP5zqQeaZPbqf5lmRGo2k1V4DFP4YG81qfZ7cUeutI3A5+6n0NAs5DAG14ISsqIsWg9Okhf82O
33BhioyfX1oMyzEiqFufKINFdQXBZm/A6a/9tekmmX3MjGlMxpDQFWHGIIONFTza7jgG6XIpNqv3
n1UoiwDrqOW+Xda+W7tjrBR3jvzmfZuMI0Yts3q9Ru5ErFzDNT6pplYurmj+oyXHw5yrTt0NCZSn
nRidp9RgKG5RD9B68BUrW3zk188wc+9S9VPdAd+8N++QwnC7VfM6Z+Xh2Wqgnz2AeQ/Z0m0LudCW
n8k2pQBCaVDguJ/s7xzD+K5FyGWYcjE4Vf7iaV+owvt2QrdCG5g5Y1SmQkWUOSnlRCHjCmgfPoSm
sdJ+CcomNuaadbWS2tBPfGuDJLTyY9F15ftSrr/yVHfgJ/5JTB9Y4UONaAr1vDuiIZxKhCdb1uxc
1S/IslipufCG7Ksotf1shjBGm+oEMI6D+NXYfadz8x7xdHti6nDZF7i8oaGlEd7PC5kuaHIe8xfC
S3+4t6pR+FaAf34VPMpS5Cg9oRslbQGXEa8WajxywxfoQ5j5eb8zPhFtCZqMuDcCIeKa/8x5C7ez
K7HSw728QI63yNVMlJl++/yBHXwrERBN6mzj9GytPVVCE3R4tOsfgPHdoTeKBeW4C/G8Fva9+cTc
Za2hG6P5PKVJRwENYOUM3tI56xGbz0AB08GEm1RgaxV1uf/qpbL1cCYypFfdxTs6wW3YRevlWTAl
Y6SjDqVIVpj6PBK05nY3uzJNP6n8bffuKZZjYNfolbAWxvTI2Kv4AcTq+qk82I56zmfqIOQNSHlN
Y5x12VOTqH+0dp4RpE0R6mJO3Y09VWtv6OgCWe9VU7mM6Ldz7v0CX5inmCY5BzyDyS1E0G1e/kh7
uQq5xgfUtuV/MwFz13tgN8X0uVXl0u1ErT8CKgafe05Re1iRXCxb3jAPx98/WXW3a05mtPg7kEbI
SHHtsndlobxqQjtXgpDhxV5hYGMOs6U4LHYPtGL3cuKb8Uvo6pdaPT7vHIJcsAHyX9gmrRFwVk7V
PAepQRk/XnfCUVh59ZjyttneAra12/QJC9fMfIrRhDgqOp8zbtasHjtljbnpwakdv0qGFeyKAaHB
orGfxQase+2cdtYMnxoyOE8dhuNh/qkw8Ko1LCiypP0auerNmlVo45UpVaLFL23K2blbiCDg7gNs
ZaZS0g/j3XqzzhbkluWZ355ZxOzorqFpEwAy/Jt+e6dkf5IXtyaZfR3VkmrWJnZZe5QB6fP99NZP
tHsEVZnf/dSK4a9681vtPMW973NHaZqETb6IsMoYoQnqwiutQwJoXU6wuOGmftgEx3Gg9Rz5hqwZ
EzKOIkPv9QU0pT5XnTybqxk4X3NFtY5mq33wKniwqYxWbFwbW+LBNf9Lb5ZuNbIxV2kU1LP8nspv
Cqc/y3UVADCfazOyG3HniCqvA1tbmAGSH403riWb0OK7xVVaMViDn2Jszbg4zRo+Hb2k9dpazTcG
jTX4wRguoAEUL8gNFaWsWltKL0Y09GYmOjDHOo36b86HjFrAmdauxT706+/p5cHoDX6qIbSgN/cQ
ZM+rLmBfYeEJLFurjj6amsj5CdAxPEf5/A1n5iisE/bnjS1Dv1STWrJytVbSESdclBPZvtfmy8f+
fUh3Zq5vMypHyud16IpiFBkPVqJoMdHaTYwdfT+vlyc0+Jjd6CCjCf3LE4+wqHk9EZNezgB+VRnJ
GctqLkKrcj7fa+YulyL9Tr9Hwyqmp1fsl9DqKzPi1t+vSHm3nPMfHtyjawUw7Hq3hALve3/1b1Ps
2S2J6MLC5FO8AJuFcWcLVWOyPwz2IZ4iBp0tYToki4P9vZ2YXnAzLySvBz7pFTOGfG1ir3qH2+eX
qE6634ZWZYDu4rstZtSXT2lPsIUD8JtJ14ep9rpGg5bLu8SkCD0W1E1Bh4hV/u3viaIHXEGuZjuo
3GVpqxwUd71GjpreBXlfzcq7my+QWpRjuDzTxOIQpUy/RpDd1GXOznCQpu6SA1nv1UiGpRn4z9Rb
Jf+G46sfBvPSmR4qNvyXuxa3zYUU+pSBGo78Hk5BbmgL2dZRQ/w1pgx8Y+oKy+fW5Jay00jZoFNr
s2pWpMPdzEE+7KmiSiaG4rgOZtfTBEOgBS3Fdt8n3PNNQrSsaRxskBP1rvmHsmDv8GDjLXYCScHD
5jKcP6gfeNENW941xN6bbhNm/l88tDbGsQxmqnIqT9UCxnqv2HV+OJ60o1ihFWlZSHh7O5mIXjmU
z/lUGCaTF6HuCMk0pfcq+O9F6fPUNInSHTgch0fe/w/xag14SP8mvA/mC0/qG1uTDXTa4Hu6Pwe5
u+aM7+aA/YrgDiKZvw/QFVzSWhkl03Grw16iM+9EFAEkD6OdK9gkluIGHu/JR9c4yGb52CGuukOi
T3FS+cMAJcsRZKaLI9PINoCCm6oKGNtXicNTY4UbTmdK55+UjmKauwc+XTSg2Z3jVXDcb0vNPQwk
L/pqiAUNF/f+heY9XWh0W76g5468EzUcD98+E6OUiZmDsEeKskdY4qBP29RCcX6ufan9yaPhYNpx
GC8RIrKX5OnNWh/NRHZ8gU8fSCDOvloW1YxQM+eZmc8OpOmBhUgq4yuBdZ/9ty+VmZbSKiFgJKP/
SSDuCvYc3eRfuLQNYATP8hRwQM5VZM178sO52dH09xwO6BSsV37ocoO28xbsBKQdORBqvHrODFh1
Qwp6TQ8XFcfAJ550pE7SJRrIKU2EWWWfUsM3ggIiJvPlIj9Ajma8BxHa5X5IIJcHqBvfq1f82hur
nyIh1YO4ARnwq2CJLA1zSKhL/VlZcs7Kmzu+WYP2V4dmRV+LTSEF6yHiN5HQfXQ3m7zngiKo501t
eKkEx9QuHDAtUzNXPw76z+zU5mAQFCpZAx8UVK0XnlwM3/Ajj5NgVWSR6sgMPXN8ABRupGAI1DqS
cjZvlNWigLZ73pD/gr9374NrfghPcYw4uy1rG9ehHtGUEUk1rFDwG49l/CCJDCyy9hjO2AvfulNU
5ndF5kLbK3PK/ftS2X0uBjkHHUiCqoG8zbWfVBA5xh93SguYziVWR2wVdKP9qniG8MwG/Q52YQrc
Kvex7AtsOpV/lbrL8Buj67nK7/ihrRLZ5CO6/h8RroTN6yPrnevJerWGlKIYGMWldObMQa6G9w9I
NuqDGpDYEEEnS+cRlrouLpslSn2tbVMKdKeN5N/6CbJ7scxmeIMD8mVT4MCA9FuOVPj26OdzMJlV
Yu2mC+pJN0smSe5kQdTRYYCcuCX9laIxIJvaPyCvorjimbMUOl/KflOnEIXSfpiP7CThnFavr7Zv
gdX4ajfEFiWutIUI61qtKGo8FLrec0iJRo0qH5iiH2Yjv4ddIKY+gy/8CIVaSJTfvq74QanQBoxe
UcNjvxboy97EYVK/fUl1HMk3+iPgGbOb9T+IrUiXSerCLXYk+QMLyCqbW6pvesCDOvEjWtdYmiD9
e4bVnY7nmoRY0cmt1Lw90kfyJzn4YFvtwjCxkttXJh1vcgyQk6pv+4QSRwkgOdbMPHZxEXe3LwG/
wVpLE+X4Rqc4HdQf2W3+tH3PaLl8Vd9WVkP/UMxCWHe2WmsbH4xcVi4uSaCZKvQoqKeGSIp+C/An
jMHvDXwIf/1OYqMA9uG1DAY4qAKtA6yGZwRJcM17/uxtX5oul93EXUT/3O9HAiQmvYVRDfVE+aa8
rHDwRS3NczM5bZ6Nu6qe0dSCWzQHLNyc7NxXvJLDcBttwzKRbnnyWIKUdGrk8uhbefcw9e+cvne1
XMp1cp/acz21Ole0M0fv/kTYZFG5u+Sz9aN101Th3F5M8Gc6oRQ5MsfYh43Bv4WjC+f3UpWXeyAs
pyz/gFBQzqlfJ7mdHL9skQdoGTakDazk6W+2XynDjyAHWUpJguHnl0UYnuBMjKZW6QxXcr8SeIQk
35Wp8cpl7iFFy0xPLAi9IoU3W+NoxfMhdh8Wv+zTEVZII2cY+sjsEG2CQk6yVFMbMIvMntpcsZ6z
TAif/bGd4QFspe1bhoRPv6t4fy6eJl2srAAoJFcx4xsABMRLVqTocaKbvFgiob/0UkZtFToDiRLl
EAqZ9w/EreygrD6tI45KV8hfVP/xGVfi3OOxHCyzrsr12/5O7HcRlZkf2XeybzibtpUpDmjdYXi2
oqIQ/r0F3GpO/2Yk2s50xBClmJOubTbzgPfpzOSTgXM0ZTTE2yESY/2Yj8lqDCA4dnrWxu/22LbU
LBIbeo8ED5aFgtIDKJdDTTKt6VOH9wT2gNHQQJIFKLwVmbzqJCQwfqqFg/VmKW8c/zVJzyxwtT+T
6jkJQBJOlPFBkOqRTxvmQpFMy3OvaBa7ZgHxXs6O+aUo7wnIv35s/VCzkqgEOzhQOfWWjO877kab
BtRfNftXnHX8wKd3vIudoexFBGBf1sO2I7XWW2jPhCVpRGpnOLT8sIW03ec2dpf1W1rHq3/3TreY
d7Lvca4K52S3fZ5Rt/GymmjCom8f7whes6DF6lOkN/q/jFVrUYyx0u/ttNdnRpK6qNXwde/caXaL
P/HPa4oS62tzdpZCXlrmx225MQQDDdZjiZfkf9kikDE4bzLjw38m5zUPzhWcW0HQHfkGKprRU88m
aVk0CImW92n9rBIQDlmymMKptE0v9d8vcWHbU5yOz9iPddZi5Q6jIXuUBgrTi/26CKeRmS+W8Oe0
8RPtY8nNi9voICXz/m9Sy1wQ1Nof6OrDCACHILbrcqeIpez84op3QuwKPfXmpwFw8yY+B/AzLi/g
Ue0LzLVmBIsGMD7/vzxQNihKjd3sQAAW5dtBvrzSfuGO9i5b8UvLlPe8VOXseEvaSPIFhABu5YgA
Lv59P/pzz4xiGNa2S1hRoWUHIfO1rn57aeOryw7t5mSgHwCY7lPbMgQwWmoleR2L4WqagcLBpbZ8
vWtkVOTZdpvzpxX4NxQId9mekyg0NOAYVX5bgTPAj3rYvNTfRSBX5+K0VQxqBNSuhkYSUVi7OLff
C4wqeKIhIF09q7a2KnROfOnrDYn18M6wk57Y+Wvjz69ynNX8AXnPUyDUhwnoaj/PC8Zgd5HkQlWn
e8FXaaG6vx4cEjGQhLaqmqGO+i1fI9mpdbqzTncHoAC60RsdbFlBfOz8SzHH2odSUh3SshCBo9KK
bDdftk1VduyGdkPB/b+V/AHuBiRq8EAq2gip7U3uUs21X2f0K1VXZUvid+zDv+6R+1pj8z66T8zk
k4UFxuYOktqL3CbqLcBuCEpj83HgANsPcTBxDNNlplRrZ9SD+vqfWKff0I2Y5d9UugkBWCZcl4HD
+yAm6Z6+S1V/kI3HfhkJmd4Y1TdlAtMmxfFQb5lZLYSry099cCqmdUTruZlA2D7gtWvcuru3zpNT
TrbKwvn827LKP2CZmvAlFLkn9j4er4LkzLm/0CD9CX5GrK0PgH7QmRfEJdqvlS4MQPf4NJbMd2Zh
RcQuAgPTgwFk83RVAwYVM1N3blCky2rPTYMJhF5uaP5xAkt+IpqErCpCWzfzVoptrh2bclGqFBAa
pk9zb+3tvuOT9Ya647LqGJL3Ds045BnnTtiPIA3QuaGxAFWUGe0wNVFLlf6sYF+GVUcem9RdfC54
0VCu3q4yi3qvF6TO2VzlNVlEbJ5ycRuje5DgX2gZZ6SMC4KadeJ9uGgH7DdHtr5ZC9Hu0r2KR82g
/FtUr08fbke/KneXYsoJSl40pB1pmlUuHuymmgbGwMYqIqJRwRZx8+iuyaZQtpDedQrwBDAuAdT8
sFirnXuJZP9valk6qPnVNfJOjPoh6dbt7tDbmw2BoMEC5IHNErnuQCW/PwZwTQKzxrLgTRiKDjGl
sKcz0b0YSDRVenWcswljovKV5iDdvThRi2TcVumbYIQ2Zus/zbr3SrGenvlaQXLs32Qw3CT0kAyj
n8LHH6dPuc3ceNsqQwxVqVS8GYjiXTaoL8qsUw0bk2Ka4NzhlBk07amAKMpKpMKZjXSPrmMat6Af
VfNWFOgzKS262E1jq+vxL8/p8SJPC3DA6kL+ch6LMSvi+00iiOsIOpWFM4u0Q4mCbVTt7j2UmXPq
K4IVo1ixd0IyUcpneSsI110QRCSJ794JI1Twe3TmqN2tJrsjKSoU/sKFOspokp1ToAL3GIUna7z4
4YXFePtn/P8Lb3wYiFB6tUcIodjnY3YcXYexSJfb2Prui44Q3kpVlmzF7iOiJ9E1ezfip/dAjpOD
sFAaoCHFKikBZ+lsnSbcLUcoWoXmZa+iFluvEYw3ZdqjvstNhUTJH81IqYYFlJQUxGuIs4Mh7l/P
spluuI1FEXdQW1t7eLFNc9cDigtiYYGRiO4Vewyg4aLMzge5pYa3A/zyVP3wf3Xh9hgS0Zz8ge0j
fAa1k7v/KQ75pm/zQDf4rS9fq3cMJxFR5NjonR7sxuvobLgX2EaeOxf3r3uX4EHZwaMFyRSHMGfr
u3WizXU9U7GsES61Q66IeLHoX1G8ML2qZOY3q66kyYckjm1i//6asU83WpnvnDUi2Zx+uyFxos/t
CSfZ/hd8TqGd7m2p/hKtV9ceg45FKaBhE2qxyoe6EzZV91cnNt76m5SA5QLbkvwhB0zO4jEumuVB
JRzd8UAFvTFNwsQ3AO8T3Atnjr4cC27DhOq6TXMFh/H30u9Skgvcmfr6Mb54ihF1BMJQiNXSg0jJ
Q9MwJ6H3Ri2xGPJqdJ4CUSm40+o86Vl6jXK9EDFfKPcVB6H/KAVyzZnHb1vedp5oljI3aZK5t712
6pDMLwm0eiAWihfrz2iazxDGQWfR9C4t0ECSN9UcU7N0k2DfAKwyHiUT1REHCBMlUwjpBxGaFV0+
PvisKMe9fcODtOC8mr39pTs4SZOwI85lrrLHc9gRdwqS8yAbEgexm6ahIFAiqkkp0jI01FBj8RQ6
DkpgICYF8l9sasnm14aerfVCVutej3W8NjbLsWyHgMmebze8sh6YrpL/8KMr0StloawAP+ekgXDC
tEUGvSXveFr/9ucG05kKcAaFHdeJmaz35xzjNoNoWd8TrlfgPPpM4MowjrMX702g5chuMqfWj3Yr
Uaoz8kl1iAPWr9Ow5ae34tcRYK5z5LW+qEZS3slXLiNT0xb8KPTUlb63KfKf/xxJLXXMjxCwVvYi
03CmI4tEPuJk8TRTtEjjMGCLk/K09QRxEDHLQaeO345/HX8XOSDZnvVxufRkfho993UU5PScRV1W
x+S/y3W8dD1ZEDE6ubm9nqUt5N945qhjMxwu1C5o98gJZrtXmIOZbGDukZ8DS8WLafuMBiv20U8i
78mlAstiCcHmLFdaUVdhHWf4tpe81P+sYotHkRM89DkONDFrYswTBXGwQE3Vuor6F8q8JThIGiG5
l7KN43PLYhwORx/bn/VKBWIx/+3WB6nQAvrQOuflVt7gF/1+eXuOPPcLgwfIswjrXzJ5gZEUuQhB
pI6Cu8kz4LJQqBh7ifaAqCc6HUKg2avNYeIv0qpWwGPGVa3dQwSPcOvwgOOa6f/Y2gNPvrtIYLH0
hvMF6P4PI1dXtidu7RiUdkDbV57lEUa7QgFhaXsx/2cc2fGDDOSl3yuQLKlXdHFLT3Mbf9sH2ggE
+lEKCg4xwcofTaOT23VlQJopdq6MHMhnzCEmcsQYT+JmN2eidpx/fFVGqzEJtGeomPaaKVHQTA9T
/2zYsLVGq9gb5SJItOsChtnjHYjJu7fvxK9wUqz0NvPx1JKd1FceHXa1y5Vy7aEUjnHtfdu0mlFW
rVwVwdLlkTR0RKAs9zQj7Zr+PNG8H3jBZO2Lhm/esYsLLQQGCNueDWvaPOiQYUukoRFDK5UAdOJf
zceeIqYtlvRAno+4EcJQJnIutegW8Wiodnq12kIQ7QYwLOBDtZH6RX2tDfS0V6/3N0wZE0hGFCaQ
IaLW4DzXDTtSyoGo3VdodNuNPv6Y2Z2GjE1Sjw0rW+sJS1M0k9/KcsDl9/lzEoNaixGPz59NHvm+
1ffeUFvbJaLB6NQYl+4xkif3EaH9h91O0A0TPmodgP59wT4vlN3j3ICGrrWS199nwqds6K3X4dWG
4gBCVIrtN10k4XdRQiN27caUrnZ18grhwPGNgt0NDaar3MSn0an8mckkvICD/g2Trt69HvtUkkZ2
My0usBVILZNnOWDZAzy0/2jk+cpZWcKS4sFrLURiK6i3D4IPMrzx5P0FZcF4h9eUerpomCnwRQvL
pqJEYWECyWZdIGxWOHk0MUCJ5hjFzPYFC3sitbBoFSlwYR9NtwuUGu1YhJ8dyle3ed9/8b2M6qd+
ILMxS1dNZ9brox0ek1viJ/O45MRRtW14TjvxyFccotZR3lIYHbiz/ds7An302sfzl3MEAKt1yJaA
PUPaH1IptRqpmB2WgE+I4DaGdG2C2OTVrOP57sbrOuglgc5xBZ7/oWQR+aWby7mNidt2fjLd6CvP
ffkC/x2Acc/1OBrCZMqaVcOczIK5OfmDUm98nrSBhTP9un3PkCZbzRH54eA36RjNoG+2Mu389XpN
ZAOS7T3KqWsOFPbwsSYCoEPaKVz91fIsOwsuUIsi7FWjorVRRatCWIDywMR+dRhg2q8KfYhPSA5E
dBPzDUOTe0Qo9t0JvWZCXElD9epDTBEfGBJ+sI5d7T2c/3XbVYpHeiaBEWLNFF/YLCjEFnUsUPUw
6aKtu8LuqGoMZ39aiW80bxzFm0ljl8eaqP4bBtQ1lH2VS0j/dP9xxBIrM7aSJmRgjk8C6tTWcjFL
kLL924MnCbegWjDcqD+wD4qB228EO9jr+Qr7xT7ndUrmYD4lXB4rTbktoEyUiEI4Z8bWVx0m6Qo7
bFPmUoDhdHgSx3Y1MJ6YgeVa8gQ+sHtVggGhm/PohHwmfQwVF1zWK+vyRXmt4rT7NqrIHuXZgbnm
ExsVf7cwNeB+7hN/Gu4wue8gDwNePp0DtOq3qiX2+D9FHxx2tJF1XDNDW0lEHVk2LBrJU+JbBZMk
HTQ6oAsZ19/drr+6KFGSaZSCfQjHe8VMUJa2hOPFVyk2ysxKiykUaz2Vn1H9xitfceTgcVXFCXiF
8cHobe8Z1E1jLMrpUqagrhcGsPKNjG9L2bpiRRyCGLx8/ri2IeVvTppNN1S1PcE9IxnYV8Y1SFA6
P8xUV4xiy+rZt6jtpc7pqWAPEtZwvw/no1UzmR7Qc3n0gek5DeGuMFxNiz3jlB3OBnujBJoYpTv5
kih1oPQ3WkpEx9By19FBTUQ4nq8CIacbxbmINBV3wlPkFSBxwTmMEGneaxJLL9sKb3+Fg7JDYknj
uW1jkKsbvh4NCG7vVcArbS6PnEwwrX85z9qK9hYucms3rnU+jX3kt4PL2bQ1pr7eBpIjUQ6eRIoI
NyhDz6J80FhX8e+ZleMaOFSA5iTUkoU+d95rKggCqBza8I/MGcTx+uDhwUFeRkPunTKyEyip7kg7
zn1i5j/+tjummF1qZtWU8+gFE1s8k33nF35KPWDRp9fTumiuRNy4t/XV0hr0eH4Cx02TYMR8Zoft
pQA6oc+TxBzOenmvqdU2IBfTXNMUUl0pHeVGNAi7WFpf717+g1iQEStXXQyNhX1fx2YRJq1l73aC
moYDkw8sceexMRe32yljIXU4LVRTD3NUQu+A60JusBSpIgWvN/rAqSfi+of6eOmW6ZOjRduJHCBe
9O9Y8BJCMBs6FKZhmHzzB3uiwIOrhJnUTbq2Z6pZMu4z2rq6bFAUP0wB6S+KEMp8atHb55GYoC1Z
bLHK5pgojTqQLAMyjGuMCziinREEgqRbsRXkm43aP1Dhq2cVZps237ON0H9fnWAv4nQjYzFHp7vy
3tORbD5G5BoVnV6Gi0u8eu1EtlHl7atTbb9FCghe2/LuRcvekD1ClYuOpI4V4/0M8fLQ6AHTVAbr
nXb5nnnSpASZxjWVd7y7G3SL0KpQfRa3S9KeAa6XA4I3sGCeZTV4+OE+XxfCLdRxnJ6Va95q25mg
ugIH2mrMI1nhJtYe9uqGPmCnqs3NEpz1G08nsxv914LV2qft2o6az/MevP4Z/ztWpq2XClBJG/3+
YD6gzScb9P7T58gdPJvqLu0/LjFowaeh8k0yMtilE/G/PD43P/Lw1CeDGmX9QBO1ZwoIv/2YweI/
fZTTrIU3nxChK7jVG1rodcEts+4EgYJW2PjaKb7QWcq8/wnDv2xcRvUUCaPc+ng4kDLKPNJ+Vhg4
At1H0/kjle4WRoa0un6TH0PN3+OayaU3yOT0PASdtCxOLzAxodgpbhclpKdiZrNArfaVvOR4lSBQ
qEE46sCeNCpeAj2Rzu5TsAnyeJ5EbEteHOyaxOees4Yvv2J574MOm+JZeZXEmG5x/k4FtECcg4dn
5YBGMUKIeR32cJOLAwo1Qi+z5+RoiBm4SF8PyG4FPN15/MBFXC5yfvuG+yHKrfTAoqkh6kLAQuqr
7yzcPP1uF8p6g/OZ4lw7OLKXfPEezrtJtXELnT/nPgsO5exQo7Y4cxXDFpyDxAO90C5pmx/rawX7
L0bp8CS8J1yuxU9Qn0bWDjGAq0aw/agEcs3s0HbEMFQaHgBaB9yZCCK6NnB7WTA+RbzSmf44dfX6
HJvE7O6g39K0MMenA/l+p2mqzfRX9KWUP3amktegCe5WnBbzPADAD/jsfPDKicpP9y29EjqfPkUy
t+TADgDwO1qUOWbyvQgjMQxaP3aKVFRsKHmB3o2uIF2m7SJVVDooCGasTrrWgapyMc0MnwAW9Lp5
FOuMd4v9mHdoWT/+DEFsXPaPeex0taU0qvmD4WInPjqr0Nx3W4WDQUWYgnPQ+T3kWwyzQNYg5pZ7
yf06tDCcxv8OPkG8moWgW+7fLMs0nHrUwTnParC6532aFnd+cERJQJ+EKF0smkRuD8GDLSvGJFOg
6W3h9zBcaS7b/QTLobmwyhxTdlsmOxoWO/dUGqNmTQAb51Z3Loktizo+58+tVFoIZ80St3PW+xO2
2Qd58Z9dQBNMifodhiDl0OM4pJnyLVE7cqf4ktDDCer9imF0rDbityhdDVM1ktBwoGNNwk0CGhVK
01zB4xs7ld/bN0Hu7PpQK9ZAqdrfR1sqWgZhlrwfGxjoKdp0nu0HG9kpU9EMGj/ksD3Ddzz6e+Dv
EuxT9DdkBfcvJMMP+0mTHc5Sb55P2U0Uprt/U687/b5MkEL8Opxq92BtarsduB1rI2QrsB9P5SLb
NbFsGw+87IPGdXaXa453u+FUz/8c6sBjwBLqqYUS6+t9WYpv6+ImbPFTDLEvdLay59xVS+VIgDks
JUQNcg9buSFyNBgwrzViByfwSxCGhugld5ind/0HGA24T/rvIYjPNo/JEN8kAOJs/zx1JHqWFwqR
iRsqb/fkGU9Qf94i0VqOjQTXKcQlA34WX013bVy/MzcDUppzpQC4uLsm/XDvxOH92SDkgfZgPSnv
p07kWhZktf5pJGrtjwRoijJB5+tAwzzA5QppX/fbsg8mGOxG3U3EwqCUJQvm6K8Y67yVUw3i2kBs
6vTd61VIvjVfzLk6S5/xDde2pLLPq1LwU5Mc2I3b67M52jihVFqLKdU1zHsY+PZWobk0s8orngIs
Me9s4DdHpAc+OksmnwkfwPF7zhJUhZ9rhR1n8UX4xThAjP19ECUVFYFENwFnOQDUj7SBTdYJKCjZ
+dSv0xTZFBgZROc/STRvRPPDcJmIx4+uLj85f3zv3z6AVXUwZ00AlTpZOlHj713AoLCTfPaXaNbQ
pRYIpwk/gT4RFFLFgqcoO5qx9HbrMGxKTl7iRG0Q1dGcZ/B4d3MObkVsEdX8FsBnhiWF0V7lA9ah
1f5YpgVWjjmrhjbuwUEfCdxTzZxgg7Mq4wVX7xS9Q2bk7rMiozlM3iEZED9RlngA7Ki2sEi9Fn9N
ItmZMJdREGYcl+5UGipajdtI9yetD6yqLHc1Wzw4OtFjBrZcNUhuLy75DwwrcpHwWw2Wiz7bxWeH
Qt5pA2ld7zvPtZoN3MylIxeUJRYeSgyk7PNOtzkaADRgs75QDEpdn0K9oL4tU0Hn/UrhZfVKFsv8
Rjmpw4VzIbZaTzddUigaKPxfrszceNXZ1+zA4RGrCYp6Sb+gbh9FFiSYobDoYcG2KFmlcH1UbuoW
LReUY7xgUJvOkos2p3I2IPiFQ2TzOf2BbJLBbpbXK3mWxWDk0acC4rBPneNmby+peuGsoPKGtcv4
gNN5qBLweyfiAqQqqqV2r/yRN3SyyRsftpPiu+n22vl5gsSm3wBcgbdlCVgjtt9+4EAyyPmvhggR
ML9/9IIrHpO5Ro5FkstEf2tcz+q0nE1tbonvFw6vGz3T0SD4Py6uOgxVodUfFBS74ATnY9KRxiR/
srKc+1Hd3npioC1C8h6vJ6wgSkB6YlJMH4Imyc5UaugNju0C6MTOuWNvs8PDPJJ/pBCUttY6/aUz
9NBsPEBQuLzs+Oax0LUVfDi3tNbEGCVmf2Emvsr2bE+kRViC+lu/036A7W4tu/vWDINz5WB9V2K6
xt1esh0d1lQqS2AZenp9wcUW4BIY9nNQYOWiymeMDMRIRFl1HexMVaGdlP54fp4SMIWEIcn3bukh
xzuflGVL5E+iQAF59UDTloNM04MfFs2q6oCSgnmRpDjZaUAesrpguDmBuxGoD8U3K7uMZz7OeIFs
AfXizgc944R2ndmWlHHey4PPnIW0uyuX5QvgvIWftTHuh+XvawOqzjAdy708W6AyLJVoKg7Ueftd
TtG/mBeY/5hEhMFXTbEg0uQiwuQOPsgkvXbi0I+H7tfJv2voHnTbNq3P67VMuO6c/Qe/AatovDi3
u9CQ833D3O6UW9EiXo+uFtbLWvYN5lA+5Ps6u8r2JPvHBbuQch75qVLsC89ujPbM7xpc8PCobtcL
EidXdUpa81bc6OcUpz2Sizl85212sPoPazQzfQsmF0iFKfFElDs2c1iqRVnOBFbVTJdcgWzNmDO4
pNRx5NNulLB43i2zVjiARykWV5ABQrF3ettdNau0bPRTPErR+sBkDeBJG3vTUtn9tOFuIj8aShm2
a+JWKxo0F141h5e5q8P+2Vc78lebxL8Um1bofvqBIu3TeQOTbgxIu8NyAnYHi6D5SY6+WxBBq60/
cQQW3+BPyHH3YSJwtv+p05P5UPCTR7laDaRtDZh1kIQicdgZTpIBwSxMAjpGB+Wz9VS8WY+8/ggB
AKFIFovAPAph6aIvWe2DLmWuzNK4SEZ2z6gAGsdy9a4Ps9crxvXE73bqFAPkUjVPz1EcTInzQE6p
7iXNoZwj6vwEIaNV4LLgxrpqEHDFGcciTqQ7gJp7WkPShvwClrQb5lyeLQFlz89GwkB3dJPTHkKz
tvjQ3vCmqRmh8+OLeH97QGpYmWYkknnzh00YAdhcnlpbGTmMAY19IZzbwvsPEy8aSGDkV7g/lzlB
0o5+e1sFZR0HO3qLS1zc5Xm+xQAW35A3q572drHEIBd7HX5dXTiY3AHWhongVQ/miXotabYQE4O5
TxTLWllFDUexNKqV5kXn8c8L0MfYXqebd2PMMv8ZKbnsoFmwkW5sFY6Daw9vcOAOMckgrb2ZuIoV
3GISkIklln0UqCi5jGizEGnd+BC4Es6+LIO+9+7QWUsoKah0h4BxwC5Ax+avu+57eX6CtcsRGVnE
rISTTxR8YLZALkNZ7pOugXOVpYE9jQMBWP55QqXd/xDYFIPEauriRUjBkx45rAf8HLio/F9gX/I/
1hsv+91ib9CXVKpTgFYo2bUU47eWZatTm4R1vvMAS9i3slHZ4G2/Hd/7t9gpCZqvV4O4OfG/EkFC
Q6dfoi+1Xx7eEfZzFoicle/CY1nNGbuMfiba1Itsz0pixl9qLs/oZqlpmYx4R1JXwRFYPq1FYgqQ
zhk0MIIEkyxqs4WI5RZrCJS9m3S9Np0K4HQUosAB9wh2PzwUuAO3qWzqZu7uXRmp9lbSr/8y623T
9ys4s64orpJRik8fQ+/w9fGkxNelC8/rNhK7ou1mlb94W/k0+KYBl+4XcytZYrRiGIst/cX5/oTi
QQPaCpHVRfNY9yden91QVqIisjdXZvF5Hs8I/NNlAtBOfyPwqd1yjGnNtujlUcUAPcn6MHMuy5I7
3hBChgiSD4cnrgoJIOb9S8KBt6sfI4nRp3CmDzUOFc6n0yD45ucNUe2/mDEzDF+FPW5VvcFGmbEE
yT4kMBtZF3ujRCU8wuqSYbmreF0FAb6JPpTr5YdMxvOFqi9v1pkYzKcLWMOiuZj2ooH0G2vs5jQ2
zSyWYbHMT6Dz+0Hgg+phO+kJlCIIyPIOZTCe/kc4PSj1hqcFiNQIzhSQZ5FyQRddiFJ2yJ1rU/UO
7kQvyZYCCi8vQX2NhtJUIY7D9r74e6Z73Mgl2H7axzJT9e8J0eG598bzIsbRAyYI4jTEb7GLaVnT
+o44Y+Wg62r2wYB7zTKFagEXkjMMaH4AZVkGMqkj2mth9d/9qFiTBxvX8m1XvAW7X0UbBLvajmGg
ooz/0BcqjzQEw/H7v3fv3eKtqsaMCh3B/ZWJqZETCyLqClKRUAp4z2YCIBUwbU2No/OqkWEXGmEK
mQqu9VQBfxV90IKSLyi4g6SLZ9wmQa8z/lJopkE/GSDRgNcUbsOTwx2w4UJi2aaYvd8SHpSvx410
eMPNAuCQpoWLAWOZeUDi4UPJggmp/vzm8r3dYT0N/EQQZi1AvDDjycwfoKBpZK7vFHtmAU4J0fRv
iYsAylMg+LSEYNWlg3HgnbJ0yoVJ/8jpQacqi4TUiuGR2dB3cSuA6ci5rXdbzQJreln5iwgI93mA
b6muHbv4KO6T28xjfwtsPFhMbWo94afXNzyJoC3y/i04YrIBA48LNJgZiOELhtYXE11Qhof17slk
UPl6FuFDgXQlOq0vKLlnMUBMVrlYjuW7LKLbwNuYq3SLXV9ARu9Gm3qUa8S9Op6H4grmE0skDOwx
WrbdF7dTHFVQkYmNNAkJUWkjSatAsbJTle6aQ/fFmoO5+cqN3EcHJQ1AQilArAPf9For8daZhoGZ
wDc6vSv18HfJpF1jnh7cG5AVqlHniqriw9NLdsCezyjLSMkwN64Tl7fX+9eMR5knYBCgvUikkQgP
IXWmXi0taOuOXvXvAF2/MAsibd4FTv5xQD7iLcYca4dP1tZvhiHIrMQrgGUIpIMyXYiBHpp15g/1
Jt8oxWW6bhHdp8np66XVJn4rdcEohJXC+t6xjsLR82/4MZ3PUOFp534PGB6DbPltZDzu4p8TwT+i
MKq1qIlR+KQqVEAXpQK8TRdvPVmJXvT8a3Q2cFAQARZ03O33CuJtyudDBWbkt2pMYL6FByYuzZFH
bnE5wozekm9KEWJ8YPkRCsQxCHnDCRYf/gHUPjYhPpCdfkozWt4YikfAQOqYfV0XYjyDqy4iXm9N
mS68DaWxIIx4lfHcC8Z0m+y1+VD3w/WDEZ2PktsSj1ZE/U41L0cbPQr2djCvkjZYEnLbq/xufYXk
eMhglcXIP+YbVzMbzBNzY4WiQ0g0dGE4WR0cvDCzvVB305VR8m3Dn1Oj0+da5o7EFXOGg4Cjuh8L
/yS3tfNGCGKm/tC4uNjy4SHOuMhujJ9dLwfQtIk6nsWxc6glLoG7xCZcakQFh8y+b+xx/A46ufB9
23VIKkFXN0vbarn9OEmOXpZ4wf3i9yOQ3v1xhG00C6yStrEcdvulmDywJOOQqEv83HSSFh3p5L6M
OT/BKAIQZuQT/COM1Jb0xGFJoHjs8OHiE1shhf4cpKP7LvCwVSeLjiFsBfLF7WQZApC0TgeOXdKi
A9hQNw+byBALo3TTZ0ET3YeJf0EF3Jf9cKEn5DPqe6uN8a/SyftoXmob4Df9qqNsbP8S4elT+R0r
b18Bjtj38TD1NBRCOrC2uYRsyvltMJVwp/FoKFu2m5NoxIViRxlq+nsaYGqfpQB9eqdZomOlG1NT
UX6YVUvnUS+7IMNRNpaE5/Lz7bWwC7HqUCsgvcoYicsOheJUhtZznJtVLntU8B2syc3Gxm2vuyJD
G2OMts29dicPUIxF2DaoRgnNzftNaJ1ho6Y9Zf+2Z3hTKgzxmuAH5B6G3WMrq6Y97m5TJrkoIxYf
+2GRMuqooQD/UffOqyO8b0shgXvBGAJKT2rEnuLlQJyWnvR/YfHlsZFi2m6GmRASrTI2GaolE5hB
Umfz+koJOILg28/zjmu0iwcVYGS13foRbipJRx8gcX4479yTj9aa+EQE36Ui8zGcsOvMJggx3scn
tCEdaZ0YwuYDPCSV7VQ9fZNgwH51AMicwn6Ea/HjUiUbs+DeEiek19NtP70Wgg4ZvWEglwye42XQ
XgF+HyQdvmiltlBKFZ8iGJVEBoXh5Mont8tzlkr/3YGtQBC5UrbfDgy9vGvewnyupS0eZFTf68E2
54bFAj4a+80SdktsdmHq8ns2TKIsD3Cb3hQQ+GlDciz4O7BiMVvkV2wK7fbCOzlCtpWS5B5//C0r
Io+ZxMSj2NQQ1i1YNQet/hUAdtvqtDMIsdLCTrBFVTbJwni6LX4w2i0/bBweGB2JonYMtybs5HQb
EdeDBC09UjQUPJQcCz7CpixR2uwF574H45HJPOuZ3kTcQDPcLFm8kbUx9nJ0wyL020QEyMSrnAN2
Fybi0NBOk/IpOrQwZsTbDIKui7u1SMJRMcR/smTjxB/7qI1M5+BgafdXHGVXRxAx1MqK75Kc4ve7
q0QdG2Accj+ELt7W3ZTBTqcNhtT5leYsz7kMF0W07UAkNBEmSR7UUcW3fsyvZOaf8hwh2wDEQmSY
ocGFYhVJygVBAnWk32AjuZBc5+SuNyT1m0d+1t2bwDjgSAEEv5ba2hHPtJcKUHQDG0RkPtaNeRZo
yt8kkDYvRc9c+wLnAYQzaX99mBeRpphqJDG06TUEnD4WIpAUdJeAgpBYfDsf79KCUM+3X4ox/fxw
oHUrrQXU7Lizn8sMDlpEMii2dl6xuIaswWmf/IcVUabsKGI14u+pbA/GoAukY728Opafro94jXi/
p0l1Eaj+RxNo1JlqWtaiviTS+hLrm/9LejmZQbvGNf18OxGNNNg+rr4OxlETGXffPKZGv+Lwkmz/
iVwKsqmiKZB8H6o6rX2AoJJUNmCkNrAQw8zGHO0MkfcLFVJ5log8fh42w05d2tAbXLL2wJXqgQKb
wdfqWxr8nctG4xsoob7lhc2gf2wilUj2tfC+irDKi9ucpZK0ejMKQ2TZSdYao1Anrx3jgeaUtJgV
+eYFYKlqZVd9rDv7s9Xqkuim5Ns20PY4fGqFs0rrjR/mZXU1ojusqnPz1yQdjIfYsnw975ThL/n/
otsdng9qOQyLHmdTy2+dCHTOinc7oWUfHv85+8keDNB4hTGq8doFusl5GufMncBVXu16WJ8W6lGT
rzyOCDOnVp3REN4zaQ2H/NSKysf2I5hvLd5QxHwt7hzkUgK+8lXSx6tohjGYcJ77n5Dvwf1PaiQ6
MHe2L2pA8Zz9xXMzLACEnMdH7Kl8pvUsGCiM+pDT0JOOdbH8O4Hb6yz5PQybU5YbFgHLK89vGlhu
0zn8vbaaHDCjx2fHIOdrG4q20xE1eapd8d/j5dWSzQsnVWh9PZEVf3AelBxxJwDa8y6DbCja8h3N
KwsAeGcNtzWLw1bqR3bYnIbKQHe8w9vFuECW009C5HNBd6caT2PToo0D+d39Sf9F3dDFtaXKS4Aj
2CfABXgoH7hndq4vrB/8nUtjpbT74x6xL8VGqSBLwf8A8EdbbRtAedBiVLCF8wJxugPqYbjsaZMJ
BBkl8OXsJul4UAD0zPV15HlGd7HphgfJ0aVAUweNfBB0AsEZl8ntaVgHKhGNhmxkqkDdFZYyB1e7
GvKUu9JTB9C5HuND22g9jK4qxkjBv2le/z8BZzxsZR8qBuz0w96FuwomHZSYtoL7BJ3zGXYO9I5i
pRdcZn73hVaS4ixCvWkzHdZ0mEUdYo7hVJ7V27E9RqcO27WOSjQJGooTzifLnjAq6WmESLdaT5NS
2TbfPxEWGuSDRsmWjfkQkKEvZ0jEWtDBspCX7JDbrXtMWrmy+idhHLmT1V6FGbfZT0MfJZJSQ7R/
PGSvkN5MlupY47INfRH5qufVOtC44xgiYn9AOXEcIOy3OjcIKkU7Hrgse1Q/j0myO8AiwsSd3u+H
WN/KGvniMYXiRLyXivkYfvBG+9qQT1M2+6dIhGVmx0ZYNTe3GwBYWUCtGHa3N0yCcZm0NBtXJraL
s5zDrUwaw4fMlHpBtG4PMr/V3HXm+Wao3bhcTk+eqxjwh/vcfqatevn21r9PE7uDNZoVKQFSJWNX
l9rkeDEQMc0O9o+uWN+xhbFU9PaGd3ScTBHd0Wmu/9GyiqVdtCdcc7DuGBrk3w/hjDzwkjvncHwe
VM48mh3yutNI7NeLbZVIsyn612xH046jsZ3EbtX5xCuFzH+H43M18geMHAng3E3RzFUDPmjr2pwL
4bXsWnI/aCjjMSzTIdZYQG5341KwsmbbBBivK4Mw2oqzqPkZno7ptMVRLfSZ1BOz+qRNWYiOwXoK
eDUoQLiz6a9ajK4e+badNXk3L60RUZZhKJNPedAuAvADuxgsCwT+mV4eN3YMeRj5PF1rEJ4QXiOi
o4I4nY1kNCrCuJaYjYrvQ+nOOqQtxzqB7PirawNhtEPrfa+6L3neNT4XwCq6x3MLYr4GYVlaf8B8
uN2gKyRKdt72bAK7N8i34TpQnHo89d7Dbt8pcIgoKvN/KxdbJPwjN/oGwOeaXNuEQOKIoZHL/2KK
LvSS8kq/5ErJAfJWF75ghZCRe5VYCzU5yMLyL3HYW7mZjBAd43vnGR8yolroHEoU2fznIEqmy8jq
OQ49k/De9TlhkQrNaPOEBIVveulXdPd27R+QKi8venxcLJQaB6ZD5Sx7u+S+YgwUsOLpBqDpraP8
PoULEbCz9CKqDx8y74r/NmBf4E+BuJfJCoMg3s+bhhOX17nYTtbOkHteSe7EUXFsUJDPGrOurenY
nAtTM4p4LVjWYQsZcboBr7/rQNnDicAbooUMyyGn1KdbrbzcAVb2HAp5cVZgrFvRxSSum5sgSJ8Y
HQv74ZBVw5x8kjYtKGeDxPf8wXKMlbXRiXoS+x2cQ8NNFxM0LcgH1pJt+CkT5Y2Qi+4+SsgzsjVa
y2SLrDjrZJH79rZGxoXx7M+uGY7XsQ2/LkNqMfGEv4C3bMix5yeJj9xUGMQA7dfOZXvbjaqZl+CA
perOGfHEhbuS+S/0hAjSbhGsWva8KwiWoEIyRep8CRldmXL7gNuydXxKt8O4hf2oPGVEFq32fyB9
ToxElLesyoEmIp5Mv7c7gHX7GRTHt/mtYtPihYtD7eooKhEal9iDTNDPmZqmPMibQWp2eR0WxTV8
HfBhE/KyEnmuVTSo4yQxRft0u4OnpfPuOa5PMiS3wNG/F45ahRYiAZPkhXj32eMMd6FsIQnjg+n1
pg5BTJDqdkzJJ1Nnuw9x69QQmz/FFUOQN2FUH6rKGon/x+NojL5LR7X6tS7VolYc11IKK5vuaM9z
1975EHwZP8S6Dfgwhzr3Hqu8C9hpSQoVzZxz3qKYFSBw1gJtHTWKoHnvryXOXgmCpTyZJzhzgutP
EQDiOt8IfR27oPJz0UIPZyonRbdTNBPvSA5LNXWQcsT6uk+u1UndDX8y61z1u5o77KEx4Fgngsrr
LJ0C6AuqNmlJ//N9IzRwV5Hvo9tPnDhOb39IwDGuZbIGMN/zbLwqmh9oAj1VSOxPlAbljOREPAQH
9GH1usSOUL4SfUFLtj1godAc+KQTqF2HZV5dZL7QDpOC6sObwXrW+1Bfl76903GvqwCGELGx9xUo
PhcFm/hpFkT+PFmL8hPShe9D8UZ5mUYM9S+WLwncbWyp6/tMX+XT8HaW4y8k1fXax5pIvRere70x
+08RdMjOsp9peTbgb53wOmgkt1ls4t2Y+2ZKHMNZDEMHAe9dXm8sCMu58BRONF8L5XUTcuDYy9o8
yfzKzmouRscDHZDkF2HDbIzmbgspYh4iSMYZgjkfHvdB3rsf36leX9kycwKvmgMlucKYcFwtevJE
hYcDuXUrJ+3Uaek15ZtdMacd2AJjYnvCbbFtnC9B77p54URl9zHIFzNn3Gs7iHN2uanjQbrFF/mn
4sMfVz0kIxcoILANpN+WCNud3oVVd5W8Ax+Kr0OipLsMj6GpkXixKg/4z/Jow08vPVgBpnQq/YX+
Xf770T0zQN9kdCP8FqT6a37Zvz7pcj8dHlj7OFE7wdSxRaTQue9ATplOus6WO4m6/aZ5dDFXrOgH
tQczsCkyBGwJ30PQe0au4vxjGxJYpAxWgqtr1mxIzQfElswxZ8beKxlixAcizugp4cXlGQeCkjyN
/tX6Ih3SP9GlWgtRxZRUKxfbwvBbNhsfsLOhG+/KneDQ8sGiwiT0/rL9yewuCjybxzXlezCLFw8c
Lc93CJqReGPpgjuYKPJDpyqfY9ha5bmYhgyel117pqaZmkuDmUz+AS8xUlHtQdzd/ScfYCX+YdSv
ouhrSuHoTX4yXKLPrfEIUVxEsnySkJRh8jVka6aIXrB+igICDHH2u0X5aWf8XGHDwpMQ078cJt13
tK3BvNVTF+tiUKU3V347xChOl+lYnIWrrDiGRj6Qi+mM54hLbMCYSlK0A148SOXq/mpbJmxcQpfJ
pC2q7nXmRUfe9hlGekNtx1jC57OzwemE4iiJBbyoYHbiMKLOZIJz2qn5mPT0rFiTqHj04jD8UMR2
rFlSH6/ZGng8VB6Nt0bwtjbBDvYsHuEw5Xx/PyulTYi8JXH08Un/Pj3bkgeqQXfiSmxU43wrpHJN
EMm1UtnITq/X1kLNpXkIejFU1zupfuQswd/P43dA9TzzZttRVGzMoBGbhaqlt9j4pCgi4syg/1o6
bW4ln0V9GLNnxyvSmC3nuqmEgk1ZckqyqkJtdN2jz1YSfg+sFgCTS25fAbawNVoFShywwhu2DeZi
gd5TvHTHHg5XM7j4u52UfU4paX+HWJzhCB4/fa4dlW7aASVRsUaQcDJWEHQ6cB6jqpvFFsY19pXI
RZP242yeOfbaVPA38vauVgnwlAjiPZLUR8Eythmn9/omcnchJ/5xAZJoXM6NGB7FrSKEG2+fk0L4
r1IfQQz+V2ZfQJ+YXo5Cgz5fqw3RGVe+N9l7/yLt9hcD8oWJmTNd040ANC71ZDimGSUCUkznLso2
6leZ5HjoQt4uJPJpqObMzakeQgVCv+u2t/ORt3n8dLLnMj2oBDdZDv06WYoFUj3nmZkrNxc2e5Gf
qCgYuXZmtPDUThI7lPVe3MR3iqF9JSymZOwEL/MdM6PH6cw99b7+ntnoiBJQaT1dlsQPV4hb/AUb
luarNILKRc8DNP4SY4gWYy9j42ONYbLqupBPatSvqpDw1WDhwW9vTD1oQfJUs1cDOxn4EFwDJFC5
XrRAfqnlGFrV7vf/+nlD0m2EgNPCLCfRQr7ekO7npisUN/g5vtnFCIYM9KtNneWmuPNpqpWwWWe2
4ZwaCP9HDmcDeg8Z6XoJSeBhIz/bVi/S6opmub6UYR1uzWuk5top02Up8my9fJVc4Q2czgiu5mGo
RrNdwnGHWfvkbEQFlRk5VNF+XrHr6ae6xQf2XEDxodoT9ZkInNPM0YNEqM7sCUsBklPzKSxIqOLy
oBKHlxLITHU8U/rm0vUA8CXt+1Da1OcAvqpItepY9tEGCB2Oizbp7+BvMA2zWnEFsZxL+G5QWa5V
i8RL5X9xttKYolVBg+W5h8sxItQE94fpEzt8VrHItE1b5jPQqDiSozwrjE1MvLlfJGEYXysCM8+I
BQKnk96llJ9yNetCRSexpja2SeO7Dx1sioa8SvO5Wp17ZX/JlZAIspkDEb9HuZ0caDKe0gwRtqFI
alTMe0c/57lg8yuTi9lhmhceSyjEdydYtvD7mK6lFg4Tu8g8P/QZMbRulIf74gPuTB2EEZfXKRjr
aDTJvKRCQPw6zinxN43RgQZtQ5zpv+g/2FEFbYHFaEVAnWUNG4JPzfVWF7Ct1p5SZfFnxuwDWWMT
Hxtm00AkqDQHlh2+vDc2odMXa0gJQwYlC7QIFpLjtHe3GD+ROuFNWL6+ELjWqJsv5/+fK/B2hJbC
L9j5dm5Q2KQ+beRHKQzSzTJ1IyIVzXb+MN/bFEuXPHhMFMOXGXEye0INkWVhC+URvZRPSb+FPUNM
zrjedp/m4dqeqPzGZumsbb5e3cYnEhv53LTPIzaamLaJmuNQSCg7yQRCBcwsyG2RTvlhWfQ1L5R8
rmmNZ/9tiBD2ABcxT0tFl6si1Gp8kwitZPV33cRlgpYVROGC9VmcvGSQjFFGb4fb+axeTw8L3EgC
I4aJuaRBBxy8mFBgdSZsHHLw64NDj+isbsXNQxMzvsq9qPzHoNzOb6/Ut9o7LSgUgAX9cPblvMLl
lqvYgFID1OdhpniF1vG68oxdr6UbwBZ0qvC26coURljzH8qAAfDCyrkOCAFny1xRZ8ZL9GQVdM/m
81JiD4Rg8enSwq8tJOUo/xdBR1TizdEYOsUO5rrYNOfKl0GZKkbZi90/x6NyqDJxuWvK2xJus402
8TG9CluULbphQt1IzBFFJIv1e1Q1FBTy9gJhFR8bm2udCJ6N8vWwfmpA8ByFwUpT+62o8kBi2mxL
NEyK5UVqMkyXl88KWi/b3jel1B1q9rVpcq7hDIW3BHuwqsaIFhad9zo3m9P+rFEJncuuiLsYxxmX
apBCY+EFc72sbLcx75sdYplO7/QCO7dBSmpo8zlQNegf604+OYBpGKh9otrd15w80hqCSbaW95T6
av8QMot0jQcSj4DZxbe1eI5tAaXZRavOLEmRit3E8xPbhVfOiCFtexbMKrcq/2AsxnFelmxTH9py
nxDyswm8GUmWICLm8kiDAax4g6c7I52rtTO6OYKM26JcbA9TpFdXyqKvSQuPykwqjSgx5OiLeaxG
fyL58HuIxXFrsOIvygDTl6tHeUTzB2ekm4tTKQshPNM4ZjaGahiZoG8WqJEAmtQI3hGg1tNucuTS
SeEpL+LOauC0j5K0oIQMPAkcfL0fUGGpKQTFTr5VtIm21WTFFMiYhfyomvgkLASe+O3nfuNp0oyq
VilGIWukMsXADTq1VfB0CKugh0BrH2Cho8wytm0NJV6NhnG8d/VGTIJmjmEeCZmm2iasiIF6E1GK
+GR3W18Ctq0IygTXS/nUinxvMK4nrBTc5rkIaD+H9V0zwzDwL+bcCREMVaV6VUgSfhmHTEMhzico
IgmVGmJkKrmKpfGxyv4ga0aVcHcfk/5wF/ZvRCSr1KY8sdySxHGxe2hfWgrATuYXajLTrIL176XP
8hgsl8eOU9YsBYF/quOXiqWqJij4NUkNye76p+hYYb8pL9kzMAuOkTAYCAe87zsgPngchXNxz7AJ
0ZRIh3M8LK3FFw61a4iBzOHNmdIAwuz1tgWEXaylZpnazixBCvn6lxuPOJG1U8i47JhxQKz71Oho
v26WOt/DK00MlrZ+RRagR1KO3RTbE4g02yBWAZZxVq7P83nxfK18n4vhg7ZK1/Lkx24edlmMzSB/
wwKaDGmXIUMQCifW6mzAB+0WwpKebG3m9wIcRnlYmz02QhJxikfSLf9z8jRuThroXn56sE4wmYAZ
gmx9bPPZ5MvyXafAyEZ7mgMYZRw5nfjbqt3r9EUivN4RRM2cwkWFzn9yywyNlFgiKtHWUb1tEU/t
VHdZsLyGaYfjrYX7VKc1zzOES+u9l5bSvqKOhuezpOpM7TOfJWXI+1ciuAbJgFwPAwNrxKizErOz
RHUWnXM3Z4RXqUwQRyLOovQqAu0FV0L7SsjFDbveIuU0Z7OvXsQgcBnNFG6IAksqyc2RfJ6SoWWR
UCApHYGlhUwtyrRWmxI70rMpfaCYLZK6uEq+4/6L+CqTBwWusZyupAsjKJQnkiQ2nX/W3g6wOmGy
HbP5kinHKYRZjm9pYytCaSUCOeAbdmEEUgGHqRwl3Eh9mYRwj5v6MAOZcsIeIYlcguZEbrmKNOz5
3ai1zB5iVoLIQubvtweyGVY6R3pA2pDA0HJ1ZmwCf+HwsTvuz7eyNeXUNTm7OVW6cVlY7vFnGr4e
fCoTSZOLJNWCcZS3BmDb0hkc9DUYvvr9we2xv1wUwJGfxftw4/o1YsqBRdbzaLg9rg/UQqQ8H+oL
8hrMe8HhxZQfNngs4ddrVW6ZalG9f/PUw+1u/PpTKIddHw+WjV8vEHEvQK/3LvXsxrSzkOclutx+
i6YQcgqeUEf+Uw5QJqjX4j1dH76KOdnKeWPVtlXuLwVr93oOtTmah3h7e8QODYrWouIJZ0M6Cxdj
MmxnLpQ7U9ikFVjh1uKTXiqc6TFtLf/4x2Yey6DWeqvsT9Cb8GwjKoXfVbAt9WogMW6MWUsmN6AG
8wUpSSnN2W2vVbU1U3ESLqa4lpT4arPMg/DCByXcisP+cAPafrK2LTm1uZoRWShy2O/2HAmQ+fn9
4Ys+Px6uUuNB26TgYJhhElQTQYnNpAdgrP3Ot7vphEbRzbCFIkltlTZ3WSZ/BEAWXhRMtHDxLJ1B
itjwyxJgyp16/8Cc1vFbItT6DVp+u8cL2jbfy4QrlDzCP68hPsG9sZCFORVGPsGtf+bmmKpaiOSL
Rqne0E/gHCrGJjMdila5jQUSrYI4b57kXFqmAquW2iGarICWQEznkan6Mt9fQ7Jk7tbdJn5PBwhf
3zU2MnEB/ZX3mAk3B4Wj5rB7PTOZ0Di37Xf2myLTWwJzuIwznC6Fg1oLKjXGDS3jmriYOPKYmqJH
jWxk6hV9F81EzrsQr5mHu3o8JZ8oO1jsOztn7y3UdejEiFa9fgwEelP0/T8rlakdEcc6r6NwbNhv
IRlZX/3abPoya21qn5q0iJVYv1zs5lzJ3y8CQj+0ONhc+QV4naGVSL6fJUfJBxclZMdEhPmqQz+2
x/4+zYKIDdl3wHbeQAIOQdpc6EG7roT3NTPbr3h9hVCQ89ch/I36otHjpZbUT75vmjMvVs4XU8T2
tVwxtZepGL1xThhkVkhCgY2KCifziE7aw0vZMdHAAQpBAjfz+jSCT5ihxBVdEkrBs0qWBEi3LsPm
C+1U7iUIeVW/pRn/Q2oAL8Y0f2iWCM/8aljyUclSwGoofjjckpaB2wfd4sc3JqxpcOyODwqQ2xYJ
z16G2AH39oKWRn51udo0UJSFKDBpqp83Uoh0/MJjL/qtDwTw4wq4cLsgMkPEiXg2hBJ5sy86nKmF
wWJ2VRDkNNg1yX6zYgPO6n8Xwo+84TEAd+QymVA8o/r84P9vK7jI06sNq36ik3fsBC2vSZ6EKdvX
P1F29e25gCxLW3JI9uKy1VuB2C2ik9xkaig0WcJbjCptkme+iAQAPq1FSm0yTrf1Ciknls0t4wxq
3Yw6QhbUnMSiWEEsXLUJWlrKt6VLmak++srQbV/kI4+Jp5XejDIsM60yFHIZffn2Crs/+aMJ2dO0
URhW+c9vDYAgOP3eXKRHfhEtO3MvBN+jy9p5lhpporlUA7e2fPcgG3tZYfZUyVrv2lLvxYZVFZ9K
zkKHSpjesJ487fOqEWJkX/o/ETuZrNJIMOk7q4hLEUL+sYYRCKWgD09d8SPMIyoPGKfiyKPkpHPo
+Ueyzc8+abyVSJBiV8VIfJ90a4ycdCOS6uMaPfzIR1oX0t+vsLkrbx543QOWpLnednV8/EN/sSsB
c9KGt9zGnCHIAX1nbinknwvQPIU3fAMNkEslAiLQjYHwBhRma+LQfe19W68C2BQ5ntdqfmMc8t/A
O/GrENIeNO5Doxt4ksiTyNNOrG9/9bo6WYgz+NAoFeuz/reH63FNsGwc29bSNk/9EnRNbNYBXz3r
17lWmA/jtHHzplTY87RfT4rl7gujTp/l45trRltprhiItG6Is53Y2+1L8xiaWec8biwInYfGbjx/
WbNxYcf3owqwf6vYgS+0zym4bzYLkJ0n4vW41u6eeZoCrvBwKinTexqFPf1yZtdoEpnVu5bryfA2
TSP/7w64MlHJ9cqzNTn6R0ZIOnm+4KHXXaDagD849uo/jFW2QHY5nDvFIm4GJnAFgTSPg9hg95/L
7q8H7GNNtCtZ5xrc/zDVm2necEs3rYuOglZ8IRQKySVeDyyle2jPUDJcnF2R2J0jCe74Pi6teOZ3
5oAzvAn3Uivc9gUPP7VgBsDVOFmy/cNyQlKzlDBU5e22PPa1UtdRQB4ZgaUjyobYXW1MJT+0MgT/
EccQIvxGBfyf73b6KY+MjwhPNDgOqPHyNer+22wThKEfj1k7dI721vyvyZS7LvSB67TimRhZyE6x
7m2OjD1xQh1Cs1i0JC4yzUUPzK7VKqL22aHyFrBTBu/bask6/ioprlq0Fnwa0cFuwNDEam2CwgeV
x4GegQS7szWOJR4huTDhNrGO6tihkSfLAns1lsXiRBjRvKZf+v+3ANG3GV/HdyvOEtIvUsf8/n9s
sbAulMRchRKfIm45Q58IbA/6lHtXd2J7ozt2nd51h27SUJ1Sy1SVERrMEIx+fTQ68EKn9xwAWaZo
DGUxyaClxhnOIx5fmttcQC9YLoZqabzCKGZXXrMOh7dBhES5uKrwP0tGzkYdOXK7pEZr2D1HM9h8
X+KgCqhZyWE5z1CdBT9Rlz4AR4EpfDrgV466ZDNb9KyuQhvSQLSwPYtyXzCOE4qfS5Sbj6HFkp4Z
2YqPzIdx/3PTK7faKNnXwbGcGYufptnYz+YcvNreqAIHx6bkvutc3r/37iPes+7ORfm4EewEkoiu
GNdMEXNsGYlzUcJBEVDVxb/nzvYvCAHkp9k7T4ggeSsxc0MBStb05sSWy7OfBA8yP0Q4kbBT1xpO
Bz2akGWEI0Ksua7W5XEx0ORZuEkWxRTSRrOhm2rQs+RsIb9GDVCsETuSmPeHqlMYUv4nKRT4S6Cp
lRyT8/FU9S7LM23BbQ8jHrylgYktRELHVpwUKirdUH0zNVBHttO8NIDBiPOxGtKqm9eet98MU41c
yqJGtdgo7/uslOadEREzmwvCKKGJbIjmQ+1xyRzPL7ujbc0R2VI97lNQEPtdJaLXC8jHvJnazywG
1F3NkJkxczsSc3W1tNMZhmJ9WbLQ4MqSpDYrRUH0nKjhaSVU+espA4DxuNcnVSSvPYd76Rw2enLn
oVbjyDgx5+zYDb7S2fVc6Yjhq5wf7LCK9ExlKeshhzkUXH8ci42pGopJEJJRbml86ByEHQ47voQa
4JGRi/va+H6bcoPlX6C9UIgMzP+hTY8VQhxEeE/2UfsGNq+v8JkchDH+3gmVnfYAXpuTHJbtpzZp
k42s2anD0+9WyGPSUlTzFQhFuDvbWZRRiiLu3yjchoyrWhaUh4TV+w7FrRMaUjJY+xxWDZ6oLwud
N+H19uUCNFC4fjXLL1wi5ooX0qWtl8SlbgF9HhLuVuenwTp8b4/uOEYqdVw7WoZuXt+dhoHYz3bF
xpBUS9wiBf8ixEKWHvWDNwKGwPcbcxJw4WIxSNNyL5I3PKrFDNLvFh7QtN/yjCk3XVyLdMy8KJrE
QedleDr/SUQUaPVJ6mlNSiVJunOjzkTwyvwTuaMvyeQ8YNcdV6j7DdpY48nDkenDXoZAgq6/t5l3
0Y8vhfGvDf8CDDHdlwxMnKRzH85boLqNnNw53/ZUz7GDEiqP/ooz51XB7ppkewlwVTzFg8Ax3J6A
JJTEsEKa1JQA8d/6gUVn5B/HIwAjLORx6A68c3ynR1O89pAXDjs5wv6pE4ZY9HqNw8zsG2YhKmJE
X7w5LAznOiAws2ebJ0SLettIVc2OeoikZdEDwBOLp89MXzn/yhCheSzkaYkqbb4zw0ZXwa7ysMSc
gla/zYerThkQqynKkKxluk34rwmgew+3rmSE9/pamsvRSJROpfNqlMgayBMurafYu2mZqwwoB5wy
x5IivzOM9eM/NPduvpv88dRV/McxuUKeJUH1uHj9RMo4zgA3dXGGG9x+npmUR2v+VMARnnTUWHBE
IO5AiVFe8O8TMh1Hly1/qfBLn8IVOgILa3UmSFv5BEj4x8HM4WkaWOsRMjEhHfh8ElemroLORXrB
9LrORCv23gkpyh2GkWKOYh9wL4gDam4mx9KSJ42HQioiD1ATsCOIqw/16qj0ukVCBNPO9oyNjII1
elu/6z61f5RR7SoN8tEsCO063qHASsC8800umdL3LdHenCzy0iChu5RXjAMS9wYx+HlfSFQBzcIR
guY3dfmuKoKKfc84eaWjcrKSVoedhmYZk3NnWZAgED0MqyN6EWNs+WOFUBEBoN1hzYL/GEVHpcYN
01OR+IEFrZKWyOBPUQEgAdDIJcyB/GRGbCheee7nRmae9djJlSaUFg2Fapokuj43qi/Vc1FKbKix
223s7Tws0FrmQlaS4P6ZS0anqJtiaxOGfGd8gxKt5YXQR5KrZd67lK/KPFEoNaa1lithXWmksiFH
J3UqrsmF1az6uWOLhNUmJ+yzKiq0qK95tznhmDCT84EQqNBOz7+97cqcq1RLkl+i5tbXZPpWdRdw
mRoWgjGR2pjHtzOqyOxwtsFEgsMN9XiPoer3wM+twvFnDAYZrEHFgtsAkL+4hRgdL7PEdGiOXkJG
FtaqQ3iwxTK/RIjh3+A+tF0CosEbiIdJohpi7E7oL9uqLRoH7hO/9y85qOvq44U1EU2AmaaPcI6j
Hy0nrkzYrIaQzF1AF4rGnb4dFXvmvreI/e1AyPVIcXtlNPDq799VgQo4qa70v2m4cW1+Guqm6/eP
3hMDGIXOWRBE6Kxji/nnUF2NRmT95Mp3avqL+gGlnKv4TtJhjSXwMzV742VC7+qa9uqIsyPYNKtf
VaCFQ4pF0EmwSY/BJpU1PTCH9h2Tfq9WRrzVKEhRYTzM61qpCUKQROyW9WBquIzgOnb3+7XCGWeu
PRTn0vSu3g1AlHDwACst0dRYYqJhIRj/vNWwii41DVNTJUoeobHVWlpe77wOcy2v5VTpwdAuKhAe
+LpiQGqYGv8nV9xLJo3D/PhukmDneNON5siHtVEUSJp8CJ4dRmj5aeSHrrgkWCDFb+U97P90NquZ
M76ZVYATfuLtqmRc5TqWhok2n7IXJe49QU+1kgzBkG2AmqT39SZKotL24ylbetntQzNKaENwhhzb
CWhuJAHEu8GHViCCqLYgtufo76gi4GQkaM0xbvDDOhVVY5q1fShuJ+PT63YPeDk2ZJq237vvS1EP
i1xFHFxj3YZeStJjFGhbt9bii1ZHegcs0WfisH6S4jnpIYm6aCvZ39PNHvfS5XvJoh4caxXCNILt
hwm6n9hR9ayRcj5AMsuqn0bTZVMsCF/MZzuzrWdcF3dI9tqHJHXceFW2s6DGBIvUVfdkHApxQUCQ
rDH52OG9E8D0Rrkx0BCx4jBktlZNUqEhGjq9TdkxUoB5L+7PPIRfJl15a1d2Ip57pcESEGqLzN/W
lj9IWXeoEWF8P0O1j/qr51tKGBedfV4PnQYLVPU6vtmH7JFNt8PQyM+esjv80JsQBt6VOYW9G9hE
pCJgzywPI2OwAzZKzasGl/fbJss9MSPGqchNsoklO9Dxse8S8Jy/ruTMz7E85+QbI/YJsTxz2UVw
B9nqJJzNkmchBPuHBLBKwV/Pl0RvIU4odl+nWi7XzvlMiIYtgdGXZxPEsmUXIRvKSSLVuKl7adu8
a+vPM2oXD+3MlHrgCJLBuhhNn5b8qtusOkdpXg1enO6XLZEDUuKdWprZPbs9UnvFHdiBhs1e/TiC
KSNi0Xskw7jBMB5buf42V6PuDTXGZa0WzUNN1C7anwdi42ZC+lbeG+EXt5max8n/lKw5UZsYus8m
1AYU1lD5g6EK8dd4yFVsQKSxmFh5noUMHoTzODAjLqiAmLeJnkLnWvYPWZ3xTVqKetviF0v/mvNq
SPO3El4/l/HA5WAKhJFCb0/BPUDENXYsAHco9jZMp5hKziKmdmHn2HB1yVcPQFMK+JJSp1R+/btk
2S+tb2Gap1u+8AUK6mbtkXT3gMqAczEMCbrYVHmqSlBk3w+f20CdTAIJWZxZ5dhid67IBpKD+vJv
l8cmqj654kYehcIQeXKzsrKQ0EsdTqG4upKbMK1hfqjAk80jXf+l2z4j/KHM5TxFVTrLCzdlCo0A
jcRemWWsjhZuzXcfi8W7XKmVTtojTzrTlfXijTisum72jLiAMCLbkJ/Sl+LKlVa3OCqgPSNqBrzf
LNbwuKzL/cAeZNEKhzwJ+te6OBvx+dnkYDXrvYVls6UOLaYhDxxXG5AuLu/yzSi5Yr2CX2IWSCdg
N8l6/leitnqFsUIoE3BaOUbUM6GTv1F8nc4iwjQZlty4CkGeEZAn2YE7gMVlUzAwIEn+lvPDWQrE
HdynSt1FAq9yMWxTxFcDfMaM7+tNnuwuRz6xQaTI4+G/mFSdS2DM8nrsJVk4FrtGXW/DGyfbcl+y
FquE1skRnYNkByNqk5GGLjXC+1CQS2aT3ydWDaMgxGi8EBZMBu5fy3EbXIpvAA1KTPryoWIKQEBy
iEPZ1aEfchdFIo4FIcQtVGEhVKXmCppsdCEISnclj5A6bSD9YKmTsTTSZaOQ+OACctjRQg3XnKQc
NL9n/v+VAGIUXtaBAH+fecKQXTl19v2f7yArGAP47g6Evw==
%%% protect end_protected
