%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
U9ENgEHmBPqpgAIDjRgax3vctt4T8uLiYTltXHF9Y9UxBx1Cyv/l6mukyj8D1RajFOgNEEXiIW4V
1GBD++F7YfYVOmVGBURULrtcOHsU00Stw+nEj6IJPZIONHEPpy/mT/1oJsfk6+xao9vXeDNUMs3/
4bBoyx5+meZQNJ/ZBb+KjMwwcd6p6WFgf4Lor4VxBK2+VIvoY/M0dFwH6QZlu6PzTqAkkVDfHm2W
kZfEEqoWsu/LHMZ5/OrILBG6o2XpMSjdcj4z2zSvDYLUaIy3aUCdQecF5gw3wF94PZo74/73hDhO
6vWk6X3ByNtcj0lFhDhyPXgiEUAamzg1Zt76kw==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
0CF8RG1FBKGkYDodC5jIIwVCGKz8Ru/3LZ/ulR3WlIiF4lyDTBol8HBEUrkWswBs8BRhUcfT16YX
kdZoZ4KXh+3+pZiX9qfh/KGMN1Y4zIHgXxU5nopLwfF7Bh/F9hK6AqPjlsPo6qucEf2Bc14jB139
pl5sP7A9f2UN2C6D4J5m2OzbzFxkBDBfKMQ58HUfIpHtwu+PN2tZkhQRgMXc31fnZdyMjtgcBk69
8iXV/7Errw9Bk5nwLkWj5i8ddcDD98JBk5kYG40yiKvPmdTUufjCz0a9Db1KkTEDibKU7Sqm5ebm
wFYQjjjBE3iDK1YmoPeML42VV6KROy05wgDdUgdj+pq1Yb86vzzOEYuuHokVJUCaFsrQaWfNGgZv
TTOP5+pbrdUf+nwy0pd6alwKvh4F+Atn1uhuSCMcyaLLBlFYWk1z6nwl93416nyVBYa+RnDq6H4C
JS7sXML0vQ+49fnqNDVGADScz/3rZOZUTKJln+idrolX/hnSkKbfjNFNjWhLrN+2mcE3MMkoOS0S
elC9v9BetK9ZyBnRePJj23UwbdSxawMxefEO5ynNKOS+5pScCUiUfvSC5XucHhuYpU898VWU48TH
et2aJ4crI36xhOlmNHWf1Evxq9QbW5sNngwdC5m21RKJejb7kx8a0QoYKWKdnRfCx2LpCDkiTRJc
wQ6jm9iAednBnzc0BQJu99dh6QYI/gSZM181pN4HwDuscJe6Y5nOwKB0M5sXelCRjrv3iyaDecUL
HxbFIk70Acd0tse/xm5Y8zJ986H9A/JUg1hT8WSimYyLYT7+/wf+I1S/eBvt1IOOhcg+Ha78XeVQ
vTU/BAIx/BgScLYqViPwq+FrtfrkRzb0pUNCd1T8PS9iDFs0agEnzk5NSy34RLRwA+8oKWeqRZ3L
7jw7AZdwlEgiMD3uwUINbdFtgEI9ymeC0ZIdWMiJUD658Mt4tjlHuvmOVzfoCj/P1rY4mOTaS4Qk
nHb6Ep0Fe7ec58QLwncbKYm6LdW++jtWVbo+SAWxl9NyPoIcs8i2RSZWbJrkLEbx15Vrv7TTxGCj
fFX5RUMa/4p2TZCsgz0kPqVsQlRP7VVDCGThBVSTCf5Rl7z4akrQ09nvNb5U8oC44KyGES6I8rGY
6aXEnDJDbJK0L+WheqCj8aHtR7mnG5LNlqCFoQ/tR29vFVMBDZSjvAktA9t8wKKpIVdqjlAwPd3n
S9cPj6L5PMOus1T6M8kZ0c0iRHvOiBDdu3LyOf57Bf0SyLb1Xj9PYuHWmawvd93ryC9owmJiDGV2
sHgyH1/eZ34KJaoLFAw5w8razQMzdDLQ8iqKQ8NO8cIBIQwO4e2jaFgdImbHCrhQ1u0pZnh96v+q
THzxXcmwcxq5deIA892DJ41P0JtDvA9BZ2Wa9Npr0KfjDq3LSh0AU/JdTcr2pod6LZDpvGkiAnIa
1MQWTNRjst/Xj/Nkc/2UWymJpsL9aBY+qe95jRKdEn4SADNpjqLCLGGMN0wZpMtfikjfeLb2KMuC
L5r8bVvJ8h36bs1Vvrf+uEhw/J0lPm8rcGkkql2KNorcjP/bg/5tGSSNn6EWYkisWM1XT1wuhl0Z
tICdLMYE/jGIrwmb1gMMzv5YjaQeXbIrmfxypiHmw0MmWW8S4qVln2oU9uu35Zvknf4hIzMIiUob
imqU0LDtRyFipnHvc7u5lLK7u1ml2B2g7a4qBirrV/tfJV8CSYpkbcZyHqGgwSxOAVn5WwN8le+R
0/ifJV3PU1Y9Z3b6zzUAkNB+jMeTZtWQqYV/nuQeHNYppkMTK/V+B0rGkHTU56PLQfEWhKMC281k
376Q7zQ/8u7YtOszeXDxGbw1G9q1UWdvvtGYY6V06KYar9wAFexC1tCWm5L6fv+2lBG59fcoV3Y+
Tw5Y37Fe8ZN8DvH1NiGU0Zatd9uH8mBlKGHtgFCqvcyyKpLyEOrjREvkHOMSnhx6JVasiCXJfk8E
LF8kl1NvwFRZeaFvalkgS83mBafrVoPGlx0GsICDFtPPFKo7sREr37SjWqeJAVN2UXLGCJKLCf2C
h8X4FLOoe/7Y33V+H0YjcG0uttw5zkTLuQXIOoxG0Sch+V62EUpVZie0sqa2DV7MN/Ebqq4ZWQzs
r63rM1dZ0N2ef9dU1o4+7nQ7vVSkN+MiTC/bLuTq1b7oPuSrUCNgMTbTtczlMboDv6VgBtRkwFma
9slvUALXTofChl1wRATj1rw+PUjiA9sYq7y1r4w3HqvK7HCh/aWbSC6sLZyRzRSnmqcYDkFDRTdp
rokRjRPqQzQfsiFsM0nuh/F/h58qz5tq3mqBplmIXGSuR5IGVPIQWuomwzg+f+0Epl/PK3ANa0XX
kQCAIt9yD0kaTrdu6WzqIn1nJu9WBF6yL/XL4Uek6sXo6/TNVEE296bNyG74AJJPG9O2E9mykmfH
v4xFV1bR+5SzLh9hzYpHBLAgZzBMYLiHnT1LDGdKmsma9vV4jAqFSKLaRW/oHfnIUwCSvA3lO4t6
MkwibTahGVYGJTrPIJSV6zOV4pPHCxhfcwvFmqUVg6a5XYUQtE74cRUC03KPOH5Hsalw4SRsLM2c
jJF6/SlpzelihgR2m5rvwAveAxeU9lcqMkQejqZL+fXfBdXj8creZRYYod8JmPlb8c/nAOi7eivZ
UUM6OzXtju/s7okUWTFbhFo6GCnScg+VhqZaCB2OqYfaHBBOdMKdhr+ibWn6ZDDFJcY8TleP9juK
v2+K2S+eVUpBnH7UL1vB8L0G45GzP1BLIPK6XwT8UGLyU29f7QvRgix3jE+mTVw5w3+056GTLMwn
/9kBCkK2kg+X14je2IWfr4MMV9nReIXQE0jbKDN6iAt+gSP3CIPE7p/VL6QdeLH3kiaOY1Or7hxs
htP+WQdfsN/2OD8H78FkGs4aG+GukS7L3s2cxUWdgHlcE2OZ64rzDYVv3DJCQZ3H3P7yYHhYuC+o
QlZud/qu3ubBJ8NmvnUmgRKaXA1QM1aoqlIcig4nSu1s//ABTKfVRbjs57VDNPgWGYTq3gPWwOlm
9R5q5P6KJKk9uuZsURRYPjFILOytxBrZRFDl5aE7A7ia7j9VxdqOytPTe9Qx+XFaCHkuUdwQupUi
kKyMTHm1DCkN2VghGgdN3vC19tEg6INUFvLwRAgke+nLWazn/MBUt2WuEiL5bovo8AxeSMDSAy/B
xK8Se+XHllfXvmjkW2ZvcrAaOTzz44ivq7Cig4+JNypwdM0hMn7XA5w9Ed/DczDaVJLK85V+poY1
xUJPmmLLxQI9R3xEPmeqG/iaTr3oBOt87WtLDx7J3/U+8aMfXvrNob+2dws7zMr4NCgKNPmtmxOd
i8g2ngh5+FJQm5ZPoJAm0jupDxNfbzIKGmMSCoIR5mPvNLNC3xNL+Fl+g9PldEOAG4CRU3hePLFq
ucKvc48iktWSkoD3NnY8r3XeDec3Cz/RtHthq4zchlfi2z3T+zTRlj2bA72NHnZ7NzOT0+BlafaU
oRb5MkrmBGa4UZ86C9MA1VfIGTjKMRAyy153GyYHgMLsAF2cJJeXiwkdLtSY5uZDFUN0mXXBfj42
dpQTAgIbeJWN2DN4/qqVk8SOTxeWbqBNU1cL/SwtxB813y5P7jZTlZjz9vm5nOQntAZqCT1PcqtI
83AQf5s1g1C5JRpIMastSnit0zv2Groo9X4ySL2GCpDi52NqOszw1FsL1dx1WrRfIeX8jQA2NnWj
sQE6CYBHJrpPsXq54KUE3jEnzvheuJx05kgKtfx3/a5SU26wKAyS/jqbWn8kLuMdgCEeZLo2y7p9
BZHse9gXQMtzLcCkaojv3+iyWo6Jg36e2Xu3/D5rW2Q6cPk5aQT/wq0KSbFmB0bJkAuXHjGv2JIK
uBmY1pZfgc7x7FWEtDiCMLSAyWUMSkmllzpXEjbsoe/6BWRcclUHtNQqMf2GPsGjf251oVg9sm11
tsoD+I1wS9AdyCdyILLdxSxrVErjNr7/6/aTIg3STU/yAFXOLlfS0pf1faRVzcH/+L1f2+tykvEV
5FsjfnCP/pSMzxnRHoACsJhWCd+2P9PsG3ft8QasSvzBZAmBG0y3IuaQR/Azsms1mASXrPC64Lao
3sqLUoVl9O3LAadPAZxaJ9ydQuiDExiI2thOLeEsoCV+3TkOMstsP+dyOSwPVRw9+NJtoJLmDv1C
4Q9/p+GLLe2/E6+67qnKmirahfBxMBVkIcSf01oxWToRUW0dKV2H/ydd2xV/P3hIQmkEltVIUwmI
Ul/7qHvQs6YCyH5baqVc1mx/utgsdEL5m14OJt7gkC+4hLwJY8FrepSMOVs2h3fdsW+IzcnhKfH0
rNFMpVcAkHuHYH00hx8I1sX/7ZWfNBD9wiIHmlXuGcGXyqXT+e6jZZtvmwL8/bT2ZugnUW1vwdWm
pOiRz3x5AGKToei96FiDo2llbmRI2BUhcvJegwxQ4CZ42W6/xY08ew63T74hrl6aNlLuM/6Trh//
lrWUwiYUGGMS2wIWoYm91WO7Fux2RltZgj/Zs0qLRtEUeC1KoCFYGrbFU8aZPl4WtiMumCe9oLOr
lY1ddqGQgoaT04nGR8YUz8UZRnBqcklhcjT2y8AxQ8GdRZUTORhoqM5UMPplRIWyh8fg7cNboBlK
3wVEHik03zq3HPi99r9KG45qXYWhy1WQ3Z6PZPIOTXCstQBTJnSFxoHLlJzy8xDt1DgQ1v0j9y5v
y0N9eN2Mn18mwE+Ng8fQULipHCGAZmdQ3ID+pmPF1UtYurYnR7RgkfH4UVc3yN7NjemUYZRHks1V
gQ/R7/0n8UK/k+0tmzN868V9nNCTdePo8XIbGF38YGbXKrg+N4aLU2UXyJUrk39NCU6or6Cush1h
Qf1zd+Fo15rYeR9zzX39bdn6mJ4uVE92g8ZQ8GPZatsD28t22CrSg6H3JR5jIQKqWIrAU46rKtnC
nAGDRWaZXKN3q7/Vp6Ir6GrfQpBeum9w+i9CnDuXXt+OA3lD15Jo8h1EdHl+lDCbFlM//Sq6ciGo
3s9Avd8fKH53WQmX145XSGJhWtBYt3L4Ns09oG5HY+gukwjJCGYN98bGsfpHk6HyWqiINQJH9OMX
gNfcWqcESpaLjVOFZKSfdEgncX2jvHFwAue2quFMhtSdmpen9oR90kAZqc4dyXourkReSbBN2Dux
+Ej5c5/PH/QHW7EeaJjb381P7yBQEAMk1I+7xg6qE300dlYYr69X8i0d1ZmdOBUafnsSeRO9dRzV
Q7TKszy0Z2jJ/3wZofqwfEn5f/kCBaMpyfk6Cq/b4RJEB9HJIJUYueUFDcC0JjBLSoit+DfZ61j5
Dxd2WIGY2UeTjg7LNZECgdfoA1e8oHcpyVQKXx40KKsLLfvT9tW1tBJCHEw1PTSCXAFXXZkPIQzc
t1s3D9zZHxLtkJdd5Zw9lMQ0u2FXlVtNKKhVtaNZxY6o9Po4S788DnOCDJDfoPyN7VqwMPAmAobv
GuOol0ZwONmIG1yf1xiC0YQtS7hTnjfJKMq1qi6iuy2PcF7crTyA5VWlEV1x7+74hpL2wucexKS1
TyO1KRXQL/MLzlkw6LToJfVMi8+bf8CVRSdiif9iJDm0OLU/zw/Y3HQ2IpEcoklTmzFgOfnLUnb+
gnazvnHaxhmMSRKsQaABmH335LFPuV1z82aC4OsO+IXkKgpU/veLHw/mLqrTRZ7nxNqB7o69NYdK
VUvdc3FWWIbfMhf6l0WoJrC6j0d4qY04g0gJ2H1yNDjwOEakpY4ftkL8U/P76tYkQ0jQFtOnjGX1
wOTvhZhmOwd36yE4e4y+AuaKYdeSdQV+JQCtIFgXeoKQG0yZO/kFVtrl5TScZuVQRu6AWYGQG6GU
yWlND7VZ5hnzhEljLCvN0x0z2MJCoyos3je2C6+JHMZYyJkWhvC5SljJGcPSXOvB70sSZ4lS/f9Q
P9d64hOf3IJUHtykCcHTdmwr602ECpQt66IynR9gkKQot99ilLdAzHmu6A678/w4DkN1C/+NaBO8
KLyIyPKWMwOKdphq+yx52wOeF1lHfwnt2TxqNP+x9cbO/xNtoBMTVYujcF+G0D2tvWkkdwxWgdsy
fTcz0d24R9ZzKu1bdbo3SeCtr/IVZ/nBAXlX/twy1gSg1vzP8zba9EHWD+c+RKZ02cV+uIDSLcKy
/3CRFhm9MKMPHrU/XJkXkSo9lrOggdBmDf0tYf44W567PzRkY5/sRWkGBfNEyBEL1pvrW9cmnc++
zlduaUrKrKBQaxjrrCI+tMM5yfDJcDWL1IdrGFY/YDowTWrOdZXELE5OqDIxDNz5pt2L3XJZ8iBV
mxRejfSA/nJ4q9mVhMC3yGx6zaV208NZxKnDiQBPCHh9TSVeAgJyPcs490vNY4vdaZwZO752ySle
FCBmGTmovqU5PH4VkPjgTiPpPkgP+fuIeYcp+NYJTKFve4m75dmGnQ3ndGabe+CsOQGRqn7zaL73
xhTioKayMpbwW8Glr24QwBrUDhhC0WVgdCDqB0UnZnbt1YFuv/sVVs78nnQdPu4J7JX87ZXLQD0V
wBpwp7OhmgZ0hQTcDOLBJydSOCMSQm6laCOFnCKrQRHSaoF7vJFWh5vm+mrBxtspn0u/nh6ic5CP
pI8RmcJKRpxX1sPRN6LJHAHtE327H+Lpwxc/prgWPA8wY5H4S0Ur+JEPq/9S2MPzTaZsldnTUbOI
xIXTvJR2LdFyUpXnIBkqW6aumj57/650CzinQTAie9ubcIJdvGCLK0fWzXVy+2oELEaBQ7NOvNLX
c4dK1d1AP+yh37q5KjMK8An9wKg9OQgKzlHNL/06xGw3uNKbV9S6RTNO6KN7xuJRgqY/uNL1xNM9
ILOoiowqAn19ME3LWnw5V87qqyqMSCRv9r0YxcHFKX7z5vkPLQ/vZ/8xNSj0pGlQFXP4stQJUnji
WXd1qUcSGjZTysq39fi38a/rmJYKv29pvrxqmS7S0YLgLb41uyT5WK58cLhnFl7VLurE4g79/Dio
9qXyjqB5HJlU0S6y2CRPb7Yuakvxqb/c5Yc5albt40mrR5vK7XTPeuiVxAM7zjClZ5b5CsrI3Uak
41VDb7hgdLDzS0QL3F+Fr9UlZPjn3hB0D6zrUG2lk+q/xJFMms4JqVWlPbCivfGsiTrOygu2uzk1
EqjOSj4LwcHEI+mSLd8+0ArSPX25/G4dDPpg2SSGOaocJ+BbdMfSNh2XWKQCQL6IFM8s3rJ92hTm
iDuo1WNX09qPjC0Djnx49/Lx4BZ73HJQ8gY/KdHPARZTWjr+R/Iwkex5jEH5Cr+p8mQQ0ERyjtfx
NqwM1Ywtpb85SWhU6PVHbjAYAQWcMigQQguOQIAL54tK6w9RXaawIVjhuU4I9yWCTGGnzMGq1Eyw
ibTBHzI3pnZzh60MoCLiu9Tj9rBEn7YlcSaysJflTbsU5eDrGql6Q3TZ8ZZXQaLaESo4AS532cmt
7zekiYlOgqiMTc+OZnc0/rg2xNzfEdq3iwknPEu4ad5kHpl4JaUDsV1O1nWXagqJbWIqyy1BqZO4
s/iRlTmSG6ss7OqIorrY9nFlxaJOS7HBD7/a2Lul0jP3BizO7jd9Ed45o2CfoiKVVLMGSv1Mr5m5
hjz19esdCJKPq/T5F+S9WRJTZ/mNv82neGsvut8bAYehjWp0wpdAzENOFs0K3GkJRI30a9F70mPL
CmEmQ/uIryB0xjEQjjIvjWWQ+3+xT1IMFn76FvgXlmg17eAxW3t8h2HHadd1bKnYB67OfYPsX6Wq
ZvZ5gmlX/iqsG3rhe9l1oyvnVncng7EAZDAxg0JCTyUizuy+YRgfyH7ata4xMCKfT131fHsSkD3r
DawmdZV1+wYTDmdfgXho/ZoPR2+Kzspc9Rxa6yyOv3Ry1bERbR+uRPJ2pM73S6GWnUho9xaCgALR
hAx4Ajhm8Wp95GWCAj1JG/TXGEQf9gwUaiV6/xl7e4bmQ0anM0MBc8lB0ABCxd+5tdL50PgxVNmt
GWwopYobOhk77kC2gmtNWev462xMj43Re/WVI3/S4KGAbA6OE84EFbofwetx7FaBTdD3dx0HrdEp
JkwuWSj2xfI2yKaS6jur6eKKBAzXPxz3xpLjBydmPGzomUahTVzamWsXS5MGVP3PE72KpwuqBYK2
sp8UJGVoqW0qCv9cFpZZUU+36fp+MJCW+8nfbi1k5JQC8uAR8q7+HejV8ADEx2RzFjnwTYq44a3y
2hHXEVhNIt3UwcOAZYF2nJmUhW1ngmPbQl5UdqqwlM9ImZEO90dxsDBLeoWRXkaBf8IS1XP1GL/8
fXbQUoTUb+3mWmfrEhFOjpOtc4s8OTUCnAuNfPYtvOiyt6Ix5QepXN4QNJLQtRmualRjAl6L64yO
Bap51sjG/vzOj479iSZxo7DVEdU5DkY4EJg+zJtG0DcJy/ksVAxrfm+t2g/Eqa6qUJAYrwJ/EiGU
HUrHVY5g9Q/eYilFnWB2GQyiQ4EezdrvR2oaR+lM20rtKdUvItj/o6w+O6iirwyGuEKmeHBhqtGI
ErcGk4nzh8lEHq7RToN1uLw4R9b0woCop1xKFawVlJ54M3G6vMMlxKmbKt10d39DwDNbMcyWadx3
Yu9rNFgdsimKl4/es1u/i/l1wz3gfSx49hxOQNiJ2dwXO0FlUYAQrVXqcKxCoB7OjCn2bJRMDR3t
w2Lh629ZWFxCDEDksPEFcbdtj8LRqBadK8T59vVSV6JMRMYDw7eXCZMTGqIWJ1EXEOqLMu9xQEDe
EI6AmF8qviMNbt1OVpGxOJPQW+92DIVbO1QjD3N47uLDmnWm2MOltP4gNMHZqCNA2ipmdhkf8DPS
U173JHhqtAPu1fNeObUQeKVB+hgbnMTLMHBbA7nlTyH8xNR2QjUunw4T+vSMP/nj/tPkf/cbQH4x
FUN964Y3VCfjUYOgvMPie73ChDzVeocJPaP4Ad5k17Kw36tviGfnRD1pWSMYCYHjkHFm+jBh9Cw0
PYVulu04sAxS2ztsFTansnp2Ju/nQ4beqQxKpYWU2wpMHK50CG4kqEWuORisTE/aGoFNKAGF9OvX
gF3A0Qc5knJh+jyxfHLHodKKcabdkxKdFa5hGep0JIeTODBf0U3St8ywApnFB7nf/JQzNi1TKEv3
1TgG/Jn9qMs8e76TBNrAO/vP689DyUoQ8voHlW4hNc9BrhEa2fRaRfK4OvzTwBvZUNDolplH/o/M
A4xI2vF2sEQVkIcYq46tW1YY95fVaqrFnHqze5r1y4SuwoqDfGm3o+84lbwVqdmuoDGoJV0ryRCN
iCMYKVg+4X7Aol1TKy8Ptl35CrjM9ydj500HRecn0terrcveNX1C90b7rlijAo1+iCOhPJwbPAgj
VhieVoHRynuroob2VN2gNmSbyEwtRirfSx4f8aQLwCEdM9s0Ye6JbCPcI0irllx8N87S17Hvk8nk
lfaslV/6pefPd9VObdP/EElFKVAESAC9ExWl3IlniwrrB8Ewe/dE7ZBLpTCi4JtIhuW18xthu0c2
VdnV9r9M3DFDjLch2an/k3XSMJoYU98coHgiaLZ7wD+BgNbHaDRAjE4gedsrJnFxoFo7XGecOvDr
NIswnYxYI+Bw37IPe7YAvcW6VYHd1l71dFX9Dv2iCNwqrg5akOPiF5p/dOqDYIv8vJP67AdmT0QV
L6CTJJufAxzP2dWkKXJVk6IfY7qVC3B2MzPrCNVNEU6we3RfRt2JhEMM1hk5EFT8QNkCmEpvq/ty
jB1K4zTrj0KhjxdJTwbrzI9CGeWpz3WqPw4DseWAJKclT9yx2OKO2gyHqh+bmqem0TopoKO65tzd
BdX3uW7sMxSfZ4w4MK3ge53TjqS8hVvLPLcxkZ7WuxrhKmAWXRWtxOWuVwl2B5N4Q5E1BXG+T+2f
7axfwFLCBzKAaEmZCxk+lqGtX1xx3+HmJuThXQbaGhrozBadEEriLQaLsW4x0qutspmdh7pZy6NR
5zWgUp/xYDhc70cSefRvDQAzIRakrpt5Bn90GERWymkEqaHJP1c2EvJmTCv8GiLUnkHxwAbH/NfR
4wtEiM8nkS6I4xD5fGzZ18yCvCMg3mGOwelJNAv8w1UaA2RQR/pZ5ejRgZaYipHlnp0jcy94oW/m
zWhwTxd0srnKMMFsUzxljCmE/bhhHiBQ53Sq9J4dIejAcmBZwtzgmcvplfuS1pBH8mjKWOWq29YF
WpwmL40HW3FNou80BhmcWfece9EYmyoZBTNfaoL3GBcarMkLpgL83rWZcCtvOMjQt1D3PkNuRps6
aWRnYMO7H9C3NW3ubmK5KonS1InchL8DmDti35NuLzL0ZTPCQZbvFvvtoFLV9MCwZ1457l2d7lhN
c5ZvtEfauFSzCLqd4G5HvZpyiUI9o7esZwSVJFSH+dOdQIdRgXFdHDllkZdkD9/IwryVcHRykJ1/
GyYNKal1wNbsR8adXssEaXueP7HxTg18zaS0tLKHXfvvDlveW7mfo6LUjwBfT8lM4C20UMG8D2gk
E9AqC3AxPgEy8l3USpP9kBn1YQqIl+Fvv/SVcFoK/AB/4khhKbso7IqZ7GlI0IAxvLZaCQr2a6sq
+p0p6FNk9xvKFuamkKZyKlld+mIWfQnpAwoV6bG21c/6GP5QUEXYkU66Y1l3m48j1MnpmVKP/MP1
5HmlfA8cm2cQWJuJbmEm7Tsw87L65moYEXDbBgmSSLImFtI4tceQLWp+hGjP3gJOh5aIvvYkThqF
Us8wMJ4WJbBein5g9Zy5DZw2y6wUTSTQiFV+qDx//y5iKLN4PsFYAZ+HIF8rNhbCAljMdG+ZZoOo
jgRuVM5AB52QCsv63ZOKGthhYZTdxUJ7I6L5q0LJikPf/H0P/RWXkXl5igPD77DxgCBsyVjsT3FO
zSJW4ZcbixT2VS9l1Cpp3DN77CALGrQ3xVsPtjsZ8bsT15rJGp5z8oyMfsWMb8InB7xieWpKj4IJ
ZdIe9ALWxk3eRq2w5QuRxs5rV5NO/LefjePJ5lwdDrO/znFmhIkr4P7wf9hUYss+QzdO/28Oi7Mo
PmZgGc6FQoGHT8y72ErB0WWdk9zZ3fyEXh5gl8tgEdTnA2TBsw6Uw+l4CWPCRF76b66f084cTOSB
aE9p1pCoWcB8ClE95uN3Ln/VOtkcKAek12kurJeSeMaFxDKn+BD2C6YB8RgFDbxrkE1Kn9Poe2g3
X+7z26N4gg9W/35/z51GpZp4Qj7ztE1LFhnsR6+lo9PqMwloSYlj42sQ6XOSPrhxA5NQVFBANcGw
Sp+RCopKN4hXNDSXR+U+qhH+lH1tSZBzEXHAXhUmusSxl+zkNcBjZNr9C+l9zRuUmdfy23dyrRmT
fxLdt0hnxPBELkR+loG1XJ9bSnU/oYEJuMd1Er9SvKeOtn3vIPFQXhr/pD5qp5GMFvEvZyhPBW18
Az8+Auegk2M3Wxw5R3UMTYGUNP3YSM01s0h1yJJnpCTZ2yjSZkeElxDmOw25wRGAFXnsp4PMP76b
ZOUPcL0X4urrsMbgFrFdk3aa9dUbA8HiORurZBm5OBVn0NJ/fDQyuM+aKpcKHVS3nVXs2eIfsqYL
jodYuofEI+F/PHlwY+wy4rNz89xQ3Q8gyUTkLT0AhwZJB4asNwPdOw1Dx8dyo4Y1P2awB4qcaGT+
gzATNGn1PVZi5tY875HRwvQiU1izoUEGCQTIwpj2dQ/m5mA/XAMxgZeLxHTR7KEns/bzrsZGO/6Y
UMyrT8o/qa4EX7NMLaocfgCdyYhXADXbSRbl0wfx55aoBVe+HX8v6UWfF9fs12DVNX1UvBfLfWlY
/lcpJa/pHinOUkBSG+TlSnvzKLLNdYcdT1s/uCJdFTPN0FvOGgkkSsWuL1dxMoqgfYO5P9mOx2IO
/id9ckyCxfjhlEeRmbtfPIkHvjKB9DQ2fK/nsFySGtw6D3qgDzRfWW2O00nB5VwhH9xIY5t9WPlr
0Nux1hc7RHwp6DltQTpkKknF+GF9GRHhciQbp3T5QO9rjCCcjpW0cIWVBMmxxrWwM42YGoU60gKv
VZVn4VHzgR0ZYk3YAlrOLwt5adq10Kwzo63kZvS0tltQFtxXQT1W7+FkdJYbPq4kH6sVT/Iq5qaO
/lpXmDrRGjuKknBxVPff9/9mM4AUD9ZB3N3Mk3VhhUQncZafPwA0HBPiZknAXIzQw4a2Ez0l106u
2uHqeMR7lE8/nYsfaGput5r2+85AMlrkfqHtGvi8fjHF2LKUP6UIkCI1eXvLihfudm2+hI4c/l3k
9CKx1PkxgRmLh9sEz+4XltBHUzGTm3PLGyoeYnYVSyOxdptCxCzm6GP8bDpBr3ZMChu9HBf7wDTn
LCPVjHowfbalbBfWttyXBZgneTOzeRQ+hVHdqUOcGqkgPWzRM60WEqhr8Q/7D/r5Pv0mFgbee/I0
1SsbCUVERNtgOTbVJFSbYHT7DJbQqijpGj/UbJXe8yxHzwf75MrQ1KSrB6gfrRVtd58u0+rNM8gd
uPyaC0LS/u24wQkyuu2nxWALCZWnT5IEswH5+31ajCsSSOEC7lhDBSFEnZFyGjlcPWz8jiqYEr8M
n2lmhaidKlmvuUq560ZZeaZ9l/Ns7dElXW5bQTDv1sC1mvtwBapV47bbrDJUUIB0wgzzUxna2Bvu
IW4sBrSJex/RrqmPD2egptcFtLDSEIpuAZ86x+Wd4bb/MBFIb6Qn2XSPGBfKOOchf4D3/9z3tlKy
nprxlIF9taqHgqFOxwYTjWRMLRAFMYYwe03jVgm3PpZ3HdqaDoR7gwuIdZ9vlM/0xLtevJOH/6ek
XMmfbWk4F13+MCug9eEgZ8foUoDt6sew7Ie4+8tB94kakMlu2nr+ujrCR5U6mADOZZHCb8ptKVMB
IFPdVjOycnZPDUgTM1oCiq7t1CTQxcmf1K61H2TnnFbxaIU35cHZQ44cbkmfWNvgueh5FRAnKZr+
5nMrbLsIOiYGVWgP+lhXyHoxpbbF/Y4VWO/LYWC3JLi8oaXeROITU2qfZFH9HGLxMhqSA09mc9mQ
zFaQ82Iuvhjgkxgb66uSjir6sDL5LAurQb5AbRGOxzOvc/SxyAT0AMbcYvuB6BX7PPglcwU9Sgzq
3GXpcVmUWqItTCU6G8a97kBNZEItmdsXPIT+GH95nI0MHQVQD9LWLIjImrVia0wypdzJ5TeS91qw
fU3qYMlpcJP7l5vC4r7U8mcexVO52ykxbFFiOuF6Q8XmeFbNjIEPJdjtPGuNhf93Nh82FFKgr6sr
80qzHoHIUdpEWksKXkudeAJsMDDpnBXLBOlTq6oPq4cBN1Gn7GEhoNIxx9P2WZJvGPERt8kR+5R7
1wlo4sOVxgKAXjdVfcTibcEAGG2LRBOtP3yurd57aeMnNTma/dllYOIX8JjqiDtgL2U/5EOGFbAQ
wa2VQhkP5+jaGZn8KVR5Do88Orw75lxn1VUofbOZzR5mmTOmCAtTkFDG4RIknrVuCuHZ55T/19EK
nnda6b2JI0lBmEzKpOPjCSsAV8kicdaMspRI3xlxeQPL2eD88viG36qCfgfv01qsLLBymMaWkEi+
5k3D06MCmRLSi327okwM9CdL9YCpvrjJO36Xh5FsYBAXvtxX6SoMgQijGeyL+sGsN+Htj+EoP1DP
K5Zr7VVmz9PbYZHO86gr3c6Fk1ED0VdEwx1b1xgT3gDkI90ArfHRDnORZ34T9RGVs6APgHCkOPUu
hL9yJm73akWTKr3npSsgxSuGGDoNr3BCbQk77zrIXelRV8HC06jxH8Dqfo4GgsY3aXA//CaSAYJR
4cI42nf66qEitUpqCnjpkjNiP/YZQnVqV3lKm87Qoh0hYkgimnJfJWa6vVJXWJC3des3TlOz7b7y
07/M9D41y5dT3rxy7yYQMrA30fOEakoQV6ToMltEylcd2uZ9HFbSuyctjM/xHu+4rse6HYUTM2Kt
jHCzEV007mmynPGEkwlEPKBBVfTY6zNNsVLy9FiYIhaNs/o40xAWcky00+53Rt5GWB5wlJwjfPIs
a5sKZ0suwGOebvBYvFmgoSfVJSIPWlhQvNgNH3YGfR4FpaVaPGOIX1uhF+Zeu9yUa5zgENr2qRnk
gFOj8jpFniVYT95iD4eXJyJf4eMomv6YcP1BnhcfA+tXdTGpvC4od8u1VoxhLaXIMyV+Ib3GKqgh
sSOjvKgfwkaftZV2v2P4ZRBPZ+7qFYydDXMKOy8ZIIikF9FWig+MovaXb2/zvtDE9rEMbfIwwsdn
QDp3HHwGIQOAn2QrRhNkUy6u+kDpFCBG30Lu7m9PMarHwbiAF2B6js9nRU+2Y9N7CGnZF+igWuxU
bSxNv5CP4wzEx+HG591ikq4JHsKjDRozhcaEoyRXANef1eePlCQjWeAGVZIWs3KFUwsML7xJQ7wD
xLsZD2fj+sXkgPD4GM3cmjxF3hezFTwi3Yds/IgmPRusaZlr1SMT10y4i4V6rSiYho1jkbu/VPbO
H1OCoCJgrf/nx84N6N2IcO8U9QhiBNN0xBT6l5cTOKpvCjGzkaF0FNumKa2RoGCJ6ZodVmy+HBz5
4qB5xO39DPuKiFS7r271vDkkAuQZ7Zv53TDqbvJjnKqOuuaLCaRp2aiiJXzm/GwCnMyzdfgp2KMX
0Iq9kJVO2bvTRNs5h2YkViweNWe6ubCtyOsRdlAOVCCGFpoPDBuao4LwIbXfkHvBxiCNoF0htlkJ
12XQ0jGS2+wLaJDBYwwCZzwY+XqoTc1mdn8aZHuWii3AwPmf14caFtxEMuQOjdQUKYhaNc6V5sgR
AnkoLeUkcyFxnJC3EEozobXVj1Ca7jtUijgw5SRNBdLjNrXgJ8KWVIvOFNFL2PwTGq/Y3hYUsg6Q
BSU69rKlor+WUx8oXoyxT/d8Kp8Hg8Wyy3wPM9t5W8bkCIz3GlwzTEQhct1FLhNwCbygzATyi8Pg
KYrSB2qPya2v2luccPYxtpNMWt7O4JFdox+x5JTFiihOYul5+8WX3xyNKfWVd9/kOyY13USpB4ak
UtnbNJLnK0xrmua3PNIL4kfLv8joQdF00UJYJZQ4V0BdCZMACusx6uVur7+RtFA7jUzeVAjoaA4Q
eLxTY1KJPOs1cEzwZpkqd/AWm23valNN1BueZmq/8C5oCQ5m7TwhHmHLGIuMdp05HAmEvsgE8U2m
qGS2XKuY/ThQDCgAD9zyXD7p/deik5+L9nD4NH1my5GmJHS5KUUFHe1gxvmGRXgQfCny43nuAzDa
+XSM8SAi8VYCC00Wlt8TQtw+mFPTbRTRgj2WpktfFMOLJFY7lWaoW7we3Su/IrS3hq8e3dCt7+4z
l6nZ8D6+Ey9/sh0Rv8PXwN5s0Q1trQfwGi6ljp4d8XQkITtl+lqrNokoCHitkdaGMeG6mAmV1H6x
7G1LyKApAmdoAVYWQJnK8wQ+rwTH6h7MwWwvlD7S980hSqd+ozZYinI9QEOWAzQo6bMzWT3Ifr6a
aJfJ2JilxMTsHkGJS6QAPG3LkRqVR/LkmyR6QAvhmBd0ubWI3EZ30BLKFwQR/fNnv3WGzqETiPQt
j0X+ZlUT4tb5aeDE71PvnU1auzrdik3k3B32F7/c0LmmtlindSVQYca1kWlaxHKiqSKS3H/QGKnJ
AIn9GbcN3GaPZ7iiFMiwvPAcYunfgKCRCMLEeh3yd2e4w8yawwtHtyQZgmYd1cfUHmdx3UN3VfJP
FLqvwmK2BUnbjNm7QBnEWU5Rs6SVlIHYh0CEco72vZQRNAPiXuHyl414z0s4QcZQp3GkNMw4Oewp
HXuNzcWmQlJnU9e+fulpr18rFsudro0XOVNv71zR5sPN4S8N7K/rfEma/to30axm4MvlIS7V7iLt
5l4QngmbzDkAyyALZPJ+D1Aq9yVRFCcIYOAICWvWRy214JETJv4lZHEd32tpy/Xhc4vfo8vpv0U+
L0oiVrz17PQZJb7otdeRmjKpCILHaA4srt579f8mw+cJiH2c5PWK48Onehj+56s3HDx/JAtsBqvA
dQxl+Ss4xY0Zjxhssn2izeRlXkUgqJ3Z5LBjbKgkJ9RSXr9CqQDSbzK+5ZkvFslzihoV3aVBRYQ+
Mf+0iopTXaZt609Y5RGjyauNY6GrSh5ogPwi46+nAo2757cVjFmawNavP7G7Rn4IvV+PCIVoLpmg
HSh3O1WMdwzFdd7gVO0OJPpAMWrUj/6z5xAeAfNFVxDSpMVPmRofp2c+7wjMjtpmxlgBvdwA3Dko
EYOxDP/X22LRdWW0Sn5rSabHvnKi/dgU8ESNPlS2m1DO7rQJuYRjd/bZIP8h5NvKaJaM0syUKhVc
1p9rJdEvrV6/dfUI3ZbF9CABDkL4HryCN2zDK5j91dLa8ZvMKYNZiTziiONfmVfI0jKTJzYrqbpv
KUrGypikGwKn9AaKMGUXs6Z0kYAQaUsYPOxIzv2V+5fZohynNpnn4FPJPKxcFWnEaVqzO4YGi2gN
no7MXTBDTTTluSApelgxrEmnTuIPeqejQlcts7C1BQ6SyB+w5HuarKPALs2HOYgwcXQ58sJtKixN
t4WrYubaRdlPDIHHUu/BN9fZbxO/52fQRiKCObFrMN2ODXg4dYbrHEy+3Q1v6Uo0MUdZRh9OizrE
kD1ceuggCrIcdAjFOqrv/BKQLr5jftFbWdHEQchcBuHyJk0ScknT2R4FzqGB1Ma4vmpbndcnfHwy
lEacIMIMz6Sf2+X1pjk8lowvRCQIrUgpMCqg803yUPEL8rAX/Xp54atUx951PaFZoOYgyxCmSHhR
BH4ZmS2rdhOYgkH3ogCTBcpqFgtHoAUnwh0MkjeLp6ZGascgEM+RmEU7jFO/GgnpEioEDs8Orpeg
4NqupmiYHokeAyYjXGfiiWIChe8gS63oW8y4ynjOuH2l63c4unFpMaSCC3Ofyrznauu/BZMjNZLD
QQEIjm2LANbEJvfJR72eolif/UFQSSL3nXyYtO5odmyS0PyIYviC8Ekgs8t/k28dzszzcBZsP7Vc
aclQvDM57D8Bvd7vFhdNf0zHqLZRkkjCf4l+x4Y1h8io66xaG4bfCTc+LU4URZvzyoIkYEL+z5M+
S9WRYiEuklIiIOlwOVrLH8L+hz4Kc6e1S/yFaCKq9limmoXcg2nQ/H5ui3ovSQQ0wFwBCNNyD051
oFLEYq1ZNXm4e83GEYQ403l1IR36kXU+F654Uyl+UxgBDykM54ldwhq/spMsLpycX2Vp7MVP2gsr
d9JDKI/BVjkPTRC0H9fpk6EkZQaARD6klnGN74aNVQsfhZZy3JQF97JehApWALfN08jXM+veoSjw
0Q8/r2dx6/1W6ApbUVQuYA6hhmx1g2sgYHaZiA0W3Q8D+6ULAE1QP5mJGnwR0G9vEgHX/HGl+6Vi
HnSNf0PGiygn1LtHnBbhrctHg6fBjkRQyTntl2R8zISOQl03UixbXHOG7b5ovNB7NYGofuSw1kXp
DWPMBjI0eA0o+UZ1zPFlSmfpVFRbCNGcPp6D5XodO6APcKQe/cqq27xB4E2E1sJLfzXIkNVrtCLO
lIZ3Af6tIZcQRleQnFlhk2UYqb4/VClYEX5AzPnwvp/EMLTr05lwFvKqYJLkHRI1VanimiYrSxxD
WFzO2LiANQg6+cX3VCBz7r820Wq5VOsp/1NsfrLfJig542VwW1yyQkLy3ByXzJZ2axd/nIHg1AkO
f3kCNjIzKj7VQBctBWjYTTEvSIXyzbs1Ak7oWX0heM/QJJnBBvOW79yqS1Sszmk1BkCH2GDL1kdj
WjhRDt/kJ4UAtYN7+rkan2X6n2AWn7A1nFPnZipx5XZFq1jgmUKnZs6DhcWxXjghNErjc5eD17Ou
DmmFJ5Tat8QrvpF1XS0CbRKvVhA6VK0ra3pMIkOg9gPC1bimRozhwMKm5mp8V5dC0NcUSHHmQXS+
sSz2/ZOGE4qqv/kouo88aZdI2jWtxwfVIGQ2ANb3GOzTGOdboeEsVNtTHWBoouRh/mnvz2Hp6aPU
u/bCzBNw95GffOtVSc8cqrq6GVh8Lz16jCgnpOm+CwwdtVjjThxPmkFEVhxecccNBScAEsdixEZT
Do+iv61E9s9lZJEVMQMQGVnO6A/Bnwew4wHWJgt2+v0nM18hvfTjvWbR8Mi+LCfednzY8t6tiwys
aa3ariEmBRWg3GIeipS714tt2NxZNWaiNP4AlvV+nJ5TIGT7o7gkGGU3IaabU1UuXFbSGI4Gn2mN
q3R/CGgzRJe9DhoEDDTSG8XsbMTubkUOVoPxChrkzHq/JdeKzb13D8Lpzq4qJpDVRuUSMiq6OTfo
Xle8OjA4bLUgFjjSJcpS5AznLfufPCzZ42iu3EYKWWZ2sxjSsCvol73uTCtuYGBtx3G/t256fPr+
rBIAcyv+4he6Nvt2Ys7p/X5l3+/+mDvl3yNkrfNigGU7KT1TOT7VVuZliZd71DiqxWp8ohhnbpyH
uP6HBs5purUGmm2YR3rtObDkkCZJbkf0unM9EZfJ2F9jy5kPpJRWga1riW/SDYAeO63CGNE9sQqs
JF8wbjkgJKOIHjfzhpcDmBEINtAhD1NFSl5+uwmOJt3TU0A5W222aOniyRiGF3qWsN1OvoZDQRd8
Eg0SFWNWHNKi0uq5pBVofWnH1huBoZjQYoLFZcId5LE5fCktX9w6jPhn5X6dAUADRtkyYX+Zb2cL
qtHKju7+EnWuQDBTZnj6Jov7k8le0C9wtkqimHKpPnWD6JmyAj/ftuPEO+5gQnMC+RoJkTs+VUye
5agnBXtTrqDN9kTFiDa+stdCACcN1Jdz4ZGFpR7coPs9h23IVCej3vdK29xszshVBdh1Fu5kBCwa
gAEhHdDkz9e7Q5Hre4zIbBewsmcwB/xmE4v4XKjWzwLsaAbdEvYounPzgIwLGV+iofIcd2P3/D/2
M8qblFGRU4GocTwmJwFnTAMg4LcucPdoqhCt2Xv95LOLYF3BrKGQq96NT4Qbhek40op5mCVrfC0n
SjmB8pxH2VH92+g8Nvt9bYRZoZqNXFFGP0jqSLtLgG6Xg6EihYM0Dnw+WW6fKgOQc5lXKeOnzFQk
rG4aAr/QvmcFMUM/Try6g9R6xTAi0uNaxFfsClgzlH8CKrD92UKdR+hb918W2pOw3WuGAxUMsiJC
Pz4eB6WG4fkPMhEAmYcnCcNHLhl/yCCIzR9sD9WK0pp9RY384lzoId6jqrNLLczUS/oDKgZIA5pO
o5NwUaCGrgWFWU37FD0doTWIVRqERbxd0kZztnLoXtMum1xCLmmQFcwCp5K4lMCM3Z/IXtk5ZE0o
nitSH+zN0datodyLaCCGzjfiDo1fpL2PkjjNGToVQpy6YLzVOh97Xve4DcuHY3vhpGkZGO4oxwvz
gFg4Fg/Tn/VQBvA7T+XT5v2uyMPBdiYkgaALe0BvkHMHKLVkumVFTdl6AgB5VcbK4F4mxQ3g4tP6
nCG+U8TfxKN9W5vsd8Zxd077Yb4XtLfRwjzYUQaW3waM6OUXIYyUir7gncHJl4qNnssNHbqMmccq
L2qQMxi3aoVmp0uybEN2xEUd+6dBhrJuW7hthtycEZ4oYh7OyrpxGNGsvqmfc8N9g6e0eeYtIjJF
mLHriaVcKpNqR5UXsxOb8CDM/qmHAtt3AJ2nEikLXR2B5AP2ogxCTj/c0XSEdTYs8+MNQswTkxji
J7Sx0vuMudbnGJP+MlVguPDH8Z6TnQmLoXIt45tDcBmyvPRpcOvkpJJuYz8r08KLXawOT9Jh/4if
d8shzG1O13NKIp2iaceFPGuGZ2Q9p6zT4E+5Gzt+usmu0AjG97ATsLAXsTtxahLVMyx6l8Rd0638
wO6cQkKMdZ0uNgG/uB0uqycRmiy4HyRdzO4Mgi0w5EuxY4TxfdQik3r+iZJRpYSf1VBGZZN5hijS
OYGw2k3a3g4XT4X34d74L1s0KKddfFwC5TrdsvPb2ZOqSM5p6Y7tm6/uL1YWflsTXlmfOKvk6A1E
1aAoKFOfh8y0szZy+Hun+96I2rr3SGNMLLc0EVvU7Un3D3fx/H+neyx1Qp/JGUEeIMrvkAcOVZPA
q2tMSDJ2lUcKT7Ds1v21CRZnQFiUqOEq6M6OavrRI5u/LJTz7wWxtl61MKbMuPDceipDAQ42xwVu
foLZD34L5BUmyfob4DtZiWRxsJDYeJ02w4G9urWrtQaKwX6JzPpUszlHjPweAS9EP6nlKe6WX8Au
UGLlap6ZVsSpocJxW4Sxy8Yt1YED9dfMXLidULg9WlVXKr+LbUT1fC3pBCQ54zyu8du6uAXf/d8q
/IhSfefh0kgya6mH3VpnyT4esnTsp4Qsf3CmHQ6UXWCY6phMFS4zNi6p8UmOOU6veTfDJNV/M01C
jRIQao+wLF/e2ZNenteYWALwals4sdtPerfSi+eC26JQrvUft2EAsYOFJ5WsMGtZeXVrmUTck510
i7yl8QCx/+Vl44QvFgc4HYCxShjNs+kFDrzrpMMN0B4pfu8epr1/Uq9jM7RFZfSmzm7+BGZ/NRle
0jdkEEZZVprWVGC0TtmbxDEhM2BZozTCUcpm53c+uFFSfwZD1hA9ybjWODJXR338uoI3AH/IQl+6
uqPU8eIeVRq6yoVPXXok0AnU9RlYs066TaNutvEIQqCqnEDYon0T4N14KZiJ1K7c2xUP+Vzl/NNk
M4SNsJ4bkAh8ieRyBVCP1noOOY8nMhAlVrFLVxLHteyCNixm8ZSdjiTAOXJvXY5tjrZmEfGVDrZB
szxdZV67d1hRKZZaKX2r/2R0QKe1QvjchwNFxKQJKm9RVVRKj7nmd5gM3ypyrQoCZhuK9DQqNhwD
4GiPFnecTJFX3sKNU5r0UFMgkrt+e0RE/gDXg6uvaLT4mULDhF2XiJJz0kjlzOq+aawUqeUggv0A
pICsBsvnCM+IjkiKZpPrabgZnQtK81PNtxidBQ+MVr4DVcw92ZDNl7Xv2eq9iqFYYEFhTANwf1DK
hFW1nf8r+QsU8AcOIeM2z317z9G9wwH3oumLquotNTjpYLHS5Nrf1fsx4d5zU+ouu6TIE2z5yx/X
fUz6SYz518LAsVshWUdD+iW/nnhMfd5OScPDxKBoXfgiwL0EAHVBhhxC2EAUVqGcDCcDK1ViPbTL
chcPoZQyjCCcg4xz3ozzo9ZAyqFd1G7sZuGadoPccVIc60iu1I/aZSNRWw6Tk4BQIR66tUHFVUOd
WKWVg8i8A6KEgoQ6Y6BuYkRj1Efj3T0YzKEi0/YboyLOVoODqNFQ+Wxdqq8sDgi3ywu/MJB3lDXm
rzjAq0iForaWONEW5+JY6t0I2N22iAMY5yGOcPxU1LuQjYYaRr3IcKZZCE/D75dZ1/8IQg4CpCRQ
YC+S0e+mNqtg+LKmNIvvONod8gADtoOJYe/BsFY4ajoIWyfpYODY0EQMN80f95w7cjCbv7VfpH8Y
Jq6+FNHeZ1ZaJaOtYg0OY9282jf4RrfcaY3vuxqRBVVnWdP89z4GzIMjPvbeh2c9KG+aYcfyvl4k
b7RTD8BTUjS4obbS36hMEEAU2UEp44dqBPJDJfD0PTBHDZjFk4qZ0UcWu9bznAabr3tUlEmZpnyD
s7WqtlxClpIQm7xryNA+vvQ+zt6NjPc4tuJoP2FHMVMg/DvrDYrBJjxDU8XdLTrBhKSkNBGpEv5+
OfbsMfVY4RHBfIwhX8/j1ZfF5jAW3V01DKniwDxbyILRx7hkIt1UeZatXTw4mj0xnv8M2SQCmJJ5
bOBnFI3G2zZJr1ulmGvplmt/I4FEU5LXnp3QoPkSLtp+sFf0ecw+kziwDMYMxwAXhp2KYwS/Nsmx
DMyl4Uien7ylJiAAZ3BnS2J1GCoTLAuWy9VXqANJfIfklgFCqXJS7srXEyL74nYFXqpxgSD+t4Kv
teQa6llh2UYHyzfxZ2Xe+8Qx9bk8N0VuaV8WZEbklYT2WbklROlSoqpFcQ4OG4tfInhooqbDcpMc
6sHtIUl14JKtEQqgrw4Wv4VGj9DUSouC/123oAlyQ7ufwHQ+1pcUJ17jp58KxqUvBxhucSRIIUXW
CFLcnFg4/2lIZB5/knJvptxFXGk6UiQpdKz0o6ue9q/PyIiu6DEIGeliB5aRUkfcA59sPtv07J4a
aKqC2wY2BeRasJyD/W/waC4PHZDrtijadkX5uKKcMN9p7Xqex9XfxqSYwjR9Yu9p35+ysERf4L6F
jjGEuNuLeByI079kjpt3FOJyingvoXJ6lz4utaWgAWwI9RsH63AODpqFpEuLK2DGRwcAybpDN6Cf
pnQ09ngLXaDmsQhRJLIxD70k476JV4cw7MXlSfcczIZDnM63au66hqWf7fg8sLYfSEVzHRhtkiMZ
AEVlp/4Vy+bXQ01l9+ZVo+FzdhLU6a5YaAks20hB8e/aPC28vs8Opkf0nuxKams+K8MoLq2LCXeP
lM5AC+utLcYT6hX3n+yZ9Sv5ijXQHN/7pFvzPUjBgsrVkNvZe7+zEH/Uh3bSN36XOceVQYDImu5A
W/K+F1p/YrNZyKVR375m4sS4v6nLQw6lQA1UvCHFgrTXniIHOXBTf0yrG0uzKPAHYVw95io9iqlK
HYAeeOcdqLRKeV0KJ6G1smKbW2eTkjUB06vmnW8APbmC9ksFHRA072nmvM4Ya4sAtCBXWhBHyBEd
9yLBKBVAYnV7e2x5MRy8AQ5ig+C7rTmqCgUmYJUUDKt7dLkk+hOHAGeo7+mxGb1fx5yYhsPdNVEy
C8AqVNXsIwcx2yF7QdFMzlD4g71/NWG/GYmtHX2pbofzvUnFtyf1crcYKurlB1KbcVz0fDY5OZkA
Z//1wv1H43ScxwM+76d+rNWab+IVvOrfwoOR+qaPe17AzDZtMqtEs9MnlWpAqyYUp/+oTekvsGCA
FAsDogwwfBvaYIY4jxgyg7Qut8O+kSX55nmuKDqlM0d9Q5A6xW6nmm8617kYHwRm/JIZ9jZrFG6n
5m3pZigPefxarOsjmATPBAg7eXEYcQdCJJ1uHEKyos1IpQ6eKY80th0DWXQCmsBVSpkJzuNrLVDi
ExWtx2w7SSsS2eDgI2yisIyKW0nawKJV1gajfzZ/gnO1zqvFW9AdegsTFALULl49wGNS2124ULDi
iQaynJ8eSFLWm8ywcMcpEInK9sFhxohTYVt15+/Sia+ns/6Q34O4vjoITQafJz8ao7+apru2tpqQ
kwtz01WEXq+w3tXpZqYm1/3U9WTK1HZPERpFuRcNy0HYKWOu6R96sW2QjT7qWxkkUngVeea9JlF2
zGZc7t4+G1CAUBWJM+Y1leg+esqsqpcdqsIYO9iDifxB25HKqUj2x0lO+DYqFgdSGWWFslz5xzfw
03Cwyn2oJ/QIm+O9Agj624GRInBckzeNGSPC+CeQ0/FURW+uiJ/Ysaswbd+eQcWG2AkrwxS3VdNl
KmVksVD5ixHdLGPmNNSgdKq7EW/FoR8EM7s2zhNderPRXZwyRVtacPJJ4mQoe9zaYsWkDM5tB+Ep
RPXCUHOVKj8svMX+ROGPsAZ09NGe1y0n5khEm+1gsWTyYwA/7H2wz/EKuawnT8ZodN1J/XHdKCCx
z+TgOkAUbsgBkUoCHrGL+iR1SYg85SH6yQLdJkxE61nS0IkIw+uGJje4UAs72+Ot8k8rk2qA0beG
VK1YtP9YVH9dJtklFzVPFkIbU3jh//RRsnlsM5TxiE0LN5D7TcL/c+l3kqIm20kk6LcLaXCpqWAh
knR+FgY0vMrxzWOPhzmMSdO4F1Gz+AWY+/3MPGWZY81edMQ4vvOv5Bi3wkUWxZ9pohzt1njDP/6R
GlcYq7t80oHiK4Xp4Q+zLcM/jVUdiNxrFc5HyPNTOuRgVY099fMTfFg8DLt2N+mJPYj5GaeFyEht
CuK1KqzmCE1PE2Ygx7SaPjBnKeAPek4tsuJENb5NbH8hEg6phoMoXo20rZMa+9N1zxHKYYoIXPhE
B8sbpz0YOAA4l4JACcBFYm9YJVUwu8fnEFAWPvcYOrT7pW6DmHkHmFR3oi4PXQmDDl7cVtrviLta
pEu+Nw2y+dinDlakEMhjJD40NVveFbe8RbNJjDsCfVOXQPfqqLGxziewDxzbew7HQHEWLZ8J3oY6
woAsEAUTlqXoqe9/G3RwgRWqYot86s6bwwHpo3hrU+2Nm77fcZaLXtF7HuzTxGp66JZCcG8Mwd4u
uWXPEjPre7C94TMJQtjTkNB4+tXnnsCuFfpsap/EBsunL63CnzBCULrLKidp7HlA7EoUhjWxemmm
JjcuhQWKRBpofRWaOIwJRyIk2YaTwmAdaU/mdnkchbv/JAKWUP/1kls+dh/VPUPy8cO29D+Bl8Zy
Iu6uJPjD219CvovJOWOMTp9FwcmasXbyQ6feWfejaFyK9uwM19eIuD/reHjAwxbwqcGH7KFNJ41R
gm9zmW4Y7F3gAOPOuu9zDKH/+7MuzqR4F9y0Goh01xQb6vGzjDD+WKpO8CxuBtek0fF3n1WIGbsU
Xa576VbZcWJ83bZRVXOO4/L9lo82AONQ0AqekH9x/Q5hlFYnD48/wp9ivFP85IDKq/InX/AV1gSK
iOkJpc4CFVr18SYoCuUoiDnhvrnUfMy4dT81bXX7HHUH+rMF9HChqrgPZ/i89LCyKE9eUC9meJcu
twlMHvrSM+Sjfg7OwHIGV36uH+RC8HYGRiJmRkLTU8x1bTrx5OhkyxwikyMGbUgr7gF81p/oPgR0
6wV7s2/luNkN0MquRfyU0FPuhRCEzIOOYP77oK2Azg78sQ34yYSXJoqhV+5sfVbj8574k51vcZ40
QbUFm8vnF2axKk4PR7l4v7/BKWRbl5LlxlwGpJB+eE7vLtS39zrOjUGr+798YWZuhpcD9o7ycEx3
pkPPpkxxZTQJk4wYA+rGopcqPdyyKB3NA9bJUtAmiTVSzuC2Y/0dBK5ZYY8toy/D4E1sFoFabCHS
COeTZSn3cAc5Wv09y7DwcmGMnV7dpPXTRH/FQ0rSfAbRyhd4z/rmn3XlDgM+filhKku57rOKc8Kd
NnrQjDVLE1mHlADtytt3evqihoY0NYAejDtbRg9ZR3t094kQNSPzKsILRgPWXeY5RO33KwiKoxNY
5vZBZNgHOmJ24RnPpKJLXjr7nf9324Bhat/JGp1cUnZ4bthluEgsuhtIgdTprRD8fchiUU1YurfW
53QMJfIx6dLVFCbRerdczXUF0kunxvi5yftkv6hhXqndnjVTV4YFZs2EG8isYOBlX9OqJy8FusTr
rsnL1aw3eSC98NoDqE5G9Y6iedKjQr3MWdB/GEz9tSYEDbCcOinJDz9W76i3u53BS1nWs8zf3lQJ
eu4Bo5WAQ8Q1lknpCUjHw3dRZD5z2mwS42tKOnA9BUHynM19piwpnyuR9JSU33vPlWB5BGOukWJY
R0baWBPJWZ3Hp8NvVaDS7/Eri0JO5gGcvyEvGQHodkKtjA7Nr6Y/SR8OWD4s92co/RrhfBhQUwul
4eAFq3fwAMzo+khbWqlbsttRLx+9kONuLmWkYFqHMBNsZRVvmuQ8MbMVo4EdkEmJyQAz1iRqGU+y
qxeCP2xqRvs7+/1o1CQlxEkvlKfiwB3hOc9eLt1b3OeRsYV0NBUTL92MpxFCghlxXRsjJcozDc8V
FhKlTWM1xiWZ5f4gh9qV7R3i6j7MHUxpjbX5wMBfYh/Cq0AwCxh3JU1WaKDElTEbwub4WXSHlhKE
XbqOO3lfhokGVsIAhNt0KAj0P7H/qToOB4TIjgbLvptDdgDaBHWtlIYyGc6DaFyMTLUZc3u5Iwzw
cs7lp77YWsoBMLa8fsvmgTejww0BPS66xbFwUZjHKeDw4c8eddCA0HPRNv3hOoWshamwdyyefyNM
KZzHtFpLbqq2XshvPFulBS+WQyu3dw8drzisEiXq+RtCMrMaGilNpN//T5eke4Uq9O2i7DJyHe25
vMllnE8HnBBNsUtD0bTZiMkG5Hh3w6vU6fQu86w4ZE3KbOxSvfy3452OMq9zL6yHfDhysixeM+NM
GhGCbzHv//xHQ+qUHCCESMdwS0mCpQSpOxDqj9R6rCZpUurp2Z/S4Kl2sHdlUxo6IWuqo8l3hKM0
fwFq31Q6SJP8LrUqXH3RyWOVFyCBXaYbxSoB8dJMkMn9eu2LcCDN38A4OepVeKcUR3XAnv9SVjas
4bCaRxqcZ6vZE+nyNtfeub+0aMHYaUOL6dkEFHg21H+xp5SE+M16ToAO4t7PRrUT8dTFSR5BAzRj
Crvjd9AyxoxeUEq/uwI8pCXuu20p8thtDW1O7aY26xBAJM682V0vA1xT4JrOiaIm2vuT+iMpXQlH
DJJdeF+yDQGHVR9cSUPFjS6DkBisU9ynOz5mfcrPinzFzm0qKC3JU18LxbwyI0byl93UjoO+dTD1
gSbXxq/3XqZVz7dSe/ieCkWf1aEkaG+sXdc0d4sriJx4dJ/3pCg+6uLSEDtTncL0cvdAkbtCiRcJ
BRTiKi2B0zaePGFCz9uebRcm6AXe3HI4M/Oc8xnEXh8Ct/ZsUAWcwAUqRPuB6ovSI9m4I7bA661W
/1iNxgJCs0tJuI0onVQCN/TRFYiedjYsKtdfuGCZarAVljK7+N7Upy4LOHkrRzFtL9hcMtNtiB8P
DkEE7VPpmBbGeb4bgfVLf5l8FeCHlWbJHJierUILgatuclR5fD+XzoVqqYGlY5Xt5xwZxBhQ3Vc8
lpsE0S/nOiykyUbaXJvQxjhE0QGlLbfOkFmagSt0Klu0W2xSLP3hqzjlSyPTLqvLCPi4t99Br3Vm
TaNGwf2Ai0fBamQfK6yJiYodL6wng0LGkmeqZ+REM182Y3Tb/DPqM++KzfpMp+gz4Gcl07g++RRq
kIq+AsTA9MIR6OqcbtCw44bUodnEY36vaJbpocj/P+Q15MhThZ48rxkEvgb4H2l9SRDmODNqG6nu
qnqr6AmBMdCAzWNIJTVudXSnWWQyaxzVAF44y5h2n7ve6z9oPM8t/V2sUGXCMdqwBWFy4s9VSUiU
3ecuoPhYYtlVbVXqlRQ/T7C6RK0X0INU7t9gN3EbTXz9CyGyHRhsxg0fyf2ptSfstB/0nMhTk5sw
mTwvaT7moLRsPSySNbWxUOuDUdksIYEMK2+lXiQS1n2SoGwCkx+DPQwAhrv2VZQxqcRvD5G+/HP6
Mp2xfCUrdWT8qWLRv6tEFRrLr7DZcKlh9YA7P1REVlk2aPyrSmUZDFkckHl6n7IJAjsFI7TGPEIk
vIxKU+v7aro6KHUOOvcPxXn2UKuC/aPKQAloagnJh4gE3PV4TbFMIaCsBg0tAeycfFL45OvbDRIT
hQMpyUiUQ6uuLqWeAWF5HW1GpKye6ECwpqZI4xnPwdFQcQvra8gTrzqNynbqn8jxxpTBU0pW+bhv
mwm30ua1jLaOO+92QbVuVfgJ23ws+/fFmKPnLseIY8STirdgG4aDbY6FXMwa4u8BGZdAb/wEA6le
nLU8UDzVy+/8wQ1xzVXDhiSepkcAgmLsLsKx2K9fILISs0wCS+qYn22NOGMwErBemPqXurz9h7WT
bgkKSnZaD1RJmgPVfbXHZ/zVqUxHJyyckM/Kw6Yz2DaPckSF5TWb7m3aOYr2jj4SIkXNTo04Ym9c
moJsNPSd/ZaKo5mGRQsPAqfGkxmambgoq9TcJtxS962AHHoeoCVkznlj0YnlFAcnVOaauE/f8R1/
Em7jsjo1hx++2Tl4nFuS1NwJg18XKQDFmI9BB8oEU1R1f2Sm+NZ8I/YTRc+k8rUqML5SroQV7ILv
4FU/JZLKRIiIh079zigRZWiL+3rYn2p8a0FbrycWQOFJfV5FdZZHUGtJaJPf/2LIgLRFic2/ErXE
xvHJ74NEoMORaiSOWaxFvZqYH77BfpAZioO9VDvcIuMiMz1NDTEvWSDEV+XU3jiFqsJI2q3zDnF6
x6YcO5OfAajtPTcl9sfJMDt6TBlNzrDOrn3a1Z8rm7z1RRfzIvYYeqd52I3kc7Ay0hOx1H81m44T
RjO5WCXyDqCXn8M+8yBxEBjy2t89RyvTfZn0wKApLizaBnFLPcTVWaRAxgxwQF2zOEP+Cg5fu9RR
nIpA+CoGTvroh2Kx2U5tQn2D4U4elZwqJMzhCXhoH0ACsqPC/31IPqjDVl2BQ5i/MScAn8SPMpES
kKgd/P5qfkKT85j1uB9f96WGYPC1t5E9gPCyzdyI01FMUUZat335aNxzhrk1Z1ogamP2JSpYGHgf
hPMQMzOw0YKYRbInbb81UOC1LSCk5wsvc41AorALsn0sKVCAJZUei4igY4dAIES5bxG4nFEKKJMe
k7QaaWOkrU/Sg/t/xIocP7BfVsrLrfOqfw/Ib1ZMLqptrDmxr4rKjog11j0CeWH9Mo5U515mdn2j
TcqLxfLzq4t2vZnFAz+RyvF7wjxgHiOdltO9ZzspXF6LFOcid+5DlavXsSKCG2NRKA4W1kC7eCj0
hSBW5tKSMB0xyxt38JzHTGgWw87nD3AU+B4oFQhKt3HIIlPIVPUzxDJ/x4YDf6TfzDF7k7Apxny4
tgBiYEh0fFnssQQgB/QTnOUNZW4eJJv8OH4kMlGODm8hNY1NVN1NNC9KPBBREhESSD/uoGgerLFY
FZIZHsPZ5lievuSYgfsOfnkmok9OvJQL6Pem+fxmmVxRrMhu9Rd3Vt/a6OemjFZpz4gEDt/BlEMc
OUR30/rW7z2Ipg0s8sa+CTLwgLCCsC3I7SgtkArGe2HpNPNWpjNVek27r16VyhKC1rq7aX3eptQD
o5+wbRUY66h7TfyNQHBp5pySDcq56WygzJdHEEatDptS+/QiYT1s9D92uOWdAcqp3e6O4QpubxsB
dJoeO55K+/JUk3wUUruVSjCRMuw/rfzQMdkAxFzWO9N370atrmZH8ublV79QRKpAnAMyiB9tiHTG
yfRx7frGj0/l+sBNDqwMWIGDk+08b+tJ+1iDso+WP+jCcKaly1s59pdKdfZ7bgUp8NXPyw+BRZji
9e7UeshmNBz3i1tsxjmS3o3+YPzrDeVFh92mYQmZmn8vzM/SW61Q12g7YmCDu4z/H0zJPQnJWNDV
js8Gb3qlqV5390GapVK3u6Khj72htl+hbIqNbC9QJ5fWulBjvyTmatA6QkKi288as4DThd39Ebsl
yGZ6FxeH0PZWMNYSw01c8SxnkvFiA/nfk6SArKWxVqT8EPyMS1O1Oj99NFLREl3WbPrvyTA3qIDz
+yNvE00JSR2xEgxqu99tfTjUROflbPCYkASWPCvdQAJIgDDD3lmAktB8PpRWDkGXKCdgRMCAfXzp
zPanxIWTUsbX/X1rZsWuFafohZaMWqQzpqhPXA+oel3FS74ePBV9KlXLFW8+lb7DVutIGOUlmfTc
T9Yu4bxio0k3PqQWKzjf3aEBA3UuzpfFHk1Pp1hhzQ4oHejmgngu0DWM3kGFACbalp+mtlTN/Opj
f15J+UU4GSjn7D12fp+lXnfI2l94HHvKgoGGsXTPN5432QlzVqO6T7IzGa/9fThiDTYQBALMvhdB
Z2gzai9GhZX+UrkEyPFhp7C4Q38T+fdYo0+LYhEn6LtcwA6hOJOU0rGsDe+Gtq7uvdaDbslHIOQG
cAMmMbfQDJP4b2hxgw8eU+CslxXF0AGD2EEkM3OJqpIdLTMZE99phJmi+nlLOCihjRIC3IgHZMvg
rHpr9IFJJl29GUHCA9iFMLiB54Ld8P6smy9RlKKdveqA/AaP5eaYsbFT9BHAapYrp9icHd8PcpeE
EvLGW5dhzo2Bhypf6a9N/kn51svvU4NsBmrYqpQ4Krm8jMVqN2J42pPeutKx9xCn/3T/4hgg+CEG
+VIstuDF+B8vVzYckaL7XWV6eyzNgE6w5CjH22mvA9ctF7FKV49IST7RHgdocqLTnYytSrnxrZN9
kHxZt9hbG/WMv1yIewGQwH+BWf6STXGQunylP8vNeLmMON+ZJG0xallXZqsX2QUzXlt835By4iPA
EpzfQB06pdvWVurUhCcli91YLJF5BOt/8HyZAVNTN8MovUj5wBjI6cVyuQug5ataD9s/3ZmCAIVX
eDE6Q8KuJT8vz/VPFemUUT3uX29L+tTJjK5YhWX8HWVPZMoO3OMTE3fiYhEMN/qlntlaMJGqepYt
9jEwTEwVTDtee6lZY3vtrRzE1pTKCuek/ruUQAQMHPkcxImi6YhPgzyEOMj74tjjYP94A7DtMk7q
7DLFwoKxgqAQdzLDZK7eQrd6fH1jancBn/0WO6lsuERRV8jxhneFj9KqMurdBhN/ag0sM9tCIvZk
m+olpgLQhBP+44S8WnoAhJBfje7OVKWesV6Dz7kPsurmHASeZHJvGrzWuPw5Ws6kgaRUB7QuLKy4
WnvuU/qkQvWyFBea3PbENQuy3Fu3gsJOyKV15vRphUBtJt/ppmdaktKPmJfFfLKAOH85zTLBNEg/
gOeXUaDi7gf0nnTDp+bGid4GMJCHcsBgTszloX4uS2PgAgT5M1CphTZooaHhpVDP4SscvPtu5t8e
lrD3nqn/aIxLSijq4XkiI6edBUPGKJr71Olgnsj9wO77872Bnc8HE98uZwU+gtiWJUrtU2uELxMb
XKXcxTi9eO17KsrjIH9nIZa9osS0EdbtIzQZZUOvXOZwxrNokaEuIs4GxqA7dYi2QZUfGXQSGL/z
0xVEAR6lVkUVvLSZb7V7N5Q8RqJDi3U4LCcO70sLez9EqPt7/EjmEm4BzhxdxiFdooZ8RRcqPMJ9
DG1Syn8IUQyXPfe8P59PmJkDmiXiKB63EG/otJizQ6Zv6wRA1PCDFvEfXkPOEadT7wpDvyqCYPa0
7Ni0shIkMKUS8/ZfES0qpIe4ORWqFfSrhFQ8xHh731GPVIzf/cD3rrBud7fUOu/F66qCeZAvDp05
EDNi/UdIERTXqV6mWFzoi016BZolnMMqqiDtzafhaKD6MGJFevBwglPwraBeXteFIRFTl6X3KUm9
WrM4iynN77hoebiFW3bYhD9N0nK5XyjY0Ogv629gqAdt/wxQc84BpssxpL2t3DGI020uF1kvpTg8
AU2QrLzrMmZWJnO2ZRR1LGGls513BnZoJHsU5HZT1/UP61k0MFrm3DO/G2bEIadeJVxgfhhVPpuC
QNU4aEC05n8xU2xkWDOwIrKYCHRqtu/M00vgFERekuj0MahGMabLnmZGawR4gHqWHn8NmCvDlzez
siUBhPVB+y1YPLVU2uFjKH5ux7yvi3tOjgyyz84ypWRunxZcezXgGbvuwavBsuHOw/0mA074DurE
XLd46fgrLrlZZQ/kdTfi2aaLcblOXjxgpJovlV2Wd8vrc/buqxbHgoSkA/W2y/57lFUFoBihgCYt
YIeoIFPEcHdQxBJ98fZFdKHkrQ+v9lZYDMY4msnzgwFWwIOQjNWPoUFDkKRfdoDm0jYetmasCfCw
yCS3tYTSTav0dxHTRf1IvKOfhEIe+GYjvWKN2BEsJ/vXVVrMI6FPryvR1RrRtD+ebwwdfdQ3tQLL
sokwH6tCcHNWRlGJNWbpY20FsMl9UIXdeW+yCW/MWXMDc4GsOXF5PnYcHAMI0hbNUZvvrV4/zWQ9
YvG7vlImQciEM6uXZX+DyWqjUD0OdCFw+tbLdNfNBd3o4sgRIvpAp8c0qWoJYRIefVHxXB4gV0OY
+8g8ogCHLthd5pLbU88Irnr342Vk5ycN10yx/xjwIZCbHTSdpm08bmclAQMkGKcu7liYlD/1Me+H
aeIkmOpJc0sb+V7ES477qlObRO7eoYgi4Til92YxfOIV8fw5F4fjq2RYx2ZL7LWuyqtmFx7SxLx3
DWBWU+ECuq3fHcEhsnWPBdB0/EYtMgmzy80VG4pAvBQ2KwTdwb8AfiTeG3ILpVNxBuT9aA5E8LLd
bnndukxIBSZluY3fzoai0IVC6fT2wRtvcyFdBrpNN0ERbARLEzW1iA1gJZzJ4W5jHI4Trm3LOWlW
N//qQS9rO1qhsXtSpnwu8D+BCYUqZxhZ1+npB7/8ABOT9zbBzhjq6umB9JcPO3NdCJWqjP73uJDt
lgzddeq5Xb046JClzcSG4C6GyryyElkBXg3S+131u7XRj4xUOmGd24bTjDiwQ0J4YICWEw6ekVB9
AbSrtFwyq9YknonzErhBFr9y2iOlvdbi/SiQ4P2n871gibAB7TMvrHjV9m/zRxzuKxTnCqFgQSFk
DnvfU2nfla7Svn/CmT2RHvP8JIm0IT/KcmWbldHgN9T7EO4gEwQd4lMTqeYrnn/br9M3sY0vEo7I
yuWJsSksB+T34ARLSehYrMCiBg0zbgSKSTIGW7x5AXosvtMZ3dtcxI0gWRveVsgsrjzIZEZxulFl
TSFGvpNDdvHXosd+DG3j9TZodw/Phoc2ggkvVpoA2xfgX3EXYdQ5I4U7nS5q3OR+KG/4leuW4SV1
sUt79a2uabZRkDWS289OzQaUYDj3bQPjOkGYpboFYq5KkKFN1pg9aaStUWVpmx+oVFsnvgCKha2w
nWVNMOZiC4IMTOZHJoj9GxPIKSKzY03ROQ9wuX9vHx5JfxaXpxAvQspfPc0tgUC74J0h+B7mQQFD
3c+eDPtpX4hQ0RQ2e9Nz/7NrGAhrzBee7lQHCJojLINrDwA2ihVLtGBQDZ4LsAsrdvOaeicTSiua
78p6d/tRiQrOtFGxXWTsVI3I0lMTmAt89Kh3VU6AoCd/faIfyii3lxWQw8HhiZLiG3nUw+VrS+qR
rkxPJ3DWFAUJL4rQvuL+odfE1Id/fIFGDMWdsJrMwoxX2tAIXfwLhoqBdJQAIpDKhVDUoCbPb4y2
Vi0EKMPwF/g5mN2G1U8wj6GPEBxeTn1c2LoyVrkRKJl3tSBjTF3xmq4qOcR3TUL9la50Wyg/KcLe
nrsc0cTcywaZi96c/nrXtgr6tQdfW1UQ2dXkkDqBZEj4mhd/wWmmycNPvTHBd4AdzJZxJ8cUoVEQ
TQeKvQyzOZUEsl2S2h39wOwaU/Oa6ZXSF0Y5MV8+AaQM+waRrwFyElfw3uZuHte1o07AQAyDnGRV
kxeIW6eNl3bYtk0d8lFVjRsGS+z5tkYREIoM3NdAu+lbnhfIpGxs/mDtmweG1fL/THtSv4YSS2IP
iWM82yzp3X6v0ty57zkqdPvdg/v78jSw5d+GcwityqoMqA0OCuif144qu87dGp96BoyEq/lhirld
Ponh3pM7HnKs6lQTyCm/dPLSFfA9fe/NvGOkiWfDKBdBTRTeXLgkIK9csUdcaccEcm0YxtwLrIVN
cdLIS28KDzlWp7YL8P0d/S3+4cK1QWyUt/gGXkpAT2903JrHnBdgnNY/giBM68L/MQGwW7Aj0BJ2
1ZPyq1hk/QvjdteKPhsfehBcQCcwVmyGKzLsZjYV41AAa2qMqX5l/68gQQsVFbgbw2y2KlWn8EVy
NAVvNzAxQK17Lk7N3wziymULbEs4943WLwk557LwWQ7GfAsibSC1Fc8HUUh4A9/CrI3qQ3u9pycW
zHv3lP7cmVCKidg/M8rMeOZdpau8046F7USDqNqOGVEbxdin7rvQDw3jRI2av7/ig3a4BtJQR4YY
SXtP/fzBGUztBv5Ujuis5oJMKdLyE1/HNXqXJ1a7sfwR+0c7Mfv3TSK56s9gFsKJR402ebGJn8cE
zndzHeB6pgC8x8iA35IfEASH78DeOA8JXVCmnGCkxQyNYnpmOPbmMGOiTqg5EtNCsj3XkSbiA6BR
ANpMwub6XBiQEdC8Q32gA/xX/f8LTrgWT9X/zLLSSen+nMKxVTxcjPU5wa9vSzdgYqqerh7Jteqd
ljVfsSxmZ7xj8wXC0HOG/W81i6qP0OuSj0UeUWVUtKWkI7XTiTLnKwkcqrVi7yOjkvx7HAHiJD4Y
VTYjuLNABLoB1DsLiG0QQpLBCQe+enVg7QyxFFI6dQmXyvTjZnaCbLMP7tdYXNQCLx9XM1Uqoqas
nfq7AA08KreLw8pzLNKivv2Dq2FBKSqd10xAS6FLeCAyGEVMkfsVevxHwfQp1EWL/4EHF5ri4dol
wDOq4rhAH0XSzKlOOIFC3j9FQEiS5si0tKFHEJY+zeyMeInqoWv+GKUjPCRnBSBg1DtW2rjbca9C
EPCi+LFXFbljcICbDjO8+X8oTxX2oB1BQsrWaFETMcfCmlt08nqM0NE0KlQ19yOOFWI/NOhvmHzQ
GMIMNNy2E0G8G1Gn6KcW7MNkI3L3DXOuHZc8G+djQrHVw9/CZqlNNagAFxPDdLeRRsVh+NnMTafA
znRKJsiY99jyy3cJRIvKOxct01fLYwSQfHwgj2h3pIgP10nMF9271yIumJxEchAy3UOcCe5WSaSE
HsBuZFzPQ2WQMtWSgRUr209/ROIuZ5pwPnh/CwA9qwKytZUWm/tiwhWea2PluIQhOonS1pnG/KI+
Wsaqt8LGgw/c7aNQeuT6EhC55lBnSCUFDc/0bKfJWUiENZykDqDI5OpzrXuaAlgg7kAyRiWCXqWD
M1V9gI9wPU98CejidYKl4OE9MBpUTYQJSwTY5JBk24cZjiRmo/OELOuGGPw13EHM86LfmKnESh0z
3Q7EPm/xd3ScsrADvJqCKzBeR2jEqQjwI9/N+DJr2SbqnVpmnyQM1Hy8yOfw8DMw1rjLclj8eh1W
wuf0nxb7IZwrGYAOBOZncB/B4d/h6UZTvcTilaX6B+mJZ/nPK87/2isLRdaXALfXeCNBic43lJv+
vTvpiryWqdVd/qHG5vqX0oqc59nnuAS3YcHMarR3vuUkALSU+2uUFK1qY3jzJraZM9RLv/h1JAiy
hRlaJ1QI+A/iz0z8roSmu14lWK4ny2cud3zlF6/y1VF8ywWs/ib13kE1vJbiuG0hKzgtUEJ0QJBd
y8ViO9WvGPbklEO0ir6kWHSNOHyYN979gcCuoy2REfEhT4cstE1Zp93N2R+/nYbio3py4X0+VwF1
budAya0OzZgzCiEa/hPy7NywyABQmxgrOJA6VlDC92fGjFtf2SCMJtb1Q4Kl1xMRqge8WiMuiS7y
5aMMXj2X+0Fnvr2e+940fdEntARR5AjXR1oj7LbZ3BJ2oipAbvWGsu6nSAvF03FBwMQpbfL5vAml
lfJueuk+d0/qBYtEWRSf3KL3gWQyTpfiTVkGZ02qHTh/41GN0ykCQuuCwbf71+D/CXh0kU9IxsgO
0pzrKYO9oh7oJUK0xM97qfkc4NPhDumkAj4u9WcT8mJ76iCT8k7bfscx+CWDAAFax6xUjxUgAlmK
cErj6oHhHsoDt3rJbboe8JPYcm6timZC9CGO3dWShYZyDTWf9nKrwTVzipOj036Tsc0c15Xb/dN5
8yiekfU/DhvAlog/JpbNpdwYeLuxfYYYIcjgEM6f/C7r5QcVtOzW2KutTNBI59X5TYsSXqG5Odg+
bakAHkE9ft49P4Btc9fhtFDCwCdeQjwlywydlTiGwBSd229WLRQy6PmOqQzRJIL5wzSslPsSfxx/
Bppb6RBGvoYcstG8Z2sR507LxZdjZj7O7wMco+w8mZplunKR6vliMckBqqjZIoSzlcO4fwCyS7jc
KNwuh7RnE1pirImhkvpkRsImu0x9eppPzxfkf8J2QNskji+EzFykg2LGUlSmJR4aOo/Pw194Ntah
dNc/rewwwTC7vD4oqIgtmoW4G/JprLFtVINK2lNwtNWzFvIvr9wufMxm0CitJ/MElu31KGR6B9PL
RqR2273dRW5NsQ69tStLCGUMPTuN68yol/IcpCAI7e/kXeXQusG4Wcojr4t6s+PHA3unpNdgTDmw
s6V58lsIAWJKGG3NR+p3u2rJt4OPayQtjyC83EJytjV+v9J4RNMsztk5jLxVmt3U3Td/KvZca66d
XJ1rhxTDrl0FsTrUwwtOjHCkRNaECpR0UrpnKFRw71gr2kg8AGSQdTvUru4iaenRVuyz3UClfzII
eT26dXJcTNGu9f4pXKa7t7dR4uW+FCf91BC2XYEHdm//9NYu2sHcIcgIzlH9uCgsM0h9wqhvsprx
tN1LQBTpMDr33TNbdaJAK/Jf9INq+xN5Smq42pUadIByPfN9QcR/pX0m/ZTeQVWN5goV2ZQt3i8P
cBMPEJ2UQie8+QsLhaClH44y6QDJ/B8l8Ct60H5bEoqh30m/+TNDtzkW4yXTY+GOsVsZ7RvDJfR7
cuW2Eaad34L8zPZE8Q2Y2h1zfvm9uv/7E0ggXj0APttncaEjQyFTL4VfBrnXK+DG29gm80hwEckk
ztZEXE8pfZ9VHDf1Agt4cKL9z+a6UCBiCEQJpLpyLiod1UYlgySGOxEOM3zMT9JBkqhYa8tghRq/
LIWUAALUQT6LqLdYzrPB0Qa9+BoRNbxZLj1HA1SHSLLbXO/r72aPKkSD1QDm4pfyTfOS+eCUB5vN
B9y+yn3TWIEe5X1/VlJTPchLDr4sC3jvFF7LiLfE2cDY0affVQPamkbCDE9oic/TFdO4e0LX9BNS
+4AMAWvzxlZNNYChQvMs0//hwHEmwy82o7Wz1Act1RP/Y0jp2ydY16UUbcqB1kihu/o+svLxHTyr
wla5HMb54DVEn3vUfI/q4o3YXOe1vgm/fvk5hcCnpZRxqjHkbujcxkCPGeLrUC/II73OQcPzIZKC
mxkIU9ywvMjbxITCl05yPK83BVPD5d9earp7Tj3OliLNLgxTi/4iNrJ/FhUw78gGMLsIkHbGv8jJ
QaaOGPZ6Iica+0dVHEjNGccByfw8PTq528gA16Ar+DGxNB9UzmelqNegBDgebICseFzhVNtE0ooK
5n9DDlC8BoYwe1yh6AE0U/flYSA/o5htmy570ocnqdrgpLIQPKXmbyaCwHCGe5QQnXUhA9PpXPKy
exO/iaeQO8cZZyqx+AELnNfts5ldUlYhPCzpWpJMcvYVRDTmjkZ6LYVv1OYT9EA7O5vLhgZSzrUG
xQAMvtsHN/QzFlpYwJxfQSx9Qcu00m7FXjumiLRqcx0GB3k4Eb/x+36upQpeAOjzZFXgIECWqFOZ
iiIPBMqfmETZBTGn3cZFQss1trZYD3qf3wASWwxONJsz6i+J3GKsGpMm6jr0GzfwJy1yHCXKRIqH
dy2PRyzIgbpZwTxbksxCC5/QzSQT3Vt6PkwzpvcEVo9nJLYWLNdUvjAxjTHrgItsQWaYjcZc/if8
Cb2Gbuog7iiXpTKkjy+All/Y/ac2yedfZOZsoabhkXQ+83E18hE0x7UHtKnh4SOqJMslVsvn51SQ
2ULjB91GcdEIFkAXi3AR9UjbtUQ7CEkSgrubl1MCe8KUiGAy607eWwBF2nArGVu1M4Pq8oDoskiL
KJSSiPjhsRuuDqSKCKrCrLHQ/6PYXzrhLGuQFDbPuTQZi9F1WZHY/DASpXzliou4ezKxnPMS9BJT
cKXVFEjrPlRTlRoUCM5Ff2LdtJEgvIsZXTOzc7nqPhWlcMBrsRjSXztzOUJZav/sjhRGS/jFBRyY
iVfFoUf/9aIN92Pr94GAEV/cijqugkS2i4HzRZv6H8F1qyNhLjHRaFk0DGGlhO9ZcO2Up2KZB1dg
W9M2+aZQn4G+GXU5EzMj5wnZ1keRx+uSIaDqMEGkJST8qhKX082hFvWdmfXTyPg3GMOTajeUWUyT
ioa7/2YYE4bSvqa1ZQwFfXlSGqTbBOnHr16JIeUR+E1l6+evelhAS3rKRLumODXfF1lP07TfIs01
cznw2lSp2JO0xDCb6Fn2WFko7sqdupBbJG2VIjtZGX7kv+VVewkJwMU9RlreX0V0z9dmu6t6SyMG
ZSJMw8jskzzTAKgXbC4kU1Sl73MrzmUGGbLhhQPlf0WHdoq9eGERz137iBuwayRUSya0PEg76Qzd
CPwtKXtWmDFQNThA/lamt/74mBIp6Yh4g1MwjhtOgYm0MYGPX/S2+6Aw00jEicfA2mmUjdhnVCU4
zHuzQOCAWS0+hDs64wMlzuyGBtIiYMLtjfietba10OxVjXqtv4JfSK+frnevsjXKhpkc336fZJq/
SYJg099pxHuuuFqZXV6fW+ttAr47uHG0buZWrQA5hShh1H2Wo0tUaNnBO8kYKEz6R2IfWrFTjfJw
rHZOtdeduSVurHyrcY1no0wAVUcrbCmsRJm38Req6XjP6vKZL5fMRvYCLsb2U1XQn3zsEy1iWQpU
EhxG+lNHbx7hJaYEF2Wt3FIEeK/Y6zp+en+8gA2or/BKlvwTT5PsvldMyc/koOqD8eJ6vmxijQYm
jC4WfTIu/gtu2MQLzgJ+1p1GDaNV3B0/MG0H/PTCnELivPjUwI89q1njAMLy5xYZN9c8BlvnUlrT
W2KyOIcUkQw4mObK08KofAyyDZWS3p6/p1l1hR7y1cb/1w+4jyxq05g2QAvh75nfWqWby+urFtx1
Tvcubvr/O60RmhU9TIZaLkLg7X0x8VjfpeJVwcEI6Q02LiLP69jnNzn1hkSx99jHFqPm2/sYgOC7
KwpxJLszXGZbu33HvVfTmzenAGxoCv1Q8d+6MM4otSaV5PmykAzazHz9MXDD+3rbIMvGGFywoygE
UyjTmOUVrv6qII72aNxxTAuwSEQCvKh0MXWJaaEpBJVZu5vUwbcPgMa0AJdY5nxTrPWObE2oPh7a
MSbVz/AodUeMC6/qZRLAdsPuDlixB3Zx6pQ4k6/h6ISKqauRd6NaSB3xuu5j5dirQ1WEYVipkokz
a+cwk4orgFL4X/g5WdK6+ggWsvjJfJxflxeL+BML90/nFFvWFlqmygN+AOLSmKp8EmoQWWqzMhF2
fCzwCuIjm1x89xP7tcGJOXbchrYLyMgHmYt2JqhkXUGyJ2T/L+Wr2XV5iUw6bqCd6dCDru+DVccq
vQCIeuCM7ZLCqfFOJ/rbf2lSGJkdMaX1jzIqzS17Ukm97F7y/S8AAO14xk1ezoIJ0/qA/T01DMnT
YflpJtcu2pLZLbumlCcL9z+lPAGWUAMdQaBI4JfFycYuj8UOk2L9zCNNRHTw/6PSOPZZ+qgGbZca
4LHg+c5U4ZuAqDLM7Eh+C3h1NwhPjeiGiNWZjQHsC3E/49Hi0jYKr56ugniTzOYnt7BzBD+Y7u+7
xsgeZAmLZZI1IC0gsZmQMvkOf5dOdMtSwh3AyjLo3n185kX7h0Xtac0bFMlYJEovg+u9127Hskbl
4G7C/Ovk5HBuVYQnGmeMvNY1oaRfHu0Pm7+5k99q2XxO90SXy00bLBKp5l4NKeAild/ex1q78A23
JLeKGTJw7z5H4EGMO5Z/9MOS+rSH6c/6doGmN6RMwqzF2aCiIdcRkRVf1MqQ91zYlIDTiJoa+WXn
ZU4h5mUWWCA1/4T1H6KJ7ksGps8ggNXv3oyI0rzwBQGBB2BJlJdVRsiY4SXdtVtQf62Lsbu4ekJj
2jkF1NKmOF4pDmHgIgAwB/l5bke/crbnWtz74oMF28u6owjxUKLvAX0BPgFtIwG/07FlP4gAsjEs
3V52XRCBabOEdXUG6wtUeIn43/qm5nM1QSbrq2WgCKy2Ol2bNS/bfeh4pS9ZNF1dtn+7nWBt39YR
iNOKb1Wvpa8JiZKrzfpafqTFBDv4H7QnAyAZJKGyEXR/Z5dFa02pmzCL+CZmIs7gtJHJWAn5gP/E
S8iEBmXIJ1KZqSrZKc+hw6NqGPsY9quJalaH+nOFWh8T2V1F5cw3LnKIQC2SzXczTrWSdhuOxRIR
4mQm9sruMoXmOBudXbCWQilwU11K9oG2TkGyGFghvUa+fZ0KLKVDSE3ww6LrPzi/fVlG11BPBmoS
uu14iCOwHCJixQz0xpov0B8ddPsMeARa6dhh6bMRWRkDG1Rw2Qz4+sKVdeBb5kuu9AfGDYMaWWZl
G0nYEWo/zuc2MFarI/OdGGfErq7t19dfPbrcb/fo/qk/UPjJW2eolXsC8OP9Q2iLdUZNO69sNEdL
+VjGZEhMHZi7QPBpVJcf8VPRgWcJj+NugcacjxDDv8t7xY8WfBAMnfehWW4mMZ1HDMzILZH+RqGT
uADntI/YdPYxOao5wfsPBfAXcqT2cbiMGPyvfNPQDzHBmbPnYNkukXS4C5s1tsCCsIFwS/rOCNGq
4CZIBhpJZ23JgtvjmQn0vXehFBzG+U++ZTbWrWqLhbKOYRishXGqQp3OHOo7cJYoCIXJWZDN0f1o
5vZ7UUp/X+8HtGFlmL77FC7bERtZyz0AxafD3ZKYn1kVhR+w4C6s0vzGGLoChcFeeFMVsNRRjN6/
8zUNZfkmxtLvjW48kMRb47mtnMqOg1sHUzA4riUXXJQDK2wf7V6fcq9ESJUqa20sIpvhmyERYPxc
kRJuNEsjk47x5V7zvP/JE1+B5O2L7pxkFAD80DCG8ia3d65MtJdjSrYJoSKMkyibmdH5mudt703r
BMDuiJuGnaywcYxajMgT0AtV+LSCDu3UpLIJWP7u0TypScK3RQ4zb4uuYL4S3J5su9UeheOBty0U
GQTDC6HB84Avxv7DTv3zWDiFbUndttvHgk9gX6QAaPisIXRQyc+g/JnC9ckxMDWcYkgghoodhCEJ
KX602/AhzgFn9rT90qQwdu9ZISipRD0HAFHcVafTFpRtOmaO4CLL8E2wC2OC4G5AvWHVvQYsfKO7
hDwi7scq45AE4ogIZHoXwacnP7lPpM7c2GI/ISWKR4Atgqs2TJNpDaV66vpg7X0Klf0qxOg+lFxe
SjnPKpSRO0Rk0DLxil2anVT9cxctxE7btvNtijuWSmPrFKA+0c6AZY70CboOQtTGn+R5UdmZKQXN
5P4dLZ0LgnSHLybWoMogXYEe2e345MHCG/9WgGKsMXHPb1OVhLtaTlwNK8/r7mduvoeGQRlxtFMB
WhGtDVcpsOamriI5HQAMamJQRi+LyX3vLZg952TQzeQCHjB/fe9xI/n7IBF8rFJ4+DyY/gyX7FU+
1fQ0TcildPyB07xvLClioFBU8O4wO0RYXaZu/gJh2wJHc3yu5EpefdO0BHgcW9SW709yeUZbCv7N
qhKjfZLlFCowIa1TaxaqPTN5/KVv15wXTVoJOMmsPB1RZPtjSqOfXYpT0suSMN8WFRwpmPgN2uPt
BptGAYMZatQAXA0RXCpBLdCTeNX8VNopeme+g8AtHxeHjTHXqPEFqnQZVYQvic+DYNmIbm4wlDYx
i15vdTF965yjdso2pLffPGY72vZ+ypkYeDfiGhKNr2ywnoSCE7FPZ56vzXGoTwgpLG2ekQ+WCMeN
DPpwK9QHrx+A8N8Q+57I4z0qS02FIBlHbMManSus2pO57xY1RN5YKGZhe/ebR4JCi7PJ4kFpiu2J
Dm0rSPMDhd0zfC2xUr8HBVZHvs5AqpiS+uwCTIk+9pKsyXxUbtxWDMIO0S92ahsBz1TKZwi5Rwtd
H2tWk40/bEMKgAHz2ewQBpUdYSiIMEZVL943h4fXpPYPQClrqADRj/nmBW+yvZmkkF/1BRKm6JXm
kAalhZ+7NbxkiXPzNp7T/5ZLeiG8mT0btQglc4mh6Odr3De16UNCAxtFUVlYZKyfCIaUAHGiLHMp
y+GcVBwYaCASfGF5MInKseykeV343vVZyrTIcwB7TglusMfFBjMq2ww8g0c/kUrFhhJwgDMZ9Xzy
ZdjbsGDfdXY1cLgoLHVjhiXfgJWEPC5qrEQZ08AefEpl1BcePfY8c5/h2JybDBzDnPDDX4VJDXK/
2amhylt3Xdg+M9Z3nRG52kNT9sAR2NojHNzvPAOXAbvkzhcV7lYCbNGWEyTh6cQMrLk2YtDzp9o7
GxGdQEryECMbAz+lKh1iUR4oYueWVygzX7J5Jf8ZVLiPWbJscibspUas2wFWDppGw2hJBdYy/BUl
nDBcDunlUX1x6ZKTylb8Ysj01m9CpH94MMh5quHRlHsMsa2/rp5HfFBq6tW/xb2nCLhR8rAVatSE
c0Tg4Y6qVUmq/VZuDY0KXiFJV9xKDoUZVL7KnM7sKsRgbGsgaQ6DcmyUCy4fS07zzfizQprsROOy
54yVmWNqbt29QmVKYvWFQfvjZcayGC2eIGV/KlabKo9HhSVzGsGK6aAGnZ0uAiNoGyg+/4nR/Upv
WhJ970Xu1krxf1wen29nO4lf9sfhtUh7C0KE29GMwKdP9EQ10W63EZiClKPSUH8/DaFEotaBdeba
E4RNhEMwH+FFUMPNtop/0+1V1r2oK4cekL8bwCFZd6M5uPQOIzFILXVbvQNuFvuVCyRiI+Gn40lG
is5nM4c1wP3sGowLzKTRtLfGKGWZVkJHRwcSuIy5+c/n+EPeD774MNJ1k4a82YSs517z7X4T9Qah
I+RnB4O6F4y+gb7hvFT/TwrI0F3OxJU8SPcjjlUvXkF+avbctsZe38PavGRU+GER58N4BC/Tyx6z
BlJcqr7v1DiNfFBcnuteca0TbV8bs7pciHLYLSf0p3ypj3WrfUeIz2JwoQ8ZWMOnwxKQv5R+jPCI
hzVWyshiFzCYSSvGTRYHBnuNQseIowKRRpdSKVZ1eQTkvkrU3C7ng51YlEMhVbs4htEHM8JrR4vb
/IGmoRQ15sXk8sk+YYYbnWJecO+eF4JFcTQeAzLcX7Iiv8DoU0Ir6L88EnE+Iu2qk8C5Y6PRtGiO
vMD9A/QqW9AnQ4z3dUIvLrA0KQZ9BS6GXAMvyjXEOjyGk5szVKR5BQC8ilamy9XvLQkbwQdL9W8w
j9zKd1F3LOe4cZ3fJHZZHK7a/s4O9rDgj4Fj/wmxqg5wQxckhVJL9VgpHf/7AOXt67ioY9xVMR18
QJjvJTGeoxz0Sv0B3HhouzifC66cUaPxsdX2eV7SwM9V6JYo3DxMxQyOTUBfPeD4fZryqKOvVQQH
u5hLDCj1+PF8LLSO17PVX+2myROZLH4LRWqRJQc9uM10rtEaw8Pp5c45pNhMU8oKBk0FVO0S8bsI
OweSOpg9xqSjTVCTg/FH3ABFy/tHN4wf9oUyhl2bCxGBETq2zU3dVi77KK9W+s5SEdw7rZcGep4O
rVZVEsYff7diq0qtg5HZBGrxPa4xo1hTWmhi/mRYpz0kgPrEVxahfYclbmtpPPyZya8Ag4IIIcPW
A5/3+IX+qLdwhCEyx27kf9A7iU+m9ZnfCd4dUhR/SHUZXfHhkqlgjn2sFnUsy8JF7bHLtF7EkDA/
mWic7+X9jSVkYFY9wN1XUnxu/MMNPpiEp0TYK/QVpWuPhp85GhwHkTRjfgL3ik9iYoohQpA9idTt
+5xzitxGuwjd+aiZaIg7LTdfIl0IQVhQgUemb8e+x9UhNM6t9Db98CQZZw3/2mpPA24bqMujiJTJ
RwcptKS+Sn3ENxvFsHX9amfEc+rhxEvgvgwROxT2q7Ukzc8CUrX/LDRiIUc2Woax1ElBhmM9bN1q
9TqdV70oCkACFqReUsJQ/YW9tWYEyjE23nO4vjxi5l/4YkVZWkeFeRtS+wKbDXsGoO5EjRdqCjWq
BupZd+o+HkztCjuR+cQzSoWJiA2FbjuamWukDHwnk69wSusbtkCJkvhisu4s82YVqJM3+E6sNiju
EU3a32DIGwDAgV+qgERHYJdX3wBYEVz9NGXr9aiBu6TDHFRWgPgV1NV3vBeleUBbMyd78JpQSdyz
4vy+QSBELdX6mVhlM7myCzQSBLqOyhFfX+64bsYid8FbZ92cuDw8+TkjWm3az4svH02orrbsVhEk
usgtbRcs5X7QevtNAKIZZBmmIa+OzD2JmZUdsj/dUFjiHxA5bGp6qrP71PwDVE4zuhrHR2Ggi/EC
nXZ7LYCJZdom8MJ/hVpNRWxYFRb9UP9r4Bs+H8mwkFTsh+/tzAftTCBM7VOyR3L287Vd+Z26K7B6
QjUUBMBsg/7k6yEPmCwTSHPx47IkIqeonD89Vb0gZslgJEffjUToPk3OaB840+5KDVhcfbpKGtCE
nUCIm7EJGZ5XRMsfAN9jSuETTSbM29hajLEqpESui3YYIpq6Og3uaNxWgw4pqhU4RYxAL6w3wMpE
tyNrXWxf6IKC+Fzk/ZNoOgF+vu5vAX3SIYffRpakPm5HJV1UejMGziaRgg5vgJA0vnHfW61Mp7in
rMDARpDzIWkWeIC38Kct15bgQmQNZIG2OYw33S35ERVtv4/Fa1lFxP6HXJY36qr9qWcfkkZ6JxqP
qPUNGNDLldjZnDkxw5FG3w9knm9qzVBGjgc1zIjQRAap7m/9G4XZm/dulwCPs5ljFSnCFtnTNyH7
nOnMTBGi0AvywRrIfP9PJP0JgMpiKbV1ZOWhXYzi6iNPE8anysjx2RrAUe6A6BYEjlChk/gI5XLZ
zA4izlboYOBXHyscJ/5dZCMCr9WkSYRuqaM7PCNjXqRuGeUCGiHPCrSIHtXRTqE1ialyCfB/O28d
d123DfXGL+JTwSyWeDFeWJMdfykXkQ4N7cJ2SY7JOmIz466icHjqYhgTgfuPTJDoh2IVCYkw1vcH
JqZQnk+DFPRTRDCcPPNfX6XOnK9V8eQp4/KEqQpLcE1yS3NDBbK83bXeDBjvoUwfKWWytj7ani/B
TkB9MQvQ7A9qJhJms5jBbrKq3s/uzxptLrpT+wjyjxyn9grLubIJOlghkqvxzs4eTUj7Sy2YQ4rn
6Y4kcXJnWhtU/DTW+zkAjV+z86kJJol3acrROeGRdecCuTcF0qslxV2FJ5tXDcVMhkDMGg/hQN53
dLxsf8nY9N5pBfxNqckhfFXD/zPuy4nqZiiNdq/NvnSQxQjD3UooJiHA1sUMSXmLX6Zp6GtkNplq
qtVUPsyc9bzM2DhWQXEFXlZt4Eza6E3ta/frBUSIrK6sTi2Jfg9+GY7tE5nuxD10GYGwFmXcuZvR
cieg98Np3/uSd6Nusy45Zaxb6LwL9pP92xspMnHLtkspRBphE85fnTYryLPkpeX1OV8XdMpbQw6j
nACXEgUwvqAsgV4mDp++S0D5/WGudC/ri+zWdiQTtRPYmZW80S8xbcyr1rwt+G/n2pYdk0/uOZHW
sOa1cYWOth5VTuj9nQX9G1qUaFmSzO/92DA7eGOuKW94XSa+s4aaA5cwR4IjSRUfD5qgnPEHzt7B
C9CeS50rGX0phg2uLVDColV6x8CaXZGCW49kYUlOR1XVX1hVzxaNBqoasa9V+qrSeF2gbBUTFWOw
OC1/+wmB/79B0Z4CLta+WMqCB4zQ5jJy8lp2Cr+FVrc+kTi9Szqrs5cFk3mODWcIWjsi6j3+FYSU
Br4ylhuDaZCq4y+ewe5ef2DNQ4dsWkAR82egkSb5qQk4QRcbMw4rouWYrJ5yW79+RlbTVa7BiRsj
t9UGbb68Hm+oe1Y6V/SSNmXbji7Enw2P6nRzbECCVJtis8SPe7hxQ+2HVvhCzJYRcscfl5DH9+UJ
bVnimbQN/1l7JPClN79mIsnKB4zTTIIRj31zCV+Ta9BQCvAQC4t6jVfJCPDFnj8QxhbN8+nfiAoW
Bb4lHq3ccg8CEq2wDA7SsiP+qBOue9XjPrdFa6ZiS/O0cOPP0FLOvsYEKLoT1fhFw8xtWv6mKQyY
YX5waSeDxDXJcibw6SNEn604qTOmd45y8N6PY4k6naxUQcIb3rV7anC0dEG1l5GvVqOGnglJxuXy
l9fcfhZp2p92bsfm+3VZbuSK2PhL/doIUdRwSH/b7rCBGQPM46mG5gPLRg8AL2TK5GrQgUEEiUEo
NqupaTs/zKIjvIF7NDhNC0kXocanWYcsXlaMCnQEegUID1mD8kZmF4eCBOTtFk56vSqQKuBP/A+X
PzX+BQz1I1XFc//1P+VIlv05KlsGFEaZBrLj1RMof8hc6P0bSDKQ5FGZt9JkGXWSmyVBAvTMEkm1
HBmuPBkqFDmG5k0/itEukduCjoY4FNox3XFTzTSBGMF+/xZqq3j1tqRa0um93vGgkqBRQ2uUOdAn
aGcjmGaWAT7+f10Jco2WSpbd3J6KHwI5LoTK+nbJ8+cmWAaT20tNVpG4Vio8G3Fb+5X7l9aV0cA2
JfmrbYTCEjM7mc9KS/ZmOxmJcwwWdc/8JLJVqPZyPVt4PJbMlOvkTc6C8wAk7ZRwbaXG6+r56L3T
lIpQXaw9mZh4Ap9lHgs3oI1hczQQt0e7EnbhFM5wLgxTNwozh+dVW/SIma+ZX4icR3W2H3c6vt7M
MIg+DATBVP7dxdhhf345B2nmCTlD4CK67Y3mqRW0I+gMvFcZ50p8WJOACCSVe0zWmanXef/u9fsW
k1SZjKyqcq7ba/g+CM4S9PLiI8sm6sDmN85HehFndxHNT7tL0Z0IJRysn67gl4BZST2WbOc077wD
9TdcFroyL4KN3Zr09Jb3HbJ8qQP+tq6R3XNw+4u4N3ohc9MS713F6oRIYqbu7d1FodTCVmI7yBiw
U4o+DF2EB7IVfh7wtMTVDSXVlyHl2nTG8DEShfqZO+Lq6IGaJjzO8O8uikeISqrE0F/ewq7UxvVw
afwAWLVQikQolJidcMLOfpWz/PW1Sd8Z2XuqUFetrlrFV+gyvYnG880PZzaXEY30DcGgX5xeGEWo
k+12SKYgPOX71qQKZihZuOxuwJn8lfhSzKUCKuN/HWMLC5E5FHWhmT1BVGxQZleOrm4CfJrLiEX0
uIOll2LK87+Ea756sLpxmWuXqthc9H8IyfjkmmU+em6XeynJ5LvprRvZxTbUjzqjLJr8cdZtq/K0
M2PKfUyFsFF+8L3cAwJarn07o90jdiBCOxUO1WVfM16i7SGA/fXxGlwUof6mmUUb6kFarNoLBu4f
2xaaW5GnjS+p8vzlZV7f19GssJLiov2Vjv6Hy/b3TfH+pYpyO/XoTATFRZc4Y/WvIec/oNIWiCdw
oUmGTvUhlmq0gx57cLtB+4wEaIP95LQELvQTOKTLCernVeY+wP9aKwt44hM8Z2Rn2k4zbwUgKj4u
hIoQaIxygHGnYfXjHaNlRAzQ208g+RkG08bFyAGF94wwCY0+7e0rADJJeTPX5DI8rh6QNBg9Ahzr
bXGClIF/vnMMR3vISZH8DRUUFz1K69sFMxXoLYAb20PFb9MsxCPPaZQ0VcMVRjealNXIKiD11AvN
wrN29cliWnFcNfodbcIR9Jm6VmcHrkwjtImoRIMRuu9yrMDum2VEjz0nidOe6kgH2ZSHEeImOKD+
hMJGVq8t9nqQEPoIxlyljxp9Wn5nxfGL1d4SFoOyF8IIOrqJtTtfDHFSGW6HilpbQPBFM7U5gr2O
51sJXqhxpfPd+pFYsnbqCbu4pfYQ6+EE+dE1y8iil1vmPlmS21ft5Shp0sET8CEkVvRHZ8Eqn7gD
G3WQIG3eW9HbufNxxHoQ8THaSOxATu60WUea475ZgQJJz8ZUAV9NRqe0XjG8lTAEPT1DY+Hii9HO
xQ3+z6NWLjYtaUqF1jtiIXRdSPOI2Lgu1hjWfj6VpYqhpd6JMXxZ0EBfCUY5OizSPmAKS/3U9irK
msVHdwafMoGVTorBviXFRg2dwDENCPJR8xC+atDm57XVrOM6E2qTU812bCVKJrrR//S83HgpMlOl
7T9JN3dfW6TbaAppwu1n3ejeU+YDWvQSV30x+pjP2/Mf+m3pLJEPrpeOC2sm5KOd04fEIatValf5
1DLuO/XlzY1rOHL49bx/qS4rhYUHAF/Ajc0V+b4xWhSwBX31EBq2LbEAh9gGtMXeuwqoNhZASuVM
XQIGotEpLAUreO/C2h9CnbSWmVZc1KeC8kfSUsNJbEayJC/vb6ICPK5puIk9ZjFfJpD1kenTMjCo
UksuJT9ONqk55MsnNzML/abTLbR5tCV67dIUzpVL1MXkFR5vVley7cUWt8kMZKgQbzLEJxC8PYwL
OzPoHCtErBEk2o7e8BnqXWkjNyurDWG9A0JecqiHXa5TI1QCwSbMNF8a1V3V77QmcKeXHrNoJOJB
NPVFrydOUKsaY8G7YS+O5xLRuCRrMIDoLKC3tXOab3gWLGuKXv/DkkCq+RcPoS34j6Y/Ljr1t3Iv
b2j1DjegPPX3fkI8e0j/oJQIpBGRWa0BbBOWaA5T12L3p3FO9GBMEBHM5kJvgVos1VzJsC2/odQy
7Zy6aeqncc2nO15CyoyB0DbaGhwKoe7i1hcMas9uGQKTQRnsTFiKb915hmtRjWfVYsAMXrobYaXh
Q76rrsCvrahFQDK2AMYV5mkBPIV+OrhW3+MxcXLBn3G+9DE/Izf3oUY8khvzic1z3+ymRDZFJ275
mBT6MqVTV5vS5titIUqjfumodbeywfzsOlYdI77u/eUrtwo0xOPgy7rAN16l2zQjIAkllNqmY+B1
GSlzggJcriGBznEU2IVFRxPlYT/DgPRIEnYKDm/GcitpFkPBoqF95qzCjgZ1VoxUdAj8CIUnK1d9
n/2AZ3D5XGehb3FjJ+ZUF7op/ogX1yCvqioboyYG0pZoAUJwm0HAi2Y28qq7stkN3W/3ptEaOIh8
HQAdTDeJiZOkTT3roKwsnjMIBQENysScvUH1Lk+gY8XjX+VEZIUfhgk8Ymh7BV1uOJofRJpF2w7N
/wSQtWE9WeYN+aKKEjNfjd32Jvd2oh5QukAX8SjMCOQf39PiR3uL050SV7EvtLdxz3wptArbv1Tv
NEvK8D9TSJy2pr6V1Rak2XYT/gO7BUHFx6PE3+9lJ7lq2s/pL/AwrfHbTQufSNvQSy/dJtT/xqDJ
R+0TXyB9+3kL0wPcsiny6b/Qb9Wks2WIX6NLcHi6MCktr7SdLDYrGJp4z5eA4Jx8MT5B7UXfj9u1
DCs7SaIVRczulWRyB9hsNkdEN7/GMWZMSWsgzJN1KA2FjNzCQAO5kCZ8iIefprniHvm03w0fCPw1
jVmFgSCd8uYS0x6aO6PPhBCOxNM9aELlkMD8oO034bd9FJRWjEPnDmzTT4b8tXc/jzhdS/Hi7zXE
K6WpQXOr5R7/CDb+luC9F1KOg/JgIkErno3o3QrEz4eJOlZKW3eADIZzKstzDnG5DCAuRFtKPUuF
I9w7NGXk1ERLb2di+ZOI5nIb8pMaJu2dOzqbZ2gxtOy3HvB6bC6LcLN52P6ry62Dl+8Y4AMzznjO
wUaMmd93gLPK1WoRMdF9COaN+EMXRhpmH+RqK1W8VYvArrmOlCJzBgJubedeZheE7Vvr4f1qrvwV
JxDQiuFTV/xZkDItj6vPrZv38zrKYp2yq0qSyrLMeln2HsnurhL5/e1qUmzvlJMps+qjaX0LeRp8
kGZCYkyUnVGAl1kV4WC4tzcQLKo6/anz5I5dNBswe+RlN9QGiFYf2VUkJj/yw1SPmQpG1YJoTkmz
nLUPGlyNuaqQABfey5XdMyKl6x1KuroSuCvQuJ5roSICcQcZrhrkwcJZS3+qfeekgwwIzQ/V69y8
sMDAmMhRdDhzv02grJr7P4iM2rDBewx5J/Xfe8HjJGvzv2c88gKzJQNhlFOL5kxdvlIROTLVnuWN
/gtOmETl8+pVYY+zZGbojFgfWni5CAwIsaEPf/gwa7+RNdh8atmKXmj2kxAdDc8ejLs0fhI4o/7a
ZSQ435LnzXuSwWcgoCgPlwxUBMVm77UUt1whZYdPIh2F40tiuS341eSMmcb8/dPP3PbpvZ5LWrpc
AApyXoaLpcodmapf9am1gcG8Vw7cjyhCVqEFurdUhy65DtvzmVjUcWrJzH28UTFetueNTseGNU0G
Hc6003WHFXdaXO4wORrca0ASmQJenN/+Pbh6p+64s2DnH47MnxRCcne88JntROcUm/GlEeES9HMQ
i4Hjz7vPwq6SXIuiXFO8KLkuEDQBmKNoAwRRiKSl3uNiiMQlAwrox52IUHard0GdhGg/RJMUx54z
Xh7+6Lw/KXxa3w9JeEWDQDlbKIZtRbh+8lstRiBMGlngSZdX96gPfdRBn2k1TAPfPUglDrEd6ml8
OnYlZus0Oyk7Jb9DTXahuHEAvVUX6TrM6n5ZZz7ytqnpesyim0ULIN0UKURLBhcyIKV3toLLb4uO
c3EycrwQ5JrhdcD55m38ov9TowQfbnumdlGb8HRe/SXiV5tHCDG+VKWtufADyyWcY+ujEHxL15GH
B5vYxrOiobXTVR0FBd3qzQbHj8hiNm8iVN7Zfx6NcDsyeaoeet2V63/8k0tr98tXj530AWNhwa2C
/zq36KK7fpFQCa8NcBF2eDZ9ZTA0IWMdaZZs0D6Fen69ikOuakNiUF0aZwb+kvoSBG/+uIvUVyF0
ou8eM5T/7TRdPD4vXXOogehrxMYhBx3Akej63U16fzH+dpp0D1idqzCfl1/kp6amfHgzEuaeCISX
K6Nzm/Hssp8T3OFwL8pjjwp/UIuQhMKqCHtDAeee0UMhFNhY2HTfYnm1Pz+hUEgSo88PkFhU/OAU
E8VGeQHFU0anI0Uc2FT/0CRu/PdBZVauWF0DRQ8LQuSN+gq/Bpd1euIqKdh7d8IfRlLQ8FXlfdEr
QHf2wbrvoACgJBV2QU+GpvMBudnHcUd99pRA7AJdoIu5eSbIKu5ue+gThSNFEfQK90PmzDiKv1A/
TGF1l06B/3CbBt8ElVEHlDj5jJF+w4MPIqV2WKlr22ox8e8FdmwutAKDeaL07LOwUzbryFim/H4L
5frMSg+7ta9jNQKemkaqwPlKwP0MZ5a+Rx+zIQWRnAOEZuMopC8gRB/51/gdJ3mztaqZEFv6g631
VqvwhC5K6X/VHl2fqBQ7Mf6vTEochuF/tr7hcb+HzeCyI1aLQg8JYCPreVClOr7Tr0X8U//kWTBY
F8HBf7gDBdt/B6NjaiUfDZdU8SsQxWJfPVU06eAFTYICXGlATPkEZz3T0ioUKErgjComB+qkyhN3
v3rvmx7k5SHWCCLfAqYjwBLtwysJFSnldny53K49xpjAXEE7O0Gu602VLGrbPplzO9UgA0rbjSSY
f/15REQHvahHmxJeenWejab07AlE+/gH0cXJU/5mcctaN6Jvv6OIx4ZDSqY1YXR3Ff1CBdHO9KjH
9IpB/cz/V5iUPFNUI7cVOhtfniYQVU8xPe6TEwQ7PWSuW+ZnAQIm980cdHjCnJmuaJQd6kdy5Yzd
ctxyR/JK+n8pY9M9eEE27tQsCm1kzww4+2+fiKlgquKOigMIf6xTT/RFkmKX3k3zFsdbfymOYb9c
o3WVTrjo3xQE+tptJSO71YdWXrNIOtSHIr24W5I1yccKL7GKThNAegWCEiegZqpINptqKdGHdStG
OdF9RMvjCr5BgBRp0HCPmstmaIqG/ynS5zHNjZTtFXPAj5wLhD8WVxxSKfMYV1c3vlUQGgsLgKw4
Wv5gsfmrzwvHln7ymUWPKYNTCQmzhHwj2Btqgv50Oim+0HPryLM/59kY80AApj93+5pz71iSOKYk
XFON4Fg9pwvx5yk7Afjr/TX1cay/6H+pDP3eqTaebiZjs4N0pQ7hMVgxz06ys4ZvwsShBvlUC787
ZingR8S6LYENsKBK9MsAkRF64FpNYxianOV9EmiHcwqnpUq96x6x8owj6rwaUlzNRDbZxhxa3PZO
sH0Os83URmbfByoKwk9z2OZeTmB+DBHhVAwfcGo4+ORqdVFt8TJFuXASsJV4HtKfsSlOFShtodVc
Dme1rL48D7O1LrQsiLPXtIxGpvK9U9LiUxRuwwd4xweCthPEnOsnLWaOot+XE88UQNZ4r6dyxPOI
xvvd2BsSqk/8xQUH8FIgUQ6GLRbw0kSATjaK+4zrRA1PqzNtYyLk39BhL5BTwqxP/RiOy0LJZZod
tlMxUoBJwoK6ol2Gj803EpC5WMVObhyRtx4noEuqRjfuuffPm4XHHbj8tvMV2GCQVJM4m/0AsuII
22sgxb5H64J29V/g6eZohZDesUY/R2jPrpzHmPeZfCfgUXRM1D5X1EtylG1NpOYV7nGafo0SaFq9
xaKfOG8fkRSJveYa/4JSARIJZOYmb77B1IHSOZt6pCYGXCrlxoaH1SuugLQBnjnfXE70cKCAKHli
U/ZqYYSkL+WE4FFfBjFuKKBonLqGJtvYkf4WahOHzFs4LYrKJME6xpDv2eCUfDSpJoi2393Z5Ytu
gz1AdIQiPZpc/eL5buPv56czw5nBYcgOi9qIlh812P2s3baw8kauP5eHa7VuooMyaXB2ZLd2gaK+
WHBdB4TYLLPv3AIXTqyTpg/Iq02DQTfrfMPjHOmnQxbuKw5k/XXzinaEYi+dVJS59OPS046hpm49
znNhSouhuXhpBINmF4xLrC4M/R1yCmYTrOYFEqq6foidXv+vCAVbK7maqi5XZ2DpskWHwqCFJ8FE
KwTyFWD++NcW0IGfN+Mj+PttAk5Z2nT8Fj76C7gitcFgrsySORXB3HZMegBdQg9ZpUmejnn6UuX3
S6gaXdgij+ocNhRmySW+zjDDKi/4SrIeH0npyanoKSkPy04z3WLAfmulZen4y9kG4Xm94xDkzVlF
CpQ1O3creHb2XylY8LyVlhBA3Kns2lxRXxLRPVxRdSkgbyUlOC6tAskb7r+8FQJIe7hJ6YVGF7lf
joIoMb2EUIuety8cARJMMbMQF9olIqiclG2y17QNm8wqcl2rJ0vso7oaAN9nrCagJZ5dAp+Ch4np
IHguBaXhI5qaobbaTOAuHQV022o52Y8CnONyKdE8AxfEXum/Q/y5YrIqeAtQ8YsM97LOnAcd0oBi
+f3HZSgkSFB0y+dmMtfbsb7RJTBkFvvIaTPaCwQ2msUL5Va+36xZhPrsbG6ATd+uzmSScEIPJjGM
Dh/+VEcZrBXgJku+ax7k9wlz2NPdjc9xwTNd7Uf951Kloqd372JPZYK1+Mgap5yHv56fqMYw5CjS
BiOhkQk0dcULumDzRNHgLStONqAw/oXDD2yfrv3HJ/YfJT5FcwVtDFBX04fMOy4Od7dHPni38mQO
k0Iun0b185z7aifms31Y866E6OXqu+LCNlk23ORsKgBQeRW8QO8a0Ao4WIYzY9Hn2Se7eMXyD7qD
JKVBA26iOtqbwDlcz5kTUABRMWfaY9y4hPjHKAgnXufLfAdmMgOH7wGlvYhXONepFyK4dfHHb8tt
njYarfD9eMl6bzXy/2MNgF5nkNFQ2Y71/gAxrdWI8ZjzISe9vA+eqSl3ZdZf8r9R4Hix1FO7mJF3
nn8jQmznHubz9JTngPSFnckJct1UAKFukduyl+eBxZb688fNk4zFAnY5XeRxFyNDkCh19qwmkIfm
If7mEHYm5KZ9Rp4sCwucgFnCgJBQtsWbFEqR0EeYq+2xR+cpPrXwSZ1XgdNsmhvTyFaX8hWBQF0h
e72ywWEpoqGUDYsc8ixHWulUcbC9lWqWScvnzsa2vwhHPMGRfpOmMKq+9Uva3FJR3Skj98uc+Ln6
mitKKar9GdoLIwZFyyFu687yaoZF0f4awIsFYW42SEHX6Ss5ULiLCQgMrPgtJTypmv3HYxDBC/Yi
u6GuKUn5XHkg4yaSH/m2w/pgJgrnPPBP1gT1+yjoYN1YjrkA2pcOsMGk3PBmdXNiFrdjHDbApkeN
irz0AhHmjFiw502Wh9hmzasnExThXEzBii/b7HUBthNllAN6marCgxs33EyqsV0wSYVpiIq1nYpH
GW3iZlT3ERXEbcRICE9T3CrRiqCjqjtmNQtO7oOiNKcH28YbcV6MkEQW3PtaMUDlWaRUsxPoXWzm
XE2lCH6p6QhrSLhkw54WfP7PfuUj/5KHHjgGDrR9DPlMvfGHZo+DXG9ga5vdKxWgcJmZ3op4hOBc
u798Z8cH+Sh4lKm5kXRb62E9nXUoPOhHVrAlN/Rbg3EWwKyhNgVPrm2AIS17pQmPqYQoJJ6bZpGw
bznbbc7dfV0pGQaQ6HrNy9QlSTma/MVtim13QxtmCoPIHWYzHbXM1AT+BYdaEYqDjN20uq8erqUL
2O/ym13xt2sOa+IOvgIKCvsBdSTq/6DWNo7obqmh9+J9DzkCytHG2PHbyAwBOMvXL3LVO6audJRh
wrDPwHY3xQCfy+71l8FhPGdWK5c8P7e9zoOFURmvfnjTu7WenjiDIJ5MlmfI5+W2VugEhhhf3Hvy
Mrh9+PejYGLTziu2sNgbw5S1pgzl4UIcakvoF7T4rG5QFYsvV/DtoX4HKo8lCk2akLUGnk87LG0p
MyReVd3UoQ9ZtQEhRFM7EA5iwC1dgy58bikUShh6Dy7L5hCx7EhPLLh79y8sNSEIk5ZB1WvMa18S
59LzoriKvX1mxzb399JhuPpFIh0RgzEYfS8Nkn38Ge73j6qg5pdFhlhs7xM0KgeZZ/8pTAZ/V+f1
QEFMUxfwaAxJQmEoCsdmpxH/xIVjRZdIjwwhhArYlALJIHC0moHnHQhJasIljW7GMSjbumxZQdwX
UPtatPdG9yrGBxwg8xmyhqOlZ0wSKzZrIRk9qdFZl3vOriTOT+Zzc0l8MnpxD6lFy1DRhtGz9ofE
f9fVGY2KMu4s+F6bboTMHbz58onI8siqv+rrqHJrdycGwn/RlyP5PqxiM6L7ani8KxeTaFYYTKTK
OWoBb4REFl+BaGMWQydZESFvroWyBjhHtKbSG6AX6r1v5LGnQ5jJGgDsI+rqKLcekYo2g55GHRz2
xvqTPqRVU8ArbXqGtuHiOQRQREYLgHWJmxLB8zT/nmxHEz0upZNfMHhMKLFJ4ziXe3dGsEroVpx9
VcQ8SxSYJFH2kH1KUpGLe/u9Di15PJpHxYcy2EwumnN0xuUiy2fPP2HCVtUdkza1tln1v0yJ8AeB
OvpfEinOxwRtD/vD23cll9mkf7+KsJD92nvbBDzHWX+WM3pdJuxYhnuy0bVKGJaT4GqUlBpNPSoa
Pq5PxrYUFuDREdvfrkLhBKDnyDGV+NVU1+NLwl/QcvxpOWVxwqm+kUyWAAkMJkNQ+WaUNg1b8JdA
XPuFVfWETci6XDky/vqEzxnuulYtndZi5fFfG5w8atMQW+LnY3JGSuQSuUw81Jg3YeDH/mXOeeXe
cw88MVLU8RpXJCpG63hWZRvg4REe8Mu/0RcX0VKMWSIdnybdf9IH1GklPWfmMiC3WypJKNN8McfG
sBrhbNk1EnGfX8902UivVOjd+/KOgO9nGAhjlV/sMYjiu3N4hd4ScvAeZ2UEDHRmASl06KjE4uZ+
F3XZJ9VjOQyI5T6xH1tfM3KQwIRy9A/MqdGpuI2LJ2WGyx0VDOEnOHppDp1LXYUnFvsmBsjviRFs
fiHEmdL2s6QbY/S9ROWUftADxFuUNDvtIYDiRDaz6Ic5/zXDCeeJ55AcN5JzRPa8KS0bCsyvZbgh
LubSV9VDixz9AMhfWduyTX8/DiCk+TMrrrkIPzjf3fF4s0U5bQUb7NbSDQQ4HK3VmPF23NdS3P2z
eMj8XoH3djfuv9Smi3WxUI4Wmaj7a1pUR81ztECFrq05TrSFkdMip2/B/0zqgCiJOT1+DT8wA9sI
ggE6yrQ8nzww+Zh7uiodXm5dYGLiRFLSM+p0YGfsEZ7N99/bmNDT39qYX3tGtf4I/XHa86BTgBu9
lVAKPe+NIbkvB2NOAtIzvUAcLWWhMKZz10RyRCKH72+mfswVM5vFeaNIp4WSRc9P5tcYdhfpm7T5
AWwWhvUrVgJ1tdwSVGb3u8O3Wux/+6Stdtm2g8zeZZJapcEwDbJiGchkgWZ6MiAVQnbVph5wrptV
4IQk+qDs3hXesY0USVkDqrRvpluODXLLDG+pfcrbV++jgsuWzoK18t1+t8uMApGxo4Fmu52yIbjr
BdLrlf+MDSXVFl3I/16eFd1XyPbSjtUrxDSLlUp0uCpCVUc9v1Nw/cLqYDaxY3nGuuOyvjkar3OQ
fqIpoJhPeopbvi2TESyJecqMxW6OIYNbIlxoxM7GDH6VXMhGxxIsZAuLv2MbZMai8W46IdcH20H4
JrmZ/1wTSG+SqZ7Z9q+aeY5n/gWIVIhGCDuy0/xiMpnHNSI7+kIA+bpcjzsFZZ+9baTm08/A1D5d
H1jjyHYU/H7aQJ8K5VjYhjmLdoKAsg7wfWfgFOdGvBqNkBC4mFuHuUvmlKn6CV1IlGn8P90Jz2jc
yDj/qWSbDijUvVN3XZ9/PY8qgIQfPMS3jVDfVSn96yLLC4gtt+hZE761/xo0moPDQSThixOiPnNA
LW+VeKIjuZoJDJ3/HrMnLw/PS44wdBJfH0hmnf9+pf0t53w+XXBIHTzdEAQ9mF14mHlb5+NH5EtY
wMykssm8zjYaaEYks7rSUGNseIco4x8Hu+yPYE61blIisDmARLsufyg4yovkMmyXy2RA0ziMSreN
V6Fn+4qeY6wlvaiRzRnWkg40CCnFiFwghI+xBxCybLRK/o26cdlfUvKriNaw89hiBV3SATNLkeOq
FVZtVaRgvZsuGP9Inxm8T/9RrQY+YFkNQKFBrHGN3LYMIQHgOb8+1l/i0V5oROYm/pYQN0x1zgOr
rBQttPZe48OXInmtX9hWyDXelNbOOX2jh3qYN0DP/xoNYajDcku+fGdjiggRJ35LN9SKJ3Knr3Z3
5BR4ZnNjU3Xu3HwCFIgZQdDzi2sOOH4zxAeoo4kOAIp1wWUNK4PBNlwLkCPGKRC3hbwko0VI1oe7
q1NX9e3yRXYBgg+ExTDwkvO9D1/yCsvLxwHaZ1CUnN93pO18Iawvwx32sm1tlCLrgmOEJfxplQsP
mFu6l1vlhguiUd//WcRCiFd19qwzF3N17/CMkAACiQx5O/wF9K5xPW4ybDoZ4wnI+tzn1Eu5klea
HQby3xY9EwhGWiB8FoBBZ3pOCrloItMb7tOE6Go6R5721zgEGDoKDhs7o5+QwCy5VNS+g275BQdw
EIGoo07aVzMC1PbN+4hLzh0XoHykhM9WYpf0/SbmooESEvnOAueRxWcpq72mvBOYCdGDV9T2qau/
FXqx9yt60YFE28eTYA6YJMcAiOoZ5k/KGzovyyqY5AFx8B88IOp42bHg5LHfQuLtWnuIzyh6tho6
kgra8nFGOdb/vjuYm1cdv5QWR5bXHhnJwhRsGsSz7P1tkusBg6lIsY7gSlMvjnUEWKJdEMZL3lIU
ACXdQ8Zc+dotT/9kggXQcMvHPcF+ZXq+3c5AijDJGnoMJfVW/pi7uKLDsYLgtkvnnIGEG7KSYyux
lXsJoOV7crhAwd7ChZhfz8vUoziBwo2CbuqGn8FuA9P88QI7J6tr/IqQas9W6YgL0rGrNILOA+Cd
ix+DKW4eX1+UMOlJ5k7LwguAWMSAfTQMJppyE77ppepd6iEqp+uOBcuN4INKagwi2/Di8YQh6TC+
5tdPGET+vVlGzB+QTeOm6sOqZ9QKL6VREvpdpLZT68wFBbmzRjwJPz5UF2eUGqjfotb/F3l46I2p
Z9TeHg6PVu7n4x6sciXgb4hmG9KfQH9oqdz6J3brYorRQgjJCK4F7tTf9d+3DH4Y0KKWXMvVSBNH
rPZ+qkOS+gs1AGZiLAvoNOMidL1Qj6BhefyPCsK1bNXE1JZFHCLj4kcKXj5aT8Rl0szTxLrYZ3A4
6LiOUi7+xHHUbwA2JrSqSZtI4tB/DXjmKY6fMAi6KO4zln9hSpVV9K2o4oxA0GEkLUsQ99WaQEQ3
PtZH7nyXqxLtWNWqTt0P69mSsLFaVl30w6It/nTT+zenDjpfuFENntDCPgQ0/n9IKaAeKOaWpglM
QrrhP2cXmOqwOModp2LGMY8cICKYHIYvEO63oUp3t6Om5bMeM9DvlMwKs2ovMb3oZF2Fc1npgFb9
nabh5l1rQiPk6Z0a7p46C82Fq47ZriNsxIw6176SU14BBMTc/FtH/BxOG5QeZ37WkBMKzzMXy3ZO
gLQ/kjbDSTgB8NhemvkSFJVJ3xvmnDV0LsLuwqbJCc247pHSeFE0CvtzN1Ak7AkFo4c36LeTmzoZ
0fhbpwicsvltbjCspu6XTLHorE5QQM3EpBu767t6dBdHBMIo3sDU8vhPVkMGHCjkRHaWxWto0n65
owwSNgPFXPJJpdE2PqHyEQOBEawpwkuUPrSnjUkdMkNdgn0p7n8ucynZED3xbl3kJ9lb/b8K45Ml
0uQpqJw2afDSvgwJzDhMZO1cIHff+Hvs36C/7Ti9QTRCX3xB6UyWw2qCLO3D2gaR7k8X55F5nb6b
Cpnv8mvCRvgF9eLJEV0aGyQo7fuQjaq6y8oxg8/tpP6aEpReNRYYAu1Ee/dY8vlP1J7EoLOnFx/L
dqxj1sBXFq1jM71bD9gv1ZEWertfV5ae6QrKzxFyIsdKGoKxaJJq6ON/KZtJAnYbrRgggGK2DI/2
CHTBIC+ndGyaXMaX/HeWZG6kSJ8qJVILXm9jClp9kTbKUvmYMXMdurq1Olimzor99j75haILN1/m
C2ZVKDPuBakZa3MXbnVO8ySiNJG5H93lVIJXBIWcAC8bu6EkBvhfNKa7R+oKux4la/sN+wxKSjgn
ecZrFGGrPvGfhAlnM5UgEItUqmQECSCi2lv5Vpacx7KwHj8SV8gMyk2o5N0ER6HtdPd7/KLzq1aq
cCRdQp7XDl55Y0AMPdkaNhIlX1T4ElzZgviZ8v8YWYaBSMMB1n5BafLTXYtsqjTboklgaph3pro+
VTU44JFf1qrbXcPsiDi2Jl6h3xjgGgylBzF6RQ8G4VS5vHboi/CF/3iS9EavWJs+fqkrzd2WEEyG
dP6rMSyh3p3nSlgKT8eBALQWPirdotaYkhNUiyVlnCtc6psZALHiKsb/wNEdtcDViaQXTVh/Ojia
pDqPm9soJ4YUIC3xq/vmaCKEuuTlOpXcw0eZlcbOIoqqM4uBcP/94kz+5YOk/ohgZaesMNUDYJ75
mo6Be2V6T6THV24Iw4vOP1QfO6VIpETp5XDJMzNeQf07P7Ytr3LAIoyhWEIxEzIF5FfeEdQm1+Zx
eKoxTUXb/vozAQKowewwFOxJpf7+wU00IZvEu3EMwnVydxocN3hbnNYmN5RI2mIGiwVgoHn0iE02
QyG8XpDj1Dr0nwu7zhkJ3x0bEPRqxOwrpEQSylZulCIfP6Kg5fiu9m/Dm2BueqybzK86Rh7Oh7gD
4j+yVSEzbqWvM8HE24AzC1T8AoUqam9JzeJUiVqBORU6dqCfKnSvLM2Q0LzbUnc0roFFXKMdNmSM
NBK6Su2pExDUMpIDhbcN7IRdDoWmIVuaeE8/0R/3++PuhxvQ1kdeel5c0ZhK8tEcMIBzlsZ1kiPR
TSbarcVTIEEf4y+T99O4YBa1AVCigy8YaglmN0MUZCIWmjoJFx7VL12Bypf6nNChx3NzbemanzwW
I/1J0qrRnnHzVz41bvbp1nWnz9w9TxlB9x7MiWizVIgqT/HiWw0rEANXG4ET1l6WJRh4XkCjjtmj
uHflLH+3oPi1MXShCv2KQ74wBmyOuSZ3h4ZkEZmDKGL1WGniJ01CnMROSiVY/ZH+IakkUZle36YY
sTKNQUNtEoa0v/oBHWmgp6IG1zP7YYD3L5xcp5U4O5rCRuVLo+zshLeDWPcY8mS5Zz2KmjrLUyyZ
i7BuYJ459go5+KpkYgOViFWy0RlRZOPlBiT5LdvGEj6KnFtJIaP7QjRstl/fP00C4zflyerd5Wgn
A2wq33RFdmqFPjNgujHCA6ntUgk5PXosj6eNRxyI5Pik67nsARTon+UsTlozzNSq0ctUXcVaoVii
BTP6M4FDrYeRAGCyUxvllylw5Ku5Y3S3KcWTCDg/DU3o9WshErosp1WnbjXn15v9VgL9WSb+uJIa
8Vp9fQ8lgSQyhpTm90YgFqiHQAc+uWrFnaXI83v14I+OsTlM7QSEAe+fNp6cBUFyKD9c8zyPhRDZ
PEQ8hmtL98dKJ2psGl0O8yZdtXVZxNoVutRcIUoffjjjrXZMHkdvzeRC+9lqVSbXs6TfOjSoJYOE
cQRCUFh5llQslP53YeKfsRqHidh4hzak02yqwU7TacdnLQhy2J+brUXFOvz2J+wOcLUC/s1UC4In
F4uCjPyCZp5ltf3T7m5uVCfHJOeBTBJJm5PWNpnkdMmmGMAdOpXcpgnPmdj4QMufTXXE3w8mNqgP
u2S62gva4Z7t14zYiKu1PggGsYzqyqca7+eoBkx5VSjYuDu9Z8ByoxwqsS8X5bTeLmRQpZzsEMN8
zppUVLJxR5VoccAxQExBquyeonDGzuDnDxynWa/I6HafMt7ZBalBGJBm1UTOhYyDLHRxM2kSl2TT
7Da061ea9ZAcCXkn3aZ9WRamLEilWHzpL8IzPbtkcr1cbIeakxe748AHQA9ODYp3u/x55U2qUS9Z
+EKf0HBCyokMVXGhLVy9MPjn5bv+MGZjtmhw+W3tdKmlMaDsgEh9mJbJ7XdLE/jyFdYcDw6fgmdm
fy3RH0MFTuweRZkUEJq3w+GpDOpQWuvNq7q+pQ1W3JovG40zrK10MNFwG8KOqOPHzRqKzaHWh87v
9Qz5cXZQqnPbYvecEKKSPnWjux7Nl9TLSgqPQNvNbLbRYD/Q6IWrdQt65r025kT7UbnMWifuRvAc
QdXV/jdsPKlI1QYLOcP1cpzGg3BJh2h5g5g2vu3Pv5UJQivxc3bBZcgNQYxKxCZo5GGic6TTjM8F
Zvg23jaoKVWMx6gaTHzfYUau2GgGMVltbchkone/16XF9WtPYz2CWpkrpGwewcQVhdcRSf8E+ZSO
UYGb11FgvACmoo8Qw0Glx9HlY6fCojWEEoVtl2/bJV+d3VrRiqoiOPacsTnOsqZYHuhKd1xEBJ/1
5IjKhBC27Rv8wvHACrsqy9HkzRxjrulosCnzCU2fAcyCOxoZ57i1D30ZABxTBIQJaAtGblP2bIiw
L8DzD2kGWI1Wx7Nzitkw/PDN25zAPwe58eKOEPtmhVglC2wdMuQZy+Tmujy/ZSeZItg1MSwCGvbs
HaV5/jOqdLYCAWM47+ZyCTKlWHdRc+aanFq+3gn6YP8W1EvRSxplxegk8US6JO8ibWh4t3wjhvxt
6PlO0oEmrJfPKf9N/MiEHIOhb3tNVUi2iP9N+OtjrUOslmKejQctyPhAwpb8R9FxLI3scY2iqA3Z
lpsmO2dz63hwJIJ3s7tAF46EMOISXW0Z0D623JiGaUxmkGDLlk0XVcwedRdtyIDL7WUG8mxkkUa9
s27cwHywWpEcqFJRRGnCfmd8u9dubUDI5lcbSKW8fUb9i4mFTDfrlRZ8ZBuAJt30WRYhAMmu48ug
CSCks72LlmOr1hFxagL6oE8Gay3j192fLjgdMh+PVN1pqXTPv5QUSimuA2yX5H73M3t4EzBJjAxy
qyrJ2E1iZK2IqyA2rKxCjP8Kkf/oOGSQgQKj9zNGjtqA1KOaCruMpekWIQgIIBM92OStLDq41aSl
BmdE8Xyew26Mniuj+kolLcvGatM3NOd0Kkkb+cVOq3to/n3qS9gW6blGtMztHIOW1gVyHv+mL6GL
+fgkXMJnFF3MNxmd4eFzAcVbg3t851ScbZfmnzyjfJI0J18JCVAg9wV8GO277XgGzHEoABblMBSY
YK9M4RMjhzoCW4rqenLRmUpQpglHmAx6jWtFYE8+aNRwPm7rpHQ2rAGohXjOtgcF7J4TbAXpF8Ex
Zbfxz+0zQZjddaexHPaBWMlvEQH4dNgV0GIWyZdTIHUOUdVed1jNCjRjzEh3GanXXTA6jzVl5FsS
nMTlwKASBfGDRfqyEiMTBR4jEX/b7Ienx+rQpbamsZNsguwAfVms0wFpgP18Tr73zdxJthWDJLVL
1n9+lt/zsnij/H9PqPCmZvZ9md9KOkgStOQOBS8VuSfkxIJwAKmntOJEcoShT/rAnK1NC7AOzAbl
Cgsdq2RjsuIJ6xg8PNuB2IMmPaYNyBygHYlTadcivHccBDHpVgFZReAEsjQZ6zFMTLtGurUt1KoL
DNZmQuFcj6qLh4ysyYjoWkdwEgR0aIAVVpDGPyB+MqeRxk58kO8MHE+FI1B9xCnBrFewgIh97zfM
NkWfPqba7KWVwtLUZmv/xXnAY5Pmp3jo2xU1WNRr/b0mRQNY/1BHFZQ5kw7UhOQ5Zm9ePxfbIFcT
shC4Iw17qB9LyzZgoD6lvqsgYtz9HjR2R4GupzbhhqmbqAN6PPtUxn+Vmki0FIxMyZTyqbm0nXsj
k1m0TSGXyc2JRXXgjWB+YN9apRZgLbiw4gkm2CciGBbHPE/PB8i6B4ZytfaKyR7Xv2mrPCT2eGYp
SszWI6u22IoDgT3HiTk21/BB72PBwBIzzV/M71mwL2awCNGzS2RgHLAwwuPCSQnM/n+pZfr+tMuc
AqYKzOKurA2wc2oGez3GGs679+shVRjbRTywiN14cx9nfokAlpqfPiyRcdlpI1ZRa4S81RmMcInE
wJFF4kaSToqgmtU77qfTuqL/PqQoDFKD8VphEfhWlHRZJtjyNurdEDo0bvXAPRMYo3iebKrE4P7W
GJwD/l3nvJ/NMupcunXSrZp+Chi4rj90LjKmgN5f8f6XrK3WIybHE7SRgn1HEtoMib+3NNZm2ePU
UFBVf6+maPk+9t14jL/1sdRgwFlueoLgK1LZW4fPPERUcebqnYyYeAWl3zMhBXFGdptb7DJA+3Mt
J54+fA5Kuv7JSPWbS3fqpN/2yf/0bBYHwewDhrbmuUq3VcmZw0zE61cTvoTToFfcfZcrmLI2BgYu
V4NHr8f5NtMPTLHFDsnHZMlHFT+8fZZCxNxYAnkx3BP6ET4Z/yGSfknb+gJ+0MEM/aFqVRHHQa6h
z5mJEU96GiAH0WXx8zFTKOT0ThD6yw8ixGcbGEl1j5Hz5XYj3FfIzExqn8OaE5ePewF9vamIas8O
CEZI/8laX/DrPMBk0LC0yNguQ8nggz4suDJCJ4qz638KxM1FYD0wyI7ZMVvzmqcaO/IGIUg6MnKQ
5AHYsZGHtDFyHyrgJQDxk4a2xZWxGNHUM2mm2iU+NPwzakh5gQMiU8mesKRs9nlFa8vDehS/tJkM
8OiAnriErjKOcq273/wUPNPDXNXG1nu4r0qC8ZzP6fJ7RC62q+8it+x7Yjx2DzEsotSg+V/eh5xV
4om5Ra9sNMpJhTAL3o04/fyU1D4nncRYfleu6D1Yv05D78VHCAom9jrm8ABLJ0smkylu3w+uADZf
sYBTG5hIq5qVXkN1YXYTHoMhPaGNXRWvNMuiD4iCpcxQ/GIvXAY0It7yKJLGoGP+9SCSnOkMzecZ
BfOAo/vme2fayqnReHtaqquyKBEO+NMJ0DQcnV0Xskt29R3fCgcA1YNysYlnNoXOwQ6zz3ZGw6Yz
dsU3bEXB+MVAIjOtbM1+5SeHZldk5tVos4Fk4tAJj0X+uWuBTj9u2be1wWTw9C/LU1PMjULWUrzb
qq1gn+0Mi6p2RCdOjuo+/j2elbGnJdqlEFUTtrmhja3yGM5JNdh2NwSPZiRf1Wcps+thrUUe1ySj
4sjz6DqFBSZxSB0+GvrdOEDZFN2zRkki2fOyrDXb4b+1fAg/4l9KQk0j5ULnJ95C6ObXrC4T1n/o
wVsgTGPXa8sLXXqLE4UyfOoBv07E2mi/B49sfo5yLPNEk0cdrjG3LQ/Xwtubg61SDuBakFS+3J9+
CrWzBMEzZJJ7mBQkvo31SFhblzUStdduhFEJV0Tl18UN2Dd1fCNGd4CbBIKkbhyTjg2RXdXPWBV5
kh1plxE2InJ0X23yij9Vod09Gfu6uiT7pBvY9D3yTjGsxsyH8Vyh0rJCaH5yEDQDCBKCmSenheHG
clkI9gTKcFJhAbYOGqk3A6LXcsmh7rFaIg52pW4AvtfP5LJnut5xFZ1XKt4p7rKDVtgMEJ876XU6
FsZV1FIKXPrCTWoz7//WSFdCC373jrYinQjPze0oX142TlkhSHZdjPeHJWsgJ8ovWf6eiNFoXBKK
voPMKQluv0/ki76vrN3l1YXnozt3DoZqBG2n1Bba5WpJ+n5vLtIGQvoQoo0+F/FvTRfclBzY1tCz
cVuCnC+H3J9MYVqqHA0d9Dg5rmahaZ9ibp0t6HSuOP0ApG2vCiB2jyolyPYVjRfZ9EvYdE8ecbEH
cDLBrjUhjzA0W5iLk+EsmKDfQOpLXoHRvZD5gXjkGqoYo1XHkFFGOl7Cg8gsjgAENjtHCtziCIBY
DNXVI5ynZphPO8e598MMfZp9QnIlmW6Vs5p9Rc15aO60HE3Gh4x7TVFYQKKy/SyZgARpxpE0S1ai
HMppRPZIC9rx6SQ2XezRvVUFCyknutv1fNDRlsQnA66qXK3UPbP9CXmRDTSYw5uiJJdxe+1g5V4m
WSswsG9Aywp7ngBXwXxIjngkL+dSA+wCzAoMC/iRrNsxz2gqW7eKGIldTbYL14mb6MGQRRZtQOdE
fhzQnvg7CZpR8HV/5U/yGn7eNuzPpUS3YXJBfEf78ydSsmj2qLBzcflPo2hDlVbGDA/FD0CqxDVu
8UrWyRsG+IENyIEq694GQx3sh1YmKHl9kGMmHDlqrveVm/cyq7MypptFmaOPOuqfC6glN+qK39yR
0mhfD+EGCKgZmdvqqoBc+AGs1fE4f9vwTOricotB6S1eKV04KmAiOzfNEkBGI7qVSX+gmUthoxSG
octVtIfGo34bWvxOtL1wbWrqdTghUgJs9jjzAy+PALyd/Ap77kaga2iNg/CwvpABkEsiB+JLiSu7
9+nT7aqJyf6NEbOD19WJMsLsln7SNcO3Jsxq7aONbj8i+vxb21ovhyYGF5UetJNOGNLLrdM2f642
m9emRriyJWAo0dXvgs+JXDG5l+zTfaHOVaExRRmOJPdkatpIWuCzLorPXp++G4RsRXXMYqkktrXG
B0YQZmsgjCEg3HYrzCw2UVmAjnIiV05b4hZP1ZVBjUWIoFe3YsviJ5cBK4LfTH1HRTTjxcCrIwlR
CO5tDzq9V0VMQLVks+101eS9ygQygtfuOU7HTy+49DbbLI27dcE2v+wV3dNxSekZJsQB0f2jStuY
6DGK5xW1k4S/vvDO92d76rHESaiahXqIWKt93C7bq+Bx72li+K4SQWrNQzghmc91JMmHPXRsoJTv
1h2TXZ4S4a/kjCQiVWZaJcl0+3iMroDOj2WFSKfZqc2TqysCVIlad656+R3W4O7VdLsoPyMGhPLE
tcdIgKDYasC+2NWLG40iA0jFcmIraPn3XBgioZQ2dhibh2ElN8aMfw+oPDryRV2nL75Ky3sPjsBY
zetuYfpUMR1HeYuMbUQRGyac5JK3gXNt/+VanjiAtbMsPXFT/80Xt/+xwa24gdmBOwVD3c5/J8pL
pb5Ol2O6KPG2PxZwo8iJJBxZilXpaiOFlzFlxE5GRlO4QXaFNI0BxrORrWHYrW1k3KTJbQW4o8hE
KN1IVBjOWDgkB269hNm8CMRhnlBuXPIqbASORg/FkY2gSOuLWKvF6JoKVKCaGm8Ol8ambWmEpNmA
KIS5rms4QFU883Tovq3nH/DL/geqsB9zZgyYWbTG9TQQKln1lijBITHT/Ti36sN5/HPHSa+/GAtX
EggKUPwswlKP3D5Ab2lej46HcLB6V+2oab8CtviZzN1Q9F1Thfo+mmxobPcfC1x5J5lTxERR+vCb
poCSmpiVlm+wsUvEUVBi1e7NnSSs3SbqXGvo7O+g3FOMYuehgQvDU/zwVyoB9Zh3PxqTUa0WGOKH
uPz79hw+u//DssrbPgDlWPz2tOMg+9KPQVlvsgp5eLC2mQ0bjJLYgzwOUzyQXB6lddCIdu/sGc1M
q050AzFIIEJDKR11m0+smYw+c9JbjeaBY3g72a2+l5LSj3qLHOnAO/ZeA96Y07VIB9fZdwlRVirY
/ksW9eRR4ZMn9agcE6M0JaXPy0iOngFHjmh5bcsdZ7CcdY7gNFNlYfY1/lcImJj3TGgEKaHnwSkB
VzwR/502nZ0idSVynqfaHlCabwl0zLnE9dtvr0YK+mb8tihXthW6N60W4EZJdXL8Nv8KLvmn64Lx
//3EJ9hVqRMC0tkNzwWyQhZ7NkbIYyXKWVQ9MP9QIGdi3Z1dkSeke9B5+C3kA5+Ax/uUegQo2JLd
4LDVuFb7dJSpTeziMqJGQnzU4KlGsbr7szeVnWvbZIlPrUPPnnAYcqWwJtpye1YwNxUGDAQQdEwA
hxQ0wytElZJxPA5T/mx6Auc25dacAFUsGwxp0JpF1CrrH36zvPw1d/rWgHVbH/AlDyS69R+EGCq2
QZt+4TtTpTiQXopg0uQ1PoUZD8y2QGACPBlqvfxlNj1G4geG/ZeFc38BxfGb28OqhxFnleVIdcYX
guWBVALypkrdDsQDWE7IL48woeexpGSyOsZyPTHi2mkbAMXx2pKNgA9lN4ZamzP7Uc4ZIcsIV7ew
Vy4x40rraCt/wMQGH5d2gsFujiEKwkuAvGJIkKD2ktm2ug8OeGZVYszldROnwf8K+/U5okBKEbFP
N+txcGor1C6aSek+KafqUAtgThqwufg7vG0492qrtsgDhTZY1XEnEMRlZUhZ7v7KYT8bMxA9sSyN
6xHZfdvj5kYqyM18K1+WY/yILEWUoENW3yN1pSNUJmgahfUxk84AhTv0F0ow/3CSEAvK7V99+ORO
V7Uwwq+3gvfS8lMGex2oB1cgZ/htPoFMBhk8yROV8NUUFxRiLxQf2BvVYhLrIWrolAkv//QOXS+g
Sc3DCSx5pOKRFP/NpLkFkQhH9HTGbiiEoQ8b/dMHHJJ6LHLUIdUzovaVi7WSxDj2f4YWfa2IBBgb
wHXtkLkJ0G79mj5Sy1S4prIcrpoOotYwmRMKdEpGVt9twQXoMuLKvBoeSEKdgS8bSV3a+m+KoipR
2oQU2DZtpLngwRX+nKT9NoFgRrIYrApTfubOMEb67im3rlk1qwzLqIGQdGg840Ug92qf+tPGBM4t
PgBGyJBaavZVryzzQcbNQvfEk240jFnOsmTncfNQLewE6yU8vfe4LvQf7hi/qoUTOGsPpAmy9aTJ
Jz/vElN+Eu/Ka2DjKhOR03jJrQUaplXJg/GQCisuv43vQ74+9KQco1ghaW5MYPv9ooj8jomaPR8h
jCG6TXCcIFMYN7dCxYrw7DJmu4VSMmyJUhspffsdqyGCl2GO0DUWiHRcPBE0pN6eMQqotvWd05j/
jANHjKylJXg/PTC4eczEbBnN6P2UgtRG3QxrczsyCr458eX/V3Bg1oPT70hlNEVhyPXbqe5tU9kL
oiyj5/yUug2zLgT6c91cbVUQwQ+wiQvqwuxYrayffcwgI/+vxKcoOopEHLNWrkohuSvdXJghAD1i
6BotKXcRLYIEOrJN4f/YHtvJeRfUiW4XkT9XP79w67Syvkh07SwnBIwdC3MmDsguWBgSzqkLeXrj
uNoC9Lb2dGArPY9k1mtK/yVlJKd/prBqKJsR6IrcdGffAI7Zw6xG6Vkcep0c+xCBQAJ4tbZ3AhT9
mPi+6gQ0oHBY4WrnCYAQOztiU3919VNJ4uldICcf37RNlGgrczT2t0gKwtD9Tv2FJTQX+/cyeVFT
yvz4ablIIeouwgjyauASrH4v2YllqbLYfieniDLBqVvXbZMlcu8b6Qrj+r/G5O+dJDDmcVHwolLP
vVe+nHISieXtrqbHhe2hl6JWa1cpWNvF1DEj1cQH6DIWs/1KJRXc8U83nF0tg6KjoCqarIRi0IUe
DBiYmefYaUP5e04/Jox41df4v1KM7jnrfp5z46P7sHKawzN8lFn6p4zDQzJNOM46QYoDtxWtZnVd
thd/WPPxqWC0Ij0q+W+I/yg++Fc8B6dCVOVixCEXDI/6vtwcC31NWBPjGx6OHR0XkQePENY3p9Ag
psrwL/KOFfvM6YNLB2ZITtLsmIAUYO6eUZzJ9gYewuTQa6B1qAPhSUrlKlJDDsxp0IltiG5dCkeW
4nGERHjVtaoghMGzzBuzq74Zua+S75Q9Jdxlt8DxQiZp3cR1NDq0FHE+8xG95jT6dluO0fT5QWeN
78/jPETllvm4yPBHo4QrYYtVqUpwzJ1LlX8ziL1QKSJVVswMnkFJ9vFXvZIS+DQfG7ch56pKJB7v
HRMsNOf1xzgipoE1fzjT2hmPaOOUu56arGlkfAqmNlr7lLJqhkwAF2uAz0hTKaXVnrQaNfpMM71l
TOXPl4XQQxn2QVhb09sVvCSOk746BwoI1Kf3wAGU/01vfxyLdzJpCAI0jWo/CnzwRY5k8UM3urzW
0KBPy2zwauHXN8TJrAfjFe5Y7Z8me6Ca5r//eccrnVMynxZXdkHpwCiDX23CGMhIW2tYEia9BoRt
zuY0EaJTAPVtJt7BbRzT50GNzYjI/bepdukd4xW2AL92nBpH1l7memei+pCAzO6w5fbLmQORK8y1
h2hVRzXMG413ljZYTPCqOzXJ6MATco6OqhWg3F55OBHiYC9T/embF8CUIim8yOub3QjvpavkPWWs
r+WvYgHJYCCW93CU4FFCnnUoSJGPC5aHY8ti40gK5w4EOXzBBS2LsS/33/M/Qlgxnqdij+//BYog
TKghIc9dVaDadwnl/vqZ5jfDQv+Bg6j3G2etRZJ6+H4uVkyCWQTkWT5/6RaZV7W2WaU+24OQRLhi
8bdtgbjcLqpnbJ9jaGgraegHDOHAmAP4Tmxm4HRX7mrB4k71kwZccXCzTYvheweSXWichGL0urQo
Q2ihmKYKSBlYW1WabZ4eYQZCe0j9XWs1IlPQEJZxCvUFQcrTTcvY7uMxoXdGNiIFCgSofkXCIo2h
sgZ71ap5fSSVKXJcyLsS6C1PpSmp43Ubexxvg+VLDs+pWSEtCXTI7Um5ir748q/fanhCpFePokrK
BKquYeFF6MByf0NWzh7lYQ3AjjJ44wv33jO8fFirOkQFMf14PLAjCalSB/kNbWyt4w4ewKz5xchM
K13hAJYw8TLV7PUNMzeyk97/Hw44Dlw9zSmchqDUwkH4TXc0HQkZg8xUigGmzT7WkTAB5UT7GNm8
N1OO5CUUYPsecAy62QkeiYGlMm7m8oXXC0wr9QmoAjsr5D1JF0kSQtZf0oeZLHgVRyFxhTcrIAMa
z0u4E7FTCGLIl23H0OK68UqJwRmsI/lZa1kq5ft4PsY7yhK0tfoc9JQ7g/h+PXzNz1wi6RNENwAh
STgOeioOORJEHG9ZUiA3NiWw1yyUH94bX151QcPLH744pGkZQc/EE5QwFyew3vvqX8y7HGrIZEop
21RvHmY0fNaKtpUnxtG48tqhgkceF78KXuNPf55/vaqC/vuH1vHcWt0hiA2r/SLFmUm4PvG10akj
Nk57LyvDW0UJ6dDSe6gmlukAlmRcUIRreoTpPAK0skgGDGacvQKIXxz/1cEtjpm3duoaNhwKeU/8
fhvExWZILXdq5ePCWlz/l4y7LAGW+e7P6cPkVgzwlG5QEvdS8CzPQCnt0xlmcEYImnldwrIeP5aV
As306g48k0FJwYeOAuBLZrn4Ea0gs7e62ylDjQSrfi/A5DJH4OoaHpAhkCSlweFdvYNLtCxXg6B0
fdTQdaV+qJbpTapvqq8ZuSVEGDIqJOk+SmOr6F5TcEdS+oc/DBX5Lj5Ayq068wa7DrLDhL7hwCZ9
2U3JV5vWSko606sXnNIYoedKuP96gDLL6bfBii92ODXerjNo8FLNUAOWtprzRJI+g4M+vFRtMxFL
kTv0wKi7NVTI6dy1QPE+OutdsqoIizeYMEIA0NZvDp1j6H6HuS/PubPcXRt/IJJLlZELFdvovkvs
wQ7aTPy100FrdD+LurIbegEBZFh9za0KsUIs35YfnllWIf+vPszGegorOeQR8HteEboz1BvTZ+Zn
NUbZJ1hLkiRKdJcyduG4bHETWtKDrpfeGZ6p/vpleP4bLHxuUrc4BtIPtYKjNcbMZA/0tmNxU/l+
B2RgHKGsKZ7sa6tj/kfuwDPvYTBfA9AcADhgdmnWPmohL/RtwJyHHrLzGheIAfQNMaGoMQmVjQ+F
+u+MMeXJZIlJlKb1EGt9hZ8Mj84nTN760rUHyDmYQdMgYSTXmYqp0QCl5ewOkMkc53o1TYNBvlAm
zfVyPOL47ptDiwUjPvNxqRvq8eXpn/raYITOS0dBnxwtgZaV2h7XWB3X11VBRhQ/fcivGsBCAqIT
e+TX94iQVvTwFNUczm374Cmbwl1d1MrWs0PsIQMxKXG226YjqoQGda+s9C/sodGtg8M64FNz6kWx
UtYIA1t7XlQCfGRjMBoMu+dO4gkWXr70ARAOutH+gqnJBLKZK3T1kJ5l0ViKs+wcfjPjKXIt6Qay
tQF5OYq2AEB4tyjYROE/wUkMTABHzBru8gahN6VmkPnYnnKq4Qa0ICYC2DvI9oxtf/txciwtt7LV
/s1hzZ3Ec8rVhSeE38icuSx7RDfwVmK3lakKb4cCPJO0kdQybOeNLECEkdDqfFCL+yMlUGWdLXkl
vWAUkUVsjy5tyiLxlK6bohD6Mm9LnHYVSY7Ml5s0chYqrQnGDH+sWLHa2m5MBtDvp6YaHtYRKlJZ
vDbl6sGdKRtFCsmoYqfHCmYg+aZO4vj+jknTdXaUQYc4rLer4Brm1tMCYEw2sT76ZGmHQQyhRUGe
TeuvPPJal93riIdwlwlx8uPGL03FAxPQEmht65wKdac30Neur6wg1h3ZxDWq8PCc1LpyYeaG+RsL
NbIsw5LDB11Hv1V/PoXzOl9nPwNYoqaPLUiv1eqr+2xJszkbVDwPQDJ2MrKgTEuS91iO23yQ34hz
aMoQMQlFhMyIpKpJzOhCWa4Q1Pp9TIqTwsjtYE/5pSEFLzR3LED5qkBbvw8Z66WvzaxDVXwiZMNY
lBBmYkUMaRvYdjZORTx1yi85xSpGANtPlHLZD3kcwQNg7Zm0hKo7KiprRAjymCX1GqhKB04OunvY
0Lv+/6CDN8VmEUo8tGegNfTerlfoShZNR0b32RSfY1xOpEJRcvijf/k/LuXGD1ngE8if94CyVLnN
UB0bms/8kkWai8z46GxS5b55mH6sDSr6oQTDyzXGkN2bRfEVzYXnUyYvSOVjq7y+9dWn45eWhNZA
BB741/oPng48rLe+6WrlJSvpvjS/ZQrZyNU4xDxgOHv0HLmQ97qvKBP3TkEGqByKzE6WomkRH8nQ
QMZU+iH7zwDXhqTxWfgyryR0ydxbNB2XiI27Aq4LkvHYp7tUiFPBxBVet/yoXvfT5Oe12qG8DLRn
IEDH+q+VbgzcICjgv9nRrM0WrJNqfyum67t4lbVmjQulZhlvfwI4XsaAUGSpwL3iK8Tp51tawPn6
udN1+dPIuDvoGRVkK5xsdkMaogsShmkFGKL9wYwo+zANQ0wxbkMnQkyY5MDOYmDnAUyVYNo5PZNo
+wCHha1WlXmO02s16qgVBm9mwC3C83Ac6Fw2aMF06eL5H30g6BgJHuNQJhrAMtCrbx3yq+UyN/1C
PBLdFH9XCUe3vL/msCWStUczuv6Q0t6qHCSvvFuDM8HmiUDCUGVL9FCzOqXBEqja3hdDlrpykDyh
qQHjoueUNFH4F7B+Q7zq8xEMDUNxFF0aegXSGHuCbntXoVIzqupwznlwWe6GEauLLfvQdNPcrhkR
NCBpqADztLwFGFTX77T51pjgKjqhzbdAdX0Cg+yjg+FBt5MjycchuIy1n00WwS2Wa2+ZLcs+Kamb
SenA9ejlYkyBb9iHalk1auWkhZUdDlDW/bDlbtXYMksYjr6LpRPI4JfeFr/lV+jtJuac4ZQCAKt6
/q8kwwvcodGKO/8y5JAzXvw8Y7JDDZ40bJEIEJpw6OmvY4TVmkIua+juecZL6pd4ztdVMGOVw+H0
35ljtG+rsV6GIUu1eWSWJfshVdq933YzBovAp/7sf2GcVVkp4SeYRZy99sIa1UrVI35OcgNPus+o
Jefrip0sKQQQ0ix3BLvLGvfbitz1xZVX+h3VyRKSA5ANjrP6N7KpRYAwzK1ozHrdfnR0mKbNSEsK
0nqMfy2pCbgl46BRDUkIsijxQroLbYaDjecLUZK6je/33URHdve2qxTmp7pxqVzPgNOqFrNs/9OP
7v+w7RBgsL2N75vVtPlY8q9QhEXOJ2rQuCtPPcAO6Q8pvuX+czJ1pXv+RUOw6SrKnwK8BRbCim1Y
8svLm+gfPFZqpmdxaxdYhbGBG3sGRcQDmAfaYALrGwubOJnBg/kjLwvSqCEeBe46fSH30HOOTyT+
UXjkSj8qO5sFv6Fa5/1fXP8Zg4b/hqAsebYTYUwq2kCxtg9i9YkIdEN3LwNh7cEVctue9aKLeyXQ
XUgjUC7MAkAydVrigFUqJpvZMAis7uRiwgA6CVHLhqdDzNlV4z6q6J/mplNLjoS0uTB/DnFEis92
G719kTx29pwjaZroQvBy1V1/gKA6i+b4/nix1wDDpcjn+yWXyP4Nb9sBi3XD4HW3ndVM0qR49PJQ
j6XF5NEGURsYBTBNUc/wZ/+Rwl7z+pte3UPE1bmCZ0UhBMgGNqwT3mxxlOKK83RJQ9aI24jhU2vN
/dIVi+DTCTi+4NJH2cvrmUYuzsh8p2JDXJyQ4FUvRFsk704Krp8uBy8cq38R/v7r4PZ0ypT/03m4
nR/laKIqtbqVgNBRyTNpmDH3j/MZUvLR9JyyZLp/CJsnIEszMLugehV7Yd/h9sd0i8cOqdP8/sJE
7DaH5gA9p6hP0Hf+9jHyDgr7K3C5ntzIRZ2o/3DJjSjw0T182rVxgFEqt+yUDg1tMZiwBeju87Be
8eFqPTsoRJj0f45jCtHkCzbcBxG5T+KnfuI5rnB8wyaNaViFcIUftKbqxI44PlJMMJkN9S/+PQUB
kaIlvjalQMFMHUd60m/aLSa8QC9n4DvvQHoN2per201J+HF098dyFr4+fDWcI9E8uPF/c4rwKRgp
lvLhDu6fOogBipxA6w/lgeve5liYAFbREsE/KVXNQrYMqbEwp1HPqTLktbZbrn5jEQNbNngVivu9
IyAHNPN/rPWQ7X86Mow9QvDqjqgetNn+fQfUk4zOIquX9pvYLcOE58UPQSwxzWRWT3jRb4b76lJw
g/2qjUJfzwxvqJ8pVUVFqSzpweEPZ9ePgetJcdkhI5HG6zf6OMysodE1OgyD0FHL4ofq9qTlDRU2
9H+wrnxp3U1RNQ8xVFBqQY4OIQMERcGjcF9V0M0CjRtfTcWetYWsyWpyesxlQ5saub2Psmornhgo
EB5a2REVDrVCn+/FsAAtxyzv3SFfhCCakabVPjH6Wex1hzHJw+bQFEOQeRjmJVvDHNxnYeWNhxwM
WjgUQQApIJ2puzLjI+N4x0I3R5MHVTdAGUPXKAz0ZkFZBZMVrPUgfyxBG2mrhM43H+OfDZTpimK+
CJjm3G5X+oKaugwoy5wbi0q/uqTI/AJPSJeUFGzZ+AeNO98AqyiJz+ibuAS4+Ip49jPRlrZgq8Ns
M40KDcBdn1Xn7er1Y+7jk09i32CJcTjEakjDqp3VJKiv9FUcwhwR9rGLDW6z51AZkhDKSBsEV0yR
2l0jvo3wMiv6F73rneOkPZdJedNvxKQCd9VgCePfN28GFZBtqevRbREMPAAar3sf9QDgycIKf8nH
BaBMHskNcpGnsGkv3RubGcIxIEx6pRKdD1jjDfTY/1QuVCg5BM2vd1+l6BgfarGHGr0iZ3KISFzT
lpBHN5KHPxAVA9ygiUb2UdjBcDQkV0RargRlwzAWCPsaWOmIzpNzsybxCUblTk7MWzqMc12zRsVU
jxRp1r5V46ygVxYr6udIti0dJGbm4vqblA2T7VmmrhU5aBFKa5yB4WM9IMRYZ0u8MTJJ8aXW5DAe
ELDZFQy628xnBt87gJGLgrBxtrrcMFAYEoHn589Q97mipg76Dt3POPLbjaQZF39BJig/SHGajTDK
ASnmwBLHFDKISOYjcXKf4tbkQ30DVhElP/RLvkD7eBeZSZ4u2XzCIQkijnJf6MXh6kd7C0uTw8xC
ZRYhsQWZIQ2k0LnTu/h98czG2kngXWEpHKAGAlgeMFuoLsxRC8p+7oKipxwrLy/o+cXh/GZd0Bnh
6JktDfh2jnPV2uPPYmjOXEDJ5Qhi99ryk4EKW9ntmgBzZPQO5hIDyo8z9gAWMx6ELhJ1RPF4q9gK
r3JQPkBMLwhZDRr0ewhH5y55Eh9PrMiQqbwx9Ni63HmUVgLblV2kgiMyI+OKK44RSGM80emS02GI
OTNBFEuAFVYAeB6zwwY6Zm8HRU1cKbYqxrIaeObo2L56V4Y7cMrVXQFSg2CF4ab/Ef41ivuZCKZX
2WKwHNqKRPouUSU4Qr0VVQ+rEQTwmju38YdgSn2ajV/RK98JVRUHHukYje7LLCHrJ2EOn0ciYty7
zHBnCI5t7XX+Hj75yPKkQhX3RGlSXdlkGiSb4+VVR5Jr8EOvs3FjK3hxt36jlKzuaQhEM0m9Fmwl
mGhk4sl7hVjk/Vctsj+nL6i01YqdFALadFy0PNO2uqaCjpanKfrime0ODlLsHeLOFaYq94zCZAiM
EiYu1vfqua+g69YCZe3PeeGPxiTP2y9XjfmqdnOWMNEgmh2W8ItVqoohFKHiRw93YIKk8rHuxTjI
rRnwgVlPTdKqkwGqll7eCZ97OO93UH8K8b2zAo5FvBF60/CrfehPEL/kgSCCRDocFdQjIwp0s3un
HRe7NCIKVRdfnsSIxZ9UVUkbK8fmHnglBXoKGCVZ4WVWVDoyFdht6BU8Ui0nZCBbPDqDjYKAc+Fb
jxpEM5VxWs6Y/WxCCMApvqPSTKBmWb98N/t35zBkdZ4oin252DRF08JM0lVk6cs6l7vfzTGGb4+l
cXyPIXnYuIwFag8ETvrk2DOYwDTg/6vpXHIqpqz+pXIHTdhtkJwwzZYixjotGy+ShKtfzJsyYuQx
JIqpsyxzIJkiODwBr3JlupArgLmT0vQBBuWR06sK1kVoX/Hq4Gqx1RYFq2GbHUMnXnTpempRmErR
oPUZV3qnd/Zjr5Qjx7MNsS/axU0KPFGE3dfDmwE3XWt5KcWNWGm3xYD2mrZiclYiQ0EMSwJeL2Vs
h5sIv3avxyc3z7G7KVeRQAZxTpnodiH6bGLAq5c1D38YsrtkzFJxIxLpkRyjh3FVuGSjxCqJGwwk
axFmsVwQ0+oCQaz0dSF/BEjNo9SjEJW9TpXAtM/2HHtNFMLt2oSY1UQqORPqiFyWQ9aa8OAP4Il1
5DqyJwXEq2vDP31XEUHE2cELvKwyMErtseU7LASr6LsZBJBspVau9veh/D/glvdeJlUW7NZEn5oT
lTmPChx2EYoZwAXOFI/Utkij6fI1oxdqSdvwEgkunxETp26jJuV8ntDQoGhE/SZztb9fj9j5M/Oy
CfYeCFjV8mH+/Qc2ZRzx4OLq+0/X5otjHCIIPowitKjBgFeIbjFGNb7+qzLB7wXHLzX5u9CVV0DR
0h/T2TPg0ft7mkLOojDngA6R+pcAjgDN0AUgJ0ZMwaSp4k9AxQMqp0k5q8456qZYiQPybNpdqrFY
6etQw96e/gc9ZIQMErg34uX75SEXGv9jFsvsXfYMHML58e8Ps5wb8lOW7DdAxhWFeEf8C2G9JZkU
GDEKyFow7xSQaAcPlWxk11X/10fBo91FeWO42odY/zB2ndwCjamzAD0C9Kyi5F5/AV2f+wofJMXz
S3Yj8XSpOcJ5c7iHDx/uZieMzzO+Jzg1C3rqa6a9cDxHSQ+Z0aRSOseBhMvpqHe6CrT1m2GHYwfZ
bzltPUlvIHqrs/b3GFNDdmaQgkS/7gCxJz6Vle4KEx+BOvCTMZe1JFoT2jDyqjULTv50xIotLqwy
CaJi2m3v584z6SVJh2MuG8pIqYB+dxtnWWRNsxYRduX3MgOdGFG2GGXW9/8OsIUVMb3bJJ/+TC+L
L1RmETDW+NnXoH80n/bNz/P1dKYlZ1NZB6s9RkIAOzep5pre2z8tB0A/fv67suCo0U60clXMk1/l
/qxnAMMK5yJfMLkfG8UstJLxnyY+WgRpFGViH+peJCwAKT2Myklg49adDRkT6PW5kGb+OwcZFX5M
rNxs551REsn/z8YaxWJQiZRth72x/imDx+XoXboCrR14ZzXr/QpEFFFcCE51cKzNYUbtq/STcgxF
TKBLYTSoZs7J1ehT46pzWa1hdtnaTfFnnaR4OCxGvM73K/LTfdIs5xpdQcJwC0QF3+ARb0mjDERu
IuYrhDq6/FrxR0GobWbSlUSDjjpImtLXNCySGEwNehG9NcCRkeXWUf4XldK2/5wb8Mn2P5RITQnw
eh/xwGKErCcA6GNLY2q7fxIdfpkXCySuFD5tvUaZpekqQp0ffsl2znpFqEJ0WYjf2hwUdIe3M4DY
MH0oWgdsEK71b1bt+cxMGl6FUEug4r1wSI0qsY2xiIBUYa31WemCBDD/hxFNZrryf2i93e0xu3Ts
jNpWcv6FNx6z95Re9Hf69jizh4gSxUzZSZaZJ5pLipur0A/EadnztZLfi6k2s9BbVcTa/WZFhh8H
VMkCo/rIxBJeIPVYngcgyyeZ7ydJL0ZPp8EZ2a9Qp24L19YeGaq1hHRfEQaD1SFraq0uo7g3l0uF
TqbTXxIGr2MfJ2Sw+I8NEaI8S5RRZQxQhExqzw2PWWom7gL9g+nbzG7lZ159UgxIq1FsBzhF3To1
9e9I91MIyVh2EQEUobQ22yetHmU+j3o+dM6qG/Cs9Ztoe4rajKlDxTJlQ3b1oP0hljau+1/C4pYq
Xu24YIpMP8EkMwj91WHXjRaER/w/FgshTWzy3na/xxgLPRovhplamDvhAYb7HN8l/EldAWRdA8tH
O2SnPzoiDeA9R4+cIfufuj3MkceK9HMS0+OJuVbEYDgma0ic238muVMfcmzZ0Vcww32RlGT1qlh2
5m/9zh6fsKyyd7owke4GN30dCdjhT2SDIyAWN/QQ5ezL4Om6Mhhv2Xz1Nf8/Vro6VUB4/ee2Qx+h
iY7vj0xJ0m9m/pdvbnz9AyN0MNDDW02b851stGFq8T0JI7Tsna0rAhRvTnDq7aE++KJZYbcvRTWY
98ZDAHFRth/PRLG6YOSckxV70DO4uhvy7HSerGhROh//+FU80MQKcOBVQ1fCsGoMu7QX5GVXokzP
R1SMFt1h6xJbDGPTKenk1BCEyy6BugB3ixqWQAHilk4sn4s2e35NQg+llT9lont0wi1923gQYWd7
xYxFyV2RA5iR0XO201RK5w16hB7sv+4XRtH3/MVlYLdfBXEpZCZvz1A1oit984/EccZE4PCYrNOH
201Yobms4Q908AmbDbzJlIw0kR/VCYUWPkkLaP+U1gdL6rpDPxP8mw11GRlI+uOYxd3jIS7VQwGz
BSpmSAM8VxxqbsUuQ/8KhEdDUkGtMt5I5jXBuRWMJyyjFb9DIfgzIodnUSgSghsOP5bzVdeylcBl
dRJwN7Vo8U571e2Kp4Dts106qd8h1Z1eaeHG4IBQKjFpthk5i2+KY4IwmRBcm/fiGJ7jV5Yp0aiS
la1nLD87aR9holS3xCQpYCjdEEVehcWctuc0U8/nsxSTORv+yNCexaPCHnzvsotSSGlrlSWCD6SP
CmxDejOXDpiar/xuEvm4ADvX1UtFLWHL5nqHoPXbEVNDYNa4HykrXkb1iDZTQiKSvqA/csbCgPrA
M6swMADdFN5KjmdJzCk6vr6Waj5heP0dU/nxRXFmkDwwCzBM5wog9b9+cArCpc+P1nK/dxp6dcZv
RSOFYoiryuTP+hWBeDgxa/cGkWdAf5b7bLIX3Msb7hTEhm/LyeSExT8zHkFaU6sK3US2KwT4PIYy
D/Y3RYVGjkUGOBWrC3/1zMFrNlSn2vAgkjKnH04shNW4Y8E1Oh5KDFy/LOeczTJ+GqfrtGC4goMy
L4v8hgSOjM1jiwUVRfPPxUYx5CsGJZXqffbPJEcf0OlA3PiZFJaip+Qt8pZlC+JzcVJcGTBFLkPi
al4duXScbHDISQXaQX3EZoDLEREFcfqbTqxStWjgGtVv18g3PPwf6LyuHFlMERU6no2uNLUZgquI
qsxRUbEydP7P9O0Gw8hXgPI/h/LBsF3JEno1rapEmj4Y5yZPXktoIFNpH/tUKrLZ7UJ34xEpEY2B
Ul062wgo+elKycUj6jbsuRZGOvZBPKc+GocYLHxOjoG+ebiN+q3QAbqAP7NGYZklIfKoFvQF1q7q
IWZzK4EjMwhJe09UL8urN+7oIpil7JCQ+xYvDh0WzFIl3R92EjCSWSu95YpvzzNn0L7LFlCZvg6N
5Az3mjBRFBc1yDKohei+VILO+iC/Keblh7DRahXc6X6BewEOJ/b48Y4I2AN4PmHgDS9VtmuOYB6V
h1AVPZHjzNWM8Ff/Svl/RKIr0MvzfyNEj6QhGVftdilxJgUb0xFkePA1ThVsHwpNhVWNCBi9WV0h
izUizz4CYfWjqYBeydkw2n5jLeh16pw4Go+azz3/uqFBTOiDKqq4XX6QBE2D/1JJUENgmwU7675M
ScpecNyCr06i7q2tvjPHeM3wXvyFFk+CT8QnwP+SNBHSYXXUO2GhvIoKq8QOaOwRLDVUpzsaJH5x
HC46advGi8aYs2Nbp4XnXMyNBxbVq0+2lqV5PHnrbTR9EAxtrg4C5a0NXyqLWAZ8HHUQ4i8s3zYg
14tW9gfe/U2QdVnV0CH39BNins3UZxBrkb6Mbyisj+r73b6IghXlnv5nft4xTZNchtkF2HBfsdqN
rJppH07BCx13UIglRiaTkeV/NASNQvlN57IBpMtA4R6Hk/6lfjvYdZrLBZF4klj3ZCPwI/QR+2PY
AfgM9DRzC2k2fenp24It+NhCx436/MQCUbnAMtJinSdurp0hhxnNcmjxnmrvIPsDL8BFjv0Ghjte
d/8e8C9D5WfTKDJOSqOrEBn9kWKkjMKojVE+7n2KjG8uvS38QCJ3+a7LP453ohe7xIqATR+mPqDm
NnYhFNhI84J7PPIunMktCOYHImnwAqjXnhB92n+AWWOP4g8cyUfvVhXUe0w3nh3hgvsoWhgGpmVE
kvly/PxY1r6fh5yvnHe23sfUTXhcxSAqZH3ELEfwdVWMy0UAtYwLzYkyt6qNFZEMXhErsRetAonF
xjhlc2RlSBMtJiXLQ/VYZpMoQdU7lKxqe9hfXhGFmXewBSQgVHhI+kykEemrsz0fN2YNReLiaIBg
n4WVUohpAtaa0bwafWMeLYYprQVVz7upfHUo8gayniWT2vzUp2BlfeY7O+fGAASEEcJV8o/21PPl
RU0z735N7TwWRCLSx0KXMdb+2hIvaClkiK1qeXhNkmVshVWdDxib8SsTfmFrmzx+gPSr+WqF08+K
Kb6f/6laTtTWx5tDZb6xYZ8Od5YFx+04dMFEu/+WF6DkgXvitBSkQeVCn9t5k0xUXmb4kuPtD2cf
enf4y2N5+pIkM3dYifV4J3SwNKX4f4Co+erF2l+q+jQHmBBbHqgbmomjyeGiFCxmkDgfBTUZpl+m
cryMg0d4bEp7j/MM+hTTJwrc5oYVzatG96DRywgdd6i4v1uuqOsQUo/CBgEecnD9oL17K8np/IKu
iWYgLKYqbhXsk7a9I07xzv00BSxMV9b45H/MTluiq/8ZMq/2GLrd4o0Rj9IZqqfsnpLBIDJUz4WJ
XlhaAe32ssqlHnbVRHgy7Zy61V9hsidfmhUFBJTY74V2Qxn/cCz0Ap1MEc9+NaTE2q2O2GDd7lr4
ygpdOoR5C3JqXkn50CsKLx6yIAtIiu4K/7cH9agUW57E0tbggzHpCtOteRnpGvrGjXyt4PKfbdbA
pl8bnEdiiKywD+PIn+SQpLqKAotLueVinyoDlksVzYRirhSp+hmOt8vK9sK3IEPYdlGO733kX1mV
DWUEn0c8N1rpXjZ9CzKlLX9140qsj4LSC8pocCX3qU9GgK4aigrfbOYc/1lnk+Leno4UYH5lgyFz
0m4H4F6IZcYawNiP5dZbjJkeUtL9fR9tYW3ZgLuRV1+GE/uvjc363f6iAd/XJJgWPeDWl1ec6ZZZ
sKZTcNdhxruhYlGs51fdI8N5Fq391dMkswvy9HTOrHC0i9kf8SHDvtOYfzX/Tdk0CBEwCgu9/4C/
ICZU8ittHjUUH0ScNinNkfy1yDQM+Qoyh8VcMFqWFlgnypeiX1keAVM/TpgBT+YeAG5LX3kihHSD
7rW74Z0CwlWZ6fH1fUd3Ltifa031MNhXfaRWuN8ypxJ+DOWQErGyECkzHTn+To/MQyUpGKbgyL4D
3ANfwO/gXzAXkyPXl+dA+vLOYqi+Nrig5JKdZ4vp+2knTPyeFoGYRS7u26x/2PoMKAnLP4HCyNMY
ip1TAj3zyZrErOte4WUW7HgjU2lFBA+ANslklxW19U21HpTjXdAsPJwBp9OaV2OTw1neNy/0mcqU
5mcn2dGt1NdSIdOonMLBJuJk+FdYZqmb18wGmXrYTgYxom7NhygSP5mWbN7cVuZYRh3dwKU0Cf/5
4baaL12+K9rodwzi8pwOl6F41bEUNeRCp/gj+NZoy0dw3/CBSyWiQ2m4cAcOSTAIL+C/5GV6/cEB
2GkKf5O+YzS3+hN1+iTyEK1QjY6xqBdjOyfyb4ixvDm9+z8HlBBfqFA/6lUsfQnd3TLuNTErQdEQ
PW/aNRMtHIk/jKBwiCe9HYnRFAlLtES2mLIgBRAyVHCMyerEQK4G5elbqluvGVZqoNKlkmEB2mwv
waYkSVlVD6MzxiWfrFfS8fdTISao0EeXAC6y1JZQvoGnYbRVK90qpiCjbInHvSuqw3qsliRjoJf9
49FXbd8XsTyS1x3+zpvGJR3K5y3yhgTJ4193d1annsbBkOzR/RXo0uD/0L/pKqUCVt8tAxigUptg
YvonnmcTLg2f295OwFaQ6JrMTpynFuN5Lke1HBov6b35dRoU733jZqlhBqkCPQr0AP3/FOyj65e5
77R7Xp2BZywhBID8n2tvxEmgt6TjsqlWUvChQ2+uowccOlZZNxPMaUHBJzyTSF2rlXOPMm/f+EiD
QyaULCf1+j6wjW+YiWakHJuZD/Q9ifkhXZ45QLswNVHcHIbpoTSdxf6KYUYH7AC0olY0CxvY52Zd
u0QkqWE9Fgc8yZLQD2oO+igRS5tq6NBeREd64zU8EffiFE8mnF0IqC7M4dwELFmoLXH6qS080odj
jTjB3DVDLkm+p/kX7czwEbj4vWbPTHWsZg4V6T96wNwvtSOvZqYcS/3OKaErwg+SvLVitQEJm2HS
FiSkrcmwBuxdJU4yO/HaQb/Mjtpd1djElJ2QBXpaKxSt3YLg4p1BLHWhOANt7MEdUQg8cNgvKftS
eeCDOYAuTL9lYuQuquEXp5TWCXCMuZ3VBeCu90E4FJZjoVhyS1MWNSOVng29W2Klo16/VPjiSpu7
07NFN5Hy5LBWGF3FmusSI/2kn+cbwAUHHib1a9r8ATVZHaFf1ZhNtAYvBwbBCscHdU3h5+4P0kHP
vMX0o8XbsJwbUmOrQDWjQ0aikjQGjaXa87HGRFplBkpIxJFbb2I22r2oULtlSiPDYSxjLgXhQMMX
gZMbT1lf0QXWoeoCT96wS49MlODk67JH1ss2LCboC2Mi3pRKme/t8bfiVvCym9EAAK75c0Hq6nui
5pFjjRcMDEO/TezEKqqAf87kqipnwsUcCNJUNNzQ4+409ByeLpZJmzhtLx9eNNMAbJwbukk3kLY5
a2SnHWBF43HUhsavVVbCc5F4UnLukXtEmOwJI3C9PLKn2VQQn5bbyNhARdKrER7hm3Dsb49aA5/K
T20MuZY4dR44CsmE9BnBdMuQlueCZJUdrlv6wWXpHUkHXLkfRt62AQr0wUxoPIgdr7qhXCrDVU2K
LpHAXgwhI+l9tNwKGhi+mjhBEeyPw5xgRrOeaHEnKrBKCY5LT0waRbHSyO3snQTo9AUnOdIj9eM6
/f/drJEKIMH2mN88gt+FXLcVpUbCFV3xw+rx9WAJcMEYAY990TO8HHIBaMxlkWX9fa7A7Loj6gqa
CFDfdGIgFQmzYW0HV+G6A41rJIpEpNAhGK9bRbRtqejM668rapNkleTtHvNklAa+J3LyT9Cdu/vU
4IjdnOuOd42n/bSiw9e7SKR4NAq4dGS83JvwY06cttifUF3w0uAn7ETfU2Girkpw/r6GLtA6gMZz
BlyvpeFf4A+WqZKSaWrh3g/aXEQSabprukvIDxIyPdf0DyvfbVACIbS29JrFL9qEPCuQkEF/gN7k
8gZbsi2XkJ5dAjD2BHeW+IK/Md9hN7COv/4kE3WL7SrEHFBXL71uA37uTBqVYoUYLUfL7XB9f56I
HKUE1knI4FLbMEkysz7t899/T/uKIeeMlSVc+cxGapmfxWJVAiqLCFwDctBs+/pZal4nZSF2M3os
cnnuxFIvXJfTThgxhUcHolaRZASyTBEhAj9jtA5DXZWAfOppN3Ky/lKZXu7FkqWdqPSWcFxNKSbl
THDdfkyYwxntkjQg8EIbxImnDvXlYzrSHM0CJp9oTuqQ7bc61kdLi6uA46YmkAfbikNKXB1SXoXE
oGcQsOWeugNhR3brOYixoGbX8U2af0l6PTW+DrL7yjOXrtksKPmWa5kIsEBMkSfLMzHq2hx73mzw
Uu/kGKBc/mcRZNFvxfWEYeD3e1Jlm3fOa6MO2sWbN4enWnE8yeHgXrVYSLlWkGFq8VAIgIyQCdQs
zop6a7VAXkAWzKD86hBs/rcNXfhGOmqUVKe0C/WMtpO4dUzY8LOBLoBL5ho+asbKKjG3nFw/9Fir
/MRyiHVvpwpbtnVIH89VGoDpNMho1Akgm1BYXAMvIUul+JKoND3CSw3/MqdBlHEFSpPfqMz0SgFM
o3lUncOzt4YLV/fAUWVpUYPSYfSsBI6rDd1aIJaPxIbn467GwXmE4DBFuKKnZXXGlO7K8o93hnq3
4bf4u+HjoKN2EqiCaQBlBbf6Z89Q37UfojIjdQN8uJ6YOwoHunHpTutF4NKJ+RjBpwAw7/XDmTVP
5OJUMdxWMUsxibAhqRRy/Y7lNexyewnWUzAUxRGlEIYQ5T5Iv3UHG951HS9HpTjJgNm8RUzZ1LUz
pss+hHpLNsTJ+6OqKoaa3iWyVhSS8EGva8Vy5O4/Cx82NdRuxvnHfhsywer7EAGBaKHNUaLWJIkj
YlM1fWFgqSIKw7Lbs5ugcv9YFhwAmaFg1gmChalhwtGIjaltFC2RI10kUwExd5jOEGplOl1UvJmh
D5AXAx5qJxui9LIg7g0tJDEbVg2n2WbQNBjZH/ePGHOKjDWF+sU6LiNgd9obNjxogjAo3vwfiPsS
nEwjyw2fsv5QVV2dXiVqWxqX8Ts5E/uB+UhxogYyMmp62vF+yi4t4H4qLdj0JxV7fYrg+aJVPLZE
gx0W7G0kAZbDBn30UIcMw4pCYk1PcSHUkH9rE7UOk73GbXLtHGsY4i+nemL6ytCB/tMuQCB34P/q
3Y4Rvig9sTGeB8kOKn7RrCL2MW+j+TGdU+Z0G7JHYtw3TnUXYUpiBo9cH091Z8gmhjR/iFjJFpx+
baJXr/XSpI7i5c8c5uKa0HMrgns1/xIbGOFAr8argZh9afk8ByUS2Kjti5O/uk581TCl6vcOTmhl
Q/LKKsTlv3KNvTO3mtbR4uzT5Xeh4znh9fzsrl/YldWcZSz0HsRiUuy8Zd80D/F77KdpmLhVNl/3
iPN9VAy4lYXpTPPNtJ+88VoGLOqMZjHanxWksV4mhaq/Pwv8KXCFO05n9hsjn0TS2qPMGrxWPbvK
U4NXDS6nBWkOu4AWv7KBKs6QKhSKkc+Oa7kEApZMdlq0SgMi2/y8QCPeWg0r4YPZJB/9g2nsEj9O
sgQIvZK/o6RdHfADkNq1cRtcZCsL27O2mzGrIo/mlXs4K+5JEzGfVr8t5VqNz4uT2VfxDOpkvKJQ
cJYF+QZqzFtFgS14KEQkq+XUEozlBbL197o3bldbPokg/pCNGDPNRyjd4HTzJvWodooOe3iTwvzx
eGZDL98LOpGDc9wn7Yb/F2Cw/aSoHUKXRZVQVZlxeXhKr4X7rx/te6B7SChhpdt7hCZVdNbor3m7
xaVMzKBw9ua8f3SPFXdME5bupHkJeOD+IMVEIHJJkqvfDZzBrcr2tcJdK4zPnCFLV/nH0YdFshJk
EmvqeNvGTD5WEPuX1lSB0DxHnoj6/LPi7sQmnFqBW1Wv31kgqkfM60CJe6ulVCTcF5xy4tBrAtfd
0ESRu5edMMfV0KN7lOXeHzh+I0/bBQx2ofPWvP6ONAP0Lob3KeRii4EKaVuPy3frZM0sbMmEC3I5
f1xQajx8Y+pikMJSWCYys40h3dDn5HrG4Tppe8tCPhTnG1mqEljmyQiC6aCHdwV0aSdvCH2z+wZm
W/52/df9n2js6YY/9xfOLVrL40JHRhTrU215DEg0oQD+sij+UrvOM49/zpIih+jBW5QFemedeh1Q
ISu/ZBcktysglPMZdEBLvnFnnNfZ3QlcA8bBLocg5nb4T8VDSWti+vUHP6jci0cygNm2hfWvK9hU
+pb1YvBB0Nd8stdgQBIDR/YvETOPOMXgW/TAYymvK0PCxxzcXbZOU+buw2snCOWTH24+kVgjDoTL
XJMcFKmBwJVdZdiZCDzteE40VupSM+nYv5Nu2mfKJdVsO96xGLHe+v6sBfHxyi3/UCaK8lp5TU60
+5QYQWiiMyVjwoONYZaPg5dSt4f/WxkxwYuGN6sv4RczCaSpnnaobseLLM64mJ4DjSDiNisIMP1v
LxvAy9oi10b4MmXpRoneOCSJhsr7F8mBeU2QZvomLFPq49vLNrXfckR/W9nSha91RZDvJRayiWs8
2QjOFH76LgSsGLaHNDHyRQD8POWhfk/ADUZkse+kfQAnJFYAO9KhhXWIpup7BFgWY31pK4umaKLu
eIK1x0cR3xUp4dAQ8RWDxT7WTroDBYbovIawEPC2qI9Ct+m0MMFt3QmASsa9Iw21KgQt3ofaYnXn
D3X+8JXEygK/5mtJ/rhbcLpmvtyiUJQ1Xk+gYBufuQXAakrfvE8UNvUD88qBIBBg+uzxmfvC27zo
ZMMVp4U/7m4e53GTsx3/DvmTMkc3j1GYz3oru/IijBSj/mr3zrkmTFGyG0oYeA5rL7T9VgWqa4Uf
LRMEuszQLd94Nn199r+Oj+loX+iOz1swWqOkUY/yEvnWczYdqvNQaGn/N42ldXLXN5E2336LroXC
YbOcRx6FWBgumvC+uAh1+yCgrRfdjG6Uv+rOGToIBcjpqR4EaXNEwVnIMuh3mjw0It/DbsQK1phl
stiH6pshiRDMswYkkQdiX+0FIeZxA+hxlHhDtoZYrXoDPSj+X6tn5LVmUarQ0LL26p443OUHkwhK
uJKc6Oj2h40Chc9+1UUbajBPFQ/RdWibmQEYfTNqktpmuCrHd+s6cRotDiIHf577nvrWO7ot2kM0
aeLB4Cz9a9VOkKTOMr9LICNSucy8NWxyL2EJA3/AZlIlxXz+oMJyy34oanZKmNdq9qMyhBtScK6C
FRi7MVpAyEL0eO+uJNFFujzBcmWcJH0c87jFJq4lt9k83vhENlN0BQGe7C3hA9lP4EcFHBZKsEWa
AgBd57+FI1st62wtqhu9jBoxrdHh920yr58fkRC/3UIZXDl+lC19PaUVm6kkfpkBITVGEp8AT1Sk
36zUvbxIcPENI2lIC4aIodRrRHvNa4omkjdmgzY5RF8U+HD4hXR5yOpnrA76D9eWb3v3VHI+mx7M
RDSkkM0rpO6a702oa4OEtsg6Laepucf09vixNSkUXoVmpZGE5/8miPhy5qKsU+OdqW+BJLAYRbuh
PMM7UCp59DO4XctraLzzvCOc1+I/krlN7xSTAFyd87WLVWT63/duxg76dbslLD/xPTQTEKbgMbqy
Y0Ox10QlKyxy2kbqKkk8PrMw3DzWVu/nUjJxv9cgG0pHU61ziyMmBhFKA3arWjI6mR/fBrufiQnR
g0GvyNcX4qkgnhcQwPlbB/3rX7ndue9xkhkRWZ8I3yFHiR9F3QFn6/Nsu1bmyAom/tVD9QR+92GR
jicNQSpjrt3ePJphri7J6e5Zl1Ax1ZIAfQVJtuw1DoSpz5L/sfNSsoPXAi0K/hfkoh/XTcgGnct+
siuoDXigaSDfZl5Y6/1P1XjXrCzmjTmaARgrdsGjXGtRo7m1dVBbPzhOQrTie4Jert9Jn4qixKMc
BOtHJrbP54dA9M1dsJVCa2KHzajnbOs/WC+hEocqBML+ESmyuLumLs1xCf89WFrUhLUVTTl1Xha6
/55kBq5tH7Xb2K4se4tkj/5EmjTtXulk8skVqXEHXaEByDDJh//fT/RkydU0f+NWIDPgpKmRcR4x
jeq5epcBasLLsedxP1m+yXG/ZsgNO17h4xPG2iC3CVzx/bELXnPjcK869pPh2ZwcQckl/yAbnS94
/8ayJoqqgtc1X4hdE9o0UgWWRiKamA5L3wOqQ1FeifslQMdJsob20jKARRL1YOdIraZw9aEYNQ2T
3QRYpiDQ/g5N0LRm2UPxkxIAz/dXIZbbEBF1uSBukDQzf31CaEQakP3aZgSbyyrW7HT0K2i0sAG1
GllSAvCvvI+jUP5+u7xp2jPoVu1GoKk1aXTrbNh8i95pgHyPvvFJMBytFPrU+PyZwUsda5EhaLc7
wZE2aB6rrq/A3SNx7m7DstCbxXLVgKwZrHvygLdyCLj7GrMfjMzsEA3s7pcbcWe1x1i7U1UxPnJ6
SH5rjaptKG7suJt3M5x9rqIgqPHi9bC+k1AutLZGrCb5gN/3jgFHpQUs8MCH7uQ9IrNsBhAMA4K4
fmIOgSe01X8tKHij6nVXb5+4LthJFd3mIGkZW6ExGOTMPD7Wf72J8LK2a4fZs5Z/PnwtQOzBHPaM
S7/0kMIsbH9T+LsjkU8hGrdFK8kfmmBBYftayTXTnx+HW6CU/BAy/0MvotygNjDyW0/HLlWB8a73
Z0STnplGPiZVuVeMgZMJv5zFQLEcvKatbrvX0MFRVtQfp4F99i2An74k6OPKxsy3bo/HdfM4nAL4
85n5CNa++uGhG0tLP9PptB50lrWSr7DMypbYSVK/fJbNdmu1sD+vcgF75FYDICpqpEz/S0HgMjvr
g42zywjK0dIp3CC3MFhA2D9EdJDnTcp79dcSwvvpvtGPSE12iK1x4eG2Mq97yuiA9nfYoMq8lmSB
1Xlx+QJG9vMCVJU+eUik1jMpaLFjE5n0o1chRhh7/53Z10CoKgEncoAhMhb2EVE9pB5AAAkZGjFI
OZqCZVDsX3sRnlGoME82yrbtnCiZ2jCH1/y83qlcCwZre5So8EfM1+1B52YtGgbrgJcX4EzpOaup
ggJL3xB5uN+z2UgA+ia/0ZFJCyl+scP3SA/Bu9u7zNXnqxzqEg6d/vYamN2Jk4NGwJmZRk9tQtbY
u6mkmLB9mbUtv/qg98jHgn8zB3VteV3yahre057MXglJmK+2vRqNvMeGwqz2xi9hYcbwbK62eV88
62MD/tnS1gzEXh02NbG4MdfWPhJsTo8rZS2+qqOV72h/aFbQkEYtw8f4zw1BIo6dmp94ljzPK7oi
ni/Kbes84eF5M3gpcdp/t1lbZIs2hYxKVNxUeheMGwcxkwfkQdUU8QrpUSK+MiwwG+aarGB2xl98
/VYxTymy9uRWWZQHasI3lTXxctUCMQaOM6bFZfh4D0BUk1ksE6kpIwY2oFMfKx5IrcSVD6/C8y8E
YpSbYQ7zvQHm/gChcyQwR5/rO1MKzWDx/aP89UkTvmwM0Niarjf58JGIn3bspp5JPRUlqrqIf8Kn
EA5f1cFybSCewPqZWTvUGxikr78l1oiZE9/LlKoXq/PvjCUXPk/j4f4nrtbbKut/9Gd/ZbNzDnDC
U7BGv5Q3FQknfaglqBvlHVjyYY9Wxbc5pFPZ077eKGVpvSt3TAzz8vTilNHS7B+QD8maVj5JxFjn
tmgDw69rBm5NE1UK1HCuY2PNO3Pv+BNIt1mP2ibaMfwJlQpKBExrQEc8vaKynFPPTTqyVBY8Fksf
BkE4g49Xh0952xkRlQVkq/lLHHFgUkbKlTo8HL3ROG1752WWr8YpVrVS0OjSzx/TCgST439LjRWR
bzdIl466v1yLxO8y65pbrAdrE2MkS4ahFM0v4m3wAq3AILnIWRJMF4Es9l9vQqULOaCg9L50gSA1
8lA7Fxfh+3sCJESo44qsnq1uZzeQM6PYWgUz319/O/QO618VhUzVBpWZsr3N+0GZQRYosv280HXj
LuDpX50iU4Qx/IgV/3EEeAHGnCKw0tyK0828nzCKwEx866IHzcTccE2rCpgvpG9uNFxPdoOtqo9F
U4+Ew1KKNUz1cbPjK0Hn6AGWZc23Q8Dr9xJYvkYB5ppB5TMbrkxgiUOAe4Eoq67pZYu39eI3Slk/
Qv1khAwkYfSBmMP5gXUL9q4GqvSV0OlMeOAfAuhGGkUn1Bg6M1F4ekdGT2AXf/w24EcPJdZfXJ0n
FWfj3omtuUCqP7ipAOWOyC6Cxeai49uJqvJZaKwYSIOMEke1B0fGYtF4Wdbg4Ep6//f6eAClEbC3
vwJJbgvdmJNlPZ5lgsii2kB3sM3QBcFQ0Bjz4mfFnW3uzb6VYN5MfezBMinLxDF9ywjefTEjJ5QD
KBusbyXMtZVRPurS+fHgs1dwNUUjvm0410qliFxBDNtxEy+kTIgaqkqUGouCBN67surHRPKuygkj
iokeyh0X8b/bg3ecOvig3IzU2gHdt9wcEXBdV5K9N2OFM7NOQetMikF8xWLXPuh2AP9+dVhlcuu6
jqzk0shqcm234ywJYonLvfLRKE2i0CoUTYM08WSLbM4rLoHNmO1m51AFhBAfSl61TWL7Gw0G3aok
0WoxRhe9mLpKRyo5av8h1w26E32frX8x9beVOYqR/v7BSfKjNAvWJJp9W68dwIhtPDFo/KJFFIb/
CX0QtDCGy5ScvI1kBX3EHVHgk7Z8XiADRkO6PqnGz2ZyPbeFeKrkobgblRtWSUzFB3xgLrvQTAPC
fExohU4b30131I+K1rG0nynJlQc3ahOTwPGLKedleeTMZk0Svfabj9myWG+PFoGhInBJUcBuNPK0
Lbu2Bm8OxxPH7+sRheEDKIe3U1cGlCNTsrqQDtYp5KQtWA83BsIGx/5WmY8v5B53mU7ABUSZRB3b
ORdTIUP1u6VFc+wyg4SA8fWrVOpveNEW9h5aLAq1jsrXzMXgPkxIUYi9m+ikQCMC+bMRqoIQpeVH
KyhXuidttQyQJVm9fdDuO2KXlZHVFapvJYNUcsV+fWLS/2rSVeDe8w+3h6H5Gmzo4mHWvYoii7Qs
s5sHYnOttOk0Vuxlhg8CtqtK9yssOtmnaN/iLkeofA6XqzNFlCYi6+2FSPOqRdMrejC6qgYV+lqs
yaYVGAF7x0sE0Mq/hPPjbZzocYE+bwTm/u/rjyDt11k7NPpIa79CuzIKUGiUqQwCRcOQEjWDHmR0
XvgQVz/Y735ncyojjthQyZ53tt6OdMv6BZutqVIV3KBTYXzz+lv+dz7OnMjb5p1WfLVLhXraOqKq
JeOKsv28FVVCXOIPbBE6Jj4TqEcwz2CXtC+3Yoa4jR52qR7NUSQqrxN4VDMudC2vEK91gR8hJLRe
NoFmP5Qgk7o2TY4etDkol9Lp5JdH5NrliZYLcDgtKKyroBZThjZDqAGa3byCxoj6uXrAoYx7Qx3l
eIlt4AIYYrsy3TympGmcpB05QyrRkMpRXB4+MvPyvupNWd3Jd9VGv2J2i+2dP8TQQNovCH1fgH5M
k7Z455IH2tIppwwgecMOXx7lDJQp9JmaHGvy8R4x4U/umj+OvgXkWtweXUhK5oUBnz0vD9Rm1MxH
KaG+oSqL8lBzlNhZGP443PRskh6/55D8aFNSq/XXEh2FH2nHf9yIfzV3RlOu3FFyfTZDWVj/E9XN
XhSOCnnYtF5wYfZOGrv24mMCpOzu8csigIr/sX3jZI9B4b6FvhnhPv/vMrhzQ+C/OP+kkxrkZWgr
/HMR+NypuP/+Apa85yUFnW+ibIqbAtpxC+77S5YU1c92ecfNbJNzaUZvlVfJ1dLuLGyntggZlBJe
o1b0oDRkF/Soj2AhWG6eQFAL9PDnJN0gCoQdEpLrFed8QWzVn7GPKY8H27/EvmNKAliZ3AHYkRVl
u4VDoZw1IB62CXNda6PjOwv1zIXjJ4Dp4V+PJ3fq7E3AqaVTWWooWDRDFQrwftweokefLhc4Dyqe
kgK7hjRoBs8syo8Pa+EZmf+tI65WDH+WxPJ5BeHEXPwKc31Hz+eEJH9dINQlBy6vx/V6DmJN7Nlu
cRUYjTERI9AO4EyAJmc5bpOqt9iJr3/a4dcbi2MlRd33SNKgEMfvCh8lFY/jOXQMn25tw6dWUDdU
RUEAGNp9b6Ffb+ow55B1XSxx58Vdbj47RP8Jw7qFvJpX2hHGRM2SgM6MtSaueVEb+sMEyOM+JK4Z
luf2MuI8Isjn1kL4Aw41dBZHgDBpSEs/DxHbepGAJz/96kVr7FHRCxv9ltres248Q8Wv3n39ukae
A3XY9KRm9tezVlCcXSsiE9pveAtc9viOlrMzLh5U5kKhFUwJDNLhA7+vuSWCm9Z9WHjhU/YChV0s
lQeUrjr8G5SO5UifiZOTMSU+j1SgnF881kjCeq0/kI/R1BiBIDEGhMjmEihfKUrJw4XXR+LU6Gyz
4cUM844Sd7Cnirn2RlB9WrHNTtkOoqXoMZTUMBFnDtsDLyrujShAH+3dn204mm70Xb5p9jPYFWg0
9Y0wR+27cP/ddT4lAvofvThjGvw0i+O3z/Mvp9po5E3Qtmuh+ZZLrTLe3bMv7yrylVJf61Y2XW2e
gbWeCchbTzYx3rPob8dFHG52u6dk3O0JhYBM2dFcKCaWA9MpEi8ffvcUA+4jpnzr4wEKWqOw5KSm
s6t8s9LL2kyYPF0Hqc1/Y4iINWqXBxqoe21xSR+nhRlLcYsi7IB4O0zxhpRc9CxNJ0U08/LKLR0T
H4PGAMq81sD2Vpw3Y7mGzUTaES0Q53sY+BQ4KQhOmCigNGz8F7NhPrjyd696QBPmC1yoHxv1KFV9
AnG7RelQX4NRkYdtQsOUEG4BRD29aHVAwAzaVy4k8Na30i2cOx/2no7QwD2JF2BYd4ebUh48U6Cx
pTwCpZswubH4wVg2sjvogQI7FxAyqsuanJPDDef9PnIoqKc7VgHwOMDzenNauUl+u2HylRNj6vy7
wgJNbyEnseo3IcucZHV3kn/GX0KL2OaloH2ULoOL1SgM45suJykzD2ulTCGDbdc9yTABRi8rBcRK
tTcYsSN0QbeGjmd0jnm8Qc1ZJfjt0QMtHKIDTkSuIpKhQK+3Bs1EjXfL0iY63LUp9mFA7sHh57Ia
Z38smOpcBH9IQ311GDRlIYAiptBIE3zJnUtW8Oe0hH+7uNqnK/csKYICj85N1g/0aInU2H6IdAXr
FAfyDocaCvAFkkQ3pch2boaF9IavACrzmJm8F8RYF2BVlj3jvKfymSkwjqBST0/D239+wK8gTovv
nQuVi3dZ2qq79AFq4apIe6xcmxvT8Du6SkwtvG/Qyp9vu+ZYi+xtMid5JSyA2KpLpvEUz/YYUu8d
RcDW0Z97oxDDZizl9bG1SlG8gqYQKqdVCYxPfiSMoCl3QYUqJIUNldYiQ2NFZMzO4hbVO8jty2p3
DC/57lv5Aap/UfUxr1NZgKNvItrzf/s9UETQDj6XPCdrXBHqdmiIOxONZWelsdFm29R6Ye4mEHyQ
Y0A5lAZUvtcm4TwSAuF3KCFisYR+QqPrO2gRnjOPrQTJVANbeMY/B5+9CVqZNrUmCDwHHeW4kJnP
iTjQgxedlawm3CdT8vycfqOKotQXXfhVHJu6zQgD8UFotJfEudcPDkNUiZEeRBJxrHOS4+poGIdm
V4MCuB38Nicf+bDS1IRoQNCR+ukrvsTVi+/3e0kLluMBZbLKS6nASd0JqBK/uWkzBfC0fxfnM9go
LIN693WyI0SaQfIuhOvyf9T87eaC67EcEv4F747456ts8aePAJcEyhrg0pCZQPVrvCuh89ap6FQW
geqUke2evQjFLgbBmRzJG7QigIfb5gX0p8gn7mMFVWk2GrNHfL1cs/01Qqw+GB8/RvuxHLSkcyae
BFibUwtTibLOGxt/pthfMsweEyjeszVdCxyTXRol1gD2uhzZN69gjXc934SvBLhgF2GViyk+eiQi
pe/sgdLCwO8VA++Jii4Q2zv+CNZQxZaCjxxJUMy8CbM6+47sAFNDX+fR8PzEZ8qEw66svoSt/Pe8
xWRAohPTbWY01ko4ZJ2sjAxM625+C6Ztn3IU90BrK9DCTHSA8pq5e/pipbx6tlAsPowlC1a/2owZ
zouCHffw4GuXNAOM7YybPR+LHIvWQo2+EHXo7m9NwQNeavpTuYOlRcjXQXdfRfrhiAkia5ibcnTW
uy3utV7rEOikn/PpY+FfOJQMneWGJ53QShReXxldSqrRGa/M7fbRAyR2lMxnZ1uDJkFt/PH4W5Ew
VUDmmLSeSVjhJui3aaqZUePD1DLYFv1d1/iBmHIpLbzpMRy03IrnovbPfjk/VcVbGZ5ZS73/cWEQ
QTg1oSM62G1bpgG/phCVz2piRzLT/pkFRtVU1YASoZEp9XYZmofzMQKCi8IUjlXtrrwVC2ebpkLX
ldPCgDdY3DMW0ITIqg1Q0qylJxE4CQTMx6d/igAmc8Znb1kKRWAE9/y1zhk8o5qe0dKr+3ctoMR3
KNXEJfLjcij/Ee/JEnGGn44OMMTnsj5mvx7c8V2vnRWjnlJohzWLmZWBFPuKghDJa8cf/6L9anLo
/5DJcKy7EmFhAVMb5iq0pKNokf1FH0hLB8i7sC5NsbfTxMjNgclLOyyNhQgDY0EMRrqfBYhJSls7
KV5zuymm2v3tnlIUNw//6jOTA6Vy0wVqoIzTTOYAxqqzSdZwpO5YKEqFS67kPSz6TiyCp6FmDrjH
2TdsgaypkiRNPG7cMuq5td9Te1VVYQs84tZHjfb3G3aIlf1zIKzdSKvVhgslQTzLMgJh3fWySJG6
C2aaLOEOjrCnJU2eoWlM/b4jKefDnwAyUU9vPxRKsFE7IYUZyRIKbpw65I7Fq3yC1/1YWrmnjDv9
L6OD84fe1837w3BVL++TLe+cv5Lhj5XsixRBKWVSaOsQ5d3WjrzXxrI1UtyVwU8h9n9s3dBMSRxm
eToybMdpyF8UlKt0M01VSFkz5uajDGahHoTfp982tQ/O7H09vWFdWGpPhpFKO84avyE+vgwsxveM
9VdrYZ2MD1Zku27oXmYe90yUPeVC7V85IL43PaVV5Ow+AKjqg78hv7hORQ0t3oXmavjUaa7//hk+
XM4G0qSxkFrp7aaz88iG3L1MO7OOVAWkn+DRih9xhaZ3XIWEyFYgqomeMlsa+Gzh3UQYfoMgOmhP
LP9B6HxCaAteUTRNmNn5FTqF8CFU3rsqFMZTLunsvsN84/vNUy1Bp86kBNSFaoNCafveLshtHshA
cnyOkh5Mg0xwvoTCE4xmMfMFE7r/5lvMctspEBBp1D2bHxHLFdIIFnFSWTF4YE9LVZ13ZGJRldSc
i+bJxVKq60qowkNgLT5iHx5Mx8odn9DI88NT3yuQPk+bh1+dDtgTf5m2Q0IkQ2SIOCYsPwrsaVSq
JfqqLZIgmxMwGVMURgOew0kILQLeu3bkSAPSFebfwFMgwA0slGsV1r5xznVjGvavZoCNOCUBPldB
Xs+aXth0zS4EAvhZ1YjfZh7CX3z3ylusl0H/fNrBU3sPCh04jejsJPjGuJp4tE5pHkMyPp7R+6qq
7LG4LtFzpDqtNjb5frdsvqR81aItNZXt1d+oCmeqyfDYDXSg0JQ2Z3FoWLx32VcFFsrLiWRXFjfa
Jn4lXGuArSrMAWMie3PPm/t5o9pUTvDfB44SzYRUBDBpEm445yOTkJMibgESIewhYDZg3UKdrzw6
hbfCjVLb3PtpJTFcMc74hLcRsFaKhD/3mPu0veLcFONyExXK3IVJ3GjeeCEoFIY0GbC+y3LviOiv
UCTLJoij3AIag1oWeD875axiZcNw9vjXfymltt3PQ0TWVajjFcdPZJZOoKSdD1VdbDpvbOo4X1uh
cRPAZwVoM/TaZzgkcVFvj+RbeGd2VdMWOLeSluAHuRuQLDImgXGqS7wztKGFZh2h/E9TKkypo9UL
TN1d/UkSoK/ycrZJA9uPWy+h5fgI2kPyx8pkpidmLvQsohmMICTy7BxfDB/c+fVtFv3IGoOx+JUq
DMFVxypanX0VarYJuiQjq48zFF1SXXbElCak7QTlpPReYbLVp07RKiIlgPExBFW5Pg+LTMIh38yF
1plZ33wLO8im2f8+JiCBkWU+iOCpSxUyHRcTOpTJmvP9IfO8hKPnEyq2U28t6VbswBnWq1q7gmTW
ntWU5Qd+bF5q271b+jVtP2D2i1X992F1uuB4fXzj0ocJy2rQBllT6KH4ET/E44SmrmjEjGWMJ+st
CYVn+ybjwtTSVUg1dvycKBqZgS2SsvIeOlR6CL5PF9uhGn5ZcODhu3F6fl0+B7Vc762JiAc8V7wm
oI7O+vBmISdVnA58aN8oERaLgKXkqbpPT1XvJjhFBqg//P+rEptNFsN9DMLACd2vlMVwIHvNbLZW
zLNMFU7/5b4tbHQT/eCvgNcF+8ioHCTga/P2RJrL+kgIKaW02nj3KcLB9m8qkKbWbFRTSAFTMD1i
zFI8/QBeFnNsEQql1epMPFZQ8KoaLu4jOE8Bgvw3yy1CilenC1Hfc0fR9nUwvMTp6e8bGDBdHgl4
J5um72RSZ8o2bKWzm5eBLfvORFLG91dWKZ9loFROjtwkKhdvatECwchHYmbZklrdXVwSwcGQdw7b
J39qIt3uq1xHhDE5Ssh/ES0QwzGwPwJHwTGl5DosSvuQnTbdsESTFYJNf1W/mahOxlhwQRgGHKTF
Pms2TfPiQcowS2QcLgFq2v8CghdqoHk2wHpuFvl0gcR62MErjyTsU4Yv3MDfN4uuOvwuOSsChvZ3
EwwInOYzeE2u4Sf8h2Y6s9PHhYiIgioxIw5zLP1Wf+CCvsXubMBUyYH7jMDowXyCrLQAOuDcaBAv
JseLTkIWcMzGu7RYL0Ymi7gfxn2tKPg76Ry1WpKvRSHI8Swp70/ekAXkbI7hF16MNkNfPweBG/dk
zCuY3O4TlBOLwxA9yVS3zCZ+RACiVM3YUN2uNhoczt7h5sTSwSqTfXpWIGe4queJ1PsdJVTu83M8
Nqa5opA5a0XcICe6u4pOGde4FKXMgIoQrUsHeDxDkhnEQ5njv8HIrzwdpCM/7k6a42LOyFhFY0SP
Uc+VjwKx3km16w9ykYWcWC/L1P/sO4ewjPxmKe2orMQ4UgBj3B6UKhYuHTQI1wAQ5xDHwEW8cJZI
wHgtOQtz49WqskAk5n6S/yRdACOk2Rzox0LV1igVilhT/VGTt0y6YevoKIrN0ysZGdjv+qiQuNSB
7lbbdz8NvHFAOuY4KuEpxdZQ1leHWIn2i3jvTf9YMe3vkbV64OQQw0QN2IoI4+0MW7SMfk7bicvK
qyclSd4EPCcZpgLMeIFxSp9YCukrQuCtB+UGAv/FyEHqcXFCej2P6SluxQ60n8QSBsmC7zG4lMkK
H0Aok/9amx7hW1p0oG12gl9HkPOmfOvoFfwpZaNU15B2V4u6HOGRmSpUiPMsajlhUE5+ROAmvT/W
4FgookGBsUNdx/+7ixlvblh2hojOLkzBHuUyihKt0wf/qZs3lmeGrYU+eFPsDSKu83hjHorDvCml
wEoJh9/FlUnIc4T2zNKJ0bFFTDT+2Lr+gtrT/QTQ2ZhWBjY3hcUMHHrFIOBKQEZjZbWpp9cb2dpg
/Yil8QnmlN+a5sJ9kZBs2vR9yNg1dW1ZT1Kg3su1fZ7d4vqGy4w2EgLqlHqfv6HKziuC3Vwc/L/c
tpmMiK3V6x7ztY/GUadkI8kpOi4X8vxLmz0MgxKPLihDHc15ncnPXRMdSmwZOQTLrqwrl2RBMu7q
SBjMalO8zfhy1Vy/SB2IJJ6g55nBuTawBBIAa0qDfEx7l7TyjeOMCToqz+dB89kQwZg1G5hLF3FN
UEo2Iq0gY32gw/jDl/7gTCHAG7uCHHrbGrlNANq2hk0IbA9HjcNtcuuYDmI7lYPZptEX2ThBZsY6
D/DjMXmALMbcFWT7x7fNWAq+7vf47TJcPQzlQW5+9f7PQvS+xT97HpW0owGNZb+KjFdUlI+NQ2E5
J5teHGuyE4w83Q/PdeedgdMXRtmrtRlxSSn0kcUZgY1ce/mX9/CGO9tcR4M040RQvYCNubZLSBcN
IhhOBNXeF37dlbMzRNdMQIdCoza2Na/YlXpXTo/0CYedg9TUJYladyQUAyS9QG1YZtU9jrhrPFKK
UVLV48Z3K716ulN9Se+ZHWK6sZlbDNvrPYvH/9DUGYLomUn7gV4fcaPgte1eUmuXwVX3sCHYN8n3
P+Go3eE0hH5BY6oggFNbFZ6ASNRMgW2kdSzHGOjphF+CNi4MG21MjcVJzUDqBJaV2M9anbvKLIRz
zGqd1n5OjLaQVT4B0PgTXMuQuTlIXMpbFPeGkPSfnc50VLlxKh4AyKU4SKKSaZuZdAk6PpwWYZ9G
hK44XDTwTwl2bxdZaL1wicafh6bk1XJRnGFcjPkJH6uqR+9FSgmeilyapkAHvGbdO9nalsWYknKJ
PfIZgKWYexzD8AUuAljo523bWnnWJxW+hoO/51ufYeRPa+pz6tdCbEdOU1bXdsCM5apIJRKKFK7M
kJyoegu1Fbc18JlNpGw7BjdsBLsWsCxyq9a8idsahWRmf2EvpiXfltqU3fmuvYxD4+XwwXwEV9cM
LncINLYaGWa106b6BdW6UI6bpDgATk7df3yXvhV2GRo21Y/a9OGYJkH1+fsY93Xyg0PRlYpnGl6m
w/sPGqKK+rg1BXdlOErk6XZAF9nJchcGMCaTOwX9fCWL4MgtfGAFq+ByZOK3vbP8lssrakr19kxT
oUsSvFE2WwyobKgKogyWtVlAriWsH3BkQsoN0yM+LiHt6S+JLNSv8S//pTlQTfwWt8kWIJXbOoF8
OUlw4RDB/2wCtIRIE34zq90LGxqQ9pgqZFNC0NI7jlK9HG4KnFW0L7iddAy3wYLmWgBjgaIO8Ev7
Wuagx3T2AffAbh7vOUXAPLCIa6C5qsTYyCrzT/nTwgKeNSvvoiHNRBqFfdlvUjqyiCp4FEk8zQ3h
T7K3yirwSKG4cw0zJxvZplc0UL5WNSU7YCbS4eU8AwVOt2aV3G2k22/EWKGfiOqyxhjr4bIOcmb4
p/Zw1YIslScONuxgzoYgjrMII9/LrFSKQUXagUhZm40WeRz99xj09w1aWnhpWGbMXQqauBPJgeBv
H09oizmRcqx7WDclk5NgamMeudXLO9BKYBnvH1J9LcSBbrvULH2g9ohO3JwYWUYhW2phYwIXmrxH
OouqfQsF2MEeVPjGpN6aJsHX16aCBqpdxxUhTD6R2S7omxiGBIAG7IMxqY2no9XUVy9q436MXuTm
YZq1/aLjetOmLySx3rlo1yJQYS717jz4ceGgTq2uLxT3NWyoT5DzEOPliEYBzSdu3fAr17bdIzbu
7Tn3nQ32PKcnfxNcG4zBRuJLm9QaO4UjL7s6+sz/lztxy3sTHlUD2PJ6Ke3kKM3xIr24A/ahUDCv
tqq3WcYLZN3OoN8bi8dngEE9naOE3yCFHuFw13U60d+Enc8UlZj5NwB3Si8dUCXR1Zph1o672OV9
qcjDpAFdkTI64hN+eW1MDTyzqAdpGs2q6QvNfF56bXwbScvc9DwMSklD13lnaxTLwJzkbLb9rjU6
gGFsdXEwp3KH1ynzfPydth37vSBevR4bSUEDzcxFUxer69SrtDEJahqo8CBSTzyiU/TYQUhLW/QS
lVGiJOz7bqXG+v+5oA9iJ4fwhdIwzuLbft5o8npuqM3puqJJDrgG9+UKMjrOAIzIa5XXh6sh07qH
L0McfcOTKFCCocZn9ciotaxoWD1o/xYJK3TTPjSaB95vuyPu9+d2ivLRjxlSwAv2KHx8/3STh0QM
o7Vw9kvv8LSjF+FK+TV7acDGfDhUfsjNS3cpTy4xJAAuXl2Y2XPUWE92gOWJBstbjOiHCZ8ltKf1
zzveEW9oo/tOK9+90pXgHu9LEi2atMS96K2Ek7McInZS2LKmuIUPhq+9FcY2Dfxi3tfmP8zlSmm6
JZ/d/wgps8g7uwFWrf7sETtdPPRZsb0QGusd+Lcoqsup3B3arLNwAEKwjmU00DB81uYiPReth5Ls
sLEbmhisPGdrVZsCf7GgMQsHRlSag5p+NZackihnMbszFFXwwpxDxm57G9boCRMCRZKij2HaV1mj
BHF+5Ted5i2m+PILkoCTCHMsq2mPeIrslo96CLOmgaDPT8oGNsSF2+S076A0erBFwQHXJ2sNrvx7
+JVU1yfK+CNMquhil8vBcfvg2D0GwL06/gmUGHhr+Mt5KR/N8r8ttgBrboVTtGfXjrLaE3yWQ6TI
3nvy05T96aYCMs9J1bkK4khIRpQfmxHC5gQYsIzcnN69ji38ruUGCKysZdjMTwDg7QlX9S+eYd9L
/OyMzhf3OF2IOhgJgQV+cPvePOsuWTry+V+BaDf/p/AxdybIBj6EvzzL2LDwxjexNLlc4ikxrftB
4ntafNRhMhOkNbyPf5XjMmjKJJF6jgNg9EAoU17z01za2o4jSC7myjLUxQUfRVyiBz6uZonRhjUh
ME9ok8MPjS8hcji4hWDg1vpKGjZ+Nb7BtE0iDjFAtAHwpIkn+KzL3drOV98a1mZwsAmbmxS8W6P+
3s39luV/tX5a+/DmkmNUFRBH1edPhInxZs+6lC44MCNIO1m1hYJ4SVLFMlrX6YEUffYDe85NA5xW
dBVhN4DeKlnkFXfTljaTH1usiN+9/kyMTg9LMoPFcGa2h6+i5e72A1iwP4OGrd6GG+RihsSoeEx9
QrONx7A0MyDH/VTGOuMB2+i9gqtpxbpQjw19Lpg4Il84QzF6ri3BSE9vfKfW/Pzr887we3xQwU89
oYH0gPZu2e/c9m+sX85jeNC4PQM09rQTs5wnnPeASK2VhnrAsB0otzokNO3IrqjtvqNT8MbkZXmB
mN+ADxlxtMybgzS1x106QOGw4foCEJoLq3qCm2WDJcT5EbC6e97WiV0VsshTAS+SZlhW7aOg3VPw
VrPvtO8DQSayv1e/Q6Dh+DzrK0SA6SzSIBFV9YANZR8R3PWndHpi7cqOifiqMwudjYYUKI6er0Hd
DB43u4oS1nd4LEg1j1EBsW2gNyV86MXN0g8X13X/0z+Sw3AS/yloSMfryN6knid0SHpIQWUB8OpE
t4uZjRz/3dRbb5mvLWBC5RvOTOoy8fgB09VGP5FQd/jSIgApRhAqmTvAD7TXmOqXHzegiGElUkbc
5i1nGRl5DbCrh8T1wZvuhtZttyLasOxhNMfiGvBkskEVCG8OwXhCYtH3Nv3dvmr2ESkLL5vpdd5P
9KaqbZppP6sbHBoEfhl12j9za4RmDSdgEg01SnOhwk8BpxsYMsC4wW2bd2L771XzPHOtxis+Xffk
EjozUXJW17mtwxVb+11J6n2MEJIQJ89KTXyfVPzUcC6rDz8uRA0E7wAvvXDJpBufiPutPBOAPmnx
Y0jPNMyJbVZ8iHjy4Cy0aNsb+lmPiW9R2oEAs+pCxo9AqLD2TFx0ha3sDgO+ry1saMnuciZlOO7G
ALGmtcy32bbfVFwHa4/WgEKLEwnobvGvpcxTjviOZFCk7m9pQvPpP2q3sPjsp4r7J48D5VpTldbC
3VgwQPf28cVAlPqJknLMNwE62hQo9vjrvBEwsG21PvgH2XRjdL+UfYVVI5M0FaxWrz7g6A1HR/n/
9O8T1eutE549Wr8lm14aZaqA6Ec5p670zasAciANzXsUKZOiggQKRbKzrKxydVwbZXPuOrvruneB
s8/Wyzgitk1+Ex2LqdlcQZbCkD3I5kZnRG8rlfNGqCja9nMOggnsD4HJH/4dwIA2gtLwfsQIrKHv
b+5gqNK0F+J3s6aUKoug9fFzeH9+RpqvL094G4tfYSpKjDnWpRDT8KWja0j0KBHZHjFLQ4XcJC2f
79UoOJgb9xuzv3PvGmWRU633v7KBzjGRD10pP7Fu9UdWGaVTij4/Z12ba7MMOxUplnssDtIvXJt0
oj776hCXdiusgNl+ceAnUrcxwUicVf/F/y8Hql074MpA7iwZDn1Av19RDksvBBRS/y41I7dpUHT7
Kaat7wfNtrqQm3G4go8kDFP6/199mBfOKhZErv5IQZ7pGP3889WLDEeWBppm4GOYo4mGlkQGMJTg
o2z3jTszCy+brxZPi2xjQv0sZISE3wg9NPNYX0g+0FlcwgDistavMacaxvSLWUG4PCZGMGDmNCKg
EOCM5dafSGsVYXQgV8ElxyLXnkr7rqg/cBFhXJgIiRV1Wu40i/BvrglaXB0rRmSD9IZIcJxwq+lE
V+1T4E3iqpap2c9JqDmkCoBjBIqbHuf771YOzPVKWnSBxefu5rVus8pGcx19048hn9ypMNySDAF2
dNCRNz8/GBpi7ArvV62L3e+Zs4VMhYxSyQJESb9ZhppzkbBsG8u8M2QHTzMl1BrjoLovi+qK6W4p
VxKkmcStb87vID1fvutg1xE7m+QR6c4RGPDPuaYMAXE4YwlmLaszDAXfyFPy2EMQDD4G9kCwnRwu
k4SgmUXrKwETYxcI+Yi0bLl44IOJ/jwPZmK/sTJRUTPgDy5I8Y0aycOMXp0KwCDiMiTpEnKYSxBo
vCKrXUI0Eu6qt4v8W6Ixdaj6XlLtq/XxAbmbn49n77BQreKEiyuJ0YCg6PVkGvrD4D3jBAgDQ8Yu
I+c1oj7jsTuS4lWN8irHXi+odRNrmqHOCpy/vdiWUX+FEH5raDNUX4dOwS8Htme55pAKuUkF/L7D
2b9ArRGpTmq884u8nzLe9vsW5KY7XDjBMNXTS9q9VrX5D59kK12L8ggA6D/uJcWO2F/fVl8e+okx
t7r8y3zGblqTW8ELEKUGLtQgCMA8HE2HbAMgxQXDzHZbnioKFoz8UtnCXpb21CzpwD2sZLg6nKXV
ek5sSVo5ISNCPR/lsqa2qwGSkDvheeLtWzcNBc137BKPqinPS2bNcHX2EqirU5Lz9EHZcdH6HPRb
T8+BtCO3RcmketFYTJ6wQvkZzdDhKg4St1qJzFEhwf0MbDZR0HKNxz7IF8iSrTJHXbNIRPmYb5IK
noNFbEcTuXbJmEIaSuo8DKb1nBJ087dB4rMK4cmCPSha+WoEEQPqvF1oorGy9CQhNHgC5juZ1VS1
D4OZKFuVWjT2TSxwCAIGWlkPBRerl+1DH3GqU4uBQdSchLw1KAdpfnmz3DdL9D1jWE5MLakaTsRm
Xr1Pqe8tLeFn3/lgdYFtpilPPdi1Y7apzvgXRW58mPXImQkqbC7U0AsjxgzlQ1w8mP4=
%%% protect end_protected
