%%% protect protected_file
%%% protect begin_protected
%%% protect encoding=(enctype=base64)
%%% protect key_keyowner=Synplicity
%%% protect key_keyname=SYNP05_001
%%% protect key_version=3.1
%%% protect key_method=rsa
%%% protect key_block
bW7pw2RvvgrUjooo2We9GEZiMw17lri1l86Vx5TPb+fM8bhfhBZjEPBdjPnIvLfMTc87BLLyVGGy
EdGw1XXcMm7BrLlVXm0SPLRVGnho8My9GpOQx3winxgZPJzHcudCa5IsufXTBwdg3pnVuXD/ytON
KbbDwspSmJaFBVxMEKFj7moU3ZnvHodNdIA/6pH+lvxaK5sbexCsFTfAUyzYiz1hpKWz6cNBjnUw
IewvSkpK9xSw73ocGAHvG1I8VhULp09z/qSajT7ogM+GzHRvjQf3CFa4RUaJQ168utsrP+XsqYkY
V/CdWgfr3gKcuyuyI8u6QqCwtFW5hsUPUe0r3g==
%%% protect author=dw_supt@synopsys.com
%%% protect data_keyname=DesignWare-2018063
%%% protect data_keyowner=Synopsys
%%% protect data_method=3des-cbc
%%% protect data_block
5+zeyGWvlujl9cQQQ//EUTtuVkZUHqoTmn+c94fRQa8PeQRTKiim0AEj0KxhNKbN30xQBEoOLEaJ
etK1lHIRef6vqYMXmkwB0NZN9jxBp+2ddD+LTdeNs9qXVcVQqmevN6GowAn5nBULnEfklQZlmG2H
UseaSo7Sw99GNsF2HIvlVn2ZPPWhazLYO3eJ9VuBlYF6I/03kUl+Fqgqcw8ng0M2mb0UDF+62NLB
6oMjrT+xyt03gt1iNwavGy6s4N9DJrmenFkF51VGLZ/k/75yW3541YhrazFbIEPTjAMv2gSaJHcN
wP1mNZYBo0hCcLfQCYEMTbMQ/O6RUplsMrgf0by7A6bgDdWHS4yI12Bl3EY05WB/Hh/SGuUu8Sjf
9Zm7mE0wLVe0toWlC4aNUYrNUvD6JxwNs8/NnNQou/Gpd0a5OYHnMvzVZU5XBdyYff80EioS5RI0
cPfOapmOQ4aiRdxreKSKENWo7DK/zlHpV7yRv/xdHRrqyeiOf62/POg0n4Nvgfpdmnc0p1qhGET4
ZfE8uk4TJnqKDLvVC+2YAIde6by3Y6PCnBDd20ovyz44O1hhhHrf8rKTvxOw/W75OGUJSFDjYEnr
bL/ertdP387eeIqOE2y9SNlzjs7mmnH3xG8jSwVYkk5nFhuO6Nxw3XehLUy+jQ2Hsmo/A+E9Zryo
qLIonFOlBpkery2ye+QMazNMRday4hXO2qhhCPP7x3hRd+z1GLjD+EWFyDnsra5FMfgZfOkY9ur8
wNdkAQGODaGkGzE1NL0tAJBeT9sz9gAPkzNFUq/D442T77YdIxTH0EgRckou9pW0m4Ru+rJGswXl
RJYDTE8/KmbXNqit3k7rSknRNUnNjJUlQBAbv9RKJEX0UWlAmVkDfHi8uvyKa8wgZ1fA7v7qPkBt
sBUcAKlbQPrWcpnFUktNUXF3UBipTk/A/lmbW2G81fLEw0TOObh3bNif3r4eFAYhxZTzJp9jTB7P
sgmxm27i7A/F7BZ7A3zlWpSiRXoN7z5ehQ836PE9cXP0bmiBK//YmRMQ1L6xvbGup80jOuR5dwnJ
ZKxsQ6kfIPWmdJd0DfpjToYBbmbxs2MO+84SFOyor3ycky4iVEKmdo63UQ7Cl/7OI1wxKqaj/5hi
U6EjBkrlMLVRQhCHlelDJPzNM6tTWnuZpPIxXG/FDdXtQ+OI+U7ihdcjmoImfR9wvd5uprbX1YAm
S0WxQb4bIi5mWx0yQ1lhJK3noFhbDuewviALgihUc0ekDXZ6ccpRTfLs5q6Fr2wGM4JXWcTFdHwM
tXdh4BB46tsDt6Tj0xmRobycPgnSEVXSBAFijt44vrHE+bus7tIjNXiQQ0U7jp4cypKBsNbbbNot
7bgEOuj7GEom40aRzCHytWJs8Xe+s+lmw+0PgTr5GXnOq5v72pMjyyF8ZSyr/Qkl0ty2KjfPyb5W
viD8xFnbRn7rxOZXvaap0oOZkYtiWCjMPn8O4SxCGMMYTqRptIOK1mRC2Q1czcGLs4vLkir1iPKi
CJSnWLEWQmDewPHPfWPB3we/CjszOa6aKQpENjA6FjHHnVyrHxKDv9oNR6wlOncRGHGMpkbmLPhw
UxP0y5B7RBI1tKJcDgl/AH11ttjeesYlDtHC7Hrvjm33oH130zB7/iyn1+mzK9OY9OTC/OtWMlIv
oGs33lkQ7Jt1N1U8kcR+Lkwm75YXR2sGRB81zDpsasX6uSrzsYbh7dfemjmflbmUb0IGvVIyk5Hv
fwFbAXRXcXZE4RNUAQFuKIRhW/ehYZYr5QQBRHvwP6NZbh1oVtQx0wzWWpPV+6Me1mK9r+s48HyL
f2sJjMUWcs1R5LRfaO3Ier9h7elaECptX4rmw8pVslVSgFiK7BrMsm798s487k6AUpSMMSLw3hfI
NYJC9AdiIFIfXlVb7/KwHnkCcmnqr0tDm9w33FoR+vopvJ6vAkOOXz9cbJjqi4xjYO+Ve3XdmI5k
q9tCsQMXiXtQJhW/RvR1Lwc5GmdwH4gH9KkquDArrTd+eSDWHUmsIB8vsJHxRYlFuB61awAWl13O
OZg3z0TMG63+jm3S/kqwM5Zvd3AgGtTrsex7EmrcPMnBfIN2lAHlPGt6k/L7Hk1oKXgjIJpM8ssx
cFyQu7z2RnQISe5giie50EzQyJBzevFKOmPrE8/1K76CswDwIs0239vEQQLGJ3EL9TcyCKguFGnc
hSMXK0zDZ78+79QShsJVhyQheE3JjfVXwcpjyuhptikkDZFtSooDam/3Utv2Ll8NRdruRN1ckCGD
8Z8ZLsmEjZsMQUkpArRqgH1oao/MBry4DE1fwMQiRj5fhxfSCH9/EuT6J3tzTOakV8Sb87gcNm1r
qd1VIXLtvVCsVZkg8BHFE8PzJFsvb0pJrIhj2M6lWlJE20RDnDg7XBoBlaylZSImHQldkRC2jxi3
xVwDKDGXl7gT1n3uWJTGzfDgWLnlV/fStz8UihSHTkH6A3aJnDuzZjXwN1MELY+omFkPUH43keAr
onA4m2kVoH/vXv5Z2cOkaN12WdM91e0itOCAAfUZueNM05+gG+X3qN/vOrx582yiaA+tkGMGR4lE
nQgZmUAgrtFzEf/sXZj5TobdQtfVnl1WhWB8rvrOux9n3h5u9GJe0dZ3xSAFJ/HhOjHaGF08vQwW
D3WJAopCbEGxiAtxN52FgNx3ujQGScunfj5igUIvCqgH3IoHKULgRvq7gWs7aQyBC1miAQXEbWrq
pxfbHjOfuHIrQBiBXGQSrF+3JPDCX+I4rNuEbiCFPhEMwrkRxOW7rywJ/BXylFaPdfT1KzS0/EGN
p6cI9A2Hg5nc57g+zfWfWbHSD8/c1SIzWgl8LdMBL9RJpDURrv4F51GAfQeTqXtdCuUktXeroFe1
wsEHmS+nZfa86bcWxE7HswKuWdZQW7ik1DR3QvjEiQX7efvUxyJIJNs+xijgfclWHPD6IJSaAqi0
cv/vEXSNf+VIMOWSKFATzPbYKyPqajt2gNGcMmJQdzUZLB0LoM73+6CjIzTPf5PHNxE5ooVBkL1Z
ZF2RrNLVSPNpU5bNxIJtViv96aBlLVkSmibLeXUlO6+dDO/obUdjq5QAvtgJUzvYVYtwm027knHu
pUmmebWUKxsQQZa3eBBsGLJu6GSjp42o4XuWZ842uCjCef1hNRwL7w9SLD66Cs54Z+vp7hRSJZB3
bX9jF/acU+b2DOcVeYS0S6EG4PNmYXr3SGT28dvTO+ZaV3ZwWXgkEYe4ENm9WTf34Q9IwOx3lyMg
/erYrqnGnIm8OipZOhH0oaTXz8YPdjA0F3pWESyzB/OBPdI2i3MsE1kQn9cNERzyhGLtNdBlHQU6
pe2LHCN2I5/C+yWfGT2DPHUx7zvfB+fcQRXQOdqm13LYLC7a4smrfVN3dM4DRIqD337FlDq6RT/K
lHR0gP0u9vkIg24iO8v0GOKNB4svwaiUabvU6mGi3noyMhVbQmL+AsuSNHMl2NARJs42dWIZE2vB
uIMSCk7t7hg7K3elBcuXXCBxl+MafEzFsv0FHW/Vl4pl5ItRX1svMGXJb0C82ub+Jk1VM1b/uMto
O3nTF760dhVS40hBIBUQpkIXW5ng3iN8+e3ktS4pbiKUxW34zlpoI0EbI600bRfM+E+IO556Zx2D
4ZRqrhvtQ3TprM3tmixf7q2QKxFBqKr3bgYzYs9oA1fpEHuW9W1OPXAgN5IQ+NHwelhx7mJE6HLM
bvMJLx/mQ6MuFoLo2J1IONkRFg7bC5NWHVswqD2mFHwrqyk6Z8pR8xg4hXUAm9BDsJckU8zFyESx
ioWHYyGUrzA1Rt58izh5jvNLH9o5wTRRv3OuhqkhwMpbmMeR5l4M0AI4/e+npCpCb+0ooT5O+QaD
Syzv7s+dTiut/814CJ9c2tsnhgRTAzMm1HiMuSoYDOAGGtvW/yrQtF0/vq66yQpDMwJy6GufWXpT
/b90L+ekfJlYk6WgE3+Q4aeJfxpnEVXcn319EE78v7zzAsEXYJSXkzhMJXDu1DlFdLlqcdZ7ov02
r2/Cy6f0RHv2OxHBuEuQpfs0PS0B3KRXIhJDvyAYDgCliP/Y0Blu52YHMGdWQ6282WZKbdsuf5rK
sMGnQ41CcPzSloWN4kpI4+kS1xMG1MExcqgzdC/8Fc4PrffjrNhZ/iDSD98elpFjq0KGsKzDLAYh
nvRXf/DKikWIYQIBFNNfnKq6omOzjxZvEyTAgsCLJ9f/8F2tLwXQ0jYeIPHItD9Ifu3yuKAOvRcn
9pqstTPg1o4LiO6BI7Z0aUMyPI85do0ien2caJSs9k2aywzh57WFxy2u62ZmIIgRPT6//5BQW7Lw
0m4YsgxGpT1Fsn6vrmJKKGcQde+AZeWmBVW6kEF3XCueiObwYyzhL5FdBFgVMYrpmJaGgR5x/agZ
o24Kbvy0SEyRP1/xkSagA39eQB2IMI/QOFAyFwAe6q0+yxuWVGQ0XGdkYjAaAXgQPuO/D46IUN4D
M6i7VFbNPGamArz+F/7q3J81zeSlJUUOvj2apcPmhrW4/u1hKOkz1kXF2qhlCC2NUjHiA+s0zmcw
7U7CHUjCpu+9TmyTOe1LZHp+GZuRgz/H3QkreNOa0IT/3DRw/r20nIR9pTvjUQUa+Gz40DRJb752
30ME6+6LxWlNFhUorCbn5w9OhU9TBfepvrt89/O0M1To3bQ7H6kSSgTr0Abrr7fmKjNbxKFgR4xv
a6LzXl/kKcqdJNa6+bnUO5eB3VBd3eTTPqxbkflpPaQmQZaHbT+QbKyggoTDU6qAtPduAdVUtGkw
BWfdU6dLClV8whiZxfc0hKaHTyuGureQsQB1z26Kepf9Tndm8YF6369lqCAxaD23pNQ6PIkIp/ui
2seaPZ05/YvVqZXos/Ho9rSG78KQ/bysLNXC/B5WMw0BTFxsXhLPwMAhVl8SwjeUksoFqPrh7Ivs
THJnrs9grPWoikwNreq3GQ5Fts2gKY87r00uObcjOMPJKzj+XvbZP9djFDi+mwIqfdBxzqihN/TU
yLTiiVITZp826CZCjp4rA1NQM+pcu399pCYkF4BH7JqAA9tuNpXbiL6VBv4i35qoIJpVJ/jTaYuv
cVyh6Y1EXjisSGEczRwlFNO5cQcvcYs95E5TRlvgJDrK1s7lbFLYJtNFhpNI3YyPE1aJlobO04MY
S51FB3QsFrVUlKNhyRCmRt0vNIFN+dJUtZX8XplDNhZO6FtXjJr48tf0AlOQBPx9kS+1AZxglPXX
GtK7KSyeXiWxBRTMUBso1Cn6B1s76bWEJGRaakAXACLcokPZb/6LolzXfLuxX63gqnlEAo0/cFfl
DqJaYvYPAzrE9+oRvpPKQySeO0RGTZ4pW5WxVb1OjKa8z3yjJbOe5yWt3FKrJAlXdgovz88/XK/F
S2/hHd/NihoKfD7O80MuYTjAfz1bw/pH/EUSdiLPFQaWpM/WFS7Kp5uD7ysvpMmiaQ4aqbaN93hd
U5lk8fEpffO28F8iwlQfG4omJDeg04r5Qpgt1RChz7gcaM1C1eiIzg3XyofEwsgbzrVIk3CXhcFY
k8tH0uKDuN/S3wiM03AAEty4yv20+9BuCtPyAbaBEWx9ATFJnMaobynfNjiZBhy9gidERqCbNIh8
B9caEj7zl25rmWHzLERPuNU0Kx6BsfeG8pdypNqlnCmwRjbEfAT8CZXQoNNB41hZL4HGHJZTklg6
/dSIDY9fZ1O3XV7c5xLi0JgGKhuJkgCY4byCgJ7wqeaNa3CE/IDjJjCqdnTo9uZQ1n+IsZ+VKL05
446tTM5WSEXG6dFZjCqCqKd3WBzg43Tk8ILDHBwvxDaIFx4cYaliH/dejWarYxHjiKL+kRBa8u2t
mIDgeh666iTG4UTQmobtLm/9oMS2RKPCRw9axZ6fZRGbuVRWcWBBejFD8k9Yxl6AZ8HK7BHe3oO0
c7YW4kSOHootjqBYbElYMLRby8Pc7JqJum7Gv38zK/hRsw8vKxdKFv2pL+rwJpLLlw0oelYJLVb8
njpmwa3iQvIdapxMCar2bNs3oV3wnVT0JAFcwgcV7u2a/jrcM6F/Skok5paoTudcXm1KM90qadBI
Wa40Z6oRg5/wtSHEEgdgoqWH/D5lrIFDOKF0rqKvc3SFq2YR/0+l2TcX9A0twngyPyeDrmxFuzpW
edh2a5BwJOvKuIh/NyIIQVW0WfxWuOjvqASX2Y65TOvbhfubscz1yitsHub+W57XpSCyntld118k
JQYVe90qu9uvB487eOUp32GbrfiFZx8wmZQrZyfaLVzUKQSI6ThKmhFIvgUdvq6MPPUvVU60U1A0
bRj9rujf/I/X5eLZY1Wqkn9BXH2S+HvjWbgxGHuME8a0y6q79N6aT67U9cMGtFoXMZbwHw+1EFop
v1Xt1Bo16B+ixDqhVjXIRdG6Teu3wInPvxOT9HdwKRQu4gI32LdZ3XQ+N6n4vG6Go9E7BOPv3o8a
oE7h30eFE5CUvnX5pR4OMWXWPIOfGS5ekqTsDJeaUCIk4mjfRqM07k3F5GcT0q1lTAnzXA1wfBSZ
fQ7r3zN4NOJps6Uz6VeK2piaQy3MdTGzFZA1NmvVJksKxRTIubXREMAEbUcdEKZhM5PHJsXBeM4X
Y5JmUykUKhBpSmOAuRxI3qdjaiBDxhgd9nazIM0nQByApZeXJww5DKPPwM34ViSZoI377cJkd5PI
zBZJQu+E5fj0DQ7J6hZNiaq6cbv2bZUXZsnD/V1TKEJdRWfAYawIXOKztxfQQ1qrt1rag7kJdVjR
FgUfPul4KN1hWtxugKVivlsgirpB44vAQC/8Nbl5eS8a6ba5TNwwaW1NJN64rn2sE54kRfzDjF7w
iAqQevQbNQYZO0TnfIC34KMPh80v8VoXJtTE8hQ4iV6X5GM9X3FEypvuKG28O/YkOqqVR2bOxs1r
EBRfN7jazNCfjJK/OThK4vQ1rzZ016eB7GI0E2AurqcmTDfuhulL6NFrwUboESJlbu6LY14uWVnb
g/FfLwkTYoz16DpkZx2gullHlrAq2xtyXCbyK0Hp7f2mSvVUlEOUmuyUlvzyVeXF1TngeD4lBQKS
dWtkjUYMjcXDnw3MURqEtfXPbHCtfxKCYBOzVOkDk2FmQ9M914qhzMO7Rf4WTQKDcpVg6enp3XOG
GKXhgWmCbu8duOPtuuLFzG7LTfYkW9gmqt08Q52MGdKw0ngxsN4gOcshtMAr06xG0yWL7UV9YClG
WeotFsgA/sJxxFxVExBvqDJCOmmKsdVRIUMg7g2+q54MuqVqYSCsTJmcf0VUxOr2J2lbU7xTkYLc
xKkgWD99JRtmSQT50vP/42+ijqaFQH1a7jmHSfTR4HdV+k8+yXzv2crNJlV0U+NCGAHQIZ2L5y7D
qqhUgMHBfUO2XNGU11nGxQmIU3XJXTwcTZA+2OMR5GLEMJnyHZgtMroq9qI6RcRRv21Fa/1uRlIP
L4iiq2a94y4meuM35YSoKdAp6YNzHkpw5uL2uuGi0V57Gl/YBzqT0bAxLxOXKD9hB3P/Djza0O7n
dlO9AkaryHynPAoARH3L8Ix8vV4iSCRzVePpTdzBm5k73UsVskdwZj3hiOezPkoTgOaBrDqWOemn
JDZgCsKb4OsjwrhmG+bpGx4/3xJh++qzGWQxYvLOxJVozJTTyXyGzOIUveu2h9tKXRvG8kuXmZ+6
1e/zRVjCS/x8pJAd01TxWvcRSMil6A+c5cQD+naPlVTP53PO7zVzvioCt2J8iHYrf+1xEoKERZr0
N84/ci2h3jX2sjaGDDY/9jiPLmb72WXKWBqG/nZQpQXePhhwgRiSbeMQlzobpQyF1oJ/12DcnHAD
s7mjHI+4HJxLbqPwCGb77jyJ9MOINZ9dXU8FPYSVjCy337BEX6slqPT4GQsL3KbHLJjJKRrFSsPR
+fh/ACPbDCpdqL2v+TD8XRsEl8TGmpStOrpXgvIuWWTquM1K4t+StTJFhxIzPZjwquh+nOFMzCoz
0BaGAl/RkXvcLW5XnVaGmcXWpeW5vKaUGHgHVa/EJy/jH78BhVzH5iG5k/mZN0hV5kkCXu5Cq2Pp
0V+Rc4usGQztaR3PGgrwIJtMhtjzer8BuNSgF9A/XODCfmCvx1a8bbmNpLNO+MEqoTBTKyE/RWZE
B/yRx89plQJH/LIvAkdlnoCgHuKymjWQjZetWuaqabzLl2YXs9Lg5CYsRyYSPH2C8HaN2ZrDVGck
XWURyCX7gd3H4N7GLjwUZLVnCH+GxVnVldP6pJ/jrYVi6C7nRPmW+iCKt27XMfb28LdhKZfx8dD4
1QXlGlS7/nJMjPxohBnnJqafInOkvexpAtY9YlVEyN4br+WMTMNa4DPkZVWzmUcXhDE1zoxWMSQq
7povu9wWc8vujpQuARTgVd5BkFpUJ8ZfvqCtNuqpFupoKmiEIpEw4je969xC3uTTKCtRugcuSLsk
G1Y7i5/NaorBMbJFoyyanQT2EozzDjGaLSHnxp4u/hc+mLcAfm08sTp5GG1oGfuCwRSyw5G/xuhy
VsxD5z7u3r4TU42TikgzicXN7/+a8fJcAZ6yhAgQCD7zfgKWk02HJ3xTQeTsCtD0Q56TNsV7VSzP
lvgW874QA9xQT0ynrGH/hSimuSueJ90iFJycwoZQaA/bkzCa/B4XxluTY9JNMSUYFupF9T3u4paE
4HRYotWn0AL7t+MEHiXPTnfB3P7mxBYFueDc77X71BROT6r4uXt4TnGj+JC24+i60m2Ka7AbDpHN
Mf9HtiYZVJvgU6t85T6wVbyo1pVQeZCxZ3937ExVE7qirOmDcn8PJOjaYlhZxgGlm4lHOnXP7BwO
QSqG0GUs8n/UerCZNXcMg3WOSMegSLhaVVOCytgtsuRUzilkYwaGdHDobBAYsavz6pwIW8p1LbPW
uEMXI4Y/KDGHfWjmGj8/WYZ+H4+R9P0nGjmRjQpVPcWrB0dvtd/R8Ev2V8mj+dx9L4Lhk++M+8MG
wPaILK23mspZdUK6JmorD4J1crPk0iGaILXtw3bo4BLZGg+jIlflbXsLlFOf6+U8tN0ddK39kPgD
5os4cQ84V0OA6qykivDaK/ofyH4u5Jkuu96H0YWN6A4KBUsVTVs7dCRq5PBpvsu06r2AUq7sObdU
xlQ2f4OfvXCLQM5T4tTFQzritPXYuJvRvrx/PkiAP2hTBkRAYe9ehFGsFtufdh5oGr7EI8HInOMr
L0UM0gIlwXVHndurMwfh5jpWSM/PRQ8FPhydBrERNZWIpftCDfkIccYf0iYGDoRRfCxMCgWk+Ddu
Yj8KcqYlXhcnuV0Hvo8RUQmrYNcnDh9Alc3JBDWbYNUHKV/wkrTe/cbMD6VmHut31IVSzONW822d
gglOQymiqnSP9ZLdiUuS6DOxnnmbyrHPxRZ1Q/fvoMGimyePbsuqsyfiOSaTSiyLShX8xbga/g/C
Kc1pOU9rHjFo3ET2cyNq37nVZeCsQEWDpQuZcAMrPhpceomc5jIJU3iu12ngz3EYmxXMQ3dYMk97
Y/Y+tiA8Skyl3g2H5SUPhV9O4IABDEBiHR+gjmpi8Zk209lBy9esFVXvEpua2DSnXZ/5A+LETt+q
9Y4C327DsLLz8KE0zulS9GR8qOQvbBS8aFbMeMb9prrcVE+3CEY6aQS1LUvSvo1xinkxvkfNCFae
cav3rdn1SmX1z6HNFaQjYWsEWuuEdkOpL8t3Nj6i3jXgIC4b00dCJtj+GZcvQfPAiL2FRCeK61yV
7Ua6fE12soG48Mqgu39ejTORzeyitJ00CRQBxr8LNqlJIaN/c5AfzKdJ6z7sBDwntE7EXw2YDEEj
FpgaONgVL2WqJJuyFqjAKZ3eJp0j1ocn7qV1cmAg3LuzhqiJgMTxEPE9TKnPdofN5kz8pIm96Zia
h7OW7JM9ISJWJiU5O8sxG7ArhvHYsqjUKtoczPVpFt6fhb7t8BCJUvtXAryq39GembC0dAvrwmc7
RG1uWDvss6n+aZHf+yZDrPCpwuUeeaWJmOspsslbe1errnX4YzQhTTqslcrctM8+eX30QWmXr+XY
2UeDMg3P4luny0KfzuPta3fKUt7qxAQQkHOg9RgwPqDE26aO4y/+owZNwId/wmj21gPvNJ/WXt2D
tmvNATyL/OUWnzA23lrS2+8HrnMItoPPQvrULGhUfAY4jf1Ly3vk2H0o/gd9WjqqVWabauVWSXNJ
z9w5S1dKYCICuYNtkQW9PkQzEiTcMisSjQVjOXjx7fD4t700hCGW6wqSF3dV+jHDWxTq979P+qjM
vQ3EjvtGYqBqzDHrUmWrynCmH+PGo9hUQxqJjqNmpe2ubAZZu/VXqkTppItAZYfzwOpJ553diEeF
UO5xecLfGzoy91ZOLgOT+nGnTN/vPyk0i+qbHl3kOYA6hR9S3cceXyAGaBfUSH8ssw7gxUV0UbSC
pfuAcw31erc++U/gtnHjxH4Zztnei/+TMtGVbLDA4Vnw9uqmgLDVFO8Er+stckFK4L1cGoUeQ94K
sR7YIf46ByU7eWoXJirX0cXyz8LpdE6QRkkxBuAJXQ6kd2+BKDR5StiJJ1gINSbV7yOYftVVOun5
LNI0Y7pnASgjntukReRcuNAHjOe+ZkY8TjobNqCZhsYmM2jx2b6+SOYC/VZr7i6zqxAf0P2+Yxlx
7HIpIvz2itK1HZKeXs1Z9PrdOvBFFgWVHuH3GjEWJXIFp7qohyVERguQUe2vFjWvRuNQvf/Tq3ZN
gtM2QlLe0B1rhzMc+3T3dVN9G4sdTi8YetiE0I4pTC5NmjdKBdxYf4wrwnr4icXiRk8BcZyhckeU
bgKLW9uEQXdqtylVDuLdY4f/86ssS+Ml6T9JpNHP5Y/coLZJTPnQwQgQJPnEMTL83JbgkOO5MHjH
N2fUp32gqtsPHeFK7lk2CkBRCcc5m1Nrr1RI9LUBQ/dS1jThhFljuIEn05FvZ6gn124VkijdgrIF
4OtXKh3DDfUdqcO6bY5jzCj2bNmSZszc8RFkdTOq3ZDUrigrEx8RYL/YEfEndWFXL6caHrtYIwMP
WIAP0kGzjq1nL7eMGqSdcPvD1OfJ7F6L1h+CwSWOD+RLrJFpvzBS9tDwWNfGrYO+fsVItIqNFAYb
Au0JfswAHgizLMqorsztlKBWfaafkWnETs0zrG7e4FfTreO85e8bXwEb+Cf7Dr2LbpfP2j9eUr/F
ul4S+P93UqOzweqIlwtWrt6PvMjzbMsRLZMIlVpTS5pEPpsLWT5v0rZhA9jRVDaBjrX7N3MAzQ1L
bSNjqQTUbpqYvd/XGob6/eHBivqJmzuVTE63TLX+rDdvHWu9hfOmcaFgbO1W49lymcqjbkC8z4OR
XXOuz0juLqSOXlh++43aVszjnn7oledmfT7W79ALX4QXS3FHge+Ars+eu02xpxxdL2MujVmzz+Cw
jDNypzqRoI5R6W6hUoNjswlrkaP1JOi3VHBfS//F7O1fjplLyDf4cH69pHZhrvWG6iGqWQ3+maG6
7fKmujYt2oWoeq2DLDH2CmQy7UvM5cwsQJiwj/pr/710kkrQ2Twg6oyKKdGzIyKf+MSdL8kDTf0c
TSHEy0PXtHy44JTcfoY1MTC/1N7VGp/pEZQgf2MgYLgdmvGIFUoJmh0sKXXnVQ+o3mI6RMNDmP4Y
QwaA6fxzLqjToON7MUo9o9kInI01Tw3Qdw2jy2joMHdA/Msm157gQLoQSG69i/SbFVwa5y+VVpJi
waC6oQxaIklEL9DLVtgpW61VyM/+xVm1hXOZhGJvU08r/MKsDQBsOedcW0ENuViTa67syG2/5JI2
7xXRh7gGq6+VDtZSSmt64fiu2xt7BSKdcSxRmq9OdpUjec4fVsY+DLbcu3dI6p2YuwzdUmzMGilK
j1vqws8nJkSuBJ3/w/FL3PQMeCPc8JB4QpHZ/shpmAA6VLHtloCSDvni+J2uKs/9CYuFYWW0ugwu
gFD8SIaEuKw5W6Y86H8cHK09PmY0IkpbZDwg1PaVwbgYzQJlAsrEBuW7TVIGV9rvfKdos1DHaDTk
z/fxDUceuAlEBHZTmqMdL5I0248AYNqFKWqhwEVluJL/9eCx8PEXYO8ZClevjwpZgeXCB2aNzEOn
KAlOZ0FQHAGchOs3Hlmn+AkgR7SHZw0sUWWVzWRdtTGeqxua+XMJGwUO/wzbMinQpDHVLNMuioIf
EiCkNtCaVLaPTb8dOH+oGjQiu/YAtZWqEsUu5PM1+yYz4gQzN7j7WpAUb1NzOa4C8uHkgl4RxpPg
d22LYkJw92Z/rBP+g9tTDyRLv2bTz1b3fm/75qDk0cDfq4V341UWQzSYP9ROy3//7jH7jiHadq7O
TgS9fu3mlSovq52TlKGGajBBuZPoeAcsbl9SahYC07GD5/ZfLDGMb3qJxQlHOcn/E2qSI9mP9+re
sKwEQMhufXUooUOem+5iDqgOYGcleNEe/UwOW03hmCantz4CjxIM41DAC3HWSifP9R5EeBDEjWmC
3vhfxESRUNCIwEhN+mOqJEwRlkAJoC/BgxH8ecdeo9hAq8fAix9LomrWkfDSBjd8lyeuMkamv+8G
EY2tGDvIoIDN1pSMPSC4pv5wv13Sp4esSfBFZkWCiGGhqfquripTBTIKxFTOhGg1FDzKbiQiZ0w9
eoUQHwneLqc6McX9kYwSG4men2KRye2vaI78fsBFxjORnsov/tHhiZnIDw3Gd14TcDH7WEpUXIAl
eyPzTKmcItL/iyXgDna2WeWtsV8KGQ5DSRG1mrSvuvxBcvADR73NB/tKPCmvhmSkwwpe6Er93Jqo
Kf+JoaA/CW/g3MWjyfrb3AfhUkMX4OjHMCTc4XNYsat5N0hNNxZyvqmtpKYKocbsXj6IAT+e7f3p
gZsXZ8AqiBl9a5zraueUURkZ5q6dVleizMhRQos92ZJDAhPQUVkOWLqGku5GLs1HJZW0mGtv3UsX
fHh1v1iNx3NQWY8RaBUqUszT/z+KrcvIU1Pjj6NEzLUj/erc2anMfPwxdaEM/cj82EsQMIDm9dHb
obyGru3i1Cczo9jf3QOA8haOulJYid/6W7yB1AXZ8z2iCOsqxv3pNpqotZ0wMyS4rd/18rCU3YRf
ovYsa9P5C3wWx773hsvzSoduif5oh/s6+pGxkIRnB1uNBbMlP2Qi3dqwSeoHQXp/3A7e0f9kJ2qv
igK1tPAd/GtptUXiVLnMG0ejtDTXsr2/mq510aN3SdVCMGnMAj7KNwRuZmMLufeBLIBGh6ZfvtBi
s1iCRoIVY2XHUmlAyIK0JPj+MFZI+9YrF9stOziUoTgLMy/9CUCGbyutWEB5bRp0s1JkoVnf25GV
YMWiDVl5GIpwS1Gw9nTA/sNYMuXY/jfTjU8W6d4VzqzN8iyA3xQXLYwLSsvH4RQB2QKWJQ4xF/Qf
mluiezVBZCPCRpwIz6jzykwBYJj9WxEJoirVxAmQINgmQsUNROPHvNoQkJrFlSGgaypsb2yrDCkP
kC38m3PBHpRIJ6EbCkUd8O502OUX2PHoRVf2WQkLhZPBIH1L89KsLebNkb2NQFzsHubJSHSBqu7h
uQTRuz1DNOyrzdtE0P01TyLE8C2xnwNlrN0tvVDDAylhvIzIT1lSpyDzkd3wvUzbN713j6smO297
kvPviDgR8A3dRVQhHhEOO7ZV2LR2Fv5vOA0tJPbIfMJmFstB1k/MS2YUy3AQrRT6JvfChxmstotS
9/C+Ico7vTvokwxkjdWpgJtJxjPBSNujtUfV0k+rCY9bKTloq8Z+WeqHsJO+Fm/WsP2tvkrOEQL+
14pOMIQk11HIGTB3rFr9hkcRonbiF0ihyYOCzkHb4ebts6LIbvHbNpNz6ZLwhNbulaXR+ZJUW14v
65w1W11HrtAyTupsTOSWwdnmrU8qjY/TkULmzQUcWi7OfjJlGafKsSmkQkptbS0pld8tUMuCbn6q
yH3a7WuM0sQvVryluldrLjAzzsm+YjI5wA3DxuemM/95P0Mc6SjEBg78OL2/yeCC9ExfildfvzGM
deOVj459fJgaKsOldG0lNc6NW12KxRfE4UH2wa+STDY6evuCPPKS6Et3kL7sisYGlRkuOVyrivXH
/WFLYQsutDM6OOtJ7mgl31KQY54U/76HsarYPVzGHPhGo0pdBoGzS6cJuMemC1nw1lF0ycvwLbBc
iQduRQ+pPK6oxvcFzmzDNbT7/qxiMI1Utynu5Hb9xDToHndYC7DkWVvOSopbbq0ivjjnBGO3b++b
T04bQgOElySUcyv4r12MPDgDnvHmdyy9+ChAg7HYI4sy/bVPZsVD1hG00fbNXET2SjSabBkeccOr
ZRTzcwJ6FlFTjwmHPNn2ajg2xUwXy6SsozSrs0vZ3wsWvYihEe4HqPRUDpZAoTFoFHmSKmwO5+oK
xG40tXk/DeegN4o/dJwAbRVV29PKMC7SQ08PY6RLIKlXYNom6kMSJoNlEOJoFcCP2Mg7mJvF2SvB
6n8s5oZR7OI/4ijagVSvJw7zmEMHKlg1jYpoH9Zx19EY05I+pbh0oVTUJnHJMOpWGTAZiEGqz0na
qRwwFm9Ppd9NPznzYv7F5b1VdceJJ1qFoO59jTivZ7R1dJXLxTimLKExb//5w3BlQr3VU/39MYdr
26Mg9dIoZ3tdH9I8XbGqaU4akpbDoPWIanl4h3+tQOEGW9Obkdh1xCRKYJGF3xziKbkfrkhZApkk
BT7zMLiNE86gmscFAOq0X2hjSLXrTGSY/F0XyDGWF6TDVjooxnGnymwjwE+SQvuGojWagdGW1IeP
mEpHRDncX8EArarTtMpaHnnPV7/Wm/QvmvKYKYPaZIYjoAENpSwun02omRf/WSI3osFattQk1/eG
TL534mC37teG9k3026r7+HImVZ/VNRcWRYs9D1mcjRf8sCEjLJV0hnGgvU6h1kOmRxzcGxmOvL4a
cDwRb7eK2gZHxKKm8VwRIzjhlFO06aQV6ZW4fADCpY2EmTMIoqaUZIfffbGZhnZfVUbDbDr4+wYC
iEUnYMJPYLPaqJaWdzXROClHtPBp5wR8U3qv9j4Vibg0nTTk8sAsGnSi6C3WzFaf2Qz9BT5AbEsx
mavwYqE7jx3B1583OlYJIBH19ULJHxkSF2KyXPzw9GaA64ezVF6sNE+Nl2Kr9MASeSJxevAcJDP2
9AaEBPTclRlxTKs9wMEiv0r2bDWhArgbK6JOW8AbFLYkL/LLpchw/rnWw6NH+JCMOi138uUKEUWM
UsQFGVRr9ZcFGY2EHZn+qhRSDnGGZ9dpM8RNEFG3pSHZDCOWYKxCYBVTbUulvfR9LJUA+hjMNnon
WSYnbfLVRyqTWvz+BeZ56/uYAhrI+UKG6FzVlcnPRU0sBP/J7mG8jPGnxrKzSZvlf3FZsDto7H6v
LeFMyOWJDSEuK7ApbKkjyWAVhLdrJQkUqtSUmjUmRvQjQ+SPxHVTvsKHkLf0yO6gMgEedRAdY8RH
pBtWiGBAe35jJCeO06YYB5FhayhjUkpyyUhqWgAcu6SggsbPz/hwAulvjImD56JbAoMM1NTn3RIJ
jePAhVPmlW4V4JKRn6WvLLUAjLytYGXbw29jssDADUgXwiRk6uTlkdB0EHgee19cKDUEd+1cMRIF
0tfNY94yGiZks+kb/OAvRNYUSaDewJKFKC4pEoRfPwpg1y6BSaTnVgBt4hRxFpquHVInxk7FTCKT
14derM7eUv+HZ5NhcaAsYjDCF2i9zP2gUTqYr9oE302ENAhH8Wa8f8CY+Knok7tGdMlBef2Xw+b9
oPDWpJgokrzze5M+jUgTC3kbbpsUDAptLvDWiZZYv3f2ipE1+nreW0AjgNOp492+pTZ7X+praS51
YK6gnsipXJBTgV1I7WS7Hm7KGi/iGcctf6MsL4XMHaO0100jHjkD3oDbfDyaxIdM9HWBRp+Eyc3l
ptexMnQEcy6npZ+mCS44zJ8TTE3Um1FxFpQP3npWIA2oqGFcRacVhrazVDTIetX0xbPm7d9vkizn
X3iZ2UP27A54Sv3WxHkWHNk5XvI32bgIsZZ+95ZLBdlsjEwuS8J3cq+VxsgPuvt4wdbs4NTKMFeY
bBe1rPsuqOZ1syhM3L/lvKDbnxfmCEtAzMaqNo/zK3RO062Ko1Y+AVCd0uUQKKfsQYBN/C5UhzeC
DYvb0HvbBJUYQvb5it0vV9cNcvqYg0/GZi20547Tkv/IyJQidFfWbRZm5kmIoiIcS+46bAEcn/L5
6qg83gq3pSq79aUn67cTrIt0+AJ7GUDr7pYfPUTcltPnyUgDaB3Yr46RTrNk3hqMSvOo1hj/xoIm
bJcSaOeVDJ+UCapNxMxKRZvo1+CtGHqvdN4Pz1nuhZCniyvDWNm0iUdX/g6+A54U8Me89HQjqNHy
PiwWdFw+l8JcvK2P7NBGck3YHeO5mOz5M/dQj2FnOXwiUeof6ISsGxxdANQOtrpToTkbUoXtRRIk
s7m1uJj+DWC8bpian/0QeFDXGlqCl1iDXT0gqZ/MNQVi8Y1hhJogn1h81OxqsCopNNNagVSruKCn
xr7Xsw99zPMhUSky03TLy7I4hMAXZ+pWZPbDkZohH2jKSrNFHWf6prA6cmEtkALORgIRGQavcWAP
X8bJdaY8uopMar9kOUiO7phPpxksrbErjd3r+tudrePA0VHMvBTugbIar1lF8KzeQWrA74RJnJdP
CxUxALlfP8HRHVkLH0l+3tprSZ/Xvn5WvoQKKf0HLvCWrw+N9e9/EHJ5vMOy24VptAeZoeoSCBaN
N9fQJV327rvQsKn+PgAConlLxRouM5P4lby62aG07es6w6CyHqg6JmOxJ6gtVLtMLb60+hkHZcar
RBKPavkds36mHztRpWWg/YyFBIEtKGoZh2/6J1xyQsfh38vARE/KQ9VeaWuaINQ+Pc+uT2s9FDN+
f0UozSks9/0nX4FvN0y9pvTxCVlsN0vRsiFAU6CqQ+uJegdgKj4Fzcse6LeWSKX+i2Ha5L53ifzl
PmsVOwthqn9owjPJ7eBJe/rd3RaWQhm27UN1jwSuN7v8LuMu4wDjae1Am/60oyo2wiLe7+vRGTQ7
np13C/mOrsaZe1Zj9mDLxiSSkZUvxE8qbk7qL1wbfQErvhtNzhaGxPp2gGuXHNqzm49E+UujpQX0
JyKe5u5wudDm5IOONG2QTdqpx17OZX2jxy9zSKhfMhPWB6PzLnjr+KRs2sUfDvphwgmzqN9rbyrR
5hRvuKLNRUykYq8a/6T32YD/PF6E+czhUE0m8xL6ZRHD7ptALSp7Z/66ojrjKvFMVtcF76E13Y9h
NwMrsCacnnip/3EVSjvhug+3EEvaAqytj3tVgu5kcDw1HFkh2p+NVZisXTphm2YFfxM1E8Pbu54z
0UrY3iBPklm7vqi/SvaNegEi8CjzwjLfii56AZGJFJLHugVv6EVHiteGJYheHN3bmGfgZZsPb5nT
Tiz+Qzk6cF+/FBfo2nGVoOjl1+cWFcZ9+AYLE6Suwy/iQ4TiOf1rvG9/ilhJJpa7lWPB5v6EgQ86
nsJOmDfA6NCOW2msxKiFtD2zxk1p98Cg3ZUDBnpQGF5dE/nd2YTfFQzcl3qWiD1vjCRkncPexWi1
AC42w6PEnjZdpHJeAfEvb5KELOaFzZ++/EAZ18r1bxTWMgTUNkRLvXKVrSPfgE7csqS0yZPYkI55
QkeHF4Y7XPYgrnnGfBrPo6fn1d6Nh3bP4H9ERwRcNgFh2a2GI8RiPC3MFuiRvC/Tlib++cuBUmS4
FuphOx2njdEtKMPPp63tXrhxQDLfwQJ1l/7pUSQe+chwzNr+/BX4tmeXaoS24/0dLYOMmZUksMZG
SrEM6ALf1U6lOPJmnCXKq1OBKkkQ5Z5XPceSY1c6OelDwFl1AKlcP0VIApHc4X0qGzcfTtvnEBcZ
R/6dn8eYWvfXE9Zj0YwKDFSlDibQkaKHJT9lm0M/biXB17ni2POgjm9NEn56wi2qM+2DVmImUFnR
Xn7UDZHsqL1AOgHMS1nEOzmq2LNaPQkksTV7BTXNBj9xNFc4IAhr8SaiUxyb1EkgFeG0Av3HJOmP
ahTZuVBpuepWL/UW4iBCeml38zjO+CRgCxrmreKJNeBJOCSnN+jVuh5M78zmDiUdob2gscf9zcKZ
IK9gy4tVnVKSO6UKCRHwasdoxU+FWuRWuQyqdaVoDjLFkBR7yTOlzM6d2Kyuc3rZ4m2J3SC0fbli
ojAksZDWzLs5AS4+dCmt1F0yxelx16SOKA2A2UfJ80rKuKevHJg1H+e4oTPDjT0NCdwL+ETXuk+l
2NZMDVtrJODxnCMmQ08yZ0QIiB/C81b+yJaBV8yRWgL1B+4lNTp6VTs6ZHNUFbJDgTQZ/s/XgNFq
P1ynqIO5+m96ORDtZX07s7UcuDZuaTFpYUHn2TV0QKCHMErI32kjmG1CJHPjGviFgd/ecl/ADj+e
eClPXHgS9u8e0Dp/E0QFVFUj00ol6E0Qot+UoNsP5i6UPvbAJaplOOPImUtdPDECDgGmxdYnSuvY
3DjzGTNO7wgGky0QhkXSTPo+eJw1mg5prJKNpgGjHJMWP2hv+LPI3p1bh2nw2I7Jm+6LMEJBHoir
gcH31zUMoFQgI2pk0SWT8uOYFx21MGfMZH9a2evLrPZA/INZr1t+lbX+KcnSes33eFK/8WNfXFbu
nRsMtbUmHDzH4KZAUuQrr4G+4KeswvrNwpJY1qU4ylbmPx3czDgvA0WBDARNVld+wiPexbRuOfPN
/hVxgaCdiIA+jtp/b6TCvpoa8VJKO837SsrUT1wxECBrfGnxzkkPk3wojxPSK6TNFE1kavAAO3dk
6EAhj6+jlhB3yEVohDWFGmyciyQ2pfMSdz2zixahoe73k85Y+goMjzHCvf8rOJCAFr38SlGue6kJ
QfJ6JsY0Vn+3SOLx2fkSciuaPt5RI+V6ZzIn5d9RvkOZ8elfPo4ebjdwA4PbWaGE8f8o52Dh3jAn
JMw2yfWVSkCa3bX/LjxSvbEMurhRatQFO2SjrptilfSJ7mtgV8Q5aHj3l84dxb0kWw2SEbDOOprA
l0qT5kI+FiobFj5fLKRNtJmjXAldkm6acd+RoiUusNJbhOkiXAYch4Ovuzy0Y5S+UFFAHntunCE5
fXDjhsHbNSq94zB/g5i0ju7/Km76qurVNuAI789K/LKo22zcXU4mXMl4uGvmjepbKcnbNHvMq2x0
zXkL72LF7RJ48ZFndRH2iMR5i4cDoajnnLMRWTWfu/sl8qBaK9XGw2HwLmB7kxxMl8pF9cJYVuDi
+Hidpaq4GJchxSy1KyWScWL8zWS6MIxBxBg0XsK0Gmr8WyWK3V+A/0Nk2JGARzYZQsmB2PZoWGBO
QoP7BnNKMsYDWdWIbWD3F2vK98gy5B+6JZ1SUV4CRs0HSMIDgSKBVlK2erLu+3UUYI/5R9Pb3QT7
qstekfbE0fevfAFyVX4fUYndBE7zEyG//kKWt4COVlvy6Dwm3GmWgmU8cYVsjD8Qe57JSJhG7Vd7
hblFnmKbm/+1DR6x62ewnP40GaUEjOsOGMgR2bR2/CKtKApd9kR96pt2tIP2+A2f/bHpoZ6fuD/N
OB3stP7fGIX4DUMsEMwyNUIFOTJx8lFJ/iDSEOQv6lajXRqff7o5nog13BnR3pboqmkBjVLzzZdx
Njse9xusDzHWdl79LytHdO4XMarFU/7jBb+W9vc4RuQGt0QOfJg18jgfAhRCDXeBrvbL/JIvZyZX
iSREhSxNOXKci5ExFo+6PbEycz5Lms9DaeDkk634eMMWSeC+ulREvCPDD+zaMJn4APkQ+z8QJl2l
3EaS8jf5ramMFdn+7ekKGzX72Rx+3TyqVvRDv2mpEc7kpb+nUM93teBVzJJT7dPkb+YEI39VBoDs
jmFaMPM9w1VjO9nSimQC89TigOPzTV43oWs3JYAZKu/wAoQh0Y3zRAn2jXFlQZcqqwBedquHqP6l
LcfvgXz7ZVOj5lIbDs2AaNBX7aUx696i+78GEe/9gqeL9g4bvQv4RqMew1uN2h27Ee4L2YLHVUQO
reyAF/JQDmQsLfLL+LvYjB/tXn+pEJKG1I2puMuW+HPx46i15xdcKhjRDhy/0PE3KSL3QotoGZPb
k3s4fh2+81/nOn6H9jMCK9f8wCFuUhaJw0aaBtwsvJdOhTgrWTkqYbpvnW5Qoxm2mBX2iMbaATy1
m/ktk4+tj+cMCJlz7+eUmmA53Pexm0WcYBeLSygQk0+UXEXVVSBEmz+4CeAyMSDEgqw5lIHcPZ3Q
iBsuMz4mY/APgPxYUftf464BSCQRzYRNsWgXI8byCglb6YAB8UegHvtSW5OfOGGibTBRZ7BtW75p
ml+cIlb4xj2BCc1L6D1dKx81Y601YjMkjVNvsXgSog0EY7y7ypDS2VajB1e3t4xEUSjdTxrJTwpn
pHM3zIULrp/yEGwmFOsf0yANPx6WP6L/iir2veBfXIbP33Y81s+t0/21VR3CQliHc2wTrrNRQhRs
OqF2TwLyR0nybEXpLtPCTL6KDV0WzoApxievV/asqilNnhIA49+4xX7UvfKpKyWRG2lEDjDQyncB
qZpWV6MiCAsNnXJ6q6MnXZgAeolVT4kqJ5UNio3zV8KPY+0HVTubOJSeJ/NZlhmreV7Qv1UyGRV4
a+b8HuJmIHug8ftucsH21I9w7a1fA7GvmgvwrWuAb0OANL7tGsx8AccEi7RzFE1oQYfipySOml1k
t4wO9+7e8qtX8AIixxsdOrl5c5YnWhGR1mhKPqyMDaf0aR3ziUL53xZXbCA+hNDAk5fimaHOTeAr
BM8s6Lsv/8R5xznHexfV17RYZSpeBZtEm3Q6LcXOG0z5aqBJ6UsrUuKEPeg2Ktscix2jRsOlvMsq
Bag2eis3kHy/VfvaLMxx1EzXxyrovYt3JGbTPM/TQjsOD85JLVXB3fxgc581r9Yz6N8MH7hdyJi8
x3COUBoc55kt6+rNaDzMG00pAXgFpZNl0VrMWrffyVvq8BA6nCL8HOCHjB50/wfZMmG56qlYUsnk
bNICAyN86j/F991eIpyZAYZVB6fRY9b6fbmzOo1e2RZ4JFuQGVZpfbR/BlDd3M3OB97z/wPQsJmt
fgPUH9oRiI6t+79CJf/nZVx+4M/K1zsQ7BZClVgpkvEsGrTyYWkGSAIIHKEAbgzHvhnWs+/5aX5o
QacreYzTKguBIKJYl6JnRQd2j/Z7s2AN8TSixQfCc15FBgjFz6f2oJbpfDswuoiYklid71TtYWFg
BArZhmUxTdU4K+2dDuj16qd+HOFl+w1FuBddCkUNq/1zRDw/OQgm1Alh3g7HEgM8gkNljppm3vGl
YmQUjx8DmUGMJ+ZMOYGYTCGPB/RdvQ4InKv/Vv5i6c1KFWKm/SY/ssMfLzT5tDBADSaNIpSy9tEz
hA5VkcCDWdOQ7upeKkeLUfzZ/r9toNgyr614mF9oC47hB8CWN7bq0UHLp27N6f7D/aY1El+asJFi
h1V99KbzRoWRuAYLS+m/EJCdzYZytcgeYX9A+DZLMnG7fEH7ZEwZQzudfm+mbscUG/y4WFGmu1Cj
QfymlAHr0vefUTZOmveF8bzQLupCAK3zlRMwUoILjLqiTyUwhd9Hijgob8do2AhxGWVr8T/HQmBQ
c7gNe9UyGnORdzcY4d8/GyIiKYoiPQs9qEy27fmKun5tcOgn4DptQjLVQyl2Au4XAFk6n0AkrGzI
Vs/Teiy43cAKMW82UzB6xzsWk0eAYOtVSAA/9CVFfRk/H9yJc80OPZTZhKGyOJlAp4VaWLHI2ib+
1O7hg2vMkQx+EqlED17gWVxtmGQkYCdbAo9/Zg837ePoUO5EQPp3YUFfSjOf/8ZYLVKoKNqKH0mu
6AyEHNRthsHmgcEbwlbHW8jeqDOR6+pZ5J6FdROeBZ+jGV3GHcteMm86fKrnP72E+V8tALxCjtQr
e8lV2lOM88mQSKLhwxYQ+9HwDEscIh4zDFLXT/09mvlqelSIG/WysfCkX2qKtry9fI3HBLmnADQK
foEuCVhiWjJbwl/m0g44OxYXzwPME5jS8/tQUfRqUYY58gSbLNoZX/S0eMX2JyzAP6ktDICUYxs5
WvQuVlBPPqnJNZmbivzHhQZMw8vtKmNJ78IpDP4cVxfo6DyQncWIRYSbat88Y4h102S3Lv5W4tgY
9ZRhIvJ5JJneSv941L8hNIiRLp6fbX+DiDjZam4OXM+nTmIgd7GAkD90FLo4A1AXV+QIdQDQbLQ6
r1du8zZUeA1b+ZPcO5CbxZf/k2e3jbn+y/7v7oz9/WdG9EP9up1fi6k6xuPrGiaft7NaRW3iytcn
LDp7ezgohofWraqlUYN6U5gQxICCHV4sEdnM1ftQueniglp56HQINct9pz1q5e+Ci24kK/IxlnY9
2WjyqOiwgKxAWZwVaOwa3KTbQ+0FX2uP0qo0UUTgbKLwhorwhoc0Oocsx2Cy36tRutNAUK8+nLZd
GVneflz799ExZk+jSypM9OYHMRfZ2AIr77nJAtGOrvRKCVlFEcrHTxbzSFR5jSk9sKipD3xHwp9W
3DlvRjVztcxi95tQLZwdbbJGO74w1YZ8NfcQkRCaKfC6Yhj2PeNP3wTNLseua6D39061Wi7Ig4mX
iv6cKXnCkqjlapI3/k8kHiWd3H7juEgzXvk2KTFh98RFHiS4J/3W58UKw6qwomP+zDYWyzcRn4KH
4E1PJWVh7SlxM8MTnyhPjJ4I/0EhDBa9aoF5PAMQHB0F4IynoTLJYtwjBP5xK2Q71yEBA06+ZEmj
RAez5jfxh68IR5GUjmKBFlKTXU+Sd+3+Ok/ewgTJzo4uw1pxdTUGEfM0BAkX4aPoAH7d7WyyPDst
IDnUifmcAwpH7XDiMoUa2poXe8d6tvD+1wO5qFK4+1GMSWhkWLzRkE/n1Y596Iiu2fjhegkAi0Z9
IlmZ/GpFdgxBs+Mz/ZIvUPfzK/8bUVQVzw4NfErFPSy/9ZBVgPUPsb7ceFvG7KB0txO7l2pCN3/l
4vNVN/jHCrrM2Z9PBTNOsNB+RenSj/ZrsgbXcGbwESLnoZ77n0EwDqiSSx2vKGmvQHiUdrO7NZsk
XqBBHHF/RNbjUQ5Yzx3DHN+lWoxXjfARNLqkRTU7P8iuIAR772wpDJHe8nsoE1QfckTCW3JMtN+F
YkmhpYABhvJPx/aShKgxwlSPID7B/dVyy7A8jwURafRJj+9LX99t+2MjxHcYvW6c8uZQ4XwmekSe
19D3t7z7ZvteExb3I24zar0toWRxFE9Nh63xd+Wn8o7VaX123y5cxE+NvX887ChA7NoiZXps4W4U
j0KExpfhD3LCuhE6f7WHU05lGlcCsUVg+SBm0hs1Nc93gvDZUpnj5qBPt2xS6QQKbqvTx9kGos/F
p8A2OXK+VjBw6oDTc+CR7SDKMvtBb5NGZeKiw5tT4KD4GKuQZcv6JP82WRT+vzaliZgzvF2nLYjr
Q6BkizKwNC/E1d4TKAYi1CkRqfkDzVWvW/HcG+ILBlvKGfEk9CdFKsNBW0AjZH8OAyseUOLUj64g
P9tgzTa8e2ugMrMQnFh6JFwqEpoD+M/8OI4gl3Mtt+aoSX8sE3wl5RRx1j4+fKGxzuLGM1vl3HFl
IYGzpwvZLDmbiamdBsle07udT8/cEoDSCX4FUtpqGuJYkbPNk5va9gBtOlL5dEdje6PxMs08F9o7
4oLT7UHtztEtn7g5zkWNZvjyXR/M8aw/LKb20LeDuFZPp5oKpwxXZBGge0RDWx4Fnm/S3iawPMmV
uQUJebzPQzKxIg6f5ZuhqlSLj2sU0PDEDuqS2wlvVJJLlLG8ljxNYQFMb48lyrraiZsTK3mLGMKx
1Te2OFsPtlbTz2TrqxI19j9pVjlh/VGM51HcLZ8X2LOzsKuvKTDotDO4YwVpjYSc8j5UXZrfuCHE
JYS6q69WaQ2kDv3ArPeeEEKecu2OGNVxZWJYS89Q7YCq5MHkAk5QnDcsCsphPTUXx5S/SAerB0LW
UDv58KMEvlTyoU6FpknSW2qsdUWb1Qq+VxNXpHnaj0G7JuyYsqWgdsJ5pd25xIqiiYeAIwuTod9i
lwJHpQdLfozFta0s1hsQ9YOZESXetnywAVsWTeTzLymj/sEzzByWfPRW2pHo6nFGTieaLcaiMmz/
zWzmFclTrEh6AocIlNPRRrg3PP46lzM4hJPGFgFh2wIHMGcnJFLLirdRC847nQD0+ZbiSX1ozO2c
2l+M8SV5JNmWBGo2JOnCChfBi4J8I40eKGAqCxDkrjAZByQLneAltljTY2S9ziuJGlzsjOwuihs4
/oIZ++0me188mJRRadfA27TjP5oTqUk4xvMupm68wkhzXAn9cHtPTBdHLcaxlMh7M3TMSDvx0ia5
aBPHsI3eKNeYIeMudWKgxwMSWL8M/+FGBoLCPiOJJoiVa7q6fJ5JsOXsCnQ81rLlaFN5qhCYHhRe
nxHvSVTtanHl4IUG+f/5gXfPhegN073JA8yirHqoMXiqDeqiI6CUUq4ZGws+xknMky/0xLEKHc1i
yBKYQo6uYpRsM9v8x+MHQUQNwBpI844GoqqKaJ35DlqyLa7pVnjKLTfIYkv8duTSFlzvcKGGsvnV
LF87OFbGzLJjGIDF7GijXCtEW+tC131epC8CueA2KR91OhQqXhWh1YKC9BjyCmIaVDdduQAgZ9e1
ADlr/KYT4GYPjh0TBK3G+zc2nRuSO8H34FdF0Q5y7CzWhZCiD5P19+dBtX+g6Ut4VjFMrsyaDgoW
AI381DHJJxjGtWyKgf5+gsJ23D6seDa8KlycxsFuHWX6UvUFh/dbEAPVw4XZ1pHr+R3yN28A4wYM
kP/9+DUsw53n4qiCpMzlFgKGq8hEqg8IUl5L5WGov3uOWvI98ooG/FNIt9yiVAQwCjTmGUWukFga
Ulw5H4+eOXNjLDfBQGrK/F3msY6QeBDY/Qdpyof2vayqReqAaD/dWTJ8vfddOwvMJ466X4tegkJI
qB2KA65Fm1OdfvbbdgCll8KisKGmgW9vPJ7dD6s/d/I15cQ60u4f3f09dkxzbKLCIhqHgyxw5VA1
XB8qNvQMLZyKvR8WAwazhTMRzb99wcS3pMxTWyOpHLBDmzmHog7TtWE7L3oyRUww8G8DdPPqz9h+
5J45nxNy759LeZD8ZMcADyl04viZ6UlMI9DrdoHfY7LPEOknSiOi+LA4jLDNCsOfs7o8QuoFqX7E
7RGXOEpAFBtVHmZM1DPlwbezVQDaoKV3wWbevsuRX19wNq4lqeDcKELMR7atA5w/ofblz+k8EKOV
L7nSHSiK4AS9kkObwdwlRtJQzjDz4FdWGy1F8Ck1OAqF7J6/lQmK1o2UUiUz5XEB8T8cqhaXq6nh
ZdWT3L1Gl2dtnitP2oUTIL1yWM1tjUcrjMR8nAnUMbMEn0YnjDzOD9EY5JuivMyhFVaFtFBH+ob6
PFzzFpTMjenfJXYAPN9PQ9IlX+FgqEJzxy8WoAEf+sRhBQdBqsEvEbMCvE3ZBkaD/GoLyNAR4J8o
VO6Wuz0HTv5m7unTWihrK7l1VHrgWu4iBaRAu3Zl8u1dVAnOoUTMlKb7E/Xtymu8qfsxUAq4NZeE
0o6uHT9Jv923uwusXlIYZrzG/AxhXiNzU33e48Waruj8WCad6oLQAjdioZdhWOQXXx/nGeYlvc3R
OYF/r8gctec9pzlTcugd68hxVpujoKJH8OtbSTc+4Bl4u+Tyts9/nBwTszyZFSRZKaq913SUJL7C
cZvsCu/sF01u5X3WFnUgS6CVJcjPGIxzieR7bTvx5clbbzdzCJw2Iud3St8v2mH3+y7gLDScFtsp
PfJBiZFVdtHkmPRf1mU1Mqu5Nw9M5BvkTF3X73FGOhK0OveAwTHTKGZr0noSZStvrAKfw4UanS2A
YZHDkrO6YuXhzNQEe9vyrYN7lefghG+lGqtFZMJDjOoboN/707BOtoAojhq8jRX+ya3msiS4jhA8
CJtewMrXKFFX/91FklY4FOk1O32sp5CRoXn3rumFtIRAfynklQTDkVH+TMoMadvFM/g0pSDCpiGp
lrqD77oOyc+tCogWi0sjMezZSZIIJNiHpf1DlulIQrL7dPWrrUA8cVXOfBqCmtUx3YqjgDiDpQEP
USf/cb7PHZ7J3Rdleicq5cv2tO1g+yuu/sCGK6uSIFgh6v4uooNYcbchb2QcDaDVgSqCIxvEQhN6
U0XNrxGM3kS9TBVaLO/cfv+C6lyKsNKUMwZCyTYA+t/xksGYTDgVxp80ogfkrHaXxvNTYdhwEGY+
1uu7zloITfxkAicJWoLA4PQGNVYNk57kq/HS/LEXH68r4ptglxW6UFhVktU1ccmRikmcLm/8Q8zi
FSbwV6Aqtg1NhSLHNtcg+VXInrISNYrY9ti2GdQZhb+6z5bSDsCQmPK6RM4wxkde2MX73wNdO5tI
TwAEN4X9imVm5BywQVlPdMC80992PKR3LpmeKvxYDjAzHoXrSp8SirwxcmTXPfkB38rh1YRn6dW1
af7D+fPDaKQqYqtmrVuibr131FSDWClNv31vqaduViTXFvNZtlhiEI1O+PChifc26ux0IUBqv0lE
20xsSoO7jIjhf6RI1P7aMDPhR5538dx1z2U6J4CCM0SRAHfCCQB+LIcBkt7JCzNAx+pkB3lC58fk
yZ5z0gDQKi/yO9lK/3WRS4OYq+zNB1HgZYVgic3ODz3txADoSKe4VzuRurQaSln22PP5SnL9BYo5
9dVZ+E9h8cOrG39rZNi96bijIjnWaReGg9F85iOe3VFd17YI+NavP1OZ67UI5fbiniOcsoNQ7YhG
9YkpNQHq0+qSDZBJFSCEt8CZUJSoQbvkQTgOedrFb00CBs9Ufgh+FzaRMHYjXYsemGaLVzCBr62E
0rUpT8xyWDtf3aVWSzKjytjAiVHVwu/Nv06bGvu9JFZn98uxt394dU+U/kSZ3bWb4ISZRt6r09q3
dfBlt6+RN8mQ8YjMzpC1VDfwaGgnjzimvdQoHK4V7wnXvaLGaeHbgR5zW10A6sa9+o9Z1G/AYg8V
xjy1RYIeu9vE1+GmFsR1dr/yTYnrn1iRdTMuwG5mczQpoFWMlnCdht5yVNGsHphi6gZGZW1rBHpu
Y2MWjE1qYsa3gtWvVb6fvOgD8j3/xi/MQtYlZBLBRzfLlh0ferCMXow8NKk53DCBhbMIkwhcVEAj
CAyr0tc0mHJvz6VeIntZtiwexsdAmQaU+h3+MrYDYV/okTe4BbaYRzed4DKWztmOwDXlhzU5aEYp
bRRVlEpfyBc0y/i7f3eoEI8FDXLIqARG6vbuUvKjl9s9tUst4v0YX24MOyquQfKl+jkGUayhJ7oT
q2cZn2iDXZ+foac/GbNgYZXn4iootMDRZN15Vt50LJnp2YISzWQWro2qmi9PU+ehiL+aXfcY3F8e
CE63sBOEUyjr1n23WJUwDfU5CwyOOS6hxKlASHqjbyj6wLBY3SVDm6xr8ovVbshWuwQoTNBKS8eX
PnXKTpgqJhtFqdcDP1wFmSmxgrJakpf6dtXhToxPP0hq8+aTz6wsFyMebL89rz5FMDIpsHsLm2+T
icLZEeXW+fWsGEbRjvCqWirjySkqkTgPaqAJjOn9rFTK5/krQC606hJeMsnfTFj0LMCneHuQPFRQ
5wW/YGf4LcMuhVDjdcGTlI0npkwJ1GaLlY8btvra5CCUdd9P9MBxBHptaTWPw6pQrvTqTIg5M1Uz
e79eMYJI+1j/53NSnVcVIk+Sg8deQkRLxvqWoMpVPDjDZdICPhcl3Syx0ajNsyg8s9zKxnBGcecP
uYkUNHkd3eo12ceKcUjhhQ6yOMrOOQ9S8sAwinOTO0VoKa+JmWWxTA0Hj91PUa+WFXiqwHuy5W3t
z/FOuFUstpINuddl0LMQyHSvLVsmv93eAG+GaQ1yy+Lr3jvnILl4IOGdqtssSMSj/dVyw3Wmkaam
lpkPNEM9/LLyIKXECOqSaCyGSAOLilxYKiaJ7Yswzxe6pYEx8KMLBNCdndUd8dQow2nPHxKMwZd1
/guJKO6ID0GYUHsbc09WUij0mPSppBjPhvUR5drlOVXO3cD9Qzv8zMBs5EcyqW6DYAOEhK6Sf3CC
fweS6J3yuDTy4mN1gjDT4pQI8p6bWa5/DSeDn4/uJVALpW90WXXTqdOxY/7AybB0vGliyGdCdzMM
a2kRkHyawTOhp/kfE9iQzitQYh+MWJ5K9k6QGDE/gDcuKPDyyLD4AEbsiggFdP2oR6DixZdG5PTT
MqLnTzGxUf8ar26Ioh9abzQt6/T1mXmP4Omr0vfC6gEpGMlRVW101oZ4e4H+t5QxZNn6vuILj5Xm
sPrkhSnqbTgdmxi582ePtwb9IKLoIxhWLHLBgFxTO7lFyJCXx+yqxH10ohygOXKu71GdcFQH6Jg0
jmg/3dyLPlkDpPUMeVfu9c1ltWIuQfngEHwodVTO1ZIJw+D/oq586WE17U//wPBYT1FIwPz1CrP3
BSKUFMkeBSrdwFxgKPNPSvD6AJSWOPkWBHkJdD/JSdl8ZohfFITgb49rGz0D+I0pBifr2UjwyjHm
F7EtD6lWqHgrMrVaodLEa+8EMNjcpmWIumeesd1E/frJI93zyXqx+sZQwvRQjDz6pYCVys6VDmFs
1jqzSNQQ+YdHfQUk2yrgtTLpIi/sKjm4HqybCirFWwmB8I6p2l1HqmdRoXwwwsHPZB2ctjFXrO02
QGl/mYgRdakwu2EFbd8TdVjvFFumD75ym1ikuVgIt30nAytjsV9ZzvRdmSArGD1X8dvLsyNWQWWx
uaSk9A1PQJNovxpDvXRbsUMfH14LsvSnZsiaDSylOJD3llsDHhXQ+YrIYN4po2YV75Z4HaquN8IL
1oxV3PpQsFh9W3QJaJndcCry7e5X3y+zetgrptNX9H31w1Fg42sT/njdPiDcV+Iz1aysfIIBzwnM
SasURiWQFobzFRqDt4xMl/xwXVDHWZL9KmgbXjZoQ00CILSTZ54B8ePgSuOhC5FTnjcmvmMFlwT/
ENy0pnEL5wpqDAZ+bmXPducncw+86konRtMC+3jCeQHqU/CD08I7zxlb0CReEY2PMW33/IL3GNnn
5NKGi5VO8Tkw090sA/G3swTDLzLOJFsQxa4qePRgR62+nZ+cYUik6Z3ni3m9sZZyKWjeqLxRwQmQ
nn3h1BEJPn7CKTkvAqe57gI7w+Fg1xCVc8LJ8sxDl9ZUWERipbd9O7P5hpFNCXKvvkLME+A0h7rC
42FM+Zg7ibinvGAH7WljpdJDsOR/zRigViHuf4nAVTPFRLwfwsj+Mg7iTj7TnTxX4uDKXurJYLql
87amsqdmJhufSGKVGCrrJojyqb+alZOVJpw072nF8SL9CdWQw3iw8t3J4uxh85v4RYhq8S/Pc4Ep
MwGY8OHpwnEUMIGeT5htt+/tCLINjtg1UOCxzsezqMuyISc3goCEs5oZFXZrbPRrfhhrmXl8hS1k
padJ2z2Rz3qNM1Eo0nMSa3qBQr5QwKll9CFvY+z/WE5N/lM2s9ZIGz+PUiwmq8VkSCiaPqzRoQh5
ItXs9XfotHPaBLZ4Qk/ByZZPfJyzGOaqoGXTvx2BUai1HFJqcwNP8E7+o8ddnyFMsSnPH9ppqU7y
Zu9Gqggzm6YTNoSwaLPkUFe3ix3evf2eo0dR2ItNK1Ty+KytW+PKECXzbM9NSjsS0tnhUJiT8MYL
PJIMY7NG0fF2qae3UkdETcbLVAYzDfWbAh7XkleCQU1sP0jlBCoap/f29IijzPVeRUM4JrDXKRzP
F8q4er/6Lis9D8o1G/Xug3Yw5whDy43Stbyugw6VoWCgvIl4p7M4SGo3QC+70zjfozerteiX042B
PyoY7fIoYsuexeIn8EQQtZLk3MrawsIlXQtI4tnLT+t8B7ICVTgShGp9bsCyl2GiWLfb6iFuoBYk
sm9mau4Kf/zJ+eEz81s7nMCPD9lVAAj6GoePvH5iy5aguTzKx9pvHoikXWqzzCqzr1ECO1wH5ZdH
rP0b2IDihQOTNj6FhCfizs8sfU1uDjUgzT/PuPWJwU4qp50WH9xOM3r11CqSFeOdP16RJnFDlzHk
cTjJevVfpjzsmERmhAWo4j6WqPbh0VwFyXeePZe8SYq03JOXOwvvLQin+L6fJ6+gawI9GK+7wVdG
Y8vYLO2VklrerAJcdLWpTSoWpLZl7nT8RAkYUFepg5Ld6OtCvOY9vuo5fGhMn7/6GUz7ulV0lDf5
Tuo9TjmjY/vL6IOD15MQVLIm4ltfBj1+kAW99yZiCNrjtiQTRAN4c6ekoqD2qPrnwTdS7ZWfIC93
s+P16+FV8UoUFormL0Gt5vY5suOJ/3EqJBu6F+mfMyhNNt+LBeS5QhCgeOmLgLrC3ZLNNxcS7kJF
inQoYvNDcUFn3w2nMEh7TGHqSFpV4vUKDZjRG9TuK8KiCk2aOywEQKWhXAreEmzqXn2UFGI96AdY
Qq8giW+zy8M85xtXgYtaAWYgizsCFYPBmdqngfKeIVEn1ZnhOuaBDtV9kJjifWSowGdXyhaPSCEd
5elGm8tlHlQuA+i9MYS3TrweHf1cOkLULqv8zXu8jBDofLY8aWjtxONdEfR7boooYYjN+cXxB3EX
WVcPSGA/yDYLWCE07uN1M4aPM7njBWr3mdR8JWQWGf3/z/Glb2GIxf1rzqm3/ozBrhPB4hpK1dve
VZCc5Xy+1kiALGy4qANCKlH4xH6E6XuhSLsXXeuEV/78g7c68qRIFdNrtm8K5q9MrXbIemTQyWim
roWR5JrsSJ0ADugjCO8zcn3XacHeBscY5oTup0nMzGd+8KJTGLDadQHUXzdgIlYdSoAhgXr5ZsYn
Udc1KL9omNSoS9W83A6rlD9g3ElifOF54ENqr31RLZHZuWYeoHtp19tMaCUnu8r2l91Pqg+pk97j
uRft6PIaloiY2L/LX+XUVDcMeDonADDOGcV8AiX07f4cIZy4ymzlkhB/CQYngGu6lpFyAEbnOu2/
5+gi4ky15Z+18PKNw2G3K8VZUdSjDS/EFDvfTJFBpYL4R9JkLs5tEHhtmgPTSFeABh8vshuDiLGg
8RS3HkFUlZZfjiBFWCbDqVRAKirQQ3J5Gxqp/pLLWx+lGkeAkngVjRa3+ETAd2RiCfilM557uSh1
tqIIBFDYI6AZrXS4V5xFok79OCqs1HTdhDCExPEXZcmbj3P7CsnT7T+1YjJtx1cnzf//X2TnFyvJ
oDT4FBQmJYpjfb+RVXgF217tw+j7tARAJTpiyRsh8XqEo3CEG3jbUc0lgb+jjTG2a+FBDi4R5ytY
D0dLPbYjKNn6KpWKp2kZWGoTw45Ax9Gmr0mA7obHJhOahHPEvfYDv5iq9qOCY+ZPY2Bcz/aRrU3Z
5UjeHNBngRPh4yb0P3uOup/fSRSVhfyFb1npWP68iiAgTvp0+2uABr03pC+kBPaEvpoBXJ/R0+wT
owQbGPY9eitgHKXTR8CN6TRb5dcZgEnMMSRZl79Dn+kxuY2GPxYo480hYoa7TyDpS/ta1N4Siwbj
20vfCjYaUSmuCvZHKq5Mo12yzqsNxm12Lmr/cxwYaSh6kk/VJSXyDbHVUNHE5ZSFTlDbbXpkGu6W
zLVnp0q31BGLRblcvdDcfULUDiAiFNBRZrzG28AIo+LOjE1y3euvWcQ/w1214pSkEMgl5mTZg7sm
A7W7Wqv85tdB9nvvXYtfzQo/OxkSAgZqbmZ2O4lGZMNbcbRFslJyAiAR33+XgauY57vzo9IQjIPo
/XRPyVL0q8fADvCbjxRMpUkJWWMEVv/fHRzyBKxX1O11x3evBnlt9EWfjJLknM+Ii6BOEb5OJrbs
eDuv01HYcnY2MuDW9CoVojHEKKGY6qz8tzYBHPjxtioJ4rO2XxX5DKnQ8Cshqw8kNTNHIR2pqz+K
QQ1ToRhajlDqgtJUgMN62DmetSxTTTocXo7r08fK47DP1kL6MGwF/tf+1rrWvSwbjIN8Mj3fAxdd
5CqMC8ToX9QXq7I+eiigIJfZc1C1jEPcipVdaQkV+uA++BrlcXS94khkuMDksgATRWYAtmepUAYw
Bk5+jq3ThMj1aCrhaMg0+haIcrb9uFaI4SjI6ANYwK4an/Sg9PWJMJ4h3/rZTb7nkaucp59MHwyh
c14JqW/54yOaGAVyt7yVG6uA8MoFtYl6ggXKKe7D4fpcwyf6lYtLHjwHBzzQ7zHmDMumw9tG6HTO
mYS19iZ/7MNmUNUfxKXpuzKtHEg6HvCm2oajhNyMrdx5u/Ivx6limPPgCmXAIFg0yKqXmnsbN1rh
+XPSoGVckE/Ze6y7sDsTnw0QQ9IEcdRKuXgr1gDVVvAsKqvr35oD8Rix6JPj7tQtaV7Pc+V2TNRd
DECIMcs/EerSyTHOe2Jc1/L+2u+mhgIjKBf/vcOyiSxko7QqvCWdsCJsSeW/Hl/PB6jQ6j7vzaRR
I6O9VFnLVse4Nf2yzRa/TM3WWGnFyEb6Wa86j3tXxDOsMzkQF7SQs+MrzrlO0RR6n2gJJULidkbD
xqjSg0uFJvCq4Tz6VDpjRzEPjz8IH9pTr2QdtwXjKgv3F2oamQy7BoVUhhtupQwVUf/Osq+VB6PH
Lvp33Cz010i/VhN7uJUKPgseC4AGCOzFQrccpoXJuBkIwKq+ThQDhdYcczJySKoElU75EikF+Xjo
PLAqH0IEQw6DF+VujmRCeLwIonm56w9OJ3BT72PCnCp47QgDYSUtKcynb8xW/WySDp4AVuhFl8hZ
BJCVTrswKXFGiUSADvCogwcSE7OHx0TANe5bb60BG/S4Nl0ZPechl40zUOORr2u3zkRpEcCyIREO
uvS6EeOO85zuHBuBODNTcvWJAA3mL6+1uHYDLNue0WEqCg2UmJJ5G/qkXnP4BTYX3Dwy1f2mZgQf
KlDwgvwhh00R8qaDag3srHrYBqbuK9uhIuncRO2WgdwofkUDrwEcIR4zgiz1Xer8FKXOMSVRQAvo
j5MQUdkPxfZFYs+vxAEF7dmGD9PQuXHsn5JwJ5q/b90ZuunVfbYW0AiiNDdA8rpRHoAqviMiZr5l
smdGRe8xTI4qsQqhvLk0tEQ6SWbGvaw2UPSNNTDDcHVpvCIPt5dqLP4uZ6O8dI6Zdjp96F2apgst
mu76Vqx6q6lVFVBJr5wcXzTukzHpsnZqEd2HHv6ZLu9kxz3jjFRBkQw8hFSzwOtvV3QbEX4zFhMi
Y+BCaO9lHoAYUx7am2xCO6ywMmH+ML3QaKqCVPeEqgkXRjT/kxN+R4540SbmQKE9bz0mV5MVtlc6
vFPuCHBwpNXNvFmPVctL8TAVLSzmC5lZG/HLhO2neGyq7ZPG19+2qBiPrKTe8Ch+UHmGMoJORAzY
n1gAOjiGxV1rTPi67RJ2HXKRdSylbFQnO8sDKnLitZ77iilsIK3h7fxlFTQnlpWaIjdBCJ4FKVkG
M0+z+eflAM/EiH7gZWmt9U85d7T284wVqms0o8dP4Y2YpofbYolAH0U46bgu1TWzM2jPxbyLAcjo
NZ+S6tTvmSGs57RE/jJzcN4WemfDSX7wUPCp1zIuhQ+rNYSFG2XEtieDRxwkmNGxyD4whyPHkBTH
AntSdnLzZDGVSD9DTUaJWkfj540/JxReMel+oZ0ZqqLEHi4vyIaATegQkQVd+HUh+2fkBMpVv958
z6VdyuQScr+1MojCEISpHN+eQULdk/8nFg5ZWx8x/0QU5wa/Jd+RH7o8WcPwpaYvv4HN/49D/heW
QezbTHqhxDgACvE/XzMH1kwPwcqXAxSuYbEKvilC0Hmczsvb+T5EbG+bJ6NtZDo99oMiHsF+Mkti
8JU0/2/iYj3tuaSHIDwBDJIJv0POPO8i0okHuaKWmzc0xZCs7DAavHtNGbEKoSLlkvKh/ZmlvGJH
8SKx9WMoBRDyViZ6v8Ihbjf6pEKwEyMi3Kal31990g/cGcMInd6QoUX/Vdeq4biCWs471SUMQ3iT
Sp2hCjIMHCPn+si+KJprhnE7AWP+M3J765Ukv77U0Xq+dwgPgQ55Vc2FTpQ94iOMv58Lm8xb9IX7
xMlbukiyhckrn9MbEuEBJvIgkNx8RHvRSI5hJ3TSVjOV3pqnuhcMkWfVOxgkTczcimHJTm5JM5HI
qXf1mspEeLky3mX5oMuZzb5rCBxYQG3JlHEKzhs/09EzTVKM3i3OXXHxFHquA5NOFz48GKhDj0JT
KAmCSJwBLFGk6UAksigTd4Gt/WRdoxHqaf1CrZnVOwK73rH1CiLYi808vzkOEv0sHylwCX5Yc1Ba
4PKm1kpBG2qY3egZaM9WNocxUr7NERhKchXeGjH8v3XSkMpGgN9IrZuSuH7rScH+BOAWhsg7EQ7G
9lXmTndYVKMJuTUGkVN/IMmjBhVEHhwhyre7wdPm46sWARhHPAUcnONCHzUHlBhcmerYu8U/yntq
xfwH7bsDVvKNGeewMBNSu40cZypGmCYtHay8mlakVHbCyy4xtiUwJk4Hxb12Svxahxz++PBOB1DW
fcxX+8mcgSbZH9DV6VFYbqqO1VA8VieUnu8Uly/fC6kpcTSGnFzSdy6C0ssPAa5n5Xy5kJltXxzX
a7F0sQW7xZ7GBsejHY7NWDh2GkXpasP53ZUbBc/SP+qxnVpJWbJTz99egI4Bascu8Hh6zIT0ZuuU
uJzpTWqZ0bfScHOUGdpUwEwzFnOXn9lpVxRtsZm9mgfIZ6CGRIMoqXHs0XPz3FAouLMU5osmGkFe
l24T6siRtoCoVcY8PGpi7jcismoRPy6qvUq4PAP2rCkV86DsmVyy7hyGDEw5WqrE9ysEhbxK9Rcg
88Zdn6zv9l8/TgnXh0Ia9YOTmTPeSnuZsLWX7sNarb1VBRiCberlpHEy1oVJ3+1unIx1HPnXT8O1
6rtlYOoIDMwPlUlhMI0B76tZ89lvj9VH+rnwm2lr4ELk586dHXjEIBZhUYNxVA0FWpNwPxDCs2lW
eW2d8a680O/z8Nu48BAmyTfqFqnsQdcz2Ug+DCI7A99tiKIId9d3aLz/kFhUW96h98RPoyP/JFMn
inr+Btj/5MbF/WTaM8xHpH+Fm8VmMg95Y5YnK+73bIee+LpZAvGMXJ01F8fxKPTQaBwFXzdVGfVE
87lVJWx+kEKy8G2A1Rf7TZFp5GTm+A4PFuiVJrgnw3yq8xHVSdLvDnmbJLymQuY2xH+x/1BmYaA0
VsT4CAI+YOEGSR1yoItPeJjTV3f8HHAnVlBeHJyjaPOM+syL4Mi+4Cxa7hP8ba4+NgJdUDsdm/lz
gv9ZmWa5ZA7Gm3id7++jD0+xRepr1YEsqtYRF+hluL01wLWHAVOt7DeNqQT7h2XHDLSw2qcVDFX5
xbTI4ChEOnpjNLVRXmL6aLeTjLF+mwK5MiASa+ZrPbe3w2lzzf1Ad8YRyr9jnj2QH3Ot0DzLzLQi
pcmMncyLkYH6groy+ek32vojxqSDhbbSTeSzWcL1vwLr20c8D/9auGiu6erwQL9t38PuLNb6qVUJ
Tts5iV1guW3r7SHS71aHn4rq0zQDHWY/Qgu3DXdclrUepAWG7MFSynjvE7iU73ATPIgSiHRK2LsV
1cCNyLv8EqHc2w8a7Pd4aod0s4rBtKL9FwBFkIdrXJKflkIRZ8G8iLxBf+DgAZGLcmZAmdBM/l2h
kqXpHtIH0cf8/ZhpsR1OOE89UCIQiX9wP02Rg8Wlc8QG2pukP4ydOImH3+0Y+vwBkXZXdeRZUGp5
N+0UZdYlX6ggUiHabY6UdhGhob4kaARSGT5lbgVNvqYxjJEPWs07nJG211toOTbF36GNWhDDI1of
Tjv16VOxO7DrmoWigO1Vs8+j1muENoPMovL5I+3fUIaaN4ofWh+X5CyBtfrwFRnJ6CliWHVgtL5c
/5mtvJk8/lpuLHqiNlmtBT5q7RhfsDH0y4+4d+qNFtG+BsUXZUexbCJam7TFlyauUoOYJr8ybwRo
KhyCKYo+/R45S7qgiIyhoX73r8KMNGXVSNRK4/N27gJvv6UYFU8Nvv+3z44raSA0N6QSRtgIQTyq
x7yN/wLdIPnuItro9SQ8ImW3oo+PC+PNyOYh01cpJw942rT4HXM498frMScRXnqKnS/9ti7cMFxJ
7ShAWlUIokZBuZsHghEAQA601vGNGvhsQl28gBRlWfLO/rQa/2HSDcfCttuqvxDx0I2b5Twk5dYK
xwWfkpMncaLUsty3A/S99WVviQi0u5zG+BhF9DrzsAxQ1w8vuhQDswWykTYe2uqkUclH+bpOmCQe
0r7CtGaEsbJOvf0bCQ7rhcXDRbeILHTgmLOJtvu4Tepa4dWznauMtWQ1VEKrIktko0kjv17YEZxe
goMrkerTCrUQfROEqw4lHNgrtFlMCO7dxS1I9QM+yFkcoSZmdVmEFXxcw5qIk7uDmvuD3f4009vh
dO1BZsiVYiLx0eEm4/Mx1PGgOYx8KjlJ56Btv0V7JN1oBi2x/1qtP0qQuP5+/diNdIy8GTEm2RJ3
HgxGNX4+NrPsm4+H556u1MAtEubzZzaPRrx0Qixly2tLiUOHg5hVXFMaijdxlUeJdyhAldd9O1Fa
AF6j+l//gafvuchgLSfbduGjcYj5Ow/u/KCuq6gZoKtDjdZg4DpQT8an0RiPHsuJUk4DRrePm5f/
yWlFZ5cmIelPPoBHYA2mHrnO1Nd/ml8lHCdkYoKBgJJUF2EjCs15hS4MbIUO34giiyg/fQZw4biZ
A5jK3EmEG2v4RTlR1rFPFBOnFEH/wYM9oIvsPp6FLOIHqXCfXs/6HgfxEBF1s+IeqmtJG/G3hYey
3v8zLehxgsFV4aNtpxKDil5UywE1udrIA1JLMukGtwq9hRR/G81wxIYByxWj1x+IjYQ1m6G5Vx4X
HE5TlMtGS9rGBPrzQdfMsvSYIUUIClxq7i1uO4NCeD0BGQElNR00BY170VzdSrzkcDkSzb6D5JpP
yj8tpcvNYH/DzAHsz5dUhQIl3ds1j41i6CW7vJztBHfmb6KArqWKASAurcR58cLrEftl1YTJJ+q0
BGGZu3SQSqM+uiTAx3+BNcAvRk9tVdDckHvRWqJ6GcNxZF7lWd7gRT9psjvTgeKjdlBiyOtFXKjl
3IqFQxbSZNr9sRxELzlBRq+804k3ap9FETiFM60QTFyYb/eXsKS7viLLUSJvHQ8KDihTAmqAyZiw
siT/hSs+5aMxJKB6wUiSb3AhkJWK4J01vxfg3/9CorZRxrYrUxY20L5s/8PQ2K4Pl1dRrSW/5VOL
5IcnAv5CgeMg5BaVCdvyMhGiPw8LlGA+GGgDmiN67I022eT1ow3wwbvFr+a/EfKDe0juSmYvnLCS
Jmo1GjZEKxaShAtPHvJcsj9Wf5VRrm9YWS7JUiyN29Nm0i45ETrkfz+a+XSdSAX8oOAOBHKr6W3b
XULKnlzR8hM/GLBoS7gkRL3IeQK61qB3tUQGrMD/79bzVPo59fnA3URaKfjiz5Fpu7L7fEQa7P5C
x+RYynkQH4N8AcAVl/QA6/jaiDohvq4+OSyK4MRGeje039IBiMWaAd62rf1LcLDha/RuIWQS3WD4
ci/Jd+vFoyon4Sz4oMH9wsXRbxZ/HPX7HyJDdr1K/9bQR5cF3hUX2PEW8iI/AqXmlT6sJlpQ3VUt
fVWbn7sETXFbEsL3iTFAIORPiGks29pbPkcDVk5R20aEfGkQDlZ4Q63KFnsn0C3utuQJORKF3nVw
XUYARlAAD7qWMYqK4+2OJJPEoXYMWqLS5zIdKvFe78bzoja2P3Cv7LJy9VQ7qQYg3unCpqY7sZS8
D5gsPsj57NJ5yvY4bqC2tAkcp0YqxmNkHwDGX+MqblwQPz/9OoBNFHcfBbFKZRzHIEd9oTnL3Iko
2gC6MZ09e1cjvLH9sX2jqibPn1JepJoR+VEtmJWXKcOQL+VjXblRwflU1QltkTt8TdS7SSmy6mtM
6T6XNG3X+ET7zDKzr3EE9Eb0N99LxaYp0iZaL+H6fbWq2ikGm/Gxdfsr7K9mw7Wu62pJstP0nCH4
Q3qYOA/SUXI/osU1HotK7B64SdCMnjJCX7jbO4gL1t9gCo3LmMYq4kFO2piZhEfWs2mwOz/K4M6Q
JHFoe0xSfkRO1NBky11kqIK6lvhtC8NN1wur34SdRyIBusjq8mZFg5WfpPSsn+6S8Ukcjp6owg49
P3OgEyYJTKTMMo5GOKcHAzN3RtZcCICPzcbELrpgBJfPu6/3ytySbWjvchtplZJoVQEol0fZ0EmF
xeNhBuB1gw8pbvYs1H9UMUzsM/+iV47WrMspeIs30lj5shTA1Exlf1N15Hm7OF/l49AjgD9oQDdb
qmuPkAQIjPSac/l4HB9WFOhpZPGMZbm2hH6v3m6jJr4oHgP5C4QOc/bVkhtDJXZOapHisrtXXxQv
ahPWVzOXpNkR+LeQwCgVkXcp03AWmqM8/hGqJb5PNfjyXdsdKm4epapaueJafPK6JG8NOqMrlIzZ
SNq7x30Ba4JvqG+HtA6xKuT+GSG97z0FQn5BXR7OVMQh4h9OFJ4zVKn5O9KkRztyY6Unw6O31NA3
7ZN/tzDJkmDxj0j7Yr9mATlRqXRyHqRZTn1rQ8qe/MFk0s/oDBX9wg3UElVRXarFB38FtvZNTF6o
H9Gr088gZ2z6Q/G/KEOi47YeBSPXZB6EEE14zLOIG50VleapgtuuU6RfsmGLU4rUpGLuxKu5Dqyx
Rpj2/egD5UkvwToFGcJr9oo8cQzsPa1rOmxvHJg01qvlMRVYjwYVP2VrJD4ounoGIcPeFeo4mBim
1748xrFzNba2/pgZdJA6wh4/AHvuDGLnMpmFIcAWMos4OLPpF7+BiotHxwsYTjM7OBjh0//iSG8Z
5hBJAw51c2/dB01whtUuAXj+4IalNV2nRj5JaMIM1JIn0geccrgR7pjAr7mvVMU/tu30aTb8OltK
4ZMz3xW7Y8/uI3DdsPSAdJYfn+1LV4UOAX+R8zhhutC/QkaFjPwESHUhU8QbK8gIIWySvjwonKsQ
Ays18hZIiTMWiOmbg5QLlrVVvv6WLjHTzDE4i0ayLFrhTlDVsgbqCugZHQZVrJq1XNJXwOl9KQCs
ays6RLfrivB4I4tEvh2dzzek6q8ZHBsr0aGZBFM87Lua//dVfwwyc4qseUylb0uRG+Ae6/kBq/g5
7K9ClsE7/+WJ6RRNHO8GFeeKjuOUPMw42YNd93GOpNJdWFvXVZbGuSm4eVfB8fT3WUk+TMMcqCsK
sPPm3zLxEVOdBPq+bxeM27zhqjIVto/X3wGQYG1ed1ffWyE9a3OQRnW34kFVx/KgrP8bAZxd7agF
SBvBXz69Vs9RFy7KqkYvNup/WEenZTvTPzfxy1zs9syna36EO3pGuvOJxesuuPikO1GO0WtS8hgM
2Iug9ieApRlH0zjHKrn47d1orB4a0MQ5L4+pFMh+dmgk/RrYxbJhlsW0qPTaLuCgXWM6ViDyknez
rLuWevBhUB/0bd7O8fEgmKg30C0HH9g3pbVqb9ZjvZr0sVIMKJj64lGNbbZOq/6MYkOwDKsyOcXL
lo/w/N+Blo74/uSptPOEN4HUK+Vl91LxrEOvrzoc+7R8qYWRK9IXJ26HvHIxQpgTEWkPvDtvH/rv
/D5SzGjip2qRv23FQEbeE8np7ut8sSQ7IuImx3zUpZQfPcaxzMWQhDGtU+/zbBG2IbbqXG9j5EBa
bzU6W1cEZ3Vw986v7QNqWokY5H+6JILnrlumfhSBLslRIFFPy1TLC21f9xlKZlQBSZlzE3HWjKuB
1xCRu8pLaw5xuIfGCITA5obk+zi495CCIJsc6NviLds2C4yCVNuoi3b+42ZR7Ez+7l7IMkP/ohN6
UVfzkWnQRc9ynkUt9IvvOSGqQwKasDaKkHjeYf1yT2Slt1MC5suxQPVLqQA2MXWLlo11YTqP0wTX
DlVL67VsGSqgdt2+nIQmcV+6UkoBt98AvGfWVnyrpobvzssgrLmmH0rX9jVwjQOVNKEsh38yuGPJ
Jcy95OsimENAxr5xfscvyVRhTsFYz1yRMKtR/kAqQjZQLIo9toHsvNWrRgJtwN2OX38RktqD1ewY
mVXqS/QbKAyY1iSr07PQ3yGr3Myzi3c78Vpyt0uJXjoOUd7ZlaV2B9l0KEmpiF96YWktjo7vZlDs
txGLcPJDtNYZqdqV2iV01OfTitCoGD8/1pk/R5Jf/VXje7dOZPIxKoNFE9jKNxSQewqeUqsXrO//
78BEGF0euA26XqDJ4iDrR0PVEzb9AI1dwIj+3nTLPCvhN/YyRWEXnP3Hw6MxsYY0GsZUJQBwugx5
/r8fX+LPtEJBUdIjMJSeGvr/7nvqHn4hz9Q4qrVbL0cv3gLKS2zE+6kAtRKrQWPM9sExD5LGlDsD
vTpb8heev3p9Haml4ZJMp7xs3HUMKS5fMeptCHyXoqc1JD/ih7MMV/Tp7GsHCQMuwa1JdaVGeO91
4cCND7Z7NpGR7k7+GXqWil1/ImWouPWB5fXUsMxAwUUomEKZUUnd4mMGo8hC6ESsKQd1Wrs3JLsg
6b5SBFkpMfQH3ikowTQ7R0S4jKR0w1EL46FydoV2UZEnmtEnet3m5eblJulTFzVUEIFvLotX7nKv
ArnMfE81ZChF+N2j0lQMUG0RBJkVNC2CeduOXBYa9TkIz8IFoV/XpuD2Pefe/EVdwaHq+kNwG37d
8e0N7dqJncGOnS/FPU7r5sTUtvBk1cxRUo0QoAawl03FIORh45ok7tHN3QsL/1+1DcWZE6W9ykcC
J9u32/gbY6JtKm9q2eF5amOoTfpFgHbaiVSG64yaYsFVBkcSabqjy+xe2VEsxP6DYPP52kpsMxS0
nge3cBwutL3VHGH+gzyqRvzttAMx66yWgwobsBy6VWqPePf7rR//UB9ifUbXSj6J/riXJEBxJyO3
BAsWAecLOwvwI077wvXGuoe2OFRGU8P0W5anbpxElzGrPXAfb65EoFEGc9M3mhyjk2bWDYTVBgZu
J9X/MvfNT7t76OvN5Lx3683b2F3ibH42jtlsugHQ8bSN3r4vd8zZ3kkquXBqAhOn+nLTYP2UtsnA
1AlBi3ZKZvsqg18YDlxSrOUbdEHd94a3eBTa8zKgrWhH4bh0eGGxL8MwB9tDve8VlNVF/jYI/k8T
3l9vj3swDWyppiZRWd3WjBKPy+UzoFyY3TRlh5o3heS+z9GD0ETZKgqGXfta5yCK/RLcw3zD5Muw
BEZexQTJPDxudddQCApBUjGBuXE3t/4M6V0iDp6x/7pct+YkrKF2CpTL/cgT/CgE8L8O02tTN3uI
1gyng9wPVQ5d+GF8lAJsBXLMW4CIpSKvjozEljZM/BY8X9RXT9V6wu2OrbTxOGHXOrmTN4VrcGHV
2paT7Ew6q/abY5ZP86ZR/XtrL7XZMhLlp785TvY8UbGDc44grjzo4b6LujKRJROEcZT8HMOl30vx
gB/zYhX0EWHSIP5XC5py/OuDjAVx68t4pMtPPK+Ablk4bRcReYILVBQdWaR1BTxU3QRbox3Sh5xg
idg5GQ9M1WknuHwcJeMUI+BC7Fmkq9MqcgS/elHzX8MYkJhi0MXgvSBIqVQ3yGrBIhVMmDgQwKTB
ASgPOMCNN5Q/P0w7lgLUeFBPDO9nGjYuQCxuPnuJ8yA2mPliThm+e+O6Wx4WgIjvnCt3tz05A/iV
yAT8VBrH7zj3o2lwFiNaUaGMkVh5HchiUJiEm+cSUhPQp/ve+aRuJLzwIHIG/iV5Sn9rzZ1Ek3tj
81WeygwNlU0VOrlzVXsdG8etSuYEMwZUtDuuN8m5oCJH78TrsK7AHJ/toeNWpNWod7UK0bgoBUsI
u74JRh56cTOX1UWJN4M55aDvgrnWna+QW7maQm60bvPcP2Fyerd4xvRFGxVG5ns5/5F3xfrNM5Ey
9UThwU8cxJFJwWlBBYvljtfHI7Rr4r+9z7h2WHQvCSnxef3KokcV1hHEozQB8pZQCaG5B7UvFZ5/
VBOELZ9iPYwggtzYPZUnPicY3MTNiCW9biYAojCycebupgWrauaqJ6fPxchb8FQIEdtMJDiqhapN
iOtEkutC9umCDcGJairYlUoKUfJl5240nHqTo/GIWGLudda6jk6EvLJ95g24Mh3gtkccDWEu+cPa
AnhtK2BSKyGmV8qFVA9mySHgrzrXkjwNAgS5WpQWLG6324SfirvgjhoCAYVX5nw8R9vanqyqcAX9
0qcsHT3Pm41exAKQhjQdrXQ+Isd+2/N01wE0vCS2SQQhAY36/Y/th06CnzlY8eqDUKgR/FnJJ1XV
j3fd/hhGYLP4+wMbhckt6Fyd/kqpkMMPkmaK3VFxuW6C76J14qaJ4M3DSsiEv8r4GwPv+ShQ4F0+
fQ85kt9w4RDzvHcEluDm8TQhfNd5wQXselXVnEWaQw7T/dnrAOtpa4PTsz6kt+nHaK0TnMR0wWto
NSzv30nLGz3cFnKv9CX35F44o6YPRXTnKCuCEbjt8XBvd764E2zZa1R8R0+XfK/tpj3WjHtdLqUt
1cdiL32YJPKothVTLh4YxDsKXm5pUz49yqojKxlLOvddn0nTAvIKOUM35PKsfFI0m+2iEDfVe2ir
LkbzVPUVqyD4SiW6Hx9zCCg/0h7okQWLaIQhXbStzyrQxxRS9MR5f/YqZfVH6a9ZERt8IEFojINQ
k5tQ+nYBB3De1hlGDoY+jTojIoIut5cbPEbInT5wmxX5hQWGfRnTN8yjYN3+yHGCzqdhfcRoU+i+
pTu6x/2vevLgSAImZiv2MZDAwbamK0U0WrcFGoKPQtzfLfjVn5Ls8tVqoJchplBHxkVcUwSOI6T1
4KOu7rzDimvuvNyWtPU2Z2N08i5tLfZKP5INslZ06HqneS07SEHeN6KWDZZIGys4UgxiAXn8QfLG
6bn2WyiiOIGrC40nZCva6Sshh84iP7uKmE6wrJRge34FNtP8OGGSUjmi51jobsytEBjw4OIgYzTp
ohHt8LMj3s6E7AUeFM1Qv9y3U/WqgCQKVaTn4Cnp+XIey1bSeIMPl2G/tFHxhmvCX0w0rxgBIrl0
aeExP+vUvQ48zS7iF7+Cijg7ef4BKOhxr++MHl99U8fuLedm3ASeqTZ7yi54e0zibghQEvz7R5IK
HAw+8yMgAXyaBmplmaPoejvLZSVO+/n/RR2IJ936gxOzr8EvdrR951c7b9bAa81hHS/cOXxwdgn3
iZTWDsL2z2FP8VEido6XnMs9jCGBLD7Yyo4kEydyVnz3ltCU7mzS1xQoe4LOjVo83Sqc9lnR17DQ
r64ILAEjK3rIewP2/xzoBWrClh+FzVhxNUMjBfwRee8FEDtrn8RK2JEjS5v6z8lAE6ftpEb47NTo
h9teOAlXeiegAig3L/uD1JGZ1sOJI16MlWJ3UdwdkdHRW8dzxoXsgPiG7/Ow6coHddu1/Ocjzgy1
61IBBFeZOq32Z0FU7vVdVDdcE+SdZdBcF/z1fIlYhQhsyWvf4WmdiPj4nMUyNWP9ZzHAkNskeHRY
W8CADCKbc4fSJz+wUxWFLXiJz+MGQ7YQ+1mTyFGrBNRcxlThy5Bwe6Ke6W5CC+p5I3NxzfsP0S4u
Bk7wxhAK2Dt+47vsxzo+XfQWj/qjOQQ/PNlkf7d4nIemDahdEOxnqEhmuQ82rHmVgkSaRsIsqGeA
JbVLdr3ooi8FOcoxLTK8pmqFkIi2OqTNG3na19hZ8a04nwPL3G3m9R0/umrZ+FbeC87UYc2OH+KP
69HCL7ZMKuauBhiu9JAyaKSHxMDT/9eG7NmYcyJTwHPpnjfvjC4andcqX5SZF7WBQdAFcd0mpwsX
JiCKQ9xsq4zPn4LpZ/WNrL3fCS0pd6QRtTaKIY2V1lI/onk7GF73SVphYwuyBhqY2N/tL6N8aFO5
cajZeZgoQUwBpmbgJ5caOtBVpGC2h2Prt2xGpyOxs25cGCtq/wZE1E3ZP9SNyaNh2lZw1t4IGNXg
179W0ZbOT63UKlMmdn/sGVg40R9tihyw2RQhkqapaJ87F+GRz2IP4Zj+/+sKmJh70/FQBmjBoAyj
drs/WaUyXjMoe0X5ZMRET1rLikmM9JXpVvnqYBJkDqvTrNx9+RPSkiGLJEeRazuUelK34hqUHdHn
ciqhTr/1QyZWmmAbTRKgn2duhBeDJFe/t7JjeQ60bSYYfNmRfANZ+2cLm7r/bkEDU3TDqjzy27nD
ePumt9yMRt4wcCIh8cElTqeJ+ieFxcJTmmHZgknM+4SHRPBzyqgb4okuJq3KNj8E6phQeMr7BmGG
stIvj9oDZRFY5oKA7+GT57swl0GHPi7gt3jqlklxP2a7bos56mBTT+61TBxRb1ZEZT5oCmtQbWQv
4P7A12W3BRxc+B/yKHGGGIjRaH2Zi8rmRbii8ZN+bXaWqy09XEoANgn8F/DaEFDzE91bTMFDqvV4
Zl4BFxgaTrp14Urmrc0t3m51hcTqFzFuN6uDCxEt7F8qEXSKdzdA3HlH6I7uJHOiZtIBsrAvXmQ9
i85JHGbXckVXQtItrtKtg23JsPOOJJDl1YkQzKDgQnEFSjN/FPoN/uYeYqDujnPCVO0nvrzcoMk7
yRDYOSifuvXlksrcNpby+IS0BvTgmHjvHogMAeUdWgF/3COTc8DFG2eyqmdiHIa9y08nf1yA8xMe
ZqzOIeci6VC96PqehwgDFLgdqOknAVir8R3Sq6Duue+wbwF7AEFjW05cPEJqjxp1lL0p0/BbByzh
UOqfNMa7M6PfJc4PXkN0EsZk36u2lLJHTAlQm64qPyRcquXvE7VnFYRJLRoZJH0/JkTpS3irN0Uo
eajeBK9aKpUAEhLQrOZN/Ru7zcsDUJQlwTn8o7aX17c/Z2ZxhwWTryXOy23z7hb7+0qd9VX/x5tl
Fk1bcdsYD2H9/OMEccmy7dMiTU8p+r4t2Gz/WbMdVVamHnSpmUeKPPQ0r/8B1rHFyrVCix2Fjogw
2MZtQxKywwuPh69cD0y+PnlT3PO8e8tx3+iPCIYaFvRA3pl2DBe5LNuD6bGadA+AySVyV1ausQ65
exwlFa5tr6YodqbJsPTErFSI9M5ukNp3n+uPcoKlh8ENKO2Cb+RyFwVK0eIjm/J4VaNLz2/EOJAO
RwEpXJfFurBw6Jt+Rmsq0FujyuhwbhpUjFAXLVCHRrKxeICMm+y1uVtWUKiyN5bE2aCyMliDGCpe
etgczdLbWZlqins6jmy8MiZR3YW6YAPSNaMcqsU3jM54djYb/9e6Xc9DJ9InARCNkAvltQXj8NOD
slvCYqeA4Gxwx/dyXHMgBbNVuuuKPJVRBc6pxTQaweqb0767TP1Y37HQ20g0dljFxvfxB8T9g8C2
kXuv3gdWWPHSJbkA6QH4076080onOeLfUcarzQv/PhhTGdtnOhX7Hcsmi1idVNL/tIDvuymnMF+O
MY6rYUzpbXvskHuzi4FgA44rmvJwvXroxxSM8MW+VyiBToT0wlbZFZZdPBRompn1+YMQLmx9lJua
qiUh2/1g28f7UFZpWNbu9mEkA0rESVFFaLulAcChZ8mof64hEa8nchKBIlOGPbVspcaaVqkGji1t
XNxnzdjmPJEq0Rr2IrCG65HSwTQfYLvi6RhFOZ2RXT0NCzU3MMuWwU7ezgiTf8Cl9629VxEVQcut
Z2xCGSI4HzOD2+WhHb3m3+WVajde1TyuKZ1NsxIEHf57kTRXuCYguJvWLPNSqwsgqbjyynYvTkpl
rV++DadRQ0cKMfmgoRbfk5KjCpNx5NzT3dcENJjGqZC7K0BcTp8jw4caBTOYwNXWKtIR/6Mk6uzY
P+COh/grxkM8A0LKOG3QjjT24k+NeYGptIdb7NcEVDQp/J+VnCFhfD0ZHyX2EqS24lOnF85G1s3K
6EIZjDyAebtP2XlAlcUyTz/U03wq0/pKC4ry38iMh16y7wKfRftwlVtwE3Rc4eoFg5QMqm11SiH1
N3gaa46C4RACPgt6Ke1rkHaqxmPkyT8zHW+rm0E9DF9VJYsISZJWx5h4Zpu2fDHnuRLEfFgIztwS
QnhzCEd50na636Ay4KtIjnm+UaX0PYVwBIael7z2daKCnKOyCMtOdl9/s5f4vRaFzgJils1B4uTb
cLHvZzaYu6LZ8buBzOhrf/dlfaG2Yyf+Cobc+Omt0mDRwos6iatwx2F8wkRORY60iyf8NPkrBnzu
meOdfL/UjiJ+XQgi37zOWwBB8LwTrrBpaB3DBaC9uG5wgkGby4frSZxbxxmUSdNkQD5xA0tpzC7q
ZvURtO5207783Z5sVzVN0kCqdRC6QmIwLTmW4kDbz4Bj55/Zeeh3KcccgBIU+JrQ4mb82m8YXNfZ
NTDplSWMBa7/5KVeNYLOiygwOaPnBXBSvJa/sxk6kWPq8LqNMvHC3WUwh1lNQmGfBevFbVTaBjR6
oG9cLAYZBGYt4Km+jAoLOBovxDKnw4yrWODxVLB21SBacLUcuCWb4QVPzcka4F61A+doLXr3ZfYu
pkAuLhltOqE39BKqMqGGYRMgFzxZpcNNlGtpL1wtW1mLFbTL6zd78A91m37NxmSzh8WiqsFtiQAq
OzSjvbj4gmdmh2p4PkP5euV9/rc+Xyly2iksLGLn0hiYztvcv2O7sKJkF3ZERPxLMw0m7L+wA8Ey
TZi5itoCvwFgz9dNlNsvHeKvr+7yvDEHOboPMwVhnuAx/g0IQO87OKGutw9ydE1u2/m49QkV/pKg
LV8QWnytODRviOrYOT37NTMmwwr6eihjev6EwrsHc658/Jhy63Vp4MhOCTx8Bls0gPZBpDQsVK1N
6aNLZ2kkBCGwHtc5kA0ybbqHoTQCg0hdpctYyNs7hpkqwmT5nM3//Bmkx/7Y2/PCvGsTB9AMT6Ot
lt+KbVTutTKemTdcnI4kxA0ve1PiRQ7hbG0Zv4YxYORd+PnaV0np/K5Suw/B/XB9Aged2fclzwKR
myITqFqsVC6/pvptAHVOvgzG8nR27xQ5dQczfelTvss8H6o1g9WnhqcSQcoDprGx1/7IFJRpyLIR
uxu9irMAVf0mb+IjeIO8PAB8N6M6XMoPi5JDkGEHK6yR087zLeiaCaPWkefvdZghCcYbEcyoxogt
Ma5vgsLKl6DpxphWyQnhBvAThq00gzAPlr7EJM46OqEaEqBP1MdWkr6RQhFaS2EfJ3wvivfab9E0
g4Gfk9NbobTCWNencYzuj5RiAAvNI8+MDHxA7dmbxf18GQvHwoPaqKO6dcGvrrt4By7qxAWQvSYZ
yabCPot9WJvmstyPWhwsrHkWugY0rfwRvvkjsD8aMnOXYCD0Bru97cIUKTm7bcbH4/XvlrNtSAnE
CS+hPooY6HS5dIlYgzPoYZLLjU7OlbiSMnaVXdSPfbFT6SvYDGBJz9WQOl9pkYSKoU+gVEp5xIrs
Z6P/yBobsPuE72fBcdHn2N6HaLOWG/LxFHFDnnjNVP7mlJfk4pGhtWlPYjciyASmcHkPo0F4U+8S
BJEbqXkYY0uNQoKDmWmJXQnSwjaBYLxrkFsliZbQRF5qkL0X8OsvQRH6XRXK6LRLzGDxLFY9M+3o
rY1zPMSwdm8bZeLQI422xlgjQG/JMAzC2sTZcfrUY171djQy7oM5oagzr7F8VPzYYhURE8+eLqqU
9J5DDPWKtxKJDhiF7WigLBZST/czJldwkHMEizb5fMxAJ+5vbIg9wDvC2pzZIO+WUK7Ta0qI7sTj
21ePE+dCGDk/8WW2LQXy7nJIJtuc2LTqxxa6EBoIS1Z1WhHwlBEzyBQ60zI3ILWlZZevnXXA7SVL
ZWHk/J/2BqrgMCra30EmlM3wjSxZVcBBPwkb3P6fjyCdTb3sC03lSWiFLuNdSxN5by+NcCp66uTh
4DsYNMuNL4lhRX6f3rteVcBxLJq8Sy/tlx9HpdN7iLVvRDklhPppOGYM6akLpQB9fLaWuKbjpHUO
tOh0Ae4ANce7DN20+v3k7WisEDE1QfR2Sl0AIJPHVboHSYcd5cVaJWG4Piv7ZNJSLTuWElb0frul
WfQPqCKW6tAZU4Og9rImcHUrDUNjP3+9Hi1+dChnAGxfjs67RMp0UlQWvj0W1wkX6es0QuMKd0qC
5+FOjPNqXDzpwPycFH+3eSY1n4KrpvW/ca7Gep5GD8fWorhQNcewuPphO8ZicbYztcs2mjQe+BEp
ftrgfuRxeCNk8WjzTR/2eQuEDHzSw8JSM25rYeLiJn8nQxPW6KByTW/QNPnsx5ON9EhAx0CaTKQO
IBcgfVwD+erkfHVx7SqJ60xYSocwrLMuHTuxVvjYPWK6zuY5f8w8pQHnNK5G0Io4RZYEIuQwZErt
srDBBioILW6roTc3HMslhhWt5zkfrzE6kdStB2tLwGW6STzHK+kkn1+3tj5gYnNWRCLlM2pVyYw0
Ofj6LesCPD+Z8iUApF0bmwgrnUmCNmzpxkkOM4nAX06OfTg5xRrqR7oW1ZJRWR2w2gsm/EDHAIBI
OWN57cLkT95m3SUhxeQLSH6ZjGPkDQWvOdBed4xDxTQK5G4MMzntBsK6IKK/4OlmhHAHoiC8O5Sw
rEIchSSW5To05QnUMI7pUMBKwSZWJmtc+5VE+QxmqkG/x+PQ6aA2gfmfIPh8Qb5EKzCUbGS7gqNk
0TuzTRPjtQc8OTO1dzdcmyvWNcHakK+24htbC3KM3m+mvkGLBnp+IUt2K6i9pi+3qRrabVpCJjxx
ea5I1yA3nhFKquXBUqupP68iS89I8CDA8z7Ebv43/6wmKX3eNYv4HJ+7kl6vmHRqghte0tXPXS2k
/mJ2rHmThDnK3xkGtyBs206YJGJD/V8bNrC394VhvkfMA80ET7I58TWKj2YX9UW1m6bVn1tKcnmQ
YS3fsJIS9mGHB791ToeL4X2Fet+VSgItHvs0q/OdTLZo3P5aUSjZCsPhGUYMZ/AwQEMQ2GmeDGJO
Z5UBVLVS6Q/ktXfDig2q03da64vhlRQwoV2GHuv8ay7hcnuzoW4t3jBtVqPZYKjrNpMvDaSml6B0
ZNyVtOMO9kwX2LTK8tOjI2Gbs6hSXxCYJYtoBYMqHJ+ENfh/IW/f7LSpRVncMO1u6tSJLdzEaTpb
XlL42/IZBCEABFYv0BTIZUHBLM3pxoJrjnWrzGJLCr0bB8/ENm29gfytDSFvHLHjBXXg8dmRQaiZ
JJJjlsXfGSjbwmbMLisNgFBGorlUP0WtyFpKXd8oz3UqnJO9W8pG0e3er8bxlSy1Zk8RRneYwVsA
D7wWlgQIO8DaLfBWE4sGVlzauRylpWuUjG5IsooWi5GB1ySnt202+ba073maEx0u6lvpmVIbp+/1
5MvE+ZuslhAfKua7m4JrI2wu5bEVWkSjHaS3HDL80ziGkE/MUknzNKcsVeR+2xhe3GQQAkG/X7VP
oDSMW3wPfpFm6hqA5xvm38W6GmncI/D+exawC4YOfe6S8nS8iENm44qZvDGQOINmgtb5JkBdtxMR
x9Czlchl/B34mskSfrvgR/DZSI4LuxCstCZF7ycaqBvHIagVi659Lg/3iO4+VbsTKrC+Z89y8S/9
64t7+hinUA69VTJFiWScLqyCq/5c0q1aftWwLfo/PTjnn/ssIWjHGp0Iv0Fp09vQf+P/OPSp6FSR
PUKE21SKLm7hR9QURb2H9a61vZKony9ysvlVc3nX/YYtxRtUAFqgqMbNcrFO27q3ggC6OpND134+
sRCJ6qvNeRBW9a2WhbqkBam89oHkYUG/J2PUh42sRblgWRixu0NBzE5x9aFCnLND5f2r3zDlGr9l
v35XxNx/1SzvynAodnvBeT0Zonr1TUn3rrO+/g8YZj3bXwA4vV6Ngy3/V69k9iuihFfFMahTZ8O7
TRYEN2E8I8qPOLIpV0yJa67jQ2xXQMcDkThX0ucpmgnCvBZ6vOUxFKUsqdGIBrJ992V+eKm1p2+2
LqrjXKkIaKujgAlD+QOPr0xORrng7HRYI7ENCHM4b3InaGrM9EitpncvwydPfosId827uIrEUcAm
/GA5BijC8chVvyFhJyc7jdJ7nUyLSWFmVKtqepq3NZAa2AYaR9PJXd3lDnw0cdHpG5QzbmbLfpWi
cgHgPb3G0q3NlPbTBOOAGF3o5sQtsyJjUJAO6QrFkRhrHy1dPO18ZbOde7hHQYpf0h8znn2SRR8+
/Fsb2mdrh8g7nkPNWXDk7aF1QHzIJr9VmBIiGfjWk8eeWYynYJN8aWrhQKhkSHTe/gkFx85pijU4
xwmyhqNUur5MZQJMSRTpMAXI2hzWketc1I7U0QfaDCp59x0oaY3ndnT/SLdtIOCZwYwen7+Z7FkP
KsnZmjZ4WyY+zEI1y5HrG9lK+bvyZYvnDAxzyeon9ptGcDbwz9yB3dhLe1mlURwTo50x28H5PryP
eI6bxwy0Vtj5jDQVmd36sNIg7D+4u19d3wDZJqSVo2FufKb8Eh1I2zOeZtPVr3x5EmFRgWR2m3y9
wTWcOdixaOgPFl3NqOxOV18I53SPXqMrqzqhjT7RE++3wL/ZjRaIFtmOPjYxY+qXH8Uy9UMtlkv8
WHkj1iUY9mFILFEPVLJjlmybXDiXhQK+cLcm3G5erekasaMYL3Zcm/ZL8+a28X/VCljb59TchJJy
nIixqfqm4MM0+TaqgOxzZvUV9ZKIHGsQbhJkMLKjo2yiL6Qf+ljUuFLPti0eCu/zIw3dOfuWtM/H
V/2VaKIaKIxWG4P1/z/CodOdRagtBOvVt0Qh12N2EbWy7l3hfYsLyXkEXozu5OXzXYrxwcaamA0g
PRMFLGTWI4E7xZOey0MBSWk3VGUnnx7/BdodRJNzvpqgAJx0kFs749z/3HR0ZLyFc1CldDopVMjJ
AcITdN6BqTFNL5g24k7N6E4YwtmF8KGxWMa9wpT/on48b3yuMQKw5yW5FwP0WLOF/ZM5VxCRg+pE
pTbsPQsZp90iPc51KZZcZ1s+AcaIxhPSAUEZDKOtsnCHSYY+4rBSyZgNboKVn0Ax4AREUH8cL0uO
DToJcldMUvk64XBbgOL1cqT9XH6poLXOpIhlMSMh0Pt8jWRfhpuWQHf9ewGelIgZGNkofbamkYGN
TrR8tvIUfUSaMo8UMz5ZYmsuk6j0w1ApQi3NTDivYnLiZ8Vc4qVtceCG3bOuMxg4gUmEPhRSZ17p
98aq6UGz3Z+xR9UE6pukXtDGlQrDY/JnPaOfE1BIr5fq1vgfmdmB7NBljqhISYoiJqNflpMiuPsm
KoQHJf3zd2OH9QHIHd0kCgIjgUt/Di1WrSLzCgbsEHb9USdqIwqo47mC8HISopv0GUNNv+dYP/g1
sDWTuQ/cqhE+0HjIwMR51wZ62iDcR/0Scz0Cjc6GKfGbrlRUf+k8F0aQF4EBQuVNlDryXYcpnGCG
3PQoXbyVxjSHMTcnQAu4/irxevW/GX9rwMLzhnnvKxw3KBFXn4rlg/nK2bcdfGN7SnvdSiY2FDDb
FDYAV4b14XL/TOpBLuG2hPmCf6IXyjRAjyS1si0zRHzOq33iG9iQKB2vy+8YaDdTBM78tCPweyDD
tTGReA5d/oASTrAi00S9JGtmPXxgyqm9g6UvcY/soORgDiAvmFCbxg0jGCGqKshmfe2SZNMalqcL
UA482314JzAFWNfEE0b+y8S4kKOy24rWFJpK4yIyR0MEDR29/kDVP8ic4RseqGKI8NArH3hmzWmv
Prid2zm/uh9/T45HU1a5puHeVme3Jn8VbM5g4LiNOlzni5AMS6oT7oaAaJcbUHebIh7PDha6rm2F
8YxHR94KZrydA+j7IZKLva4dSq8cGLj3hLCUtCDWpsDH9aZlJz5Q6UYdXqmyr+Ylo/Vsw2NDJktk
mAQH0q3XAqRtjnbtw9TtRvWKDHtg53j8X8Sie9SWHlZqQlb52LA1W5Frplm9ImimGxeqpFKOv43P
RoC8kCxVRNBTvkZqjbroi8OGUnsUfm7XwQ6t6g+8Q0ZEhtwftIUnUN4OPZ6hug3vdHKCQ9WmJJdR
QTveppqaHFgVgfJvIUZ/dh3KmEAEzKxkvL0U5oCHEcOmrP7Q40RJI6fcRRYF/0RLI/YiD1z92lCG
odwt4uS46s3u+UtyHGfwmxFaeCn4cO9qGZgbvSDjW5Mxw/Lz1gBOZkHSjFhPNMbhQDIZ6YCHooHM
ZuO3Nmjm/hUbE+Lr5IkUu4XyHcpxOK6miW2HVGFcu+0I58fbBRDBWhAEbUOxOu1lzEDmdpRwHS19
OpHGAKh69GQnjQBVKKKgSb9z6rM2UyB87PlHDOckpmDWyMO9i04r9bwsJ4xlAS/Sm9ZFv27qYz/p
pZHoqJFFVifGrqsn6pbJXGrOyuEF/z0JRhxPTFq2QKtyC9/F7jFUB9ByhcAWtJa8Md9d6YLSwhBy
gNCBhQlDqjncwQq8aChLhLc3YoUwBnz2XXWLftRnqCvCoc5I9FQA5Ix0YPOiihKy3nvYB4LrweeI
wHtDuPHtz8JvXXet/wwbK/LYdzveYsJ/nuDupkoscTGW4SqEzOuAzk/qjsxJNio/XKef9/JmRQev
n1BtxT0MKM+WDGMOwmuSCgHkwsq4akFOq3Mm2Es/fVgdY6h7Zw80CNJLQNHLZ9S2kjySyzOXdLyi
v5CyunhYRsEKtBgY1thMAyh71HFunbr7FkoGqbtGiUaZfoGeXyB4NgPGLD3WmHmysEnj3YCpEHzC
HVURaJOB0WvfVsa75y+IeB79rkM/V+CT/+zWlct8qznbEWt/0TKt20T1HvmIp2c4nZJ1R/A0oNOg
Jzp/evYGwLqP2X3J+B2GKEQckJhq8oAcTvAOoO7jt2eOrfLoojwXLNoIt9H4JrzlNxF9J8PoRWPP
BujgjFE4fMFO1ksr8k3qVeVvXxbM2QlutkT+aCm44PJrSUu3QqLgQmz9BgTS8QyAF5m72oVEFkZt
VqKm5USBKW7mxAOPjWDeXG7jc5lXYyCcajEOEkFHh0lxQpGPSoOQgcrZOK1gjZvPQuSRZ2jGsmON
j4rHNgZRXST2aUaOb1eIPyx/ylfAMDt3sufjzYGglejStpGwsoPPR8dQgUuuUzdObsXzQXoy0QqH
aBuUporo07v0xFY881pUI3qfP9NWCp5OtjzwB6ljtRKYLqieniRV9NpTGBjfn4Qc9Ye6nImnBIQ9
/ty8iFa9fhcuT6OhnMGourqB+gjeMo1a0kshdJlt4Qzj7XNbgQd4f3J/OQDluif2OvIJvJwuD5+i
vA9kTUvWUi71fKcwBJz4y9ZnsnK7YeLmilyU67/y3RiZBWhLf2UThRgl4OWeOEvbLkN+4ZshkoxZ
dU9LKk3fHkI+4BL+TVDGwhxk9+D8tzx6+m8yoOKewsDYgznYNwOHQfmAJb+Xm6duaOyl0GqbTMpq
SL1amTbRBbjbryWSzxEa1h02XSk7HDkhlogiIjCHIqeD7IHdLoumzarXvDJG5NrKRXdeKk6erChN
DLc5tO5YZQC02MvgEYDJ2XufUkpE7OCCYRz+SnnzxGlkOQYvwwwkT34uy6hOJVbmimEwrmh9LF0e
yimNETKsE7xDf1Z2+XujKDMrkw0u4Kx53WLDGr5Ydz6RPz2c8/dAD0LLM5foa++Hu9BOM3G9Q/Am
6LEkevaEza7/zNpBY1QpH8n13RZ/cDUvjQI73GrsmXAxiTjenrm8SaG7no3cYavmrlUbidt0Hj0V
6693ZcPpG2i+WYhE4IyEDL//WWjWRLE1bLSHaDNTEG0nzdhvVxWkxgZTkO8KMBrw9wvlywTnxC5D
kWCHkqEYYYy1C284cqsp4So7qpu1aqBhk7tv6nWlGKSCBENU2SR74u5NDCNFpSlcwiZyYaKsNPw8
ifWHyjyMo4D02KlFOzTKL6273y4QjPF5h1FP9IHLJHsxaaSJ9hlEieW6dQQjpeZzQhCesrHCgp0U
UEnkflnKEmmH/jlL5n31e/Ezwj4dv5FEHPxVUOzJov/y3aXJmOPxkzlLMPx/kGgsXb6YOrZ0j6Rz
tpwXFVgwViN0K+q56X8cCUvLVvObAwCIHHB5qSuo33db2oAenVDP9LPT2757ovrkoI9OWTds9//U
KCgkSpwgDzYjpv720X04ssGmpkKf60gbWJkI552IArY3spiShQs6K554zSCnW7gPrsrJWOOSKxSQ
ho2TGh4ir/7ehhmVCg0E9YT+70dEp1PC81yy+Rjg48/AjoUEmVa0OHtjQo6b2Mz1jIY4wQ2IsyaA
dd2So52SmfGsgCD0S4796KIdvFCr5lZ9ZCCnAyPARIs1tY6jwVEH0/NJGPuYd+39yPQBiprWgY6f
dhx9EssZdAbqCixfbTHODb0XhLeOE0n2qqUbH7fXE3lgugLV2ZC7fAGsJiB6M0wYdR5PhLM4jSpi
PpIe1bGcIuAtscHkfF1UvceqoXwua3CGhxF5W5Lpx7rFbarpibuIzy3GDpKCRDYfaRiYGigRJNxc
3xE1g14J6EIpUd55id+KrQ9tPT2to83Yn0nEv1LUPMGYiGg409Q/kPO2PPehw6Wf0kH1ltArRvU2
u5POtE1w65D1awnqn+i7KXuwatlfAiihymvYFdUTxVPZVb/UTtv8g8RuZ+GtYMGYUIHRR4ZaXqGk
qQ9CYNlpvIsd8Yg27IjopsjqiY2ITrsJBk04hVRFxs/FGmKEsq0Jb/u91qRSsmUEgtYG9dBUqcJp
WVYUoak/e1jIqnnKWPaqSwj3lwWpuMF7E52HLHICOEyohl5HC0y5q1EZV6H98AqPf5uR3afNevZa
CHUH2rLuwMQIHV6mhgJGgzM7xYxf0k8pwCXTzIsoHQs4WgLYA8lFGbNDeBYfTMxdam7rc3kZDIE8
PEqdhl8MemPD/572+YkokD1R+1SpuMIpluMVSIzQXNyQJY4kmAIOaSs3SlT0zrdD2ViYH0Y9Iau5
eKSEXrDKdvc9cGwkYrH6ET+h8qQcargbpZvxd8GLpXySXv5Yy4COuwuW4Lb0EMBhL8sI9WBThmnc
JdCNli2pcD4vds8591eCWrPkuzFJJmn57SAg7kVAvUMdK+9Tsj0F06zSzf8/HQOCymH9Kht8IUWi
To+h5/bkx/nu0QBDoMvc36gSJakt1jbRkvQqppyMMv4kXObWEawBheou2H55koA8jGPQciN7CEp+
+ObPnQ5dbaOvMQ/Lhgu+fP4VRo9XXnWVreMiVn7J9oD2iJb8x32X8pHMZA5sa78yFPZwRyqUzhc/
Kl9sM6pfo17v5Rv/kHhhn5p1/PtqQBHPt0jMCpwuU5diA2M4+u5ZrLf0Ce+qlCSbE28c53MNHRBW
OC3CBofmidirbRB+vZnNRUYcvWgsdkpw8GrQkSHhlUwBovHXAzgvKvTYrEkwjE3gBQ2lpS+oAM59
iuhF1xCrETdB+R9WzZl5z18xGzbwuZF5mS6d00lNwdCkBgHuhFZyDssbvhN9dFxuQ4RO7Mgx3q7P
YDpXsqmxqxGwoPoWdLg9JsA2ODIfrKXjxASzqzV5B80cliaYanRmY20pbWvMSEtc81ihtABOqp9c
6xgmIWnxX1YFHtd/02l3Q9dC71/KNi0PR4mutwOlR2Wk6L7R8y3dHYRDxAHzCXK1xw2YMgT7A3tq
fU0LlBDQ24PEEIkmVjXG+9zgpnhwPp2i5Zhvhmse4Xhdn8iv0KyFRdfNEDpD3GFuSb6/lQ3GHJpS
HuWxa/ulxuXvjF+i6/NXPJ9m1tKe1Gu6oY2s9D6i3cvJTIFJe4+p1JPy2XdeKmeMITXC0j4D6kfe
1JXCQVqH4P5yO73aoQMYNeRrqByZjVlIDtLPjUGeoR25EI4ko8Q4il2geypBnttFZN/H7TdLTq8Y
g7n9sXQx9hF94ugGz4M8JqH0MjkiQVIlppzWmvlPwvtLBt4wX25MZhxQ0eWm48mKiOxnbFm4kR3g
674q7UV8XErcN0zz9/XWgfOoHYtle0PuQxEwNXu2/U5M0WdqijhaJ5o9l/6i8dyKgsSGqNcyVswn
m+SxXUWWxbzWVq/6Rs3rtRu+gu5LiK8xcQWg47lWV1fprQVkJgE2EMcwk7XotH/Tb3moJG/QlK0O
szPjZpjJH8lNvX3pm5HYRfA9jSPo1Aa2rH21EV5wWhBy3Z8X/BecfyBFxlnq47NI906RYEya/vBm
3Osl8GvVg9h2BbMAIMBHd/mY84qJAq9V7TAGMoXES8T2nI7FsMiCTlFK1wlOPuxqJowUa+g6CXg9
EfkrYtO95wRvErpeo4wJG9BSB8Ab94D0hwb7diL3NgRF8UUtb48qNS/DwHyYCbcA8dikhvmDUdMx
4gH8csHcv7PGHoo+Bl/YeqfoVi3AD+fFm9tW6g6Y+BlG5nB+il75rG2IS6hgf7l2aUMXxPe8rdWu
kPU26ubaTW77qBX+8J0xJ/Wcb5XTI2w89tiZYsx/I891Rad+04d2QGd2FknsmVr2gTpfQz5s6QPW
FBr/8yEF+1UpBz83QztkcmoQAvbHpi3vR03vPfF07zxJTQgnH3boIthk9J6nzztwJCGPbmEn1JGY
rHbSYstxbuKanp8r5Hp2iPn6lWxFN75VtUtJjPN+e2pQoVRev/xxP5qBPFKGu++EpBT+fgFVPr2M
pVEpWBhW5rtwY929iHaffmx7DfQCgArQ6vgCOvFyxY4+V2y0p7fry6LtSMsGfb/a2C4OzBm+ZJVB
eTTPytKB3BaX+dJT4tjuX2idgVc20C+eZg6/KhNLVX7xDy2EZ4k9YxZmkbAp3qWej0l3smL2VwMK
jWaNrYlFfw49fxYfkI/jOFc+raE3vFzn1o7pAPD5n+GPCMPZOU2DSKZ0h5/DvWjmIQQ9JPDE7xUS
U/a/ZkNaOqJsEu3G/wuCG5CVwEnYrea9w41mKvdwRA7IUnH5i8EXXTIonhCdKfygxFzCgy5h4ZNa
rQoC2A2gEmIzC/qKBVAXGbV55syaO2oF49kcOH5O+On11QHdIGM26ucnXMb7UBs+gNLyshOQWs/u
XKjROmXFAZ3YR2GUqtfJYrLNVBgd8oaJ2JL6U6GHjlyN6eUPaNlYaRa+3t3bWZro+9y0X1uZs2MT
gJ2IU3nv0btpDFvwg6YaHKkX4EW0ocJVpLC3D85EP9qpRv7uRAtU3m9tUn7zLipHRbJAS4/SpU2l
R0fhnxG87kS8yj+Nw5tr3JtN24MQuwSpLV+o3CO0/+x6MUGZAJa8ufBxwHSHV4CIB3Wc7ab0iG9n
9VvXUeqZG/to02NIwyr3I7QXp7QUz8ZGgfJGrJ7wk150CwuRkpAz0ab6IljMd9+vJOuRTSwJ/4Ca
1tQbqhwI3vfgECMK8W6t3XmWysn2MTHk7sqfq92/j2eVXWOuUrW/zzX+9aH3e4jkIg+YhNORRjh1
gjE6PJCvxSqQh/n5n7OEQczZvHLaxv922jTyQCc0qk/AEzHPfYt6bhXNjBdxHzl8BBfJ3Cq+ludj
NMF3FODqVepsOi0pLaAaW8Z5tVHq963+F91JhbM8+PKT69Xg13YQ81WpHAfATB6uWOc8C2jz2SKT
C6TLZni6XHudhF2JCBBRz4dAMQx9TYUDxGi3rEZX9AKGVXMlCdNwYg8p+Ym4cDhYz2Q7L7FIv0Re
GVRw2tIlT0gL+x1sqCiGM6toGexqxXDXxCAwbdSzO7Wf0BXmb06xidownJoQnDg640rSi2DYJH6r
excColFk04e/K+Y/AnlPVdSjyFTapSlzPp9Ag3KzGo9pI7wHrejlBajvbl7Em/OtLCvWKdsXMOPq
bNq0Uk4ayfMlqimz+KwTnLGe13+TDIO5fjMvtDxqKvZ1fUMUnnYjDu7ppere/mPO3b5inswTYoP4
HISyqYuHDukuoEy1haOjNjxUlMnieC1tedrU2qN9aYhJtrp5VN/5Il9mRMSCmt9NKHX4Z/HBrM7r
2sVUsNriS9rFw1NUDqxRiOWI8izYx+e5BLsq2y8dbvgy6GouKKv/Qcd229ay+IkU3ELvaXg5neCb
ZKeCmlEv1NpZ9tg/kXBOfjVxIaQtgnopJTmo9R6jq0jGfXYx58QvHXrGneUEyncRV9qHLr15GIWl
xc1yUCNu1Q5+7YfK2eptFcNlsxNLNgLMosOayRaDBT1GRU3CYBIuc3jSEmZcLkowf/MAia86BFFH
NDgf10gZykobwhtpytThuN6EqZiKo+PZt/parGVs+GbF9H0b6+rV3+yUQ3ELRDpdwe3xj+Su5V7+
GMn94Squb9b/bY6aObUPvlqqXkA1IZNfPPSAjAcN4leXPTfyemW2eMuHNE80aYY/EKcPqmScyT/H
0qZfxqrAg1JzcwesNr10eEWWvQe+uRXHQBe6yVpzAOM7uUh4W94Z+mXiZxdp6vjPPwfcl0/Bl3wP
FwsJhWZ+j6qYWxN3imWrlQo06wRFXtkf7NZ5YRxM2O9YPvLkujvB8WGDEg7pvSOFT4AL7gWYPWTE
kxZIS2sGeY+nrPm+MIsWJr6RTGOIf31M/bZkjTvYbhvbOOuMVztFUq6cNmeECuvHf22zIfp/QuUg
WBkLLYS7PPloglidrSotkWjYjkU7frCUcndBLMy77wlPuFeVNrni1T35SM+//rj3hNndU8rEZczQ
C5gdmklSiGvjc1YAJ8q28NyyA6WY4arVajhA8yXGgiRHy6GSyUykeDYF1UWsGUwQsfOrUA5A/X7R
vrcTrcQqLenWZekJGcdP630ZmTy/qhKj8W5O0cNAGAsjeR1uQSie6+kN/MO6LvP1A1TW2KEyiZFy
b9FAKxgxc2dYGzoD8slDUeUnux3Oxfxc3y4pbbk8jOwkAW/lftbOsKGKE6Z5s71F7j+WlwsFzcGD
7oYy65msRiNGzZ2+g/jx3V04KeVTZakVjdNdoTEk2Jw/0OOTx2gMDGQ9D8hMRsDAsV6RdnB/H9zz
kB7sksky5bvlSmbrHTBUafcUZn06FKg9SPd1P7MFZ+rfXvd+5+rv2LK/bwMT2B8ceoQhRVE5rR1P
LxJ1047peSIdKqMJa1ZxcpIXqNoZcrchHjl+gh1X6rqFp3UOCEM1fLzwtEU8cfuxH7DtBDVE4lu0
TZOWH6VjYdC4yjQbIOdyGrqtezZU2J9XArlvNzujgsziaSbxDbxdbD2XmbRKC3wugs5QVkd06E1i
jQ/S7saoKsOJwKeQwOOHk4yuEm5yjQd01/TvDkniSEQ6QjOxKbv7Yew95pAqevn1F2ebiKT3HbdH
t5IJrETGT0PBzhbR5KXr7KA+hMguA7/1I6HF4GMZJ3RViIEnqDS5tC4a24ryHx5O9agQd3rf8N5T
C0qkEg8AfCp+ze5OY23X3dJ8bKZNuWP/DzeV+THnKwyv85Ewwqy2C1aHrkNkz/4b/p3obxPuSuT6
5QG4VGF844sQQGimXvRkwMoQOEX/FCEuLQ0nWc4Du+A0rPBQviWwXQbR5PjNB01SHMLRkO9uxlDb
Qj9fiYgmt4/lymr+CwvQKQ5ydpYxF/OOI5vAvcNKVT1uivvBSEIhQG0FDnG4jC8udWC61wiRA5ZU
MgyWZm2VdEWoKoHB7XK6H2bFR/A9b8bpXZI8cGDMLh54rj52V0f7VyRO0/5cuKqFfw0D1pIJxdEr
OnSFUrrpFyUop2VO0WTvVxT5wY52IG+qK6ua6SNEO5esmrEkw74A0UNzAcgqZR+bpftyhYVQqyF8
4RNcSue31ZtUjLLEwMCWH8tdpSsNhGOwWvc/EaXZywGqOqjzc/HlgoxkrlpuS/+fXDOrbipLlfaz
0daPR9RLD+4fYmBgj1IFNEnX7RWYkHPCPUeC1WpW7yUq59MWVXX2IYyJ2sDnu8SZgf9LA079vpSD
/eKewuKKp9+skxQJ4owuXY6reX6VMIeCiS39XbMXtvKRTOpIBTsqzOvc2fE5PcEsN0O2QoecUqL4
8nPgKWuLTx5vRpo2VB5GUOSoqPFLSIn9WdkWBFxKJoPsjpogjQUjCnn8PuKSXH613BiOJZfNDS3R
HBr5+R9ZjDjSUGPyhF0W4/Dv3tDi67NSdzti9KCOgO/mWbkDBX98PY0DuNv+30J+vicyM942TFsX
zE2eLeRCJPUlAybUmDWJbO5ItbwEUL4iQkB1WHZ8RpdG0rojbeuzYxaXCv+Z98P8AcDG8i9nAfc3
h4HhiR9eRVfzEzpGKosc8MIUrBDuQfKpy/fSmZwWXbHO4DMgp+uZp9zeDf3wtbB0IlEpO2rbZZwo
jiZ8VLU96k06uErx5zpHvN0g5kiKQfssCBY784BUxZtNEEhsNZevPu3k5U5YavSpw//8n5UlDK2p
rzU+w52/xxHBvcvho15uqWQzneLVoN4uE0Mukhb0G8YgNi7U8r7x/HTJu8mijsEobTQMPZgEcLLW
VWWzF8/bhY6VplZBeCFSay+4PjyY0ZKCrFFGxVLi4Yce22Ltd9VtlrJopbWle8IpxThwoSrVVzTK
7ikEtO4dffHPvQ4LOMwHlofy8qWCk7WYM8TtQWGQyKMjb2Wz+Gsd8QLYjfalvsiuxqjF7KDxA226
IV1twvaGPGtQGem973xUMXvzpPlWiWwqKuBsoS7BJIv1b/eZtiudJ+OT6ILwY7br8fnkQK63cBhL
ConM3lBkD2SHo2RCkxbhIqt2WTc8w2DDvumQyusE1FbR6+GkuVgwe7/DpSGKaR1X0cyrIGGbYOw3
5sdY6+QnL6/FfGOxIPIwakSSvevSrlBACAbXiNptfB1GrlkL/qIUXePuTjM883Voy2DchLTKkUtI
TiYX8lKOStSnnVFgC/FQpjqBjfFJv/YFkINfdwyPvcLqIDUHIuAnsMu1w+pCImFQmrfslFprLH2R
XuVzH5V17qZlxd5+HZt8Csw19CIT8JtqlflZ1mJRV8RdFTZb+xtcBtgNYXXJK/YqXc2RnHrka8PZ
cvOhSbgyLI6ZJdcUM58upRFNb9nAA/KRFdeaI7buosUDnxqvpRBrdQFR3sVFZVn9Rc2LBmoxwE/R
xeDLZ+KBmWvkvawULyj/yoYcVXte8cFJ1JzBlr6wtAOZWaE97CcRV1x20060UrtwNvDErHjCwCuW
8jmTvLCaSVHDd70i3xSOlrZ9YR3fDMoLooJ9HCMkUN02Ni8PdeIiyIRlufk/BBuXtWfuTvSPVKIg
cDEgmJTALPoHssJkF7WD6bfSncNtXuNLhDmUmhqDJ0f8ThbfzcGs5eEtfthWZktmes5dHwnqdGN7
zuT/kSjz0nn/jfjuNg1wWlejzrbIPLz1kb5TRWL0luYEgwDHQuceDUYWN8vtVG2hJuQ5ne8kQLe6
gxG0k8u1S2l3vpJoEcAPKODg5gBJPC4oJXlyFNmTbdW7rWNCsPXvz7f6nLTbnLT+fFd/Py2BKLNm
Bz5JBaskW7R1RdvKQfYbIPFF49Oeln+3w3GLtB2T7WBHzsoZ+j4Ws7CmSF3Eyj20wRmTKY5BBhew
AW9ALi83y7l+UuKPtuBReVn6EcocAOLwQqcBdNTPKoMxeJfQ6pVWRhs10JNIk3kV4eKg1BIMMi8Y
oWA9ZOSFonOyRjLOTjbD/QorpIylgE5G/JWLAWCAoZJN7Y/PNBtboA/5ZqhCKpt2IdO9dajeO/Zw
hNhPQmw41Hfqiy2erw/fOd+GsFp3ZtKwjdPZmQXp89b/g7PCuJWiASSTn2sYYuKdvJGLtygWJpVG
2VxLp95HmWU6vDKHSn1HKyivlObk3079SvUR3Cdb55yZ+uDN7neIobPokMxWMVZ+E1kECeXRNgdl
SoPbLfB9iSHdWclDQx8DxoZM6KLLBgNPQPmf/046ZJyosksMZ+VYLJoQKdObUYwvVJeeQTZ3uS2U
z2/k86gFZ4owR/YDUmcl8atoJknx9h0oMcVmGSCH/VMQ8XR9X7WBq6Dx2j0sMAvn3mGVPW28rjq9
w1Dwu3ShrJVBRlPaCzS4NzldPUN1fH5so0gqLy80olqB7RCgByuyFuHXpPys/dOMW8+jknRX6XsZ
jRaQQGG98hDxc9wxS5pURK1z1srTD7NZCnVASHFA6FX4rGHii8HT1i6/0AT6W4NKs/9EMRco31+k
v15e0Z6EjCjZQUw0o1FdZVNI/AzDONcjRy0h1+GJtQEnfSCoLlaJyKuSj3A1Rzr9IrFZsjbjjZqa
J21Q9R5Yos6wn04jbwJa23klULcV83TKsODg+EmkbSxRri2QeCg1DPGFgYvx0BUukuX+A8Z99zi0
0H84IKPLPJcR65TZVKUBtakUz78C75egBQC1mfp7MzFSH1As3c2AJ+F/FNMZI9ulcO+zd9FWeRDO
r50MVSDHj80eFTYHsUK841O3t9fSVawWOQL9QCaJ8GxgqYjC8mbiaOIasXr4ze7eQdUc3EwJQ9i5
rn9h93DTLsFhr892eLgqvDZNdpLwsIwytiKCzXKxRolnD1q3Dzg+rAP+YrKoua17XcqeuG5q/K+r
qDkiEJkGxgtw698AUmLsXMJqEWxB1xkCJOfPYDrNOix2BSgK5fdLGKWFvIpYZb/VUkCuGercshkw
Sf9Vr3iwuz6nSYnhceC5wBYbtWeuFhQUVBou6N513TmrquW0gGb5KxvFx956WHFn5C+/8Qz4ks8s
kbYcIW05pod5FvUWLuG/+L6dO8WhXufTUEYvqWmCzG7t7U2EDYHCgqMjM9xmkBdCMN/4yrDVQr05
73g48mZcb43IaX2RsVYZuHps+ojW9AQj07Bh0JtnMMoaEmbVKDGNtPj5eDMorLfCXFHA5FGujSAl
MCR9s9vsA51pQJ7+mkEMnE32dykuDIL5F4OB8w8t+As9S2QoxhEIjyr8gud7W1npKS/7ti85ic41
C83azBQrz2/J1Y7DwZaTYI1kf3ZSDcls9/Ggv1VDP53nGD9/eF9FWq2jExrz5edR6VtgvgNgUeU3
shTOT2ZJU2xKQCFhqT74HCzEimsEb8pw6Brgxf9/WSgDGtaNfAyhYwWu7CPIOwp7YxeJ9iBeJEug
9Ex35rnthJNegHEMLgypimaVvBcMPNNmvbbA7fbj8beIyyKfs2W4cEfKZNVkw7ynGcBePxsy6cn6
gGSGi47jcB5/gg3ZiXJqIuQh2brb/6UJ/MMNc54579vRu1Q0n9r438lMn3yal2o3GY4IU0dh8U4m
rgr3fG3s5L/PQmyUV5BgGQDrAPmaFb2AzWtH+mdeGHT1QwgjDUkcl94j3fGMqnjtgGfshttuhYzn
2p065gi3Igo9w6BO4/CdWWgDD6wqj18Vg6kqQKi9lytQco5Nw4nPtszxDL8Tco21vLTuvuK4nms6
dRByS4oo7EfsZqa7LMlqF+DaPLPQTFCagjl9ryvkEY39xx7F+VcDSAS9/XHFDFQK0uk+TBvRhsGA
mfOU6IMZYB6W+buzbku8TC5edRSNHzyO7OAUkCtVcEYubsJBvP8Ly6busk5WhOMElDqb2agLZNsM
lvYhOjfiVAj5q0chw4BQtSV+BJDPlMLVgwbvAumcI6hWrYQbUoWgR+nUReBgZ71xNckag4rFCE9W
vtxO6JgFEa6pd0CVwFv6N5Noc+cwn4r7S8QtLtxuEqDM9DPSJ82FSgdmRbLqUoj1p7HLWBPCgnoi
FvjNZCpf+FW3kcFP5ijSPyv1AHlBn0Vkp5pvIN7CHg5XIp1/LIDgx4aAY43ZdvBOXd00z/i/+qEf
36tNjTXFMdJcn0/E7SEmUoxc7vah3BUNvkP8EydMEswuq42LgKK22IE8HOGlYa/NL7fZDGkeE/Q0
QVILk75tmBUz1fvpvtvZnt2ijjkLYrNN6CVY3nERswtdrfkuHrmMp5G3ocVK6WklgDvHA78kvin+
27szpXuQkZVZ7IsDR09wk3vtfM+5fkbarlPLNv6phmwG0eC1z0A5+kkvrgbNR6vfAWl30lTpzjv/
1nZoKJJE0FgFVroFdhI67gRiGQZGike+/SJv5wvqzltBseIBYyN6hmGPX+xOcYJzbxIBZkG5DCmo
maOz9h8TARVORPGgLatxIXRwKP1NiuCd2LO4MXaQDPvtSpOwfE7rCzX4n0kl5Ii0RrJUgLv5SuWF
KBTvnrfBffm6ZVdpkExHNIUv/aQuP+XBRungb+0yDWyD5iNrZpru9BUBT0+8yzwqY8Um2ofE3HgC
oF3st/exdnB3CQ0RHivPlYUudRbP1aIJ6lTJnypBxLXz0fkyxTp6T+OBVi1tCkOzdpalL3VGw8H4
MHGsjwZazL6Eb/2JXTZhdiUuxmcxXxaE2nNThsCtK8YdNGdJexnOiAJhuKyOHsVflrzoBhymzLux
+zx45yG5yaBCVFLaKnp8pE0TQtVj/LzLsZ87gjOtkQg3NCYYywYSPgfiv9cw/S0oqBu1BeNv7/Xd
DwmY+Nk0F2KH/MTvqFWKBnhA4llJ6gLAEsk5eV/O4GOXukNnv2sxnSHedb19jrENB3RHZa/fRQP3
HO/lIehSZsHxAhIpesoticy9qXHSdf/mskaDqF1nVMXD2aebXTR/OxM+Wp0vRj8nQW1+AnGy7qhm
fitwX+qct7MVlQ/4kojQGAuiPdrggK/okaVzuYsUyEbH2AcyFJO/npUZR6SJBqgt32varZzGOJxm
maDLqrNcnV8GzRwFoitJHzoY1OVLS7TUxGwhMe1bOWRfD5s1KMN4jwySlarZnMAN3KGvBZBWYTSd
/OEenGBXjKRemLGiH11xpdgPvWeI3UPsLXxsJAmoaNyXuiL26CWW4XuhTrbHHCF8N4uS1KmsMaVr
1uXCYJIFbjUISKQha0P40AAUz7yb9rvg7YvrDdSpOnTVVDtB3wQ9xsSs+T0Dd0xBdLLRItrRAZNG
HD9Ka0CClmWc47Ezy70ZuXq0kXD4TtEGlcnmO4ApLkV3mJqWxBSfFsQPsHLgfculjVTBfcnSvaAF
M7bE+JUlIadAR/5daAz8tO4f0fdwx7uyk0Q1RfJIoYMR2i2EllC+MAQdBp/3G+PgpWAA+Mjy8nUl
vBrda8X1/jl7bblQejmIGGy9guQU0kbf1swH5rDVceTUl8Ax6YX0kAhjdTcBMHcfs2ZtxYr0tz44
tP5jXD8Tnp8EmgEcBGSYuMr8ltqpcLhItkfi4s62b8IK11zVjAh9ICcYWp3voxC16Zj+n6ANHlJ+
zWoAvOhlFjwvGq8cORYhE/69vn7kWssR8x/bQPRuhnFH/uSmvAioqFQ4E91+DEjEX/gfeXD1U/po
2S2gs7koloKYgQ9OHNVn9ea89BwR+Fxs9EPCnpH7+8yuIv7P0+0rHIZbJ1k9Um0KVk6m84L0JLBF
SxTvfE935vMP0qarXkokMReJyROqQXhjDcnEYoTGd6OtPK3Ciqqfxg6Wzcj3CHYlj2rUQoBKuKld
ewXooK2I3mAnB4vX2xLC2Vk3P7N8o6hLo4hcd9ZQ/kylp7ZjPPYPfj7kTysGm5MD9b6Xsqq1wcjI
7jj7TjVo7vFqS1+K4HzRDviUGyCMsxlXrh8OPWp4Ud4unHiqD8ruE7brKWRLYVNm8T00tip/D0vh
6bC3wmlQ0lL3PfMcJ+BruKvgGTsziaMDYhSCTdvLJZ/AmqLFUzpusDpqD8t2HdroNc44LjGv/9sj
fiXjnl4/Uw/SIWf7o/7ajp4WJfQx7rqksil1TqVRMsfUeTd7SMgzsr5K0PSfkPi+gqPfVTA/cfIr
69skyZQVOnMx3PSbOHaYMQSoauKpM0L8sl5gIU8KkU9M/aXAqrPFq2f0hrx/wGVGG+yJlKaJxpZc
m6GRj3V7y9XyuizeNJZ89tYg4selmlgI1qA37hXe9HZYccoKOxYFgfXeD8wGyTewOJxtLUCXqUf2
Vsm1Zr9Ggcgzn6ww5njij+LxueZOCUuBVp65H/Gpiu5O+daS7nzUUk+A3qtG7FAAc7eSoSH81P22
WJ55rvHFeQEB4q0R2d5oa562VAxgecXtKkla8KyrroK4ZAaxHHtf/tSEjy6WAvi6kf04pBDSJKgi
W0ahyBj+6Ay5mGCvGCcvR/wmQw+pNDVhT3aextLimrWgsow7J8BKf7LjqzGolatZuoWK7F5hvQUo
3Fcv7i80ifeoR1mfWKmFGU1k7xlv+ijzYHU6pz4Vq4r8bJeO4uZUiy03Mkut69c6/f+ghadJStDz
HWPdHxnQP2/AEPhL3IRQuugIt3rdDs++M58Ha+wD+sDF9le/ieRolbclhznzwNvaRWylLRAedLC4
NZN2sHO2hKo55zNF6IMwzjzIKQ7bjGhRU+crJLMAJlK6IQlZsTiSKgQ639Qgjd1kK5RdwapRSpBE
EeniLu+CsHI1ho6q1qW3sZnGsaAvfk1Q22gC8j2lo0AXUlaXIDFuoeu4I81htLz1RCZrb3K4UH57
flhtvjdmG7y+CCNaCKDvyjMwyYgf7ECOjEAyg9KxPnpAbGaUYxsO7m/nqy2lsZP/+KVMxL2ISzK2
KuQAA0hzRt6rkZUGGpOWc8vPRAFThpGCzZV6cbQ2iOm53HeU6Ylt3CCvrJekGxWQhm2M7tZ9VzLs
2WPvs/DaFs4cG3rfq8lpioLa6VpK/lzHER3/QZjB983vbNPgL6BZSz0odIPWf0Ezo7Z8tZKgwrAa
zFaFShOxNlwYUsYLP8Lq4u9hbq8rPOOQEkX20t2638G95lVht4W0keeo6Y99pdKWseL64dYi2/Q4
3YQuWaCfssXiApwA1SwhI0JKTI9Qo66YSuLp77RjgTb6Vz12H2CXdb/yHSd1qyV8ofgmoZq4fWpL
JWM+UV2Qe+oohCJnb2jcoOFhcMuG8Wh+fyxelvcgJLADoch9pmKmJ3FV4OUXS7O5/6oZorvrtaN6
7aQX50P69/FoQps08hEa45+C3ocgrnLJgiF/8kBDO9BzD8Gyf2fnjbr50hHMcTkED8zdle5SHvvT
NUwMNRuA67AbI68TVXA+C2l5ZORT3sx76kzzZJyICmsB2Cxg7joP8khOSfxJG6V/dTuZkZ+N1z1c
Wmd/xC5NKtpGeN6qaoOw1cSuPY5Q3Ci0CjpCyS4lG3zZbiiapY06OHrFi3RrfKqSizlrWBq7DeiG
CWd7gZcmc8Y7QDlc6ZhI829pb1eSZyim5xIPKEYO6VVXP4tMDXjEPjOeQTBkLDoQU48FWzvr24z+
/Mva90MV0+e12Ct5h1jEMs3y9za6Kt2bsStoA+vA77shUMmCKcKNCu9gNk/res267H5/p9mniXrr
xOOpBS5rWusmjoHZdjBWVA7Q5R45jbsdQLqNoCTONboX++OW0VqjKQLmhg3KEfNJWNJSTEY8z6Hl
RBa+f0kpEhlknzg841tjoOcMh1Lav3RkDSO6i030AB7EM0D2FHLsSZPInEY5LKMTswd5pjrddU5z
qf2yMDsFMMOJGpmDOz0f1xtR9xzP6CGPq3hbshmjKERQ3Zw5Fr9Ujn+soGkmV2Mn4WEGkN8rQVZi
Ze7+Y89/2AgrRQk03lKWhGxe22WbSKDoB/xl4WJ6KDjBqsUvZGgzlmr2z/ZAMYWCYh3CSS9FkpDD
UXUwiPFvNVAwhurEaqd6W0Zw4ByemC5wj28LeDhII8Mp3UgqS/N//GGMlk7sypIeaNxGXR85VqK7
QcrMjq/eKIv9zC3avtswm4RMn0iGEcRYJ3hjKaLCht2jYeK++JunLNnhCiDDu/ld4wjogaWGVA79
oXMk+Ci88Shltq9cW98eaMqb7cUYqFd1uPkZ8mI8aqpsN87XXK7wjXIfnynOHZDvFM94NDH1JlmD
BFaXtvS5c3KPgeEXSDQyLBOoLqlmawKKRJzNV8JOXsIWhV29LcbtO8V/ZKb0wobPJ0bbxCoPY4vr
f592+00syfiPOB5MZfm2DTDZp1jXCZtzzvhUPx3ctpPc9AOf3G+xjz2ZiK57CUP5MtA3fykbv5r5
FOlp+6RlSYfyWQY71LH1oIHL8KE8VPJcKW7CowKtV3jOYUksA1rdvgdZjJJMrf0O178lf6rRyFeu
n8rXkTp/CdqTXqnzgAjsBvbAT79DpFQS8BLCW7A/Vxt2UnuFQOo7JFJx7/3veCd5JwsKeSNs9wRi
bJN1KAjWl6P/zt3AYKp5ihQYNvvvudNwlHQfdlpiMPD69e7EPEbV03WAEqy01faD2ax+cM0whblm
P/6A+nTOdUtLTHeNHS49+kddO5IBZ3UPFM8C6+y6eVZfs3XYcNUIp8bX+oxSn+Bt34zG+KIDPF1v
t1qmhKYBKymQg+pzH8Mh0t1XxsC9uvA5uSVN4jbbOQPBs56GgYj2w8LZEnHY0IYz1k/hgWlblpMk
8G2BQXnm/q91fOZj9us6gy9kJTIeQ+G6g80j6YGJlJ0BtCpElcDfZRHiqSbeqyouZG+r9hLrOSkH
uS/waEv+S4GNK3HZNIqgleGUlqOBP+1LjZBOZC0QGA21seioWBwdmpZN82bu8k780MqDQ3Lr1g72
3Gp0c07NX+QsTvXdJboHE3LLHpOL7gDfaq36yvy6fV4KbFxU3D5tMoMF4s/l5ya4tTdzbe3yVTOW
PaFezy6kMVyW1kH/Az83ukti8XzcYbL+aHKc8Q63t5S9mnr9zdtgUPWaYoWu/FeUpUzkM1/gJAXh
5qMq6/DxILafRD16pGETSyKdu/+E/q19a7oij3prlHPa4Btu/+8TZyYV9mDo41aEiuRzQ2QN7g53
82BySiscB8SxceJDHi4jyCNoUxPFj41AsH09QcbK7D2hnzDONU9e3ZaO5KU4NKqxKrLxYqsOnLyz
8uP/Kkw0Ao7fsO8fsEqrTinwJiPjO/4uXB+e3bN+DmddRQHghfAnS2advN/cDCJzGj8MlPSucDEB
F2WLcuP8ChAEoGOi+yQObJJKReJlGlIE6Rp4HA/TYmaBWBVfgi1SMbLmRdjKphJD+SYL1/JdEYEB
yf8MyCqSCGmwf+Wpdtoh5uxg9bW96Db4i5BFHfQjSdX0UbHkw+oXzk4Qy057/SZL3JpYGHv1P/Ct
YY55VoUa1kjifGCcfIXVpGQqRgvhylHm2qFYnE3y0o4BO/CHu31LiAJt12+FfAHPLWXYhSIwW4OU
eBqEvwFiXCt60ij0tx1hRkwG2ATRCNbNTAYgsbfCXkeFItoxdnKNTwBDsOamSoJsAhk9G5WG6bRd
SEGzRCGQdaM+deRcgtvJAjzHbAyReoESZb8FvhJc1oTQanxdAEPkizVJgvHaj+KEssPnB3MGkuJE
gW7P2i6N4qzdQbkFuMFGIDPC2iBD5BbNHH6084Aan9EemWZrEO1+4Su7HZxpZO2dvbAu606ZJCBi
HZB1lr9pnaTjWd36T9f348xu9DDaHDcw8b6uVQZgz2dsMAgjmaKLcq4SgWiO7bAhiuFSyvcG9EOx
M2Jr98uxVVeiSrmomyI0JjhDdmtjbyz8OJWO7ybOvgHw+bywApnErdiICk0tR7j38HHvcwoh2HK/
ZdzzKD2jmtt3X0wWKIsi+JRgJxBBvCOXvi6xd7+3ImnvkA0/WoNG9n9uuQB276sSBGzSZRB1DnAC
xp2JnPGBYAs38R4m2veLIo0qHImmKFHLTb2KAqq4d73CkKoUOmGRaAA93z0SKjULkUv4dIeARQmm
xGc4VIH1PM7VeXV+FPazmW5vLI+677DjrCLe6ZTMC+xVy2fCCsO3Ka1OOyJt7pVDP+kA3pIPlybi
OVqD0b8cwm4+ncdmRmFAHvFsuvlU0EYqxINYChV9lpHQT1ImlhYWYqQNU4mKrPJ2oE6+j3Q0PfcK
CX8+neuPgvKQ0dQV9qqbMsQpipyYokKMkqlblFwWTuOIk+qrp5eTSP+utDtVLFNVOVsjQzQsmqG1
/MCXO958VpIal8M6PhGhdMQcvqTklYPs8Q1U9/CHv5Svu7+mxM4moOAX8j/SSEVM95836rQYpOsp
h2l1LKawtFljdWnTkaGcRmJfl4LJHLnXaH9H5zoeM8Vr4x4M+DUCG/qJTBRgelN1L3HZsIU4Hkz3
MPxMjfwkX3Qo700mChJNUawDO85DxnAMEF/EK0t7IAOIXlleFjBpgGEqFmvj/qx5/6gSwy2qc2a8
R8EL5CrY8m5aC72sub2oyrCdFzHD8PfrTou7wiMwNeoPVgX2wh4pwLUU33kth/QVwqHCNW6FkZb6
XUskxuJ9kBdb9KA8/soS/DIQW3bKcLiO378iNsQLwpyMUlxHfmAw0f0ogaZtQ6WAglfSNE1n6hmW
N9QPcz4w/Qa4rpPorXFWkf3g247Pwafh000hcbwRzdjalwtni3uTXMRiQV5SLim90Xq39jzszoAF
taFplu1f+wrGR9VElt1BLD6WbCyMVbSld6JvZ3c8YlnIpQ1lnwoE8P2jwHK2FmCH9428/3D0MVTj
8NPyJqJFa+ocQ2pBOK9VBTFq89KWhweI2AlQggBurhdB1IlprJ/gkHzwAT0uLmf6nQBMnA6nIoHM
lY/BncySrOsvMdlvAFrMfXPUHPaN4kMTKTTKzl/j/CV00JcKaiVOtBNVhcn9Avuzzp8Hmuz558+c
2avyF3hkRCpH4U4Uvkl1+uMnneg7yy4ufBb7lIBDUsK1SqDRbc+vNlamlI/AFtnnR8F2z9YpVKqd
LJSmI4gF0lYYv3xgU9Qhe2eolwRu/aVoKdIV8zoG6KCUkgbvtGIslFXRo0KZl1xNkOWTB2lLyZeP
eVjKhWzhmRpvs0+ZSF2gA5MRypdUxm7lvsrGAMGkE7WKQfGyoWQmuEESQ4hH3DsRSHlXdOje5Q0D
jk4HTblKZuSG7zkfJifwst8GyjJq4DUEi5LBNn5TXONJAyCvP1hHGBunbnR0cOV/COn9Pm+bMUhE
/30eMqVHOEQV37BhdK3TwgW/IqjbDXUCAMIT3t5gR3RtRa8sv07JmU9tDROf2iIqpGALmuLVRVnL
n2ugnkUynTf9U6dBUCKvW5GQ98WjIgC6LY5uIZHG3SE2oAuJ32uew08VnxH46bovwobCxHAGBcPF
YxQM1oiUKJim0vP2aKyYDOBYB6wf8WeOzSvLctaGViJiWuclEO7VUAsdWe4jt/S4ucHyeWqsoi6G
4lIkWu4ydxUz68/0EQoJjYqtXC9YrJ4iFtv3adgqBuKEPbMSBDv4NxJsqtObU4IuZJDiDN7HefEp
WeLiauUwQuBw9UW74HVh+auEUGc+8sBR2B3bS9fbn2K1hf1ubqnELmRUgM/DvKBbqe9CN+eVdZIl
EuuwdLpMKBmbyJ0IgmxHhYe+EVyA6ykHmAYsPowDSTWJCU929IV6jxMiHdmV5ozSwkBVXL5lVmYG
qPRU88aX/J4iqvb2q1WxoXGNlmkloCu6Bg2rhYMhnCA7rhWdVB663S9wCdLzMBeYhbVEhzY2LHyi
nFmWGksmjaxgwp11BV6Prxnc70rs0fhWn8PDWpwzVqmSijMm1+/US/jeznI2KqzGJS9mAkYqe3fe
+KknN0e18U05KMN/vE0bAUQHvmW3TuCnAqJAikclfdCrgBf1jp7xMLl/+zIElfQvTUGwDPy4Q9nb
7MIWhpghPgzf5DQR7UJ+LNf4LYR36mePmW6eKW1zBCmGailr7mAEEsebZOZi5YwhA6PuybDXVUQU
M1YDrgrMvPBOTYMZIw1mVplyjDzttjIWGL7c9OXUgacFz3D0v6Xx/9rT2N/d4LVJaGOcW62hqLRE
fVknxYprHjXhfZuJ5LA4lXUBuRCGp3c45bytX4LfNWh1eSgkGViYu86mc4/1yZW6gtjnaXiXENgu
lYQku309aQwYIE4s/MOsF27evi2yGAQ9bvTGHmIlH0yljyZL6gvgqOHbmoxpsPLLGN0hnXlNd9u/
cfbgw5XCvLmnypd+PPiSGBCJQiWbGFUniYTVQnpQAgnFrwBD75/nJxF6RKQ/u/2r0PJqP0VmRhas
tNBlrMtr3WFRyp/JbxiYVABv0XBKG3W/UGPkqOCYtGW1q8rVQ90iUdgo18ExL0GPRW/pCno3Pd9I
qM0JQR8yNiuPtVYEBJ/hHOv56wure4DF6v9FRM7z2pXV0rJeRdjBJyQup5D+rZgflLatpFVqQO8d
ZmvN1Dg2j1L1jGF5AF+7WWt/HrCTtHBJMVI+F8kA9n2Vm2HzDaIo5WLf9XDtwyNoYsnFaL9A4CCD
KiKAf2xnXDMQr59aAbd8HULT2Q67+rhvr77JX/EPkKJjP1kAQlVDYZ3e+egxzRPoqquo1QjfsHiH
w7c+ba1HfzUsUNNScrN7M2K8muumV+3Q8H5JWt0DlTAMncx0J9WQeCQCI/gXHVuTWBMT/g5exdJe
6M18r/337p2JE35GeSoyzVVxFnjChMX6UPKkagN9uMne8RRUrXjszDWMY45/P4qEVoGV5ZMsrvwV
MZ+9Ha6OOdl0qu2YWi318o3GGqrY/o32PJL3pecbkHmxgi7Mu2wUBVMsSsdEFUFPc/S5cAn+Voc9
MUqvTaGRXrtKLr13EFh0iFZIv9q0VC4uPesg1KNAjZRqHRfoU2w6n6zLWh321yvBOU8Ug2KBrEiA
maSeajZr9UpzNXPThfkQsQKCOYfNtP2NBSuC8lHI2N47K1DUJCn/a2omvhqM386TZGArqMN13lOB
C7zapOPYn3pjLl6bExizPXsaq6eSzUTgX2qaOMrkB6wpspYgroYOb4E/+lKnhGNKfDLT7AZg2uqL
LVr/Yihk9PsKfahe3SZBXJt63yM2OjzAHAt0vLscEObtlhtYkYoSSpqvHk2p6nVBNsuSRlpVrRmg
XTG5zE0XZuXzwarD3IZnwmmlXaFn/BIjkLbgwqznGgxUYpkBDMHEkjpQ5Gm5wpN5xXMFhJM8bVev
GtVcHQwNUlvV21l8+KhhIDvkfFiqkEn5LOxVJVDSL24sjXPVgNdhyhWea0/hmbr5NXuu0j65Cri5
lVbFrUHi9MJ2yzFKdF7pSSIZ7No0aqmv2sTkSF28TYlpGbjfO+DTgFnQ42GInJcnnQW2KmfHrkBT
DOKJ1TiwagqybDdWHP05i2M8fJHalmRam3bzRmgSK+HH8LAwOzbI2tZriOTFhPAgirA5CDJxCbbt
BBYqVq3C85VaOtl0AtoH5UfUR39EUpphourokHJsdYiH3+FfcEGySgy41V6tGMWssJOBO2OOhdmF
cTNUH/Kw2KnCVmaMqWvt7xZmkWg+WmHaVZe8QuTGfiIfBU6K9tLZOfnAfIV/+krhALz+iDpw0+Oc
c9vfYfvRAWMpJ0TDlZ9OuUL8TQISLVphjyBp6qMq966U/9+CjWq41yePCxspMlW9kK34sDmmjR+B
rpAAkAB3d49XKsqDTUZsqZ3MtYzWUtJ0r5LfxTuKFUR9D1Zq5nQLIRtJ/Qn2wV4mjJN6JqXAJSPq
VSffeFJI6r+9S3mMehQ5p6Z+SsqPPJiO/lBtAz7KDB48Ud8Ri1BjbTWqHYhE+NTyzwBn3HZMxOda
C+GgtugFbDniqgYjR7W0UERHZnYtS1mqSjjJ9IE7cXd5+uOUkO6mJ6AnOh8ngJ3P6v16eVG0/9m2
M/Z+VLqRAsal4Gf235cXonZfbIL7X8FGmuATiEVkOOjIF0qWxyjdROy5b2z16FODvobZQhpAAwhs
mFhBDXQameSmy9B6BhwicR4Vt+l1/zPs+UBwkg1kE+ZGBH6gWWkV+jby7s6uEdMDhocqGZqdIl9O
NldSjR080/4qDIT0H75sgkivtM5R+WeTCZiP2BVqD2XR+hRaSMYJEdHRolTBo0o348wvFifqmQ/n
a3pPNKIv9UM9m+3AJ6ERuagQGXziF4yOfUR4DjDqgNgxxUC27p5J9+ybUo0A9ROnD5q2a3/hNKHk
hnTvIPXcC1aT7Wj6RgZV4lxrVroz8EMJaR2utp2QIxPYLbNFkX5OYqqUAV3w5drYBgXrwTjPwwCo
LIaDRQZoCwqPyig5F/hROn2zbrfbBzjVdsygUmqT+187jIYdATsUsWJCadYsSzEJ/LVlXvlKMT6Z
MJqJTL556X43peBtm8Wu5LlwiDKXj5UZ30owG9yCn5lxO0fGPzkz4zblNLApAiT0i2Pg8mDbSwNq
OtMTtAGNoJAuVohfMYcD5baWKqoAWSMv4tjKICcjnJX0X0U5IpcxYsZkaIaRftBmgM43nkedkvnw
N9UOqE8EpgrFRjZ3fEuE7zo+7zL1Msf5dQBiuu+wkOXtpkCZVLnnzeXgoS48/1XQNx8hruYqmLt4
MQT1RYRualRKZfIZ6IpoXxToTmcunaEledFYfpWVDx66XDuCvcelc9y1cHZL8gUe3PHQXchUOguA
affT+Wv1vlFgPKZkEVFd+UOjFOmU/pm7p4D7e1gSTIjVLn+htwSzZXw6mzfrN+sUU7pjBJleVPfj
1A5qfTjsHFt20zjXkwdIZ5xzGDe5KuV6BIdNartwv4QgTajkGIZ2/AsX2mmjAsdpooh3jd0uhFR1
wE92jNpmcMtYmo3JxE9sp9XuXhsJUy18WEpu1gYNGFBzbIpYFXGU2Np9ySH5DriXV5Z6SGa8KWv8
9eqh1/LnMtE80UmmWFrbXwiXr47yGvQ8+6dYclnbtstNMyh9toK+u7DUJHh7wc8XiRMVEsqRNlle
kZQC5cgius5wB8Dj/WBV6oUign3c9xpmbhnjB/eYXndbl624NbcqaiNcuxVtIFlXrJNNAveBgVkF
eF1elQTTFEi91hyZQjH6DiGpbc4yRhIYifnFz1rmbm3nndaUh9b87u6510vfAhp4jlZgfUECGKpe
xnwcRbC0DRx44A3xv/mPTaUDV3YcrSYmHUFWVsjFKXg76+sNN8PiGkPyElEaV7Et1FkVfabZV+50
SxRDFInWiYlYMQqsIjnvfzX6nFm5pTAEwwHI7hl/52CUrFzWGo2vMtrx/EyE08V8ESNT7/KRwdIO
vaYUwpsz4oqN8E4gXBmCA4kAMZIZwZ4rn2oNY/HeDaE5NIeRM6f4Of3/0R1CeNaJdgDuO7skE7tl
do6MFVLndxuNbKCUQhY/3Dcy5BXRhO2z8yjllxt3B2NfNUlQrpHyAZoS/bXD4B4h8wG9yt8mb4fB
IhSlhHgWKiGN4QOxjDE7P3H46umjxT6yxUkMpj6rxa5c/Xd4yqBd8joT63yp+oOiGGMLJf6u+kkk
RsfPCM3gGHd0Fuzk0c2/RqtLHtRnBW+2h1AdhxoI3gTU6NpWhUacmRMVMVYp7XxZPH/LYY6T8xSD
WHMDAEZ/4BLP2gIHmJn881IHLfo/NgBPHaORapBU+QKOadYXOJBiZG18UtVmCbTeb3P5NV19f/vR
3AS7GBdcuFJCRz+62HWf+anbUbo6uog3Gwns4IxRXZIA+Wv+DiXEWwL5PZSlc5AB4KJIzuewz9ha
8iclruh0mRHyCFg/AtZ8+KA6fE8NDCJQC6PHW0Eo3YcgXQDcD3KGG1TZ81mJ7GhkHaTPIAa3mDjZ
qJDoJy7SrRFItyl4YnXum4KgOpvcUb70XhlY1iwtxwTyXoORnsW6s939c+wkFKD5JrJgojXqqIQf
EdI0VnzLaJ2un9oZ7YMKl2uZvMtQ9/kxmDbn7Fr1ZtwbEICvX8OCeJe9kc4ymZOCkFX/omfp19fX
40UC05IfUY+95AWFQpxDsQEXXIYEH5+6qfL7NHyrTXjE8bJ0X01eJwu9nHkXnhLbQmXvEGpc8AcT
C7c3CwtArQwgaoH7V3lPtlswvEBdq7kJrzKUJZlPJc++/fzyhCpkkz1qcbOU7gyBNtBPnzXNGgpV
9R2nbg3J/g+itw4ix0YeIpGYLVeKWKho1XDqDQ/GFEf0sgHGxYDiSgxFl3bC5V5lgQA+YgGYkV2R
01mDgwzlJ8exIen2jlu3dCiaTKvcscL7kaRk2WDzkiw1fdn8FlgoFObUWuh2d0LLh2SwHnlzvr3s
97D8NbN3pW6OOSVNh2uFs5KdRu8O5YKMgTtrLkK5ZlCegekzBzEo4AM2STY0dDUN1o07VfaZjyo7
vdorjKqIUW1J15gaVsrRFsfWP5sjytMmcGiDwiPgeXWL6PqFSMIkTmVp1E3B9EpRMP4Mj3Yu4T0z
LO5kwE/V7Jwa0xWEU+LKkAHdaAc9VESoBZmRwTZkPn8ePH1Qqef1rPPsYNa6AEVyskKRsJB5w6mo
EN10Jct6vynyn3aWceGLiyV2J4Ak+TqI5pheUvJnSWyZSagxsT1Yj3MbPsaqz2HstArFA9+8vGWs
j/EZSk3A3KpJkrkAA0ieJWK1NQ7dP+85YdagFwmTx6Xp7gFR2GQWqEj8+UF3fsG6ILMJvqGm9C8E
PWnKKNAc6Y94uXQ9FypHipWBukxZYUz7CoKcBHQdDSQ4nnjqEWG9q05BBOSDqpC98tmMA7aXmtE7
vSqf5GtdLHe4HqPu8OBdJzkocE36Vbw0mSaTgTZ4uo0Br8c+J2FqP+KEwE7Ya9mCT0ccEyKUIKAj
AirEPjiDO9DsfgZnUuXz688oQpYvaY4WIRyWdTF3usW1FlT8DWmxYGMojut0zr+Y4M/Oj/WaYWSe
910q26e7BrhC3f7lh2DfVJ/rEfi4O7+4nJpmN3p8b1o20utq3A53ym4X2J6q75JGteY6+r+BzzOm
GlmOJd7ZjjAm8lOGWJq2kzPjKnWCpSQ4aERRCZeMtRTHrCkwSIBYIAbMQREkQMfQtfLCMBbtl07R
K0pIL6QMWdrVPcDQnNzPy1z7F5iBjQHrmnPUeHB9BdgDlj907AOSBbKKKNjKjXbtz86veoUeO5X4
zPUVN1duskzJv5j+z7VO0f1l0zFpQvYpkSlcQ1STK/ZFj1CQtm1wWKI7ZMfDtZDgRJlepbV+6HuJ
pQaklAC9bWt24HqkXMJICZukdvHCsBJjfiURKgT7oSfs5w+xHz912jDuBbS8Ya3uxdYDIAnpZunR
JWX163GKHQaZl5W/DuJfqaV5kbvHQSWoeuSqsbnD8exVgA8MGosKBlpJ+hkozxcxyiItVqJbZ/Ki
DVLIBR5/zDeeoUVfCqjCARMPiDU0cFPp7nYAyXnuExkoimAHdxAGxZJNx+OZ0Y4v1SOpKPx+0B5k
xgMEX/RghaM2UBiPNAQ86gWGQG8z1zLffci1eSqofRCeH4d9PTZ5ffeNzBZ13wRun/BpMBiK6tTm
wLt3yjWXIUd2bmN8SdAh7WNf9yNkM6MS+RiisuO3oza/7rpFkbLGd3ewkid0o+WHOjIu+bUZkLUJ
BCb0BL2JQ96jpVNKActhIhi2vr6aJ8qyF2MK4bG86bSrwWMmn2NJHXIuEX/b/LNfupXNtHt4HjGe
Il52cyLjL3BPrRft7eTBlr76BvpQFfKbkOklEdH5tJeyFIKAwg6PuxvuYhXTCAmMFVsPIk/dhdiz
wi9rfS5nw5oAEzo6qEkLYgToZuo56LCRz3NkZjYZ47Su0jKNNfEbcfjDy0W6eGLxe+cHoBnuXLDo
6LAEJr+sLVrrZDUESmP1SKZxQL8QOEOBu+szkAjPoFFMCHgounQeTACdDI3B7kzOompZW0QXRcIU
H2NLEIsLizMImgrNxUAUp7E9BSmUkiHsiBtK0kXWDk3ReIlATec+n0x9FMnsjr/NFm1C7vBPHyC5
VHRK0XvIbZ/CRN67ZSU4ZY0VVgY4p2KpcWyPEmWXjt+8chIbXCPAQ3Yw0gd+kghObFdkLpUV8Xn1
OAhIPktjtYPjNStszD2v+hSOe93EZPODj+QNdBSio2cuQJph3h1dXKNqKQr4xqj0CC4Q36AGBekq
iv+L2MyLOVNURKMU1gN2ePGYzS1MDxeopzx2epHNcLH1udny14Qp9RU+DfL4lqx/SBvDhFy93Kx5
klaKLkYUSYFB3N+JlUvXj9/qfYq+o2vTi5OirQUss/E8lK9ZYIcvLA1IWV4xVe5o1WWrKUYbjRDM
ad2hEXVL9KftlGdkdHT1dDDCwI6PKeWHNtmKb2pu9Yzdy4Kda5mhCRMlkNZRv8UY9YGmkWBBs1hY
UF50X82hCfJj1c//GHZfmxHq1mTh7oqzwtgTcSTSUISiAb+XZWlYmoeXVIu0MDxJRrLBhkLfeQQ5
izrbHHlLyLmYUpgWfZsneLKoRjveVq+cbmVIm96sqvkUk+gVCyBcrnwxY1n/BPf80BJWhXm4+NXd
acEEDtBm7EsU6psH6N6BWyxgE+MgbDGIlZnHBBx308yJYXVpsuemDXC8HVANkWafCe0ccSVcS1R6
6NGoLD2NetQcWkDrdSwLbJkPKy8FZAoQzuTS+4ApUgCGYqdPEmYcW9USog6AI8RsAYkYdzauRBkh
PaOMy7HgSqRE57Wezd8/vraOWew8C4sMXDsECZgJrcGqqslzP63Ua+ESTRpeBmih9xoX4ntZtIQo
geSnb2Z9gltsBusfdSaHtCfu0Fe/4Q4ttsO1oHwFIMSis2JUhzl4fSHnBVAMEmRGWriDfR2yGxd2
XldDJfy/SQfBaaCL+T1s4WW6FDvbp5PmQY9QkZVgdzwtUZd7YDDH/jxw692goNQi3kjrUwR9B+vF
46RvGqfi5r0kL5tkgFIfbOkW7LVrIDeW4qc6hb4fE11PqfwQCikn2pFUEuzmVf+VU2D9AEe3bR9i
Uc3yZY4oWkaxE6dl1vmG1Jrw/5uA5UqZlc4xvDjAc7yIHjkGCcis3WnVDgX9eB1pjWy5fnDQGu54
LOAlHtzePXuMNktaaWa+iE4lHC1TW7QZTYSDXONdvQdwUp8H/u2k/0X3EgALiT3Z3jBXhc2qWMUf
c6MVe4j2jq8S/Txl/sVZcI4NxNWipxbnRZLxY8I8qBzT2LqOJPA3RjC/CoLuGc1v+4CmQPu7HvjM
iMMwNVu2No2/C3GhmX+4T2HW3ymfv9/oNuUl4Y3iTzIEKTwEqM7sHNbzUSqhvvIL7D4dDX2QBGc3
bGBWl7MeWjJELGpmxQvkX5xYZYGqr5mjwFSrBckBdLVn05wUm8WP/SDI3FSCnUfSQ3JkIaIEF3rL
WQwoBC+gzNLCiL5CkikP1cQ5VBDhtAGHoYWXfQ1Ym4M4akbI9/66eb/T1FTrVViRqZ5B7K7vk9Yt
OuCZ2+ANxLxLWx3xVgDrEVH/orlfPcLM7bguBQVxOoB5VOfUUqVZigB+/uFd34BIa4CSAxZd9+3R
xn7FaSLT4qCdkmCc1jHCfcFmqIrUgvOltHTGzYStVLmSgYhfeXT9OXvOz2LTCccVk54YAg+ryS2H
whLAlHvdGFGnZ6uWM+XY89y8BIUJ4xLBZro/0nFxY49CjpOpuaZh5LaxStbrPtg8H46QaXsUj1h8
qSxnM+TOiqn+bQmbkSO+R4nnh/RuPjSj6Z270Oq4ePIYW+hSLq6noqKknYrijndC8aDiDjdmcTjD
3pX3tUO6pOBnTCN5KGcOjdBvIpgg+kKeViQ9Z2EuVm869YLKPpZOpdEOKlSIjoxq7BGZHShUPeid
BEjNAchyv+SFt5DJfe3+HZWsBEOdBgZvuXRnrjS7P38+VHLE3tsfUmUCcRv9CigmQEft046Z9Zrm
CRDfUDS8tT39r61aplfpx44IxBYdWt6A6pVukFBW2aVD51hOtzNueJ1DorRj3nNuMuA7JFMm7Qfg
mvqhbzVDhh0eC8EH4J/kBS3jOBruul8Teq4kh45Ly+kGpQ95WzABJxBLsmvkb2RgpmyIl4/LaonD
XCrsY7LfoquUkGKbqW+C3HhNl6bbZfYyubE2/Qbu5ru2uEzYDxmzsvXinLoEMtVZi+K+hSO3m5Pk
zwrC+OagC9yr0OM0je3fde+Fdk/CiFkjBN9xAexQYxVie2jbww8g4t9cdrZF8lBGXopMNBzjlmVb
bYhvOzmuTZ/HTtt/ZSeVODmVi42eCUouHKkscRxJvfFdeDODNDM5eJxqscWVAvM+ONojFZhiJISX
3MVuMAV0kLTMc0BTHAtGFZrInppXktCa1HEyUWAXYSrCuhPEDmKCKbRRME8E5Gr25Fb1PsssSjjO
SfZmxnrDy6lEMfv0LZ5wxH0r+bWNe+1MwSYFo62+Hv6Hu8CsrqwPlyDejxUcdrYVL4BxuW4IpsSW
bvIms8U2TX3BLDoEKXGfK19ra97hvVfLYfPAtpdTlVfykXLlqkVvv/I8xykY/BWkouywjcVlVnhU
QgILvxrhN6zNssVzTcLELelGNFvF6avWNiH6G06mhIHUZ0H5vbZY8T0xNGmavDZ3J84UgcsIyd9F
3agpmNriW/04D/2gh+MJCERCYA2u3Zgo4/tDJya1g0fXVuVDNtbQFVPJz9ZgmQ+wRcfnI9TFF4bA
o0JmmORFM8208uQHoCTLQco2VVJJbCLMscXhhE4pxo9iTnRMCX2SKMtdugCr9XEUcbOcbCFDXXHI
Lien4XQowMklyKuOcqKZDsq1irpnpf0VT6b1jbzgmcP/0gxP/Kt0ez3y5J2ygqFLkoM4wQUPMkT9
KwhP+gbE4b6ddUJz8W3F5o8qN2At/TVV3cWFWEHno4s1ozrUq0fr/YDSGmsBqlO/FdW4EIavBvIO
xwLe+vuamkwZK0wue/dUzfczIA8AhxlfxqCIOicZ0kfIZhJBl7Z+QguofNRR2mIg4mesvF7hnTmm
XkkqRFIFD+kpp/1E/q9fzkrVrcb2F+ljs4aB+yRKl1qV+JRD1HuKGRZ+NETSqxvL4i492yr9kIYB
7kpnk+qdMMci9uvIH9FFkb8Ial3GHEQwMfjbzA7HKX5NQvETS8kDukM2Pxl9sFvqCHDZc3eFeq9B
Pc4w4TUZe+x8GTWscQY7NOBXU4uTeAhAYkveLdxMnzwWqUiWwJdUtL+4LS/UvYfjjit5zVEb9efd
VAVNXV0ExiRExw4a+dd8/mnZNFWs3Si6ZZhyQZjgQ8JlxUUblidRfLxVwiC6TvxN5YG196YZyfDA
fHqr9a82pw0DcLFMC+xlCHdU7Zh9W77VdAUUkT1NNObDZAI9jquNbTK2bExUdZgOHMvZph/TCa3Y
Wp5RwK+/R7WVs/YxHai8stAgbxI5WE4lH9/gBISdtzdwH4Sb1SvqMoRFUbSpFIrxCyT9gMnOK1Ao
B40qOjn+RDABA1dMGq2rW359XILAskzb2AnFQPhduVri8Gc4HwgCtANQxYJkM9w+mexg0/EhMbsR
oxqTYQW7qM/VHWwxa2nu2LimYOeCvBjyyW7+coZ5p66VbdU7b4CFnXILAwBmtAAiIWdmH/hui4jK
VCNqU93Dt8yIGzIlygMhhR4GnCpfSlAnObLorCg7vsvxN7NGezf+QAmDFVPTAYlhwgb3UE1AAehf
ry/zFfSfWoUAFg7xc4qIvCaWhOOq4jf0IxV8eC/GS93LKns4z8P2u+R4Qdi8LZIQ2L23liImMspH
9olQDumCehWw8mmWr1F+ClAkqEzCKvcI1jL/GSTxXl/aETKC+soI4OjPgrPaBz3cxHNZoMk0mpcU
TnDck9vaCwvs2V0wp0WWBkEFhMh/QiVBiz/0ytYiuM5PvNlc4Eq3KmObAvswJWvIuzLl5gBLwNhQ
SAGlUdDpp+0pptmMS/qIcOHckDQqV0qlJtLpN2wUQ3VXwOMArIEIm78Y89nMELbMfwgrOf+P6J4W
I0c70VxNJs6TES1ekFBknuItUsRDfPXdAIvzDh4c+ipPzgE3Zs/EDtR5YTmhhPbiQ38srHqG2FWr
rXCwQQ42LRldK4+m+bHw7x8zf+Pml1NnVmxJQHTOhfKdsAZyzz0Ai7OFvOq28HTZ+4LQ4VmUl198
329RV0RfAbyboqHCvlBkr0PHmhhRAsKtsraNNg6awlbt7tDIHpqwZcb7+pRlNB5eiTZNGz4NOrHl
3AAWU9ivjdDw9jd3LBw+eF6URcUTOmZgSWRCbsZC7BgWmiSG1FBFSmPqk0psJTXXQxW5bSQ4AFAR
CQZ7nwg3h2ueALSjH28xXkLRaSZjOkkVK/ZPsGcFyL3WYU+HZTVKANrqdoMc9U7lsQyrd4RDyDm6
5u4MzNKhC8qmN6EkrrwBADOuS39x709Bz6LUhB5RL5L5/N5XT7AZmVAhDP0pLiDB/lpDtvbDDK3N
N/DTQECJRle3KQD8m9vVRrp0deVX92JRxVsbulm4xdvoYdteiyckvNCoVY/POCVy3HpeUymJ1/KJ
GJEY1DZMDpQhZ8hDMKyk6dMG5DyE2PvUKV7PbyFLP3875tUfsp/Dk4n23Znfuo5pacwEtqkhw4to
D/CMPZRXJ6DyWM+GuOfHGik7UJzV+3vxG8OdoWVVfx5FrVsLbqewYWAZkF4v5CknfRRnzTMgfA9U
5Nr16G2iqeFRvtgQPaWfQmz6e3Jk3huV8pVwiCqvL3nWd1Z4Y228QgE9PpFMNX/WZUPaRMRaQ+5q
ChCyfO/ik3c2tZmIg9BAVEP23CosA1vzgMx1wzRy3cCpQg2n1KTkcs88dnCnCnlW69px8+y+lze2
ZB8SZfzmt5d4J3hiwpVPqy+/yvweT/9M/5u0m+0Z1MPM/WdD6D2DAtWPj0idFNQojcWG4gD+41GH
ZftaQc4NiT5UTCBEMOujqgZSCLPk9D4j/G/RYTq7XHcjWh1KTpljObi5VO8LTMlBicJrDaiztjdW
ir2GmOSF5Fu1vN/6NoVDq3FP9MHcgpfqbbGSku2YQQVVKm/PMUghrGqzqpe0kDvxxww2plY6Mx2Z
C27DcnQe/hglkfeq9vLtcMUtSoytmYsNdfAHR0wFPDA+/n3XmcVHSucoXKhy6CbpcEuBlZxb3QRa
QvgAV3MRP+BzBUV454pfo2CBAtSN9i/PgOe+uPCI1c9lqDUMmvnuPDst8WbFIsk32zq0hOfNUURV
mWDL7jyFh3PYqt+XMr86rQ5MF2/GJXJYtng6/nO+IHgqpCiPJ5zkg9dxDb5/yS6PpqhMgaZUH/09
yeMWQ5UQfOw4f0ZStu5779bK+URbdecTZN1Bkc5AIOVqZzd6QUWUiUNwXk1aTSql1/0YVqNOdMK/
RLT2jXD4fn1lLl30sne2bPj2iCgIi3fo9PnJjC8y24J8EZdzirFGg2XSYPeoVUyNMeqGOxlQyZ2G
BHTjnFUg5WtytswR3BWCfvxAQyP2LRJNHpwg17lv5Ll19IqR4hs+cRsMIF/Aav2TQ9GEviPTlMXy
kapdzZU06SuHi4FdL0QlYlrwhBbuxRa1t7w61XgeUpRLcQxBNuhCfnT6gxhMeYDF6f+CZyfLlz/9
7J+ritKEQn53s0wJup7b48wPqylAPaYRCqceqavqCHOkuiU6o2oKKqVe5COu8Cnxt0LJitwj5jFH
dsXZlR3CvuvW2kvcLCqPZ3uam+Nt2dQD/WzASPDAnJtP/6i6rEAYEkjr4Flrnn4DH9sq6M7UXdwO
xWJYCnpG4CBwplXLxI1B7AC+XJo9p8T415bgEJgj3TgWONxxzNHXujZ8PJG9hSeBZS7YN3zPwTH8
L7z/9xyzCeL9G+1qiY+Z5rKXVBsAg1gm7/E3Db52ZFuGw4AVDf9OA5Gt5KNqQh0fj+i7oVdVbxeu
SRcdgvlITm1SzlIre6j6HrfYzVwbywyaY1CTNuBe20kBVnoiDIDiXxl/O7IycszTx/s/MaPutDfN
01YzCOOcLGJCIzsf1Fd+EvYOffDpevQ4zUpVXREO58Y09J+YDSTh54uexNh3GNXsRhTQ1tBT7o7x
Q3ygkYh1jFlxPdpMvoCXNaMKZSDhEbuoZUjzzKDIJEDGXGaLTqXMWoUyp0TJjd7d7RAyaF0x5Ih8
QUYfd+jPbarmKBWlmZaZmGY3JoRTDXi+LYNOTlw9oMAIlaMkgFYnZQKF5i5YfihjIW8kAfigsyTu
Q9jFfMXuAR49ANWIQQi1F5M3GJyY3IqJ+WEurUL1A/RY+UoVeJ3ubfCnkpt3Y4EeNHemMC4Uimhl
r0BobjBaJpBST7+q4BsLXSUCdo2ek0FX4k6qNVuk2VI+uwHpXA5YthZON+MUpTK0Es0haWbQ5xNq
ok2tmzcUtLhv2zcO8b8nDG3GMYsbqfAzno7iB49UwXgoy9lGam9C6iKAk+OXWGFQcJJMNhN5PcD9
mo0xxKKcyQbIhI4LY1LS4X4VcojiKe+126rfYFAhl6Kzr/YHe2YQtv9+gcds/bqoXjFMC8sf5Uu4
TEm+7L51tITaadll42RmT74ZUGvvQTTSRvTLE1QFFuslpcdTo4iV0b+BNd3lWgK0qLqG5qu5W5f2
IY78tFOUyaT1rE/GC6MNiTivh6PypRzihAW+f09Q0/UWOEAC0/SdhIsy8aFT+WEVTPto6VEXFqrO
Hp0YmUuLFk6Hc9+gVg2QfJSrI07pStM5f7XF8K7R+0k0MPc/z53J/BjyFyHLj3Dj1I+jzdgLEOnG
KI+w6saA1/26q1ZV4RbferBjvjJWUAQb3nsNHX44+E7hZBdTJdx1KvTtDyNxB6TQRlqV6WY7EsbZ
asELFu6YaxLG7nPO0uY9uDK/CGkbImpbu6km37djhWGzLtQf5U1nnmAaK1VL31/KHTGLX+x5TPdL
7d+SMfKWHX4Yw9CYx3OAIiHaDAC50BbTyBpkwO1UFOCu+rSwt7846+K8adOBSjtwK3/sScHd7MB2
IruY7FyxF+YSgmy2revvrZVN0+Qu7YeTfZ8K/846t94eCLBHMwwclGGlncvvmZ97pjesnc2b+cM4
+df9Aswz/p5ZNxs5ou73D0juOlqe3JjymH/cG5Lcp/39G3lmPWk4VoBIVUvZB5NOrCnAm0EKJ5Dq
gfkEh6Zb/bHs97xbgt6m1JiZ+ur8J9uJq3XQC833L4K0+HD0uriYju4F4zQMvD6CRHkecMRtFdqv
9Jo0xcxnhl4Yh/Tr+HNtQswnHL3u0bb9MDRWI/RLAH7DIysHf1wshZEjOsoaU7ftVlHFDLUkHToQ
5Y0ISmeWgdH7r977/q/tQsOfyrciWoKSEMV2k46L8ihycwBRlGxACw9lRheEXamth+hND46K3NC4
j0IQkbfuwQfdE7KXrlSmnkI24ztHcm86AcGa2U3/j9gB4R5IfUA1l0EsdZne3AjRpbW/JBUuS2Jg
a6EWIzq4KDoNrKN/tiq6MYW/09a2303pr5TJ+Sn1YzaPzlmqofPbvQM+VnZr7iChty7B0Tejjp8R
pg+exDN7NBzuzAXV12G5+dIq1RpA20/HCQY7aVmyaGHATAEO/vCrRFePS212KSerhifHmDEwAYF4
M5nQ2MyXa+l3WlOClYsdRwDgHG2VVfga7HHSkZWWioFIM7ZhSZNd+Xz/Ic9z9h2N5x3Y1XsaM5xv
xycS9ImVslHUYqRb/cW7BgfXiDEoxt6cj0gn4YmwZd1rR+apHDnIq6OwyLx5XTvuHGE8LtyLN/C6
UqwJNZiERUPmhlb+/B+D1NIwMwP+wPBoTFL0Wgv3mJJYUCOJ0x0VsUp1u3eKIVx1ezkc69c+cdLJ
+d/N+UHh1+VuPwG9F/VrMCsL4SpKXlmw3j7BB0u9CFFcGbDs2T5Sr6mROi2R9Q0AU0LX4jb/rd4c
ujW7dybMq1KMPOQORYxfR4SaCpoY1UqDwjs+ydsczGVijwdWu72JEPODIzA2xBRtG6DTVI8kGqbw
566p++gKiT/OMHr9Nqp6Jp7bEWFQk34oT/dO+rH2HlmbETmoMzPzSXo1CZjOq2SEPpikSHx9UHjO
2/HxDP4//DmqqxqCJn5xx3R42MkqtlMCrCa6FHqfQjs65a3GFHMgZKizh9y2pZL0iZh69arwUp+P
BMTBd+xuQCA2rcA5O3oL+vDFL0OLV90BQBb8QPR8H/3KLel4Puu3cVxcgSS1Oc9hv+Qvo+9Z306N
0QD7cuHk+vjjYMQXM4530gWoUZamPQJDYtWlbThq0HPVHl7iVLPhZ/rUv8+Nl0lbNWYEyOb8blkQ
+m+novoFaynsxDtj8x0pAI/MOwABqGoZqJFxWxMnAL8ZYOGwIw+b0mSdzHveESMLhUPF9Q58lESd
jefR0vVse8o4xGPqcW/w5EAFtXOhhHl7+QCsNWasOTC/PEtlxgIrDD3xaQu9+iN9dB1/0wetTBKe
opTV+G4AjkYaMiJVZdz81mDOQxzN60FqTHKtuzeZE2CctCVhNkDKfxzpjX+mDwAdsJMZ64RfCCDc
6wsDDi/jtIWOlOSNYSicSXMfrBDaPWsV516H+n2vssvXeMG1/eQYA6c84CN7MIx3Vg5m8Gzg6jCv
Ny4AP6cn/ct+RgKQi46xO8Iqwg+39z8DdOIcAGjt+f0Dlza0Ejxbj5qMxNHQkj80i0rP6Or4WxGH
/GdY9jYtdy7GmE/vZrGmljEiRaMtYU/3bK+/v+EvxXMNenIXBwwqY11eyRvXVllVK9Bwp/N4Ayb/
O7BneWc3T2SjgjfGzO60X+NwAgvwtZeL+ZpDR5hEqzC0bu2l5zUZAwBcs1f5n1eRd4qz84ApxGnq
/iF8w980uu6FFBO2Db3UNHrYjkk6DNmyZrPozbfHL3jWOAsVSrqzDLrlgEyO4sBKfW2Bzp7uw+al
lCLJdGuwgBFXGZxib43LfDevaphSS0EataoF2spZYCHUo943JCRFW2iuiAptGNSMcLK+uihwmhlg
8+CV8a60hneDMJmvIYWHj++nI5ZnauQmIZaj0LOtsJR5mAq8/vmuVgkKIdCYF978iP5w2OiN5FQQ
9D7le+HdVd0AxTiul0S39oYR/Xm+zxvBfWn8LK51ocVE38XP9JaVR8F8/Wx7r/foNiwrkCJiEMM1
sa91NxeFTyyzMRrD55pC6HtWlDdje1K+uhkAwPLw1XGxVU21RJJPc5aP7eTXcsUYvE2jXEcpUDCW
qfD1/3yys82omOjwRemiAauGRdzU1AdzXMNix4W4MsFPsXDbsdrDsx7M/9cFNhM6dxcAcwyn1UGO
eJq0z0bjfzKvTmGn8m9PcYAKnl0VHRiGLxwwg4/kXZsrR7RDdgN66Pi2sQPGj84pQqe/q29BO9Xz
CCRfV15+GpfnsoaPWWYQS2SmrphARXS0qznUuI0/LGNwzWV+UVE9mHiuxSS/nWLGnV+2nwwRkvUJ
/o1g37dAnSKZ6GmGa6ccB9gu1w5pg3yYj9Tx1eaYeyRF6nP1IXLL2t9nQwUDoA5O8+qyu/DHiSXl
bzR5IWQmsyHPIBl6gjoiNAqLivo0OYrnCnODzIzFB4T4xggbMhl5tqkHGGCFbTsKb7B8t8koIhiL
1tYmdQIkzayUqpUU4GdunrzgPwKc+0aQRaPnXOCpMtFLNKWLE0tRziKd2QgG7UQEU2U1DCMpPZ4S
POQC7hcOS/x9eTzlCpZ/l8aNKPSiMHkuDYGMOvOpwUCim2kdI7n/mdGABdHegNRhJJeyXEE7V1oU
sDqZA99dQxhDi5QUNWE01H5E0kHTfyenVTjqJpLsMHPfIQ/FiEU2xq9faV0p47ZF4Ur/7GWuWkUe
zsjVkfPxmtQKmNN+1cVYXPZI4/+r0xWlXXrU8XW+6xjKWF8DFGLkuiE0CGl/9cGp4ELwyqK3i3o2
xQBw0BfiQWAiCexzquybXHgwTGR0rw+nFQmtbD+//29iQCt97EuREnPKsaJkV8qPsXDEzUW/IqcE
OJj1sMhNBLyNHKM0obhpsLC8VAJkxm/KjRflKHplqGHTJeUsMYx0G9xoKJ4DS1Mprvf/BGu0IOMx
CTZeJ97DXVxKLem2cGPb7zNoCGOCTX2mgFYtulkQmF/PSCEw3GQf3PyIu4IyFbKOPCGWyTo9Vim2
DahtfS93O7WwBggcZoUxQex+3fktYUUnzVjGBt/1UZSk6ShmN0C/1s2VKej/1/WLeV4ivtR0rGks
R78bYw59AJ2TVi1ClbREohdFk5D8mwuPj7I9wdumHV01Gm5L3QU1FzIu0hZE4MC4aDpYk2xt3++d
fRAl8bXFYIbE2b1R3rcjfnYKeCejWYyJHnaRtP0JJ72KDf0oXifCFrKdM9/KaIOdec1rEmaK7LIY
mNmBom9ekg/WP9ry6Se2tjQ+IQVOV1xIkfw21Y2w1xYRMoWYqzWgChDk91yCfPn6tRCmNBTY8VXN
EP0XdgYs+nbGReYbg86432Xljh6mlptKlObF/R0PQ5QDsb1KS1qlLAyFT89XJOoTJT5GBStpYkRr
FhIFMznLPq806MFjIyh7z538ZL05NevYUCkFCS3eRQr4A6WGgeuxpEGv0ay0zGkPmYvwZECALm5k
l+vqsB1Jv6W0lbn9+o+9r4uFZYLpLY4V/tFc+Z3KfSrEyDVN2CJJ09a+kM+H9X0Q7kjWDZj62eYN
axLSXEisnDDxtxbiaBEshbK8iP0h7q8Og78uotaUdDZYjIqulPXn852uZTBmY86N4QMUIFyxrO97
8nkOQ0hQeHwPXmfwJpCn+/xoF0X2vrIBnZZWjUPac9R0IMbwKMkGN7kXFQ91kczrQtUSk9vPIo18
SSddQu0NBUIvnS892+muGpfoKsCQx1uh0+ZVzAqDF9IYyFB4JF2CmmZFWEj/pvrEWGlkAe3p/Q8C
7UQysd9ukgE+AU4UZ/2LOjb4Bx3OVy93x9aroXBMOVA1We56L64C0d2TzzLWj4Zdy966URJicmkn
Jdrbp06tJQuQLPF62vNbjuVj6hqLKvtRBrh8z2i5k+cjUnaMdWzpobnV8rlftUgxstBA3DSrmH2r
rTjt5hpEadOu6L7GgUsNpNmjczLksK/HcZLQBPnsoHB/LrNNWzZyQDcaxbk6usO5W/8LFmTno4lx
WArmY2zvBsyD9USvmEd6M67zeshIKosMqAy32d54VtrEG+lJ4g/J7j9Uo7i17ckZO4njahCsA7rE
5hi/xN4NMAVBGrK526XN4a7Wy2bJExSWAUYsGAZMduJeIau2TmpeQyoAITFdyvbMEO3G/euR8lVj
vqDixJmTY2LocLErB1fqim8BWTCderjdPVPlF6XZYI2Witcw/nj/aszbl5ciICc7svAbPGzpXrtj
4oJCKWTPE9yokPF1YnPcw5qBZdEu2bp+mazNgZfcUWeaaYOGMcFN8JwZ8xrTuOlKw/IoO9XKjdAQ
FFHKKYEakcspiOmNBQ/hmYFKr3AEtvxa2chfK+1f+e8ce6UsvW8H2/CWBRlca2wa8fEAjtlHcwUm
j3oR+5w9OALGXM8TFGTW7I1RE5+B0TQQa7v612DYdgyKIIIkQ0QlbqQ+fQaEchBTJSNzCeu8pojx
MOOzi6yQvQd8qUCfQCCsdtbZ+KLa8pJnFq6QafPMyagMWAuPKR35cPG+eSz1bmBuNUmbBGrOYPd9
rorB7EdjIuaOxd/tJYoFEtVK0zCrQmTUR60eEpOp4JP2qVlSm/j9q7UQjDFkI2O37SNrHGBpeqM9
twmMiKL/xsCuFQIK64mbtMoOJaw2OrOze6WKpw9dbdGm9OvHoqX6jSik9iEEyxVOa5qXGv8jKQUp
hswwLyiytXfD+dxbOCCu+WL/rNLT4qGNwMvEpJUx3GsO3Tm3eUcSAqo8Scg/KMYd2pRzAjPG1TFy
uTWEpKdLqglvD7BxgaWEvUruf78v4M3apaq1of0U4sqyxMi+Z1D1e80brhxdI93Od973DpEA1czN
HERSRkFee1rSbfzuhMwotSL59tnhqINktqi8+vWgqG6VF2yR8B00eEviS0/MHVS0c2EohAhRFUYE
OKyqIrYmecaQSLWdnfIe3rtfSfF6+E/oTExWlSeb+ymLKQySTHCcpqBifS+cshpZx7XnfSE4gvt6
wUjijXBtdR9AXGGKderMS9et9poFHt2IPGdneSLfC6sfuJc9RHf/MvLyP4Y6acGcnLSLj8W0WP+7
OazCBn4KEwfOsjB37PptCfQTZSF1DMsWGWeGXVZ2scf05L6JWmQey5rjqUwAP3DOqzIj6LUowr8a
3TiVRIKEQjO6e6bUDAkQfz2X8zR1h8Bsw68gF6GO4NsUyvnQl7kz6ixlic4I4NqYMzFrir+MM/yL
9qVanT0LNo2uRwLR5H1ImJQlHKkr1r/yZNFBF0rXUXTq9Xcd4OmvcvoTOnGozomkBzKRcyWpy6X6
dfBczCwVye2MH6/sMOZPiUL90Pr38hfvjSypU6Jw4bEee9zBUZT8HU5Hvd4a3+EgMI5QVI/5V1P4
Gg3/GiW3BW23FGlthEmrNTQfmeaK89uv86SnsYSTSdbdlm0ihwY628f8aupMMibIWHAh6BIB73UL
BLzfYSFBFTljIyAJzm43lZwJ4QQ0k9nFVns1R2XvEQyoI3h8DnZ57nI+848whcLyEI9yzoRwPKEl
PdGEDZt28IXOovs7IduUSMGNntSsnT5bmRSlW3yp70+KdHCi4Ocf6KEhDiSLbBgrPQUf+q+UImA4
HHFrJ2VayVol6Xy55JXAHISS2Q14k6iF32OEK/HG7JjfXoly7YiJeOpTcrp4WwlB0XkcR2AhFe7k
eFRUIkv/Krw7B43ZNGGyiOsyYCpNvEocmM7dlt6HV7jhvVl8Xm+TR/w+K7FMgnU0NNRJ2TW9/e4B
QXBWWeIIkqXeOVeUfrn2Tzc5JXpCYFbeHweVBSLZbfQmt4rPTBOpNDOEpmTSVbpPqe/DNSOhe8b9
jQgyFnLeV3h29e+k5dQFgX7Wi5phZr0r9Av9lobJxvH3PGWch3whqcu+Wnf2db0xsuwusrz6/i8A
dxhQBHb+fMjUcy3tRmDN0vY5i5TV+cZF+djPCF/MxSsFxMvxQ2SGzDAjc4MHqm18qTD1/+6W793h
7QsDslZXrjvLEnpwN03a5WFKBnMlahkvrciwBgfqnrNwW2xfmW8rKGRs7Dk3lpvsk1Xh/YFURBZi
yWlpRh3YnL7Sxi0Zns/ro7TCd2tL1kDinM5Gkmey2Csfo4BEem7DyGID9luDhqymQE2O2gB9f7ZK
mwVPKBIxAabPC0/2ujw0O5UDtrhcLanSwBkBXitj36MEa1wElO8RxZXW44KorFAqoOiPUA5GuBd4
fWEUDP1f8wAljfbRe1bID1Nn2faFNwNT6bEUxOysyd6FR2rqWrdNTxVEvJGLYbTn2WH36Oc5EnEZ
g5DFoMS7zpqWTW9d84Zm989MjPHDuXacWzsODfu2p2KeeXjqlE9WimtQpZ0BAsW2vMp+L2+cUPIN
qtZi7zDi+32bm7yFacnCCcxBLPR64SmedttlCB+Z1WdK2fgTGjMMDBGKhEOxy8YJEwSPRMfr5cos
Qi+PSEuFyCiaPt+3IyiAhoWVu0ZfSsdNAmZcDXef5OgmVMY883gtoGx+VIDlhNI+I16UXGstvMgG
xW+KbYrynoHTVaCMDhv/oxP7wNgyRmZjkScIbtQqA736Db9PT1PESEpGrr/13Mhq5LnzN5WgUuJF
xQ7yyfx3wZts0bikJdlUueRvr1v9Lfo4DHSXVX+uhTxiwHQOjprPaSsOkqj/FOl0uydNFPTku5CL
UmsGZln9USytJ8CTSiHHabx6nCOmxfjCfoKO+M78wfIvaUrRFV8VjfMeWCE1LZ5F9gVsegE8N2DR
pOTrkXQa6wpQaQLqF5fmHB8eWz6aXDlyJKh+dem8sMWEfIcQCkjwzsWMaWFBDSne01HsZ8c7y9QE
5Pdn5CyMGiItQrjFI0BlfSZohw7L1lJJ35PrvL+vaKW/qZLsQ7YUMDq3qZvMQLaZ+TWnK7cNEQkG
4NUaVTY+wnXQJPPXWQvBsc/UhTOd9YcmluvnCm0amNn+aBuSDM82s+ZmtPlP7zEnhMn666AEFH9Y
LMl2UlrvdiOvXfViIwRawbpN5fjyg5uGBO+KthiyB36h8dsIxXCEGaWNogrykXyK89fK510eVxgp
8n2t/iZYLn2O6+PVXVJERJ/vXnFAtuTFTDhFo/kdpYSuM8YOgoY0OoldePMclj1ukx3bROa8T5mP
92o8ZFuC3tCrqsCVZG7ZJJJrXidXJgfTTUQHQA97lNYEWo5vnn0NqqHx2fAxlyDbVAfWD/hR9xMy
5EUKrfqyQAolpGKfUIwe+yU2FetvG3gduBTYVv939UjDosmowUhbJbJfPVWVyL3Q9V5mBq4fc+Us
TJHMe7eCq8Yn+LCCETQ2RPImS3fyHbmsOfo4IQCx1798QsAHOJyORJZUegrij87qTVCZweWVzjZy
PtopAvTKZsZOSPFTxLObG7OEOXwZ6bUxhA74Mj7S9smtlNqMJ6VmrSDEre6m0iY23Pi+gBv5DQ4T
kW8LLTzCDC7fsu3wkrk79n0/jjTIoO5fvsOK209LN41OJtv58gTBrRvBekjTDXku59ANbeJ6bfO4
g2zTi8YP1kQH0rqbc+g6y2HQsOaOSXow/Nd6OTjfE9UwuTKRTZ2dPSF5ggKdo3NT5Z2G+cSo48tc
uYx+iJ6Xl0wZmqD3o13jElwmOcjlpS1FXr59A5hofmBz3e9ZUIni3RE0LVkxa/WpR2PFPrkh8mqr
wIYfLs1dWRYVQ8ZrijWSzQX8YymQj1xTwarakLfgaupxKbUbp1tUTRBFjCn1Nk5l3QblVOL3mYlz
bKb/UAZ2Q9K1tleZRh2zlgN05YaS63bkgoXCVYTnPSlVzqHYgv3aDP2mfubQKQPnyrWevFjD49oZ
4lY28N+IMw4F3J/Gi/HthQ5JW7XDLDAAiWDt2mPgNWFIIboP0m+qXuzcPELc/00+rLrhkSC3gZ4Z
0VhZxuQzOxmoz33UPtjljAsAcnHMCqdxzEt31wssmHzl/b57aItMkiDFrethpr6ap8PkhLbyl70n
UEaAC/P5i715BL0ERE1wzqPjuWleOzUj6+O+o3gcfXojyb7l/FTKRZDpgLilEuqA4AzwJMGdokLE
Wd23TtZ+kZkZk67mQDCbRP2qF1z2r/Sc3tlbJTMPB5jEcvD1jsty7bm8VfB/BFlSPVncc7P1IyXg
P8kTz7ZZlyW1ocwA5xrWYRlYcjeuVK5dTh13c4WQBxC1mg44Wr0i1ICp5Z80HipfFw1Zn/XQKVuD
KtzBvokCvBdXB8wSs/HAvl++uBNG6SlIqGMyUK3citN8BQqgCwtjyjhLOeTcH3O8V64sP/JcrWbZ
2pd9BydHqLySU+lyy2k1WGjaP/jAYEepkqG9vPNgmx68TeTXmfjcst9PEDJrUcu3zHZHqLe4c56O
1kyXJKMrR/iC/KZnEA/D3rZZQVWIUzIogP243rcQTUPH6buojNpgEgehz4DACH3Eg52AEWYthQZs
T6MKssd35yYhUJIZLWNDVNP5mJJyYyBPRatxmJoMwx02DDAdzAIhurF6Pl+LGFJoJo17oyChAW14
Ol8bZea08OoOQKssuthmToCqAJP70P/R6d+NHHLtpjzIzfdteLTs+CqXpc39t1gW43IB883byehr
SeK43izRtMg3jzVX2uok9KHj8GlBIdW2XSTlU8w+cAuaZRsbqXfrQQTBX5zNwRh0JiyySYVepZRj
ZNs2yOXaUvD34SfJdqNPiyYfPzoe9ZxC99Zr4XnVinJU/Y8qpUFl4WPdvUv8LyLwqvE1GNrz2yxz
fVf+NtpyQndTXhY9tkicFrgVQ5+KFLyr0aZ/j+kEhUgQTKW34g1H2ZN/U9qcFwrgn0hZO5ROTVY+
GAlQiuIAid/3pg6K27ROpld4zTmWlERoJvdC4d5Sjw57yMbWvW5g/Z0WHU6+mWsMqcJ0ePd8D5el
ygB04y+trWljb0R4Sg3tFW0gWYukXYl21E+50FVkS1p1EMIwGyIf9ImRuZFDbQVY78ERdRC/w7rv
9a8sf2f1Fbss9W+/mKclul5mNF3MiSehlCrImaM7NGRJTjJYMM0OvDXXH/w3Hsg4shICK9XBFLnK
vC4T+U31ke4vSaRLvuZaD4ebVxPRZqCx3bHgWRP/dc8glIVBCgxrGdziS0nVYOWsCrL4gG/2p6hK
bZCwPK46fCAO+9L0zwz+T8nyLCKsK4R0y3af+518erpM0qHV4oWXB3usEJJB9+jLy/NwWXdEPBwY
E2LZOkG+fRJpb+NoZOPObcl7ZK+anUoj6VYKfWijfSLSqUSIe+a3lIW/ODttx/WkA8NTVQJRg6zK
P2PW/ISYOYaFVLNzEmWL5V0PegMFQCjaZ4G337GmG+wD15ZMa/NJv52b6ts2IjdpgsZ1bzp0ZgPu
zLtGL926T0p+WznZwW9mWHTr7EulAPSH1zDcpvNyhlzHYu4NKZ7JUSOfl138QRA/AWd1sNyzU/D3
/uBGSBndRo75mGbVnRZDKbYeCfOAESGUvEnjH/AhbmsvXFjUXviKemF/jnz5logHalcXKlmyt6++
4bQN3rlCiO1rwzEribr13sxJZYoJeb6gjdH3i6urTFJ//gjKthFWB11W8OtiaH+R5gK3TcBwbnDW
Ns4ecI40dAy4nJkiBy/TtjarDUzOItcVNj9wRJRCMZni7aYKqumax4yzDAFt+CVv96l5o2E21NxS
btMDXQ0hXI4X7LGxUb63V88Y4MJM1Y7NfDnns+zLuyO4dOQxaMSbA2NqcXIlhZkB2Gvtf18UM6Os
nL15InKQPmrr0n73mrcC4xVv7gXIJD+YLTO0p4xecZy9UwIW8ph81DhgQpP+aOn6BNgyrSvxXa2X
V37NmAntm3rr39mynh+Qy7MIzXGjZULg7LN4NHQmfjPA6Nf/Gzjo8192q+EQNoCtIBk7beyhFIt1
PEKNINsPs7krmPprXBuqg+3WNoXwbbk3wwzMygvPhEi2DGud7C6KcFywu6FGngafEaKWisptEPny
FZq0Vje3/ZHfvmPyGCodKnj4/9aIfp232Ucbp4r3gxav+HXHbrAgC57wtOVOR27eX0Nt6EYFA+UO
cHSjKjV4eoVMmLGjX76Ynf8Sc6dnyUvvFU8/N87GExbDTk3233HG3h3z+suZZqtJWkWkZLlRU7Cm
ur09KxjPN3yRSRn7hpLupRc3nXHo8CJM3slUvG2+lPtKXb1SF7QI/QADjEXm3nKH3KjRrVU8hFOj
MwjTNRZCwhbRUOHBVHeRUxqf77QRXoGhA01NReL4ExYACRCe49MZKfQz51OtVFxawb6Jy4FQQ88v
3U2le7scnopr78hFqtjV45K8xivDWBvyqu5ds6/Xmt0OxODNDQdAOziI75586qMObfgcWUbmi5of
qQ9WxSlw14UBN2k7gTE2KJuYpz73LooOuz4Y1mXE/mSxhsWIGt+hfCp4BPhehsBzOETFyIqim9Gk
Pi10bEC/XOg7OO5+ZcPoIFdjJq0LzZHsJR481UsIVRYzNnFcHYiuSY/dXrJR8XyjvCIzWRsPwf3h
ILZMcf4OChrYHHu8Es+2ITL177cz0ETItvDgFXsc0Y6ljufLMhdsSpEhrHzvoUvyaC+YWiXqG5Vc
VFFnCAVGLXiRX9aa4Zzvh5P5tJgd4Y1TKDmjtkkj2S7+R7UwBdmjEwUPCWBUkeJdXBgd3PLLlW0W
/AOryv8eMV4M6omlYnju47RVjNhHJI5Nr9/Ia5zWQpxYGej15ty2KtetzDUtkyEYOa+ccEyOsdhh
WlaGx3znlzDF1+bnQgQWl+3xUF44V2wwDfSjBkh8d8LGzAPyqQ3Aa8WXBuXWUEom1YFybMEmFK73
zqrg87+vQSRw2+z/uFt5UvDIsD33sU1/Ynti3+9FKCtcJUVxLQzMzsu+6hRwJsvry8xFkuJauwU2
O63Ey3p5JTNFeb98MAyI5I5/mRPRAKImVgJBftua0OBA2CBj+cdCl0Mr2hce2cln3upUk1+f2w8A
TN/X/Id2/pvwumBqJWVGjn22qTPyk2ZrNiXxxz/f2y7tmbh5IlpPnb2TLb/nsKLJUP4jHDFBm67S
dPuyEkIW/O70mj2vUSLJ093jhIPkJuMYBRGIqFRUXF/D5CcNBp2nZQuzHqUNBvws7ZZxkEhel/Dy
raBv3GAWEKGCAf2XOYZ8eJqOwgmhHMxDgfPd8DmgtL4jRLhiLLujVrBx/SWG/KV716MHeEQunhfT
8USsm0B400dZia/6llCbn79US5Am3zz7UuD+jdk1YZ41nNBKMocdTpvkus3RqskFgH8UcTSJMYIm
aIahDaoeRCm+41T60aTF2LGWi+nIoVaa1Vanmayqvw92MxzliMqUbtecyVZhVPOC06f78gv6UXWX
gr9S9uBxlcmfzms9wEd7oz/+7SGzzl7WNG43Q0SFhUgHEE16FMuzn7371w+HL9G5zOUok3706WU+
bKEyzKNlEEt0BUJMsjkZRTihWUpWH+M0OlbxPEI/sdQT+xaRmO2cV9PFHyN8wVswFYMb+H2+Iey7
guOCYsFFamsGW5JRz+c2DRmMn+Ms4vLu/2QhkunRjBBI2Cpc6wRNwHoD+J21gvAzZrVUfNGoNXi1
H402qioOm4TOKZsORAk6NyPk5K2sKFM0mx4ewyWn4YZWNR7rhhOBYb/Uhbi3TBjhoC1Olf2M/yH6
gMHTTP/TIAhZsSBr70+ysyWtC776oxxVKXdCMhP6yXd1gMAnz+3eZCQy1J7qHLWilHD2LIDKszUV
LPZVX+UghOnIJWoOQ8w+zAfKWN4zpnaIautvvCqNFgpy23s2n1OZJweE0dAeG2KvZ5XfNvMhvox0
bSMVXTfVBiOpQ4hVfJOa8++kklygqu2PRBnKiBZOCcW5QrRKoMxrpXrjrSFznmp4hB31x1jAqJiJ
ft/2AoQqIfoKmUkkfNWtzwhoM68+ilJ3/VSWpKrgDIsbcDO7wjlGwlw4mo+KHfIfb6YyOVLy1kRZ
Y4qJhBOZfH9/pxdvs5uEsdJpGRV+jA3tQEz2XXKgvxM5UojMUK08ex4o1zRb95tGbe7q5c7dLgC5
MJWacVwZGtwabmxjlo0fRITI0VekZzRjnM3WaVlkPZCLfKpgqBCpuZb/545QoL8gx56lIf3+aVVM
tUL5DbgjMDJwz+H5DA44IpqQXVO35bmzDEmABOcNwf5y1uIcJE6P8zXVVQHjh1ALECt/6PaDCo13
timMId9hB48aoCWpdPsZ6ETJ1bCXyug2CJMnMoamKD+fIPOdyJod1U8y9J9zl5Ecc2VftEdcth6j
Y6QrsrcY9XkJ0SIHdYF0htn87MoMefAq4r7VqbWlJzp8u828f9n5OaEzMn+gQ248VjkjV1A6PZbE
BFuiY6rV3eWYt4jx7p0JVR0vM4tx02LF2Ybqz/Y0BF6oJB9y7lErtkjh9lLuCY1gr7dQbASxtGav
2OMN+5qZTgrGVV8d9397savh5A+uw7E7/++3C4wSp1ZUoLVFRzc/3/3Rq9+XRQ3wPoosrebsUvho
HnjhZNN3lnvLYE2rdR7A/jY02+TQLdeBL1/SBurl37lsekXSlL2SngmER2Dt0i24Whs/MMng545z
xA7DTI7VDg+PSyB38bcYV4kFhWs5zJ77CoDxcQti08cmKY0eorsiKsYzExXqIxn0iIN1K90VmdKr
Sw1c+fKWWrkIyKeriNLJWLW4uTvS8AyVUIGtAwKx7q+uwLeswc7tLeqwvX7SYFTunqMCNK8BP1MG
Vu23VVDSgrJUbTg2EkK/0TIV7OzDDiScFBmwrCw71hr0GUdn5pa1rdVzUXhtEhnG3V0MXJp3aiDa
nO3W59N0NHZQt6QNdtXCcBviDCRmSm6bfFCQF1YV/TCLua/GhBiKcy8CIj57khvXf0zOZ9Xijv4U
RNQtFFIGOpEl2ka3SpkqVb46VC6f3rB0vibc5n+pOxW4yseondH0Az/pH84D8Yw1g5hFc23YjLDO
abtJwp3HZAOz0aD27QPBeyTSbnGm+2BmTddF3Sv39liKfuVI3/rGuhYtvcWyTR8MYkm0QnUshe5u
sabOn3P/0rvPaD4cgfnh2jA6SJK0VOzLAyH3S+FQ81b6CZz48l/ujO4UTSMW4t4TtJvOQ56frHQZ
Om0zPB5BjGihuKwmvcu5q/Xse/po0Orvtx5rCZAF19etTud1bMxI6JxRx+gh7tUAR1lGVMFpgANY
do/klx3K4d9E9tr3gq6+1CrcQWMtTFoxAjda9u+Oq9BW5ufgh5OknSbK5gizVhc9HmOHPVB0ZhKF
8dMRtnoKGkTmGmpAzG5WVVN9kdulFuNg3v4JtlgGIFgJx8pDp0BL+DhIt8V7/rvIaDG53QzOl/qZ
qbPtOx64EZ12gkG+x0bqQhELexmFsn5n849gf8yG/yaUXXJslCctF4qGyuJbAKHjqY6/Jw0Z9KCV
dzwrZis/HnIhLok+shsVxblOAMkqd7/t0MeRpe44KDxYeTj4KhlPh4+8v2CRX5U+l0jvA37yx4aZ
z+IAzoU/loSDz8W1WYmhzKcSsh6TGBktYD62Y5nonYIUSFpe91DDmAjctWVsLtYFR4o8CfgSf6Oe
V1Bu782yHaLyM5Wog+d24T5JQjFXeEtFoRXKDFWs359s9X2qFys4QR+dNfvTtuomLeneu3xaZc4u
ys+0n+LvCaKuIdsPKKlYWSTlfnh1KXrTnFHIZ8Zh2tyrvJI32UtK+cH8/f+2a35hzr1rrb4tJjj/
4NrtoGIrJJCVK097wi6rkVz44VHy6W/4xRrqQY8Op2qv5S26YmlTa5EvR5YfIZ9LXYo8mVDmJNn1
/gr/VOW+xRUK+sUb0t4kQXvswEgFNc43otkx6A2+eNiME5Up4NvuLDNH0A5Nh4SIOBYI88WUYkdu
tOFf52yuzUt8qNY23+T2trTQKYqPtmnM7nQGdMQrzJHjsrVwAGdykUu+bupyabS5DQwjCNVqjc75
oCLyyj8Ux68aPD36IJgiuJ/eWgERMwDs8M4u1qUPYQJTMsrZGZdbT42GG5F1SS1Y+rOglUgXRaqA
Eipl5CJqNbEUSSY+8tGNoZ9kRmgNK4KiZsiUsTYz72HvdM3TBGFjllLIAu0S1biEXUt0RppG43C/
V0wmCvt6G8Ah/MuBoMniwOP6W1ZujfQIb2ojfLrVOAJz6u0ELXmqF+JV8l/jCIcG2VIE4eH5d0kl
0gy4Hg9nphEYV6YTnteCHKCoq2AO7iA9EGANx8mVhv0ARyMC+iCDRElyRiNPfJKKz694ssFmaAUv
18pX/aw7xL4Hwqlqr/ZWZwCEd6YEqqbWYipfGXhQzmrFD7IrWAVMaiojEkWHizX0ZZblvIzyCoV9
d7M+YS34JSncN2GKibOIKh2sB4sgL55iYOgZDBOJXsBmlGYu/8fXqBGQiISGqaVMjMed6YaRogA/
/rSRTe/zdKYkyk51/rB7OsmgwUI4jbllu/KCwD82ZrfyYb9hVvo3VBYshqKOeAPKaoyTXMgiHxTV
hjmNcL3owGv6X5ZuSyJZgc9GVGtE29Xd8Vu9ZSZEUsn9vSCOTapOKGelG1L5Clh6jX/DB1Nt1mY1
Y4YE7OSSjpZ493rAz1iL8Rcel9tVp/a0d/dd034VbOAwwJvIGQdo4EMLnvt3nUwOA2xVKkAwC0Yy
JOLeZKWApgr+bPG3bUfvxpxFHhW117lZ5FxGy9s23Y80xsJjpwSb/Cpe9NwbYm4tD3IptHJ4RX3T
GL+W8USf9oHkhD6xKCeEuO9zG1PmBxqpNuPm+4hqQtvhe5ovK4whRGOpfG5w0ljYziGpPw8uTcmc
zXeUmmE1ONjnlFRdErOV9YaEw6HIScWDsCmmNw88V6hKFswhRtVxzszl3K1Fi5COriN1TxTVgcdo
s0A8G9bIx3KrtYAj4aZQz1lkwgG19/DCDYxl0oj4i5/6iqIq5ruOOBc3sUlT4WOSaw5ZXDpigFVK
SkpKV3SCii5AdEUwrvs+yU1MhLJkS3ZeSwDulr/JQ7Fw6LYAbw5Slf1/HWWj/7bWbKyrOSObvnsB
d+dF3xsZBYFoU4mHuO6vzyXSIZQ4eaivtzrGlIg8jryVuDNbl7nS2lUdOr0iT1XADnw+Qyvm8Fze
oO1LKsuEO4d5ff7OYEMF9yC3F6PQ+vJmalVjkjTFFCqdC78atAk4eGpSASu0Wxdp7Oxcl28zfPxm
KrveDdWnsgXlJeG2P1Sw+Oa7/CAOdk854Hwy6ozYfjmHFPsjsPL1trbwJYTwA+JAGz49acYmSOqi
fS8FG31JtBgvPbaCro7wNC2YmfE8TgYFyPO08EZDx4gvnA2H0g3EdM65H0ZxC7KPCO4FOXsT2dJg
l5Gqc5WCULjYYpLl0lzlnMZmeCVnnQLlY0vvktGuQmuyXByNK0T3bk2cD1XR2WyLtjDjt17ykrCg
lmsiGpHG/b3DdeBEZkI8TqlsNnenR9H33ZuQAqItsmRP2yIaLM+rfifGRi6zS2qA90yXHZQPbXOp
cnZTWCkXXM5lgcypwiHznH1Cr9HSXHjx0Ir4aC/6dz8iAhmKAyijIhBHloea4sK14fabtKfV+pb0
/5wnPK7QKzpGNdaPI2MYMNsBduGG5/Y0+AcbQe6lslU3zH3P3kcMsda168vf3vZjX6em/E3QzVxc
yvOMj6K8o193DQ6FOmRZA9ESPkPXJ0D3jmrbqbVWCyfeMy5vePS4D8othTvtn+KQMfWGVhgFHsBG
/Zfaz1MnW88sETtUNrJMPTGScBPnY0wouLDmo9h6UVQluSNbLi/AyN3iIFUg4CxTOVEpJ/xY+5t1
fZ+KkLJunBYq4DgQcVnw3JaNZ0mJdJm+mGjbXmeUYCE+qnzSZuL10Wc/Erq6569VcPfXEXd1bCdi
Lzn0Yftgq0IAMwLTLbGnZLpgx10e+DF5vix+oAJqAJLGUnVGlBFhW30248K6xCY5M3fAK2S2UJd1
Q8C3lU30kvB2DT3dBbDs0k5cr+fChdeFMxS0YhqskKR4H0zQgdDVJidn4aY3tm+egU4scQ/fUnEF
/oxZOzR2fuG1AfPJJ4MA9ygvKUEgaPATbLhflD9uMtlb8wGEBMoepJo+S4Gs2DCuXYYZkI8myN3o
4NE1mYnGM4W+nup2zFKuwn465y5jhTrGhzM76abMyZr0XrEvII5eYs/G9cfClq/Y09iSeKyL/qBt
5tGmrtPdL0mkN4vqphDZu9WoHFPE1gnvYQHVCToqWWGwwQGoo/2re7Mrd/GTp1jiSBvis4xu0zJX
/LXLUY2WPu1ASbd/ieM3z19Y4mLG4KQ5tiIqlL88KL6wh8dztBbK41fxnjiHb7S+Y1GF8Qaio9y7
VB2t8j8DGO3a3tsR9HgIulPZVCHF3GFGJEvtUXzvYlT5ZumSZnyZyvn1sXV35Zuw4asMeSlDFppr
SnD4JGcG2Rt4lsNm6ofNlODCg1/D4m/eVj+pKCgFFQiZB3jnxfmiAgmebW+1qW2/vh2/01Vqo0ZF
ORDXH9ydit96NtuesPOtCi1AVHFxph0v0O4hD0L+hikwjtkMkpboXP4+P5Cv8hCROTggj0jE+j1L
Wf2x73qQeCLgRDj7LdsIX1pCXbjDq5VrLO6rqrVr6k2xhwKzTYZvwb76HO5qeKqNd9VS76JG0433
nc/AuJ6lOIOb4s5DiQyFCzfJI+vfrs/BWpzMv+wzjtPi4w9o9uiogPpgv7uT89anOjeU9PhElQZO
Mqp2hOukUxxWdNo2MndzBA7KqHE9tPe/CtSBKT/0oua1yAOmt9DZTUCdqMfuyOZQK3HAqzbwRQZy
xaCJQQwstaeTYYUkMj9bBs951b44uKE3qdWKTZgGsyIdgorLwYFvnnP5InfAXrRJ2x3SWFgQToJo
1syhHBGKaQ/XtTC2r9l0yDdynhskLzcHoryvMbqzHnoy4aV98/zaKu+FO4f0db7G5OQhpAQgrV4f
ZsUFMJu0eJrDjnTQRgQ8yQZ0Mop3kTZOUZaO+/sl7dKQOr1nTVpIZmaHOh5psnxYL/La3jdItQaw
sPBoyVYIx3ibfQE432k+liBNe/BW9+TTVHqzOqr32PcJWqnXRECGxMB2cqN4iypLSLb5yYWLcgwQ
pRqqEStCYq1OrIDX2CNADaBahYZnZ9B++uxYZd2rJHaz4Z1M9ht7Mjw98L1Y1oeJ6RZrkUkxBNTB
xjLRQjit0UJ2xwfxW6pVT2pReZbYdsYBp9v5X10pQTxFv2Xrt70lhymi8zh2dqgAnlCPT1n6+SIi
BWpr6LwJA+of1AzN5KzyuVnLLK9DLd4/m50wHDyL0OfVTDVAJP5P2ObGafs2Q6otyF5UMJLUvhEX
zxJeWFfYh/INIKpQ2PuTHWa1dRWcRQiARqrDG5xXUMXhM6XjN+qyAb/HuU/NcMprSWmWQOG5wcBh
q2qsRgjOizahv+DyMYTyKdaAcWJfPHcIxkjro2OWD8V/jgLSqG7pCe3l14nXJs0fYN1nvShGCiwC
R1WOIk5yLGO/Rpeq0qQyWQYSOaJNvzcAt9DXAaWbguOP+5B3E0jWwi8VJqmrp0Gblmx/C+anXulw
OIPM70Gcy8mkYr0I4lp0QKk+R27B2rWoAet3t4XB51HKuMqgP/HPiw5SbJ66wBZd16TCOZA5l75u
MejB5QzbEdpJ9Eq6T21Wb5RgKsbDridauCHZDYXkiEMMRf3gCiyJzH/JDrPXtosCuNRmJ/FyeVQp
fKf35DcicXY0wSa0dqVaRTZbwfiNOK5eXkBRFh3Vwr88WxGOHyjw3qvUfXUyNinSMTyPhM5FqQqP
gNtP3C91GtQDCA66XKaWh/eqqe1Z1BtPu/azw7uwa5d6vP1aD2R/8fOwUr3SYkyoEQcLHGFFLLvx
QBo0jhuqHm1wnIM0nsDNMMIThucHxXAiqILDm8bmlyWpYnBnN8iWav5DNN+Gybtrq3ttl03S8Eti
6g8msI2u5d+dQ6A/gyb+IvTEbWRjVQSXxGa+XXV6qGTtTT5RHfU5IgJeBXMF9AqfsaQLkU/ikRke
KlO8empRiTjmRE9CI1NApt0WMkb7LTtemkPaaUyR+qsAv+yUploXvET9Z0LbymYbyNbp/h1NfiP5
Ti+Pq9y7hd2bAc3oPKGhce6KrHYPuwL+HATbf+6mys9G9Wc7ZQQReTAbl+xX3B7XQsSKq1PTTGC2
vmnWSCgd8WeVYmDwoxWv8Y6tdU2PvrDCmsyyHaxXgnULE4ACyt0BcaI3+PwCX2WQRKwEKuGKk137
iRLqdAQbs834rB8MhWQAS/qWlWzwDYVKp6ji24QtwhPnwdQq2B2awrSlR0uouYht7lWOaw8KvNov
vw2hNkhQ3NvGxrwvmkr6pz+JTFRbuyMDXT5GO3qTYlAK3plDBomBBghYjN9JdNof81CgpgEyIkIx
r0hla4/gK3vJaFeTYsyCfaLlbUID3D86daqtLeopntikIsQzWaqwkSRrSiikMYC0SFQ7k30gG3sb
mSq2qlhHNFh9bM6I4cmKQH+r9Myl4NmJlkxEGD7tP12fDs7HrRAOpwbNXq98YYQ6qJ3MGGB9ELb3
4ve6xfYWSrqsrOVPedhKcqCZKe/qZ6t03TxMpF8oMevVmkui/kMUqieKzKuLEpW3lbmkoEWk9h1H
IwSSPFrjrIL6m6N5LTCtapHMC/4rM+HM5LgjreOOY/7JKo1PqeYOBAaDEcdcrTWXluAktdelsLba
GubRlZBr7YtHG00EgSsrL9IfKLdfq0PWc3lTzRlYWec/MLhu8Bvtgw5Q16pSDlpbKL8ehqUzhLdq
2GEH/WZsO4ZzDA6zG7MWDAAgj0qjwctdaylNeDZQeb0dRsZEGq2RorJMsdd8ySXSfNb5Z6IO1kA+
kvAEMZu2juLK1AxxdVp43+mbLsvyvPLVPJiRJAYHymNXvEbYx+2P9wgNFop4d5GRRA2a+TMpkX3I
dBlUZDsn7ui2Aes+Avb6cJB71FtGDTOFnvuiPSDXUO5ULnWHDGu6z/RmI715cW0Q3kS2QOh1c8GW
Th/IYm7JUPOvbdWpfkhkHWebgNxA30Fc3QbsIpAXP8nqa4WnUMktB5gmriBlhBExF2FpfBmPbgY3
uLr1N11zBM2zHpzaGXlXTcmkQLe8INQxbJGvaTQhKf6FRslI+RlyXXCphSLOJJT8UQYNGWQzrJzp
n+zVwS41B+6a1D0D5FXSgX5+W11mHFjdP5/gZZSajPWEKnm4U7UpTFY2onU4TVXFImDIuEhb199K
3/+0S7eqPMEn1QQHbrfq/JUex56E8if+OY+vc5NRGzbGWzByT+Jh1oK/0vXGwGKScOW8d27DekSm
pGCKYGex1LTciM5UVs8MaHvUGYsjdQUZ4HpSqfU/0/vVYkcVFbR2c1AgkMmrgIrlEn5QpKI/mwna
sEcDyDFRvVr/iTZaMc3K//NabIiXQ00bhj5HkuTc7jPpKOrr3IuQi+5xGe29Dv9i4Eoy1G8Zh9re
QXSoVURZl6RhU5Zo0ib1wkO1AawNrA7qoTLiY4uSSSTGYP0aCrtsPSt/yKIyom55JordQp5y4Vq2
r48/9brbyHp3KU5CY9CvUh9QN6W/dG28uS5d0YkMMvD55vqJEngVd43HEcbVWRQOKoGayfBKGLlx
OPOexNbRrIcJhjQfsc9EwK9f2yahGrO+B3UOeCXSQTtICVpj9R9Zn01b5kr6Ko8sbHgJcghcVkzy
uDGFsbL6tP7pfqLVJmCQXug6fyhgVoTxq872kAZdfiK/J3Vsvfj5vboLgp12RDRZU90ZMPxFhmBa
jQ0dB01WRJeGE8sAIatpqeemUaFg5ZXohDRORxgheSYz/gvP36mhdxXvDtX/jhtLWXlfJ7HCErr8
Ossd55rEo50yMk51dgygizRPxSBDbO2/AcG0bYmVSG5ndWRGDnUAhG4tw04It1A9FAcwEibzUJqq
HgcCHUEzikvYVvB9QW/FycEQ8KhbLmShIYw6IE+nizh5/oTWwqcd4pYT4Jk/wEmDi42J9TkPMk8n
I6P6ru9mCaGndwKtwlHrhNWFgyqGb08LzlvjwILF4q6IX7y1HGY3IageBDLJF7j9CLUwjWdYPMJr
+v0I4m8xR1ustRUdzkdZHBdKkSqHs3zvD31Y5Wis/ZjZS7PqCPH+x0Lo1zZis+RY8XWxq3Xx4lfL
ItNUs4UinxntDtgcYlxuDQAG2ABUtssC/LIupSgcJ4R02TMpsl8nIyJqiFlICQoxq5PO1Hlpqd/S
xIKGZ8pox8w+j11M2sdhOZUFW3KcTkIZ7qIijpQNQ8Tr0McRU1iKrJa+pGnbg6VrNbJ1gjqg3FuF
5c35nXm81wjRlVmwuIvCdE62AonLjiLyCXX8qdVtNpbf+HXGBuAuV5UkNLNFHYGHc2bZhfJHohAj
RjpVddPzpHjPHs2PLPLC0eTJXGA2QSIwqMzByuoq3soubbs0EDD6I5CdWbhnRxpsBDFbwlstZ6GY
ijtNbw5kK1DkiITyDEd2tHk6pX0SXrYSoXqwXHbqPkqZDRH/3H/qtBG2wVMMAWpz8nCIz9gj3Uy4
49TFvo2oHGvh5GEwNxjlNpfNpUUiulk/xHifLrCp63G/sIORGEx972MAUwrVbu2mcV8Db2AO1UXs
G2wAsVPTwAGMl33baAKb+1QKXhNeNuCvxvfbDRotZttlZL9g+b83GtYHthzbb2/0mWvnGI14ihjP
1RzRub4juMMdEwwZtQHeykW8AK7CIefsCf0IjVdLvArY0rgaZ/TcKJIB8CMVVklIcqzVM5TbWvXk
7nDSoAfCWlFOc7sVqxQjHnRvTBSmJrl10N5uWh5G+gj6POS/LNiCCannd5np9vqpkodSeMpDIHm/
id5gV7N/BCU9n69XyyxW3P2EcL1hlYeLb+ouG4SPuruyRniPt9SnfIUMR4WHT1R0OTtH1TaATxx/
AqKXxYD/m8RhOuo1oWbTtA+H0R0C2DmcUFK1GIf0oTjb/Tnsz32y4QUWgKr4I+xxT6oMsFKYlrQ2
TeyxZJSnk27xz1R+S4LRWSIGv7XSBzXRVWshV9n9DZ9wIBi7bU7fCnGfshKvh7vFtYgaFmgZrFSa
M09ieV+zgd90dRqwo9s1TcMMrMVblJWNm1p9wJJgw1I68NY21C7cmctY9rmGMXGy1GTmaKOcOg0K
gUXUg1IhR1WEIKIIRRs/ytGtbhz0B08vo6W9DAwZw3cOKc0BJWAnZjwIuxGLSj2RZDSURCW/k2bQ
bw5myPMPO7EAQqowuy5WPZIZbTIAqGU6bcUW6a/EhAS6LEGqfryod+8WDLhau3QU6iAN+eKGu3y3
6gXzmCymKxLZHYjb2DeqrgDRQ+CoCxF8TeOdnKpCv7mgC9p7wFcUQdFIftLOYctcF9BrDpsUKExH
giEquLR6lOwiGlXybXkqE6AW8dJnldqlwTHoC9mBh4oo7KRB6xiXJyEEERkC/FhFt+89XHbkgvNW
UpRHYNeks2Bu0QQQJRJrpEl+NNvc81+RiVs9FTSmtsSco6HVibYzhvnBop3mTL58kUnl1p519TKw
eUdg/Qr9nnsD9hlifY0akSyd82jP4xFwVBiG+1J/8YzIzfZBCo1vpE1l0QyXLb6ci2uD6wVdLCLp
rJu5NQTFbXkgRK/QfnevWSVCHKANhgnQx7TV33P6BKvivI31kImGXQCqtREidJ3mfajm+UzDFZUd
68146alkKO2EhBEcQFlDrzXcFFdIjKnFkTL6ZwQS6n2Ip/mfs4DVFTWZomXrLKHYMa7D9IL5fr6R
35Ch8EE/5Z0svBIshEAsP6gFUhv6kAyc85wAF83bZcjBcs13f2+l0Tf204t7YYIwPd5lqjBDVXq6
oh2Onj7qlGoYmAh+676JV5dWwbAcsrjo27R0QLx9Xbs0qo0EEsPJNAjmPzuqQS66STs1rfUi+b0O
Qn1Zk3KS3AfZRbo1wgUxBqVAo4/M3LLiMymfWXEYeDP7d0thyvfOaRmfdxQQLrwvE91zMO5Bjv0U
JXd8flb6TiZ/cWd58Vw/Je1z3JhwxQuOHrt4ipOfJVpaZT2xz649MS0VDe3CN1Y1KbEwhchcKmJd
UPhcJWY1LZa8hHYo6V3D0pOZ0APXNk22p64AhLXaOpuGuM8I0bzEZOtAluRu4JUPF7NI39N6hbmW
7MuX7vef7uvUevyXGo2xXObaAIn+9RcPnRXRKeNmvkGOO0h4zFDue0PoH17DNa1I+8RdBZo9LRyz
0o7VmfB3f+5KPxOwEIQYze1vh4lv2g+L0d/MrUw4CGybJqfpbTiqrwUjMwj/2N5K0eSKPY5dKfEe
qI8wfhm/BAthjlDz43Nw5pCm3pzttmdX/qM/+9m/WLeuRhtyXZTA3CH0gaOLZfhmJgz7z4H904rN
VCeDW/mjiANsDnP7Zb5I3F2tS2I81KOfLzVgzJLhZoSjKTfGHnSpP3lZ+zquo8xh6F2ZcVKproxB
Ibh7PQwvrQieoCByU6pFt8Pg53rY7H52FfNd0aUUwTVW3t65v+7nc9JgsRZi3tZKatFh9lLG9Xqt
s7O8RfmDxEOT57IxBIf6+7nCMONs5jc8M+Opfujj5lcUIC3QR28Th0JO0nwsYExW2RSdA/yB+mbX
EWw7Bhdcj1TAzIDONvuQR6Vt+1Ts/yYR8r269Y/UuX8h2C38aP6LEqxc4jsA0C2oK45Qmh4yhtZ1
6INo41zgoZXxchm+1555NJ7TaPHtmeXWkPxUEB6eMNmMxhqB28L2a2uvyT8EG69bf4i7sMNy8n97
hUb3frX6v+4KTTp2UbYKe0905xQdEeXlMyVAo7u8+mC0jo3D30lmPAUOwl4M3plrS8WwZMQlk8mc
Dcmds46nNezkrPKCfCxFaz75k+ZIvwvtptTJCVQ/AGEZiNqr/0basJ1o5RPWJP3DzbPYo6uNQe+L
QgKiLPD7GhVPKVYqMIGLBEPUNBZQw74HqvYLthPTwkxq11GUEip10D6Pa3CSd58HA6tYdb/KAWq3
srbG6Z5Rial+mXyMLlMBzsNSQ4+lKCdf9vZENIb8GNPzzGKMdRhyVmsmSlJYd4LOvuDHA7AghTRe
cEY6q8+CyAaIqpKYVjjGyVE9kAzBAMUxX/kssCo5wwnmsSRM6dN/AEEzXjntKpq2Xin70H8Poqdb
4dvq6/vxibrtOmTdDqbU/4AKJXgji9DIE++Ngq+zGPSn+Rg9G2ceXVAhNiSFVg3pcww4Y9zABEV0
l30zQqCz1jysvW72TEdzwxlkpvX/vBztpnfWNpQojLZ5EvffU8oYAlbQQR+rqqiJ6eNdM3nZ055n
/SAZJ86Uz+lx1m042cCLNmt4ygwf9vAse5ezpjLbpqYrrNW5aHd8nCA6bBvOFSQaKWFEWfUcFpc0
qpz94bKcxp7aR12BpkhAHhuTBdUOfj+tW541X9kN6mPYrCWBpL9yK4vZhfC9JWc19K4J3NRMQdeQ
iq6N0S4fy23wa0ANKDJePHe7iWuNeUhFXrpNGeYDNH7sUfC6kGM4nv++w9OdnE1dPAKg8DSqS8wa
Ng+8XAn8mRHfRyplKMTPHqlb/4tV0gwWt5UJHYJnaYFkP6TLhJuRjXjqa7GhXQloYsbZx1tf9G8o
h433YmV8eUD8DYraqhvgUa9f2KLlgIto9st6LwCYlhFF2JVFbhRtUDJrrz2aPwRipu79NCYheIc3
ax28zjjJNojpEN5anrhN3H6CHMPmZamZZRMT6SipfX3q6Rjmmq+efULM1NzFPAvp4ayG+FuLu1QK
l7ITHg4+3hP1tfKZ4xRtq1QnTyscv9IWPhZ5ccay/MKgWkyEBsbvqvRNuBJoRQJl/Y+JhNVTTCB8
81F2ghGN12puPEqqA8vTqKmAlIc6X27FPkVQ/0RG6PlQiwGB10JKecub7W54aasuvVclhCP+fuY9
oGttjH6NCkCAESbHNW4dDe/A1DwHyWT9/hOehCgQtKecDMaSJN8kYluQu5HaECDX8LOg2/FSw1hn
OkU3o4nNilkC0ppc4gRuBDvmfwklUEZDggXCPfI/EnZDgquKNGdV+bGRXNiiCXCtugWqXN5jwIMj
PBKEf/a3iS0BwqG4CLYcdJG32mLz+Rd1xBXo4RV0uqJF+tj6sZ3MIV+ztykMl0DaWFE6vJl+49oK
XJVFnPk56gqspc+uqfWy/Wi1B0P0Ng4YIMUD93rPSgR+WzZPc4RZZj13vsW8yqRNgfGs27VeGOAV
YFIBFYWqVs9Bdl5mk2Q+b0EVCkz5irjxzm4rw3wa41RkH3LXpviXDqdWj6rVUjw2tzOMaywACcoS
nGKO2sZRxIQnLMCW8r4zENXwz50ZK0DZ5lfipAm6YCxef2d9JW+d8psjfOjHpo9auCQBJBXNI6U3
26GFJHn01gl8OP2vr3LCOn0ytIAvo/UlJZVsno4NpHOidpGw0YPxY9Z53MN2nSJDWzDIAg0rF+ce
0eBLrLkVxDuBYeGJ2Wz5zJ3M25jagxP9jpUyJowfwG6eZemOtwCVsToJI5jOs9nDnPcnHmLoh+a1
7h2D9KzdZfVv96dPDupVLzhwTud54adPovx7gM4lO95TadTvxxVuxEoQwgoCd/WwgAFmFkjsj37x
OlnNkz9RgGY4qGqM2Zzk8SQ2q+E7AtKliqMn6SjcWtaqRDhWmojSewtyLV9/9NkxFqabHix34ERZ
wbO8VWwGL2Pgk4ZslQGaoDBIOhBjic/UC/6RCbRJ4Tbr4mehisNALJoSMQxvvbi0BXr5YmEcbcAd
XPkhe/QbKFZpOK1/O2Zw6LgLJZXrZnk5HRdhUWvLPseOG+YfNBgCY74gNmc8iD7RVcrtOB9Nwpvu
PEYH13pDL86yGXVd7dhZdFVb6pQkV7BMnsjRzPdvX4ie2eRVSFcQ8DBUxEmTUgYElXy9Vfje2CCv
NccpBoUP1umpcB5M7u0srQBzg50YXODVH/mNi0FH1D3s6/79K0L0NhQv6QVG4TL16y+tzfXHApBZ
25N4X/zBsCFZLhugT1Q5Q/6AgapPUH4k11i6iaEPkLAAlLvGQ3xnyG/zxjmPl1BbGBnya+zlrDUF
BEjHlHFDhN7F4IVAMdTmXbX5q1LJXy7Fw/Bf6VJmwSYkn3ThyGZ7y+p8M7FmlqJuMtqRuh7mHj+e
6uaGapoI4bGF1gY37HsaGim5KBpmwraVjLJoCyIzfJc7LtC17oRm26lSxqcpvh+TwoBSL9ZkDZ9V
bk3JjbaQ0Bvr1REYWMVP+/br1PwOqe1U0J56EncpQxmJimw4jej388bWzjKafPkgNtNmjjEJaaVI
2d29KEAvEeIDTwSQKhn3iPqwjgUcVkCigzVU7wN6NNXC+SHXryCxzv0+b2y4RxT+YDGS3MZN1sBH
rPXVpXXg7A4eiNl7Sp+HLIo0v3OF1gnSa8JnrKweOwWoaaY9H3niRm4niD9phENHP9mJJ3v7e8Yu
cgzLj5HenG9QEiF6rovVmDlovd433FMz+uo2k76f3QqKg0hiBBmHHmQZiLSG5ZN25I/PIU6+9fdZ
gDTImwD9Nl7Nkn6RrgCJBIwQTF+g/hRViKtZ526fb0qWR9fV0qOkncdd4TNRYdLCPts1OlnvGGWc
79dOp//L+s+vJ82LxevUDjbjKytBHDryzRI13nigBOgf3f1JbwmAadPDt+BA4cqiym640Gy2tleA
rKg8PX6JqZgywOEDlBJpCH2SrC7Amn2omWnLz8gJQY/DdDqGP2oFGDMg7HDVt/kI2DCSpV0ZWK4r
53inoakM44hvgyLQmvlnAG7EVDSOj4JdxALZSrvgr6GTTwPXzH6j/9xZ48U5mP2qkInxc22toJYy
IcMi/RjH6qUm9NKyhGBgSnKTZbckv0nYkAu6NWiMmISyfMF78S1Rs8ghoEAGaYxhhyqeVECBL3Yq
BH2xZViUKg5wRjyt8UCpQBoZdfOfSP8dcSmYnYL/ySXAXG/FXn3Vf/HxfduMjWdCdqalRYt1Igrd
l+J92WGuK3e3/MNmeAGX4fJQ8lcNeB0Cvakx0/IASqW4W9JFM9/HLqiq8MvRJGxzY0Nr94dNlCgV
Itq4po9qyApEmM0o12BzNkx3MPz3lJNwepQRp+8d/ghwtiQBdo+cNAbBIavp3ckb0w4uqAO/r28m
nT0sFGTNcoSwsUw19MvDcClaut8+s2IzrGvcxyLKoueflSXxSyudESGB4FNhyDIQ3wmpMK1S3cEe
cAFukf7dqO1Tsy2jo2O5kNclPeYeTKPIyTdNa8aIaFH/bT0/r3SBxUqfEnSb1L+c7DR55DjJ7HdJ
uwiaCklvy55gSUg8SV5TaffsVgbBQsyGzsYuNy2uzhlfC9PYbsXyULJppkcPsptK90WETY/N21gc
2Pz78oByv1LGxOsxPowHix4d7enNoG1faeKIooYyRctuVKmUq42694snCOayYpBggAYJWS1KsCgj
AvDTmBjdAnKSwK362kq31TJZzNp8Hc0kjQobLSOuaHBym5iKy+sy9pq4J4nbbS+YNCxuySM2w4/N
HcX8eY8L3Y13AObJuKF/IRdLhTWyOFXVdGy/ikt3KHvvmsIf3c6u7ninTStdOIMnREfTvUli0r4D
/Rs/DDX7WvgDbxXRG9fwwbpq5r31Z1WcBEKYRxJzO3eJZ0RtDIajtFnRJpPbVDNxY/e1vLJuplS7
NTWEuzx7IA8HAuYcjtpEKqKvgs8LrwNHB3V28Zvv2ld8YOMPhS3hS1zTdL1nw4v45kFM4WZ8z1nV
MH568+JcCcQcisS5egvfiMpHrSdr+1AP4SR/h+06nvZBApkjiMN43sY9yGIBNqNlAoQDDz6ozGzN
apQkn1pVuNFrVU6dLGSfcSM1j017mBFB4+g2o03PzDC0Eurjp8Y1yFHiTdrKgMV7p9fK/wg1yDMa
xyGVhgQCdTb3FMN1B6HF7wNdzvay6mynfdGP81qAfNEo8S+Xuy28+HVUZRiLTm3SyX9775avB+3S
lX37m+lx2eEOIuoVkm9MocOPc8lAvD0/3FlG09ORrjufQrsNLCzMj2MYWQOW4Dr9cwEgWr1AcgS8
p4/gm5+17hS+JE7Z60b7IVPSnXfyxcsqh74FzeFiYIy67REZl4SW/vFLiYOdJuxqpCKGcqYnK6c2
aZGjfY0c7cCr1ghrfm410+FYtORNsSXiOdfE+F4hfTSLhPFFS0sAESkIndO4tnmDHSAfFE9qVdZO
yC2SkIhMRIk5jPLd+GN9SrG/hHHMCA8u5Zt7EWuDdpO9TmMkzBRD5nY65Gl7JDOXevXZyNZUjZYD
6puUcR52/KAr4QS0IgJQ2TbhBas9/JXsk4hVkHCXS1ZOg4wT/wMTATlbahjtpXo/6sZhSstydHFh
sRrLx/slIR1KyCJeIl0hdwQSEXfUFo3euhCDVWLy68GjGfG2mj6bPufyGy6vcxFpJ8DhNOUNTcyx
PY8At1zlz59Jn/+zOyll63j4RY67ubB0I5OtyyMebNqIaMqgSTye4GlaeJKMaOhUNeJBC0a7ZHB2
bm7VKXEiAadXflhor4Q0T7twhheknLiRgv4urbfw3/zNzIOdzIxYjh1z3qSAFXh7DEoxglzR0hoT
AS42v06qZLqJi1KW8f0LWUn4UgrOm6FPilSaC9uK6pf0+Pvju+jLgNwBIjvfLvjidK6K/B1Y96p9
RsnEH7YU74AlQTH/OjbXjYnkTKzlcL9PI34l+HFSDC9JRhj97RJeRf4fMEiM2kaCQbn5f5IbhOua
Fy/wWsFWnuIhUoZ/7DultfpK83b/ZobHiUrbWWB7rpMVaH0z3LYeNwAnIn4B5YlCHE73rgT9nw6X
4yHXOh5cGz0+O5QEnzVlu18ZQptx5jML8oynPvlLH6QDl9oBScHKMCn+G+EmToVRnh41D3uradQK
DLNqIS4vy/kvn7rWktY5W8o+T6hqgN6C19VuX8chNnduub6yshqFseEWJzNrLkaSltTH8YPIX8TI
ATqfL3xGDjRlCz/i7HCMbrZwQuxnLvYmxUsYSoNxToGAf9yISuziyinyja5fGjNbb7tchkVTyMWP
+tmh+YPA8BLFFL3L6mkLIIlFPvN7OK6LwB0PHNs0z9ZCvBwoLYb/sjtgY+unrKFGTlLnrn0tWLB6
gj1WneGGgd2J07i1s3FwN7UoTJsMeI5aylFTQisJuc3aOFNxrsiCk9WXORNTVuHFbe+3CoS87zR7
79ZiTqePBpCxrPuCpOmTyOF6IzhPlDJ80P7PY2XHHo884KaSEXMFGtxszoU95lXv1QVgUpdJ9OO3
1Pc/pHMX8E/CM0ZrTu/qjQAlxP4wH2Hcu4G05edoZLsK+hVxekEGduIPZsprONcSXCd9gypAmh9S
6LxGIRzO5CiwEXYBG1Ep1lUSCKE9Etq4NPfTeZcX4tO7lodTswqwYk3B22ioPffAVAgi/lLjACQu
evchQnz7PEOkU6bJKXgZnu4t/kj2zCKBfHhrWtnSRweS+YGlbeLK5YveXKS8xnbw+N+V6nlJKKNB
x8DBD89oPp0jo0z3RXzi9WB4/MSzmruYes+c7WjZ/YiLm8s/bFA/6IvC9HMGqxnYvMBlw0VXZnWu
SScEiw1SDuosoHtcRuX/KXTcJX7QJDQT/r3rDENzCdaDbpOF7xt8f+f0WVaYfoqR3Y33+XyBIwGi
m+4BCOWuEP8ulcpALO0qR54OvjIKqpLCE249sclvGQg0g+4C7AODvIrcZhfrn6vutE7ENDBiDLav
vfyxnSLyX1L4GykS5u+47cpiuhL47ZQvRWBWrLfmMBkVkbxsmwT0+f9DXxQXwot4kqQd/alKXaEB
bO4uGhTE7Kze7/Fa+6tZotq2CxLvZdlL/BzrCMTpCO2uvu7eKws5A0RLDU1UIV3DBfSrmluvfEPi
u21/LmJHS8MVK/Thyy0DrkTLAMDV7XL3xOFuOsh0u9nUuy6a0jbE2sVbkK1N+7BVIO66KrovCCEW
eiVhJ22WjqXTwvsoIzcaktbbhhlbih1Noj0QDLcYafmCppwPn0C+wCAJZ9Ak0GEsfUEYizThyu5q
9Ng+J+t+VjwgDzhocbz9k+4Qn12kbJNyrCGvvzC4cAulMXYwlA+MmrZ0riqNH80++RzL2Sx1cV6Y
b7gVqYwOMcnuDagNw02UAE8Zvqirn/TYrDJqmD3KYUcmjjJNaLeHHXHEgmteWaKV9p2dMpGT5rmy
3bsaKTvL8beNykDkwA4UWXSJkV5akaV3AhjoBSMIfepORR5V7uR2NPfVNVx6Q923t9RKH+Zv+itB
U3z/XeFhcbaWZ+W6j3IwftgCkRqITOcNSA2+BBXUlgv84T0WnngaCHhqr0xilSTaMWzAGlpjRGqD
VI57om+YobHhT/4SwCp6YOGphcpXmEX7WQf5FA8l3NmPsQDjjeY0bRuQ5s3NqqJRc5MGYFgrqxdq
QYZ2qDhIepGkH+Y5aPEhChhaOOvanCEdbHc3CvfxL7dFqUM3VYutSK7ZixSJiWMA1yB8D2yi6gOs
7BHnlri1qasUnVR872Rp9W8TadIR0AQFENgm5JFoLsXIxO7c0ZdExlcRRRx2qCYrR0PjDBUHL7t5
FT7hk009NyOhitrgN8CvWwaDfxFdQEp94BxLujfEKag5Avq2HxXXL+rLPR5dxzVbjDzvRCWqKzjk
jwzNV3RXmSsbuNLeQ9qFQCYvi9jV1hI5KBZbquWS1lra4/jNjvftPuOVM7E4CmHiDjiMNk3ZZAr1
vLIlo3KY8uZgwK80f/S0rS6v/KYNhuxRIxBZzROI7s6s87LrAgGCL8JVN4KGJNOZN+O0etUZ/t7Q
CxK/ByZGzO4nrN8/R72pImz4fNU1yoD6HSnkkwfsBoaFPk0IM+qZCK7+H3mpaYJ+nywZxHW/7a6T
aWzmxb6gHh8rVwM19ds8TWfrw8qhwy+3gVerVqzAd8qx94VcPIonOro+UTptopWf36PckHnVsEvr
WHDTOu/KaGwUvzNDiE+R/rxufsG+imj4W/W9nAoVvdamGDaU0S8ux9DX2ujn//4E7B/seahcfE84
LejJRiFyEYVBi4Dv/cZXUxk+T7npjjO4xr090G6OZ9DrV5hGcCrMOCKtxR5pA7Hc21QK9dMRw8pg
2TiOKZ24HTn1McWdospUjsmrQ6Wk+DvHbW9MiUAijT79NtDpWXAVecqJ2b1qVCpWmtzDFIqI6Vk4
A5qvAdx54HkbZ6SZNBqih2ehbxgx1tuFpzLU4iNAY+4Q6TpCKfRshqzYxBmNUWEnpdq9CNj7GV7J
uCgYHQL6zPYPK9k1VtjFL3zW/BxmZffV1/4CmJsg1rsJ+PVNLYlNvOihCcLo8uh6XjiUIeWWEoNH
3z7Zt+JCbGZf7M2UQ/Ha/GqVI5fSrVtYRJism2HYX4JbNDPp8uDm1zK/+wu4vtKD2D7TccOmjVBw
JRK+1LoOx5oMUXIktZY1pd740hy5PzPo5p2tC0B5ULC8a9+nCLZelNM3hQVYM5+CE87PlJggMuuz
T3vFGIYPjDuZUqPMEMHNoSUxQaBGSR/q57o7VOBe9y3yGy/FZA1Ujj1t+JgjNKlsnZysR5L5Ts1x
cSAv34LxOjyCPDtQVTJl+HUKRoIcSl70QKzxd9fJXaMobL3xYvqqidDLiX7X2/rcOAjRi/JeOFBA
dBYZe8ey1XUcgcg+iw9sQkEDhMVE/EzZu9aERukx8yRVHLzqxRHjCMmMgWHd0+MZj8wHxdjU5sIn
vAKevReG6FzzYIpdgfBvK+zl2zcwxLXuk73HY+JN5v4SbaVkWG5l1L+8x1fwIynvBxpuKI1hLDOk
lxxDzN5TmT8zcj+V8540yCSVgHLUoESW9jMfrrwdUTZ/SdP8hBZUS3WxcG2Uza+GG1863LOGofKb
Nc2LfNlwXQUaK84gfZLsP/v+tqWcz+5uHu6fwmJJxJk3lTacxrOPRD3u1ACus5JRnCmsDscXN0lv
gEaYAljgffEWlrp/csBvSSe0R0arHtJ3QR5i2EJ94xm2N+4HkGabG+s9LpZgBYAcwvrPuPbY7YP7
Guj0vxZ7GA5fDwEg8EGFVj7Mp5jra2e58E5KVU47p1j84Jh+pyF2jtv+khg8pTIZvtLx+WkfRSRU
Bi5ruAo2e1zPfUhxF/XkAI4Z1zl9sAxlQlzCVhTitjLah9v0k4OGQKiaX8TZfjLhJi5lZkPQG5no
S0S32A0TGLPYsWRFV/waPL+MXd59B+PvGWCF7SdcO/pGYEA8Shad5maWnx1GIARZE4DHMCR+8XlQ
d1Tr6jXib163Cg6dobuAJs1+Mbahk+5UGkMtPb3bs81whwKwvxFjG5JGYvwtvK4IFoJjyu4OMFl6
qEqtxrp5WBsIKSrm0XPxLJKgfIgvbIuHHtpY9i63YgWvYTd9PrSZJosoIXDOE4qfSoKYP6cQJu4m
cBs5MCWdVnUkRjOabJs/g3mHWJvaQ9G+FySzMUy6Rnim9Un2wf/Zw2TjgO6D3Y0ihmdiVWs4aSp7
HUAEODykQfVBHSLwh29Bc8vd+PkPUDs8U7YuGHos7DCO8tqH4LDWM9Na1qZozqwzXwNHAKK7FRfT
X1XzSY8wW0hSCGnaX7hkUpoXRK0Y0vYMzs93k6O3NCMtCQEgGZDCJTAp6Lg314BFdJdxOH3LPA+W
wVUH2Ivrf9VhjSZLXL5mC8NtRaIzFfv7Vs3q57ysU/Nb+LMZEavqOa7zfxvki3KXsRD6ZM6ajvcT
1ntlkS9+uj4bAqnbzVqgJxUumpbuZAaqBg6iTTQ7qHcn4YzZKd8R91ZklY66SxzAQGbg+yTX2Rfv
27xSWMr4mUK0tRj1kSjye09Wb8KIVp5nECo0nzhP6lartZFOT+uHZvDQIIyGcEHTB7Rd34u+6ydt
cYc9kqxRjrjeSxrgJBsyWk2S/Ze3kmZO2ofZdwTJtEagtc9SdcYt01eFy+Ap2HNql+B6tgEl0WE8
1+qf8eUHWdWKvspLlqzT04YRGBH/SrDdC+S+zpSwI3ynunSD8QC/MJUvA4Mx9bz5DVOQOeyIlV6j
O3EF6Hjd7n9oc+9hqN8swnZ6xy9TejkFHBbsHj+jbP5yQ2vxKwfVtG+RIfLaNqgFISEM0GQsqWU6
TWb+dYslCbbFKEGB+qxUuZvJQcZNbSaKzq3psZwKbsprwRSN2rVnJBxWDpo9orEgKGk5uTFx7G4X
Xv/Kkc2iqY+dVWOKI8kAnIx30Ir1ZmpKZnLukNS9pGLlFsJDXh/vmiJRx7OMQlW7fsEkI5ad9ERZ
nhJXj1tgq4ZarbRPtx6xO5fv1kJtkpsSOXIGVCGaEtuzWLZ5vtEwcEWSEDfaUhs8IEtjpFPNcbGh
7JIi5giSKmVEtwauUqummZzqh3zXnOz2IFY2fMHM+Aq11nhbEZA6cEbKpgmF0sv9XHKdsU7YyI/d
+2Fx3O7waZ9aNClWTkQTdYX0PdvREboFTpvtNilM5dhRWA1Xa0ttgYfPKJ8U6MdTj5CYVBQaz3EG
LEY5nWOFAaw52T5wpIhRulb5HGfeqmwrOmqA7St6S9iXalB3W+rfcWh3Pi3izWXLkn64Dgd8o5YU
UiRISvNMFKTeag4NHhsoHME5XS/nMfzjmoG9nBaxz86T8zlc4X/cRevWRzXbX02n3mmFSVrBHXBC
Uo9OLCcZlggKMwv4/5AY+Fm16uwMrjOfuASuC/JRJH6D2AupDr1sX2MRQnLhYLc46Pp3esqo65oh
Z+TP8TapKcTxVcMSbAX/3N9KsImwyK0W4kCFUowdC9R+FITKs1hns5fMkDm9mBbB8vYXRnUr+YLo
voZdr0KweHm5yHifAe3BlDemnZKBuhWELIhjlBTLhdveJnlm7yOtFCBTJzQ7RKXzyblBj3pAQFDY
minwBKpC/vtQwvhAcRr/AmUnwA7EeBHTvSlvyyEZXSHW95//0dn+h5owH/t75HIDlUujLaz151lQ
xJQPHetDn2+cI3U6NAFLlHe4JNyC7Mq+NKgExRbAz2mVJW0R4jL6YHlsmiuZ1CEfvjhxcPeNzwa2
cvGKAXlMIFaYTNmXeFFtcIPirDZbbbi4E/NwtBVkArTIf8kXXucn5iwQf+TibYTsD8lgoU/pS+se
qVHm7BYRJ0TRsuw5hEmJqE5CkzrecgM0dF4X/PDCJzsfi7p4Kn0/jl40zYsqz2X+jdH3Yn7E6xe1
DtfxGLeLsEVRG1LeCmnZSjGr0rr1pjdAYUPiWLvTGnFgXjdwVC06Wngl8eHPaz5rbrQvFImWK6kw
usiJ7KZg+Qpn9kCtz6ZsjlcsBUWkIMqKXTaeAeyDXaP85Oss7dwjWfqDxYQA0I+hBOLcC0A6QGz/
vT1a6HBTrk/K0YevkTYzirHTp1c8/oulFW1VoIW57qYejP0Ben76OYmw11fQaQtqMm7e9GYSymO5
/vaNC0Jmm+1jq9zQp0W/lTpzqi/3+o221YWT99AzsLIlRdJbbCYDDhDis7U4entmRD64DihjfA6e
i2PsWJw8gndK0DKyhgfUGo7dcINV508GjQD4mNN/iGT69XDnxQem67dc6iBxw+ptfQKOurGpkJa3
CRFgXyaqocRP8tLCFFWncATI17d7SpYoKC2kJYkMm/E6s6Xj7Zvmpp8oBvlcKXOL0bFwFJE8mG1W
7uiBRdnlXU5WmFj8rTriaGy1TjD3GPcnjAJsJgqiv2Z9n4wlTESfsVf++vU2AsTVuYzayuyhIgXk
yTsWyNt7/GtzWI+RaJMaEqrQjdp1ZKm3fpd8diLiwyWBF1iwT7Pshu3HPjr+KF+6n9x74lRX+ECc
ZCvy7hR+TDQEa9t6noERyemtV80ZJIrLRLiIB2HA4qPQoQ8D2SzE7lhnMTq0PzfYIv75Rpn4VXpw
oP9cFQr9JRnQ2qzdeOLcWo2B68Nt38AzK2B0IZ3I4UOY2SDFHrbMZWqAVNVZXJsJrt35NTGR4Geg
WyZXSBurJLEtETezys4P7XsJ/KOQzTXjbmxpBBlJHQrTP/FNlAxt0PVUP+OtL9fxJ2tKLB9kfdfp
oISPKbGoQsotSvnTr1KIQs76B6T9VjjLB7XKwG7nk0NwIPHg+1Wfcq0z/aJBt1uWW/NCe5t3k7TP
pABCOKDGKWVEqX2udVXPvSm2EFzouSxFm7rO31mAGAKmoHXotfYl6XnQpAimnD5Yg2jRJ+b/PCKd
SsP/j2KPgMvjQI0TlzgZP6hSxvYfsYipsK51NrbS1IxjLzK1/Lyv0JlysxIGZycHr4u6u9shYdct
4s+u3uszKxleXYk+lYZrs4vnrz15WVJpJZy+vVMdqH+pFqYwO41ereMcUWxDVjLvV5lPDYH9uv0x
Tg0AJkuj4hGqPBrCAQsZGSD5a0PT34RVAGtdQk48bqgKtWkMmPTgZKkcwFJVj3+p8SgFMq+6fYqQ
FXRTwEcjI3GZOVourRg8Eb6pRqB1x6bS+64kwlXMgOLXKdQTRoqIEsEU+OL/En88yGTntWWyncd4
VTEutVDUExQOvnfsAo0n7+lgxu1LpQ5lMaKsYVsGy8c4YAA4kfvzTtlqVx9VoVQieMXounp7csA0
gA4uDXw/TpZTZyAy7ixQ3jn9c+CZwbwYXRyuy1Dt+66MysTEiZjHJcy6i+MrX+/JewvJx4UVlTIr
7WggZqQrXxzqfLldP56v5Y5c+O9jA2WBfe5CSJD/V7EC4Y+Av6ZwL4NUyksiuHCUI8OV/LnVHORr
C2gQONBEqo2Kt1FfhGElFx+d+l8uBvmxum02q2vvYqPIEU594ryB0s0A9eS8pyv2HHMqlSrjqN6B
YS8dCw72uZ5Ui9n4bQBhvNJRzmn689GMdGDJTBJftgPRkbtehGDNVj5Y2twk1LaSpR/lFoHiDisq
sekoMpe8kC7hEGegg1LiLwDWiGS+/g+cs18taKbq2Eevb4Uvj9y8kJyXwwAM3/wgij+dCF7rB8tS
RhTlPcXqyFbI7IfgMz6E/VHh4pp+c1qVESWi6tF23ZN9sRfOeDBdp97bElyFwU5BCRBEMn7qWf9H
fE+CcWG32hHd41bsZDctiPO5keQQg8SzlkhRyiveAVqEWfBQqmnW5bKM/4Fra8fNArh8ZWhZa5oV
csvrJ66ffvWzAu3NswHA8mdKWmoGR69Mf/yt4huN2tc0xExRwDesmuzKDgUEqwUmeZQ7hYeO7BJ6
Dkm31L1rOswiGn+/7DAMUAqplI1G39aU9AqPS7QZWrGMlzLjwvCbKq5xPiYQ1YkigeL/oHRKwJ+R
OicXQqZ+GkHHYuX6b9xwDBwIMHwGhhhBi8XPdSdr0aIsjhuZV992mQ7XJb2p9N+44FOPnaatzCxs
E4K0PDFiepFBXre/tFhRXex5Gu3iUTdBFKVavV7KKBzk8uz62MoX9ebOaxC6+rkc/wqyZMHKkgAE
/qcsbEw0ERki3q7DvjZc0kOpuorITyzeVccBy4Oz/YlSgunOlbiyia8K2vkMl5x/vLgVAWCIZHOU
V4NVBu+irTvPQYjfYkE12+gbJXG5I3omGovROP3MphL+faJqo3DJNQ4PVK5cS5vhndezw7himqto
jXUBe/L92J2PevdalolPN9mURXUeteTVYdzyuLX9pZq5Of53rpTy7A++TBweWPjDBiuSa/HAxNul
1+TSF0Dicr2vmq3ylnTzl3yIrg8T8Sdikd8px8eBANnTGu5rEJMeFme4iuF5KOE+xjdBhu3V9UAz
SqNzMx29Yo0UTjNg+EBOpEijhivPNOY9f7wmZ2EN7H+xeog9MmITZB1mEGXktn7uarM6Vq2ilu1G
r3bJWFQsuzPDwYeLdRITzfAmd2Rio0L0/GQ9lJPqG7aDL5cisDOphhPpvSeZZm9g3xRKDdnmEXzY
tulRv/Jn0MCVzrcCOwxb9At/BpPebpJfsSyofa2/kS8JFUJEMIcD+0UgnU+x/pa4rv0ZekSxmPdL
Q7Yvuq5qA8S999AOgCHEev6n+zaCOSriBswM9g6NnoQmsthJM6VW+8Heox3PwjvjsWci179ycE2e
nfCYTnbgmjznCqCPwwXIwIk9+E+8tEr6ZRdqpVR8FfkDZaUaghytwDwVg3lfQTawBhhfWMsNaH6M
X5kP/0JQwxG0cAiush1uL/Z4IiarXpM/YrcBmXeNOyl49CtSB4OkkYr6MJXLDDfMswyeGoVZ6qD2
0laYvpBJVXmXSJ+iPE2g0hz/gSVjVEcBg5ovJJvxgAFyvz3MzodrHNGv+Q4VvesiXm4rIjLL4hXt
sGBXB6tVfzxGfPk3oQu8rPmNszf30UYjMV7QMpuD+B8Vk3DvMSSUFmJimo1fibtuf8fctEwCdYn1
7DTT9bKzcznQBz0oz5SANlO9vp20q7QWfE1NRg+8By5++9h5E+F7GoJN1tlQeBw9is3GNHEBOsgf
vze5ncfYvVv/4fX+sMaFzDW/NXnkLT7r/qCbMxDOl5R7GJ3/wgfY+L0By1zV70bRaKMqiCSTOspE
3YqIwPbIo9GF8U/9gAzREDspF32d+5DeQCJlTa3ItMLXPjRfUZ49/WXmBnyws3n9OiHk+YLfte8J
qxGZIQCeMdREqaaJfWdVu6o4+J8SNa4Y2Fstf9lMLOpon/7kfK9V0nnmaZyYBRB71FTcTqZcvnnS
x1JsPpOB0MgA5DEG9ORo/OMoWVyad3ykYEoAgK+IQkqZwG0vg4IYs3QnBdZdpdxhrHzdsx+DCgs2
huzu8Uhv40Zb8Q05StzSqCLT4uvLkAGARqWaLr4U3q3JNf+aIfNeAorc2uqtLIGu0y0uyKZZETO1
AhO8Aib5LHD6bvEtKVl6mBlm3N3ctRm6b9daCbqwJ+llqSgc61HGFpxOrl2GG1bg3LAxq79PuAIE
owFnAX7TY9HgHwJyv6JTse/M5Smqblb9aGQDbqqkFZpuuf5jHSSFTRdsKFMq8vjfW1zO/mzRmXFq
59PQTt0w2xOGLr/sHXygVooLSs8449tRZnosxcWVfOjouB2gxctjN5x2lLt6eex90c89/O+2KO5c
Qh2rrYnVO6SlMnnktzaWHUxlf045KVSXk3ntP3mV814AK3f61+oczijkV+XC+NOnn97YVHqh15/1
i8GUPnpmcOFfosXkXQEjHwRGVZWdDnT5cD6nGJ+rPyS4c0peo3go2vuVuT7uSlqo8baIZB7KzvH0
M7/5KtqlM3APyM1WhI3NtHBKxxRJJL8AaNzPm5/q0pkL6WkTlO/Xe+af5W9dOJRankOVhZDmcFBl
wa+GrxKIsFz9dIzuHR2SIdKYuLwSAW5rNN/JsTRn7UTsCEd4RAsORjsQBUsnHJGs2206MEcIjvoQ
PklE31t7rWbtH6csQgbuWjRSdmqmBsLqZKi48HXV5wXeiRleC2SEbasjaQDwG80ctrHWm1+RX4DY
qGjtT2C77npSm7+S2gdvJJ/NnXk3/ktqxMQcWyCtVB5d+3v1BEGw+FKonfhFahiwmrAUeTIW3G+w
SN8hj83NoA+6P/XsgB8nSatLiaHBBDBQ78HofQnvZHg/67mmCZ1dCFCALkCPIj45zRmFa7aTEW/8
cOVemgkjyLCBP8BB2HI0Q+qPGJmjg/PvPmaqJ0m14eeq00h21s2ga6nuVz7JApYynMG0jnaa2//s
lx+DQ5MmHplxe+Hm6OvCZpHOeO383m5VXs9ktEFcKNx5xNCcT/g6RHv1Vs53MjWRqhhrTuBxr9RH
FrAMCN03+FE10fExZqxg/vCZCd4VFxDNmOAlFkWpisTAl4Kjh0FL0w4Yhzl91/SGChpoY56kVbSs
rqghIMY7jGTwg04CBEE1jNJB4NH95BlH7jhSkL/KfBBhuyhq9bln0L+iITyTCfDfkTBBFloPghRt
T094PguavyPZ0zoN08PxttuRD/V7xs8KJmssdaG+Itzn2Z7pyJQacQtr2x9I8nXWNg0d2OUZxeAP
duqxJvNvM18Cu3BNcKyUZOTrNxZna/xpNYPY01BXERDmYcHy1YWB2ocrqg4JPIT9AlK0EYDKZqE1
U6Q8CTSeeCwdJwAgWuW3HxdxaQcuAxSJVm2VIkJleo8x9znELHfRf3Coo6HE7p4dCmhm8m1qP3ts
acJDKwQWKNCocIfttPvht6EUmyutkbWG8mobBGPUU38EqAkctL58n/ef2Rzo7Thdq8me3s1z67mw
rdO17jReZBHcgdZypIPYM2gzwoON1yNBTyz3gZJ3FKkFBnr4fbq4aofBPbj6gwLefcO4GwembSgO
obyMiF6S2t3jdSAiwelrRZkewvUbD4eUwty0vgSXMIHSZwKeazZgoEmM0uETx1AlYZFfNgTcj1BK
Qb5lK4yhSEk4+QVLPEV2/iKKqAn436dqj9zNqKX7Vue0BPU+EMqQXhphKOaWoRqohjqyd8r3OgnU
3srw5/QdiDvvT738OJm2QY/D4/BAFDZa/5DzJANTNfdRpWGkGEo5qb1fRlrusQIgNzOa2LqCKkbl
KmpLF122rfa168aZJBdtKLXFRHM9mU1qzXmkwKTn+asPe+KIH6a+El5/6a5dLVGFsyu8uRLSyman
oaxol81/wD0skk/Nyfox/03z4VoUpmAEwupMqgjY0uvrunJ01GyMaaoY7qOQqLhfHa9avSHL1epT
EYdjxisZ8J76/LeOLphfrxswcSCxIfpsYr3GlPfS/7vBL+Q1nXGxRrlZ203XpTVRQXL8a/eKwSW9
HyV92aQtM1gMZi6F9o7ns1RLzLV2ABe34dlaantuoJxxljCC4nOk2RBsgw6UZ/FtxGsKxFo36Mlu
raDc6k7rFWTzdeNVJc0rc0Hi60/O3qdcBXw13HyqdXsn3ochpoQPghJH406VCYViJfgzvzRZTceF
KDgtJoGJAbJ7D/rLOz4KsC6eR4rF8ub2AmyM/BvjDB8Xd48Fe+SBtBrejMLgEgWZGhi8xlnIVey3
hCrkt8JPdBMxDkPEcMvVhuQWPmrfT7Pa5fqgiMewVtRy7ER3PgqRKMS9QW4kZrxwgkiDnPK2jVq/
ehEu+eeu92pmB0uk/NAn5oto1kCD4CPJn+zBfwDFnxHm+fSI8lRNRK4jJX2EnegNznp39QaSfKFf
lgMd19G52HSugXfcBs/1/ZIXEL5Jkxj6tNDq6XNrDb8pp6F8kyYZE6oH5c9b9AhHdIuBfyXryNoA
D4l6y5RmlrDyMLdU6QoZNrZ9oqFjtxiFTyvV9kyy8YARvw25CrDCnlLDddOg4AnsFYpbglXHpSCR
Ec+8T73jSzcQNcPOdMeIt8HCU5/S1QdOXunJ5BW7orEBPrTnxO4NDjyvTpUzla2d7Sb4zjlktWd3
/OZWDKmbjOpSauhcvAJeVvkRMbw9doS5cHJ6j2fqKJ8uzdRZovY45MMo9LVgY0UyYPEmE1QAeO+F
JUGFfzN/KZpDxwh3ewlTg2dhuzgnFnyeIxS5mTmuWc+TBtDxg5KFrcy0+IVKY3buysCjbzxx+fg+
BMhl2fbAA9RlQBm13cO5WrDmZ5nxo6dKFpXVCO4N6ZfSP8roj9wKGamiS3OE9FHqiEIywBubtr48
a2nBrL6YUMX5y4ABiSUeiwjBDWoiESt2LEjP/Mm7v6YovccoFnpYpNiQw0qnkSx2FVkqI7gROvVd
Y2ahZ1ufLEu1c4ZWtJMzPr9aBC353gVwzFbFLneDapqIXTaqOGPzV1//U+qdRbzRWHn6pQmK8y/s
WOJwoXrPYhY0puqmpWqztkQBmjEgDSOgM3jjJuZ+YR1BwwlduPFpPAb/9xagZrmQNxU5DvEDVuWg
VYx7Zz5I3g56HS0CfbOVUEGQPvTELXkn17QOFjYT8+DJVGCCKolhTfURsV3zsuQcIYoZfBhKQrZg
COgj5mylg12J0Sd2xItd81OTtNz4K6HaHOk3V0+4giFwhD5oJaMI8g0ttulb6y+ipRohZI1rrqqH
yzN15GEXxNFWZCmScuePJozqxLmfzP+CFaJ7YzGJJb0guwAdXmDB0uhgDa9wQ3GYMMNUTWtiuIy8
QOm1r36vy8+oAr7qEmg1HRTncSoOCczBdpYe2vJDjmfCJPQmE5z8kRsSRWwd+npBHqRYllUJNS4f
GScEj9oB7maKLJ7HJ13mc8/+xsLXm1XM80qACqXNPyod33JUW6YVx+1UMErJUt4J7xkz5QCMDpIn
XvgRvBtQlNVUSkVZA5SQEpwmzyPxQC8uk6WdLHOR+c+Sxrevc7VSD3pd8CNyAjnRhvDst74nWUaZ
OjoxHkCssrrrb7x6NmPYKkitDk9P5lFvrfFHn53Kn0uHQMlw37DxcyGek7Y0d1W2uLP/0hL6VJa/
qyo4ZXxSFlMMoPD1lzjX98iK1O38EdFtG6wQgwy8xd/khXqEjimhBekw9j0VqrUnrPsfIamXBHmb
5fYLZSm/LxpS/XvmmlfLK8UScCMw93ZEVwbjyFGb0jdBsI4Ub6Cw5I0VbIS208OXOezaOtmrxA+L
7RBcSG+9k54fNyrfK9snzvs/lgBiPB5yoXxWa1TvG3KUVG1Rs8SoQAWYhdeesV/N3S1GPZGen2cl
S7+x2wkMaMH0W41xJi0nhH0wg4ACHTJ7DjEXerA5y3qOi64/9aCoUKnG8vFyvt7pd/2FIJYqsVzF
Gkuxn1nX6/3SVSyUP/mnr8Uf9/MY91RJ0/TXG9Fvli2VfSab5eqnJ+s78V04OG1/gjJclS87qF3f
Wup+0oF/vq6wALf3YmfOroX9SZd2BAp1io9QYRYcoFwzVO7T5Ba1UF/DesMf+t3ZCpqnx089hckg
tTkg+y7fPxALd7qrnevG7WmcJT9Fx448/6MKKSPqGVmYEpDygxCbdwDk0y2Vj3N5PrbVq4DHXMEf
5KTw5tnnhwqGjQ1UVOg58u3vyjVFtF4w0gykmR3gc0Sg/spsYGJ7AlerDtqTtpZ+EK4aBlbA+ZxJ
pXV2DnFL9jbTmjwqRlzkRaAX3sjq00ObW+IejHxsMrhkl/ocvSFMfvm3ccS+s1Ki6kGfvnAMQj/x
6+CqOYxLsV6fFLqitBVtd4MVlLpuQjzSM6cJ0DJCSeswmeGA6iuOtMdQCPDhShbrfrVzQ2f21ObE
x8grzbOt6dd+cEMVDrvurwz3bVx04LjYxmhxw/J1ZSSgsFlc9BxVGE16KTDIVv9fkWj6on0BEDBd
KGGd7uJXHMC7K24pVE+Y/q6J8BxYsp9gRknCQh/YguALAyfhRx93Xm9VzYAIUTi0rmCKIqy/CvBF
1zNz1zGhyiSgI8ZEt5k746fA62h5AlyPbG9IFXWEeJg7OYpTnNDsj7Sx9rU7wynlpvBa9rApaweS
ZNhGvLeCH0ELyOAO8zJhY57mpDeuFVieeCV/gtT/bnAYi2Lrep2QMPylV+mev07qyXxoZoY3aYNx
Vs2ZX3G/D3JLRD4X7TDFljdeTqbMKAjKc8cXNLS/r9/q5Midpott9kj0prefzyt8YFYUM3bV6sRT
LLswqg13sA+1ibECkFcwhVI36whw9sDkBzrMa8NYyoXrcJuYSvBByv50ww8S3SaFZmHh2nKKckaq
hesBFS0LNXKuzb8N86p9umAwLscrZjCA46FFUTJI1W2xW7yNbDs4SneWVjnKC/3MN3ue3nQ5cvnn
crXkbjViDlu5WKMUWc6Allf0+lDHWimPlV/Rv63TnGwOHDgRFHf/nSGooPd7vvAhsFaBdEdQISxd
vPgDVVP24WjzWjuUbWMb8YyP6PKi4/pd3bn++KDLplADJJ8CUvSthe5afad31PBwSqRCVt9dIvGp
55uljIMc9HutWI6VIsR32HTHIisoX0u9Vlo5/YfCtNDhJRDV4mxv6Jn9BmgL+/EgOTScJpT5fkuj
x3w9AK4Uw8mQYH838mYUADSaBAIgWcNA8AU09bxal69HyO9lnFPMUO3FM4RCdJFi7kr1bfkhH3ha
I4NDZRD8ru1KHtQAVC2qHZRUj6dMlDI9S5maskYQeWmyEz7091GFQJeoj2DwkfvUoXutpwub9XVj
4Shpbj326Btfw1HvwFVMrD0TYSAa18ySuyAnijIyvig7Ur15qGMrQw1Hu/bOYzmIFa5+eZGPDZy6
VUPWO1M0o79kSAuRskMhDMEyxaB0xpPE1VXH34bjx2/oOe2DkJcge2/z/C4B5w7bW6pFEMhCyyiO
ES/n1qCaTh9DyLLewwdYPPNmIbYbi1d9kBiygz8Jvnal334rtl5nMR/RGjZXehFktyJ2KOdySPdv
VejaJFXGmKxdZIIuMuoiFftrP+Vy0V7ewxsggyXnSBAa3lGxr4EA7s6Sl+KgcmfyJIWJU/Ye/hUe
Moq+ydTRdnqAtBEmRr+QOKG3dYYybtIMQnm4Oyzl1popjgs/vwpb5A3saHZdTaVx/8tEpyXwnbBJ
LJZ1uQXOucFpERHXC58kRqgHCyr33RUdSRTP09wvbJTfOpMhLowCOcOlZpt6EtgmfwS2s13bDsym
TXva33kfLLTIAmq3uM2gkclXrzGXRKQyldsMNaMu5nepq7eYIpzEyrZiaAhiNtnzpFkXGTLywpOx
0WkrJY8KHS4YpPCe01mVg4DsYX40BSbMQHzCzUtnxFuO/isirgRg6Xj51HLv/PBcTCKDiEjsgSd0
k5v5p6EM7GL2CEawpkhJrg4MNmunyeqs4KfnXA1djw5Mnd0a9GVys9RzL7C91m/vXOkQ+tiV/lh2
w5+A1ehXBwg4Pcf95gEws8RTlMuIlizh83APF4xFZQBtBP35WpWw6A3/fqXL+N0Z2ygO35aoaz7z
1EqeqM1aVhSYb7Eu7HFt+pkcySSvNAYGpxSP6XYJ0gB/XgtqKZHxoiL9xFGQ7UgzwDXLqChfc29n
7cwGROkoJ9XRH1R2GAqlPmD1nLPCh7bLTIHs3d6Da/Rh2yCiufOhbk/z8+1Dmz3xgFLyx/s2x9hX
nPxY3JtFuAFzj1Jx5YL+HfYvDbZxxTlpjLcDjjQF7yhMZadIOjrdvPSYlm7G39Cje223Kw/8Nb+B
Y6ICNYUir4HMhU6G5i42Qhb1pUSpTbkVrdy+xhabABte3sGUdKC0Yv3Yx/NdIzH2owjwghsLlpPR
TzbIX6daSc3wJg6/fy3OPHyE8LROhFbflFB7LVnwYeVezFXVS1Sfh8GVO7Q+4Xy+O4G3cgfIqlZu
6K+xyjf4PXpzmkzKHV6vQGJvtNV0ukDOHlNlKIg/OuqdKIsnxPgnPwXxn5bryMF4Wu/YB5MVia8b
aqYUGVqcDlDcqIrz0RrarejIGjEvLEzaBY/zTUQBgnKvc+Uz0x8UYLQg+Fp6ZZsslnqBXlcGLw1T
HBhx4HWyV6B4r1aIG91L/Zq5AT/UpcqKn/CHLaUakeWCKMU77Mca8/yuADrX41d4XX7yJdeFKZ/Q
6NgK0GcrWR7e+4NCRuWuTJfW5SWEiNMLvOfrH7Wf3+zurlWF/ozo2QJ8Jfvcr+FSaWfRctp7r9l4
BX2LDMAb9rzS2z4ZRXK3SA2MR4auBw30zgogkUAgiQ+ECukRWaZHPUM7Kcf/UMoA8aHw53RysL/A
gVtSVKbhGf72vK2RjdYgT0F3Bz9ntwqkCA3SchqmR1GCipPQCn2KLBiWf4EgkgMdK5PUPFwQbdSX
iim394rhGGzElly7ZLcW5RX8MllXBchbQ7bY7YAFfsn25d9WR8c6YO9syILrNkFrfitUbxGetWf8
raTpifyYIQF6segZRVan/9s/EKeQrIKveCFXq/jy4+K2vdbIluuTYmUNu7G7wIjVo4nMvBJj7Zgp
vMi+IvqgB5phqfOVKz2OSPpMcDl4IvGSNWJwHxIIas7TvvoduaiYV01lyelU7fk+luXGpYFWZDus
fziuITLO20bcaiMJveVaW3HqLf0xjN9nRNTPep6PIiqahy0bRT1sMog48nnWhRTE5PrnosgSrUIL
cvHBhjzaV0mMpDbsNVlaeFOZsgrd6GoBS3dmcTiLRKfahdfr0q6S8QjBsS8QBaZ3CV4nTnXnM8On
SOhLFAbvDjeTs3dCzF4sMYfA+h7S/65iLWRb9qjVDgNehZ9c2CwDA88pT12Iy42XbNNhy9waPSSq
kYsSsgvwpyP0L62yVGEnOvjCpPCnSyrfTjQRL5oYZ7oOVK3T6aHk4cZB3rUWyFOBgM5ZtAXY3+U5
vUdlbzi2HDDK99Y9PPuNiTukSCulUNi2tYR1U69La9lXT18lZhMO04Ggu9ZBEtnZfQ4OHa1HCkhc
0KTH0t26Rgq9QJtAKOoVOirqAoGEHpghseQ53Eak4lr3boaQudch1jCSUTFRaSmzWHqZ9a64OQb0
//W+0zHxiecz9m6O8VTJDlbw+QukIX5WwzJH5qvHPAoAc80uT2DIPiL5r1+E3RAHO3hnxYmgVM1N
KD2pxlAptVTcNg/UbqJQB0vgJJj7x0eWMMu+klHQS8r++tOrgk25NKe3vpFLKXMWUq3dWwRiLDo5
hCRVEvCsvHLbGhP4Pg+cKpNo1U9JMey9W2BFBc3hNZ83fgO+r6koXlAKUraKQraGbzTz98jmMqiN
HiLiq31VJuX1sWLSWbkCD30b77b00Z9hiK+UoeyE9mn57nDeab3o6290TeyP9grDBl3nBG6TTj8b
nhLjBqFG/qQeHs2nPf+P2Rq5SHpYbKbvULraThG/4YmxxEbNi8U9l5aOIfvOkdQMXXWO8FeR3AFt
0NYpRaqXZJCjUHpQglEBprj+bjZO4bATkfbiBSaT09PFBY0yb/fk0pYstZWU4qnrDZ1hQI3qRwsc
XWY/xaGQ8Ge97Zrtj+p8tteSMx6J2p03slxtw+ECakzr/ORNNQYzGR/AiJ8xPoH09aT6yV4OEej0
m+Zwv6fptl2dU77p6ElSl7RyQLYUV83c/rSS9XDD6UDKOYYTmtv6EBqlNJsOn2Z6VOTSNXTPuzHf
U3c54v1GkrfI6KymMVpEk57m7Q9GzFAZhagM1aWsPn9Ogp+44NVj32okDuO134o3sr6JjEXoOGL5
lgM5O2YgXj8myhkBo/77fydpq+bMLb9rGyq52M0FbmD4VozY1WYXZ6qvdbgS0KXbIItWxFii4wdi
4a+LBtjkMarsFMlmT6QUb/SL4QdgflEC15GYl0N3nWt//sNuO3Gi2ksYB94dPkZBX481QvfspQJl
Dubf0QmSLX06Kn9fJzB4IO6sL/tgppiUICvy1BGpCP8DjhxhcpSAn8GWGTV42zP2pHlrjki/w7qy
M4mNUPRU+21E0EsrsNmy5apHp+Qo+uaMgSDVr5CDfKDV9JPkU3uOmcYB7uTcwq4Sy+b0PQXNQbBR
giJEx7KZz2+b0R//8Q0XTqqwKBwp2etoSLzs/046wj/k+wDEi7T0heqlo7ImbyQSqGdoRiKBSQea
hmH49hDliHpO+Arlx8O/MyDSBvSZ+hdZG7VUfbFg6FM2zCUqq/YsJh5HW+yxgsswvuG7g1q+nSyw
orpGoyWlOz8/xANuyJIdKrd/PJZ+1EnHaaGQsdb9NAfNQ7oKr5w+E4fxRQQ6y3dwXLRj0gxbgPJW
MbH/h75dUIFhhAa+4zah6Ii4tJwVIjPU7iE1S5sQ6sHM5eX4mZnjDR5SHyb2Oh/IcFURnoyMDYs3
2YjnsM1BJsaUDotpkVQZpmTpCLg/WEbnbO0FbmKoctRkaW9slvFGIRWK6IUUMb6usui/xvCNsQko
Id6djrev/klbXKG3GWj05DESJhD9cNpT92jfLA4Sw83TiMI88y6uAifKzycr50V6+AlIGSpBBn6q
B/XZ1oFSRcGIXzILCAyyTtH6+II2TZePpfWfx2nC/XI7nsStwFHU1oMgxd3Ztq0FKYtcNjzDGFQ7
cmlsSxGLF0MrsiM01TWxAC4eLWdSe4Ro+ld/42PX1hWv5EZ7Y4WsaSanvaw0WGYUhPNcegS25C/o
bJJc3s32FkexE9v9o3TBdow3q4nsShmNmRMfj9p7K7b9cc6WJd18sX+Q9P6cEFx4R86WYM0tGzGX
XfpcqrS9b6aYxzE4wROZd2hwT9v8YoISaZtMnbtxHxIw363WEpLTaFOCIE1R1/+X3JWDusSpeqW7
jPiDUOo24CaLMN5cfCOqbVyMb+vqaHgucszmx9l9B3wmKuaSEi+pFKiz52agSorNZvAZheORShuc
AJZgJBhd/neaC5InLKBuMwCwWXq0i9m/jMVc2dToLcP6KqmuOAQGUDI1n1qpDPLNWHlvPZwqUhPB
TDt7jqrqYCuowebBgXEiVhLXpv+w89PCjI7XTkXSIjUXvzBs+sNpmrultFoHnIMXj07crgVJ2Qn3
9VuHde23pvWR0y53HwZS8g66B6CeFtRiE8Prwv9GIH0TwgtUWgat2eEA6sHXhxRXv6A/zrFx0+DU
rjLow+k+BolmBSGjuO9lKEc3uYsRWN9rbiHMo7E1isl6vSUfqKKfXBlmzisdimEHOMKU3668V5AC
cUoJoEmKDL5wYYtWDWhxVVDBc79YpeR0OLDsqndeAcVCM1Phz0ZPvkiL2sI19/w++I0/O93BqVcj
TUzm5mdau2pZSEHTqb6aQFh3NlMkbrLg6aM8F3nbd+Gh88r9jBVnohuQMwHx3pvUJGflhOBp17hw
KOKLr2up1jWqkudR+pDQf+vMEwzOo8bE/Xb1h1vTEMs8rj1zMIy15381ykI36PurIluDjln4qTGL
7ftbWfNTL1KpltfwWNQEfGlcC+wlKRsjV1YNPwuMo0pfCBJnHBRZfUpLRkoiJyDMRkJMIZd2tu3R
ng5hRV6tPJlRqG1AosUF3401Ve0Yf1s1SILEj0E9TKGP8iAtpdt3JF54Es1/XWvmPxSe/pwBr108
wlgFGWFxbBZ1r4LzCwrewG+VqGzXPPuobjhiFU6iFbgWvrdqIhfLqUIn0cJyZmyzAP5tKmB5Rrw1
i97IZcc/hME61zM7doWISN5J36YRS0oLwSvCFcaYoRgKlMZz+yeFcH68dWUqh1Fr528dBy4VFIgg
Sqh9PcCGCqdOWuqmony6CAt7k0w/6uzOmmWZOqMgd6dmL91wJBgn9/YkdDIXosLAVsZaSIOWMpCz
oRNT/d9fLVul/6xVItX8rWmbJhaSS6NK3IWFFysYdGM833ra4/6tI9Y4PYjtWaK8c8ov1md1jrcO
kQtjgpNgMaZEfunqV8oR7O/Lyy6O9MLnlRQkoxdEVv0/wRDuD2FuW/Ndy/mJQNPhXon6cnJWLVMG
y3EjD9Fx7Lj0/IfH6d/wPGRzfh9JpZxMBLbs24X5ZGY4cTQw1rbi1W9+5dtzKfKYNJRRymrFrMk3
+zpzGztOY+QF9oXX0AFKMF73wUXElTMFHcy1wsrFV8K93x9AwdovbtyAxEvwunUi1ZYpTKSe4VEd
biIm5ro07uHB9t1SSxkcCPhG50WKrnrOU4xT+Odgx7lYsE1Hob9V/OLWSaDwW8d2nlNLtrg9PTau
/nRK5XiKHMJVTplyNswt4g26C8p6Em6ptt8g6FO3fl5yK79HQzsW750+fmBEd99IGqYRx0tNYVRi
aZCix4QC4sEO1yZX+VJrMqG/ImSHismF3m42IDomxiZ1xgwU7dx4DXq4M0D4v5G0iMl6C2T8U4iV
YTFGib6qtjtnFkAsvgye+2io4SVRSinvtvf981YSN1va9JgXXPQD9bd27efm4z4lPXFGWCpRmjTq
U1SkhfcBv3H7nSiDneA7SUbhkBq9NZbebkCB67XFA1h6f7DcEhteNyKQSomF37r2vkzGr6MV5ymi
6P+httZktLbgEDNO2+qbvQSDjyGcYRs1nsqOhpY4Segw0PMzYokS08KKxoRxzfxCoZUQKwHSioIc
QyM7Y3ovlImoLHAnZstEn2NE6rV/LfpI/pz9gEq2Uu3YmnhV0/T8/q8blF4T2qpJDQzit1cTtBLd
/72SlwhVlZKmK8HAw9sUcSvKJHD/ZONjFrsrAqa9qOlhIAeteFZBj7QZd7OpkvwGxVxSM50YT4Dr
q0gAmnHu789lqmCNmJaY1IIF7K23muJCHfcZr6fkiNneQARU2fNgypFLPHOAdrp3Ov/LhG8ujNTV
zMrEZLQVpErvyPolInT7NXiMqpfq2e+WYEjoZEqmBDJRz288lsTsozqZMGrkASQVWj8Jt9AOOfE2
By5nFTe4UnLArdI2MSavcX7FcWX6iaWUveap6ZtKyheqGM8/4pKxUF6noHfGyrESPMFmrnXD2zVx
1btKzPwxErIlENrMeNVGEwcMOta3mk7whFZZdTFY0y0PgUlFjdUrI4TY7M0XOmJgB6ylvblJRm3h
9mG4/juk+18YipKcS10wGAS07lRercjp0MYx59LjZEfNEJYbWdS2m1g/1RUPb8QFsa+GX/n25JwM
3aR+1TVFtkJXTi6EtFA0cQcrb+w2KgAEYinNtkAOOBaVw9dLAMpsNPt6tT+kN1TZsYP/rfVjHfgi
K+1kbksvwclZYWE1hBqFcWR8OonRHDcxHR/9QqwvtVCQ/UsRhD8WU+R5y4uciz4dE1ytymyEeEui
MnaXAxKTGyga8PjKzptA0oTLTDhS/R2/eK1iIiCiBIiCo0PVofcteyqg32TkfFa8QopkrzQJCFi2
g8MnYiKfdO/Um87609d+fuzdprZKPaGjvkR7VPb52cmnvHRTl9xJHvdk6y2bjxcHn4xPzPilhruY
K9gnwjj1a9MCOZdLJsZQHQXYEJ5U+DEcH/VJY5DCkOf073erYGVRyyPC/c0GGzkk/WlbJVXDm5l4
XPoRXSzcL9Io/e8h6ZIm7oUWtxHXufl8/FKmlkt22j97zfEqOLnf+8QEIdr2BbPaPhSa9s1yUlNE
0VnudkPeI3i9AxUvpjAxd6jcZtd7q/RVZOExfT+kGFOd+tACryQY5+Z3iw8O4w9Xw4Rbwda/D/EK
3JOuyy+/AbKkS8W44ODom8Rhq/qUEWDfy2iZcoIOZAR3jjVUR3wNsn9Iwy7M/vw9Acaz//8hnW4e
gPAa5CIIBUkuylk2Wj1sYTNE1bO1YGDFGWFtGgUm/z/at8tP7W6rUOXsclAIRANK+oHG11sBA2Ie
qYLyPBh7m0PMx5UcZblvj6DjS42F1xzuO1zI1YNO5jK/lvewJEwEXiQHtXP7vxUpEeVcIgthvP3v
mxADBUFIlaxy2O9a6bIokM0VdfCZnLB7fBedyQJdI1/IhvF8sPWsFxPLExmlZ7thswTn6B4FZn0G
k0FXWbLCEsxF0HGWFBN4YCaZnU0ci9dkSr2FC3augmLcg0alOjHs9T8one5jP2gjVi2ZGsHQS5Yt
++zmIONDbZBXg8YpWtJNw6L3WnxyG8KnQtKVKIGEPD3/nUpw2JOicS4x6/2HhEiD3LG7MvCASczs
jPVCyEqx9/8BLjI20b+T6VL1dns3gzjghUUP5gOgv3wUTmYjhjPZVag/2dYvrD9B4UT1VQPX4UCt
i90Yt4LE3P3p6Xep+Kh5GXjsGVVqUShS5+2QhFFfSlUBB/wyAwbahvQXw+mJvtspj88SgO5pwvxb
SrnA95dfj6LMCbl4LDAKYsUWTqOC8nr5EUNCplW+2T/G5xaxagIHdnHaeWDahjhArh9YmTpiH/Uq
cFwuQ7psFXctdrbFOOaOraxXa7UVUXa49aqpoWBlfzqdLaega4pbL5ifkUDqkGIQ9+lZlWMCyOnv
zXQrot8fJ9zr9IZkpY/28bxkBshdZd5ZlplowXWza0mJ0UdVh4MUw8XBMBBJQx4gjfHQdpgxg94p
66CNbfMq8JHpu1thq5/fUeoe7urkSfsfHwFraB1ot3yCvRP5WqbnsSh6AQJzwq6mhAnEwOQ8PdIR
h29s7jlBXvO/h7mjpJRdEgzkzU5s4aDrc8U+wl2cIb3dsjx2uerz52YqZt/f/vbVioViAt9mAyoq
2lu4DheY5mWLQEZu8s798mKJ6OGlzWMGqI1jfc7Jy+ypRnDLq26UWlYvZgpk2B4qtY92RjgeE4d1
k0bbG9E0ZNrtzvJZSF27OVcEEvCZIlXfPQMJaQwq9Z7rLJ4/kYJDqA1DBv0k8IAv1EQjTV64cZrT
mfMuzRQYGGl9z2hmviiVEhZWVbgWhj4ORPOrt3ar+nXQBFUCv1or0KdUIQEIzlYsISE01NyuUAjD
ElRJjw2YDNcmMOFil7/L/hidHvbw2HI3/y4JYUvg6zPayxz8rFBbU/8Jjvde/jj+1niORO1B8SaP
a0JVkPwj7WGimQ/5ul0Ce7VgrgoHcoFktHVArlqrB+gVbDddlE1lK0oenN4uALGxmKjk/31QQ/9+
5lySenTB6WKIW2T3F+xnXwNveSZY3Vp6nBiU95dJEhofimtOex+ujqTwmdiuZvK/Itf5FlHFKpkV
AUU6PtFuXSqp3+gkcFN1hQGkcbhe7nrv2kjQ653RmXDCzmGHjXHI4rhIB8dSz65Vtu7YSACXX2vR
ZOyYci4Xe/qhJvlPsda5VEkGnyECt214Y7LmfNN9bjblckrTen8JK9+YtI2sa5z/G98A6udqnhe2
xfGSHo1aGqkfm59KXMvagZrqEBmSCZTgivFuISgxAj2cZAmuBT17K98lh2nq+q4weGhuM2ZZbS+O
/mOhcRsAguqAg+X422EGfsNAFCweP/bESL4UzB7NiFEmgQsDNV6G7bMp2JkKb9Bw0PqDFAE6cNSt
6YbKwQgiiDSPkqhKpQg448HDYXzSq3Iy9bWsWe4jxSfNqn8cz6hc8vzRWd3gsWMNPfpPSUO2CwHs
K/y4vAMVP3Fo5PJwrEd4TeUzX/Dg28oROcqQhVtMq5xp8Gi0NyVDXcSRfPkqsXHopp8mX1B9c0N9
YS1fniEtc2V9cgL32MOyOs+3JF8/G2ytZOiFk5Ec7WXYnb9P+FoZORxzpTnlg1UvjnJVRQsd5hxQ
nXnT28x9JGatybXFYOyBwLPykuD+58Wk4KTOurWq+2cz5DQlwKMK0LjeHpyjWwm2Piz6jce0eMKM
x247Rv9iraMKScwxHH/1cHyOJ2/owS5zLLzsTykrC4ekZRDz9QN0PEdgvUtMG7S8DLNtW5pY33aq
BuXXiwG9K8g0xDCUX9dAOClUxg8pG1TLbLay74GREVe9lwFp/ZXKiAczLkx+qaTeGzb2jPXdtf7W
iwPrEVbqpUjP7C7dTdGOK3vNpEXWhh8bI5nc3HaKN7xdQOERF8E8zhOi/XM3PjhrlUO4fVkR+awr
Rhcy05nGlfBg6w6uddatSoHNy4MldVP2/QoYWudOMExoDZH0IhNWHGclGgVVtCdI//X9ZvMb1sC0
Ntt6ElXmTEEArs2qxeQpbF7YkC0AFmQUGBU7evLOkLmNZpGk87znHfGMyMaMJHM/prOcvGvIoRyf
TPsQsuG8N02K/7qw+teTp/RZRStlCdIOr2thy3oCiiYft0NeSJZM0zVcoyJcgj3JjQlf6+dgT6+/
UsUXCxyUgqik73Jok2nvTVRuQcPrQBEy1Gl48b4tY0J9kvO0yY89Q4ezn18JekatI+lL7FxQXNAf
TYA64s0ozNupj0rlVMNKPKxMqom9uSHcK6Na6aDjfvs+HB+khn5Y7OlazPZyu55SdH1LuqD0Ib82
0R40SwsSE5FI49AOIN+WTyI/SZybKfUV4Q0Djh4fzWIIH2kzRr6J2L/teYXVrPfo3ojlijQCEEXh
8zAURtZAaHodsdKSarJk+Kv1upLk3JfRAtHEo+lnskGfcJD53h6aIIm+k+COeCP0ZbSJZ4/92z/7
tUBGG06Fd1tiTIDcyroa6Oz+0qMMyC7j7ib28kGTJ68hjTe0CsVVJ44x1Pa4HLPWOsbISxFbQcnk
WwFtcys50bnQjjqtlKcEcuNZqILxW2ViV4FW2OpRw4WzG4Mk8B3gsXLfxAnGe8UHXozoABUdYLgU
l+vhs7EDcQPwbUhclgb4ce8n8nXAlKQL7xAhRoo7IY3m0wEUdauQnmFfCSFqMA8VJQskoQXJuSbe
ikcRajmGqStDSEDAH68PRzcvcGCzWBP0xAl2Kkvl2lwK+SHjZ2dssb40DM/2w3EG7nGVb3YBiOk9
DIeYTQ0LZE/N3Mw74TSLMf0xx6AUuAg+7bgjmDd9pzdC7kT8py71pjTwfVOMt9wFhtkRVfKgm0zs
OaUqRHItzpKchsVv81F5E2qSXpFDwoQnXgpeQAgb9xZXQACeCQrePzGBdbxKZaxn0GNYpd7xpkOu
GFLJM82YfydCYGv5n5/K+6SnYzQu0Q1XVlpuapx+ftV1P5j19UUVAgVl6XXmfyw53joYRkIbvchR
G1ppHDwy/usyhdzrZGizMyguzZKw+u8rbs6KJFzmsfeeGyhAPzXblue+WWSDsAPw/E5HfIDujRCs
yI5QsKax7xVm4ek8BgAuD7Vja9zwNqRI/AwZqlyg5GzPpHnBQZtQ819K8FWu/HKLrGNErXqR3Kzy
6/Ib3WQi1cm3Vr9/FFmv8BEIa9UreMQ+K2/DXk4bLjrP5VjhB4da8xFc6RjqNkVvtpVIGt4Q+7yL
jwc62Zg5hdMoy7yrtwUjRt42bwr4CYAMdQBdOAayNc48TWU4I5kzLiOJiMWTZmihE0mzDsM1Ci5c
vXfFcN09+EGKgxyGuRrkJNwClIXaGDSZqeYULOHK2ETGUPKyjgl9HKOJs1hBVDkDmiVtb2UrCLBK
ogQMMdnTMXbfc0rsQRVPZGgjBbFHBW6o6UaBzGEks9idxsXdSWolX9ULCYckbgB8hPp5LgY8RN4N
n0o+qGwUgRoV2wjgCwNlE28zKPDUAOjRFtwdT2Sr6yYoW/MNxJ9OH2pfi9qX2qA6jYhZ9wHVDypl
bqItmaaBmwrxMWEQoxZa+q43YSKhFKbO1F5BYgjeZTeDKcQW4kOLg9Lj2sgGJnnEWXw1e1Fqfu14
mIRTN7ti56zxpdLtoUc1N/nkuUQBAbBZQ/k7sQLNbQmIkB4k5O9bav68/680eFQtDl7pImM/hOYb
tYlZu9U0QEA+SbviXsvE9EsIis0fYuCqyTJTLI0M4ZGadh6wi/PX5AJZq6AwBQOh00d1MKxZ7s20
uvs7BgXAhX6APXJB95h8iD3F0I36JSxxgTio5hTZolPPqIYgBHONJy00pyOpl/j0oF60SYuH/rA3
igO0Wsxw4Ch/adKQmveEguKWWs7hAYCxHTcTooBlYZd+oY1Ny0w3TYtVOKCBywO6qjajgb0wvyBf
arWffasuX3vn39yuMrff92mzQmTcMwAUYO9fCRLoDinUiPe6ni1SrEQ1+zwSIEhBeZ2mkjv+ShIV
Wvy9CLSlha/BAkozLnJsxlNPYqlU4oYRyG8vfzTcvYn/xRd2vOTmoxnVWWRv2uQnkcFbvmEVo4Q9
VtS2EqsRWGObST9RS8TX0qVOfL/LQJbAD1CpQMv7ys8E4/h00qmBKFLxP1tUshLc023cNnKfIq2k
ojZP8DXQYKv8XvAYWGM0LNk90wrNEhLb75c6YJ7ARGPtyuu1/p1sP4RCPiDIsPAeseqjLhe1qgs9
Ma2umaV6p8mdziE1O6rLz/FrbT56xRBMmFlMc3bpI78nPjS2VXqZ7pOpwIOBuq+r7uUI8aByi31v
hBFXQfhefIR1TEp/0hHv6VRTwK/XKr2cle4xIXF9XOJEi/jqrCJXIF4zIizR9HLwAx0Lbvrgh2bf
ibT2upnb2upj+I08SAvIId0OHKaQJGrY/AhaEWmMM5J3bKw3GojPaRQubAUKnRWvPWL8h1pwhHAn
hUqg3+ZV9nAxL72nMcuEGkiZrD49YgeTrRdKU88Tmmh1GZvsQ2tx9Z9biAvOPiCVKm6aV2GAIl7h
Wk+711Zw7tmfpQe/xsiendHMQwM6afoj6xe9j4UW6oMlTtjCAVQC7lvrFWbSgwu5qXRkfZ3OQ05f
A11J2ZWOZpyJr5HSuPttaV+O7ZFRcW5YcFmLgOzrFJj3Ja/p1bk73CkpmtJ19R3tugtmeD8AX9qw
LK3gsc1UbpDfOFR+O1ZHM6l0uY1sQa2rBNhAlse9PV4Uf+gByGtXqS7ZiWIh7nSohbLDnpT6mojn
dbyPK6GyhxvGEQazIxN+VOShyM7ew7wX99PBKE54ljRKoUfmJJlmjFk+6ZcFS9fap2dBv5rGaRN4
aiWcanZGgNEt+iVGhFRptB9hCDXPwP1ME+Sz8TmGIULyBnfCugHl4tnHF16J5DEtJJfHIUOPteDm
CVfsymLh/eorh5T9CkaTYes0tHW0c/VQVRCZ9VGe7HgSMfAjUKSB1dWu5poMLPxS18AGDyjt5CtH
lgcVlvvsn43xoNLjb7ZglsDM6emiOobxh1alpRMBeJ1Dp+T6GBdTH1TLkNvq9yGmulE3eWH9PJpn
sWxzFJ5JJts1ha7yy9wizCEGiF4bqgtk3rYpM7XPk1G7Rkczw+YS9lYxQ+j6PpPvM4ui3R0Vb3lV
dmND9Ht9zX/5klvpd8uEBoW+6VcDYVgzABM8fSgk53VDwpvGHrUeMRj2/3V3Io+2aPwGdNN96yK5
K3kEEJjPFWlA4Bi4UDhmiFVbI0BaeZse3BaUBMYyAh+x17HckstPn6WZes5sv27e7Kgohxlloty/
Kq2ybAwSYQ15Ak0YrlvVSCXwy9VrmqO+xMMztjBp/fY/qA1MdImskTIKH4dyFuxbdwZW30K5jv2t
erQ6qMXEqBn5qnMu/yANZDymThYWNKM4QkiqsJTIyAEhOLS8mzvXHcatXXonqA6Z9OiCpKpLY+uS
Ybk1fdIXLhTwODMvmTxXv8OHDmGM5L09c9mlbSE8awwqdKfuCHd9VmnxvaPUQYK8j4DXHHFJtQD0
eOV/CLKjG9IiFZpB53GQ9L1WeiH7KMbj/DZfhfrgYx+wO7BXvAwjK0JHX7FZ4beTJv+um2DyGYXT
c0+/7h9ujn9RGoG2dhXdUGoJ2B6X3qjKzibevEhVtLb1O9p9/O6lYI5i596IsxM3a/Lp6pQ2Q/y0
ZUgSRJlvfCBAaVjn56vZVYPP6IsWFq2uBmHriJh1F3rEBSKXBUxapIqJQ+W5sI+p8fxOdeS8h4PK
WWUI5eVyyWsb+/wmYSRAgfIkk+AIaIAkwpkkSYkfPakvDyEYw8aiZVUKfARPw5fdFX4anAbKCm5C
Yw51LbyS3uw/PQPwj3Z26LcAq4nzrEACbqvCPDk9gR726JqwD1IhnyTWC4EnU69so6N1WWtwqki1
M8XyG39K7Y9a7okJHsIXwQWT11xXhn50f6vuGcgUKWnKZLwv3SKHeCKD6ffHwBWGl+UG9zS/iwJq
8Z4MXnBoSqiimjcgs3dhXtjSlI4+psyS1FE7U+0pBjMAvrizQdjEUe4Lhen1kHVd0WgfrJ9Md2rk
EubQIPK+a3O3T1/o2+7JUNE0wFXVRmiWd0J6u1KqgSwtusKB45uEqS9XonwnhEr9SZDN8+Qey1CX
+ZqC8GL7IAneyYrXvJEEm99DBiqGpXSHato515fMz00CLtNyjfHGu7Lqku5M9zDneigoWG9WGDFO
Bz+92sMT2jAslpRsZR7vJj48tj6bi+Dy7wUe3WEzPM15wN9NW4WXE7FdPymYNb7USGcK4DVHZLip
L3UTfcekb2Pz7pLU7/XIqgHzpED8r/HB7Imovjx4Zum3u9Mmh/JRtfLloZLFXDiatXzWyzcRhI+b
AcF9BXERFKOGSDZqsvHyX/8lgeV1G9DQ6LLdYDB2279XLLDo+Zggkxt2ixaLQbGRF1xOFNB7smnG
HSlIcioxp0Hbo9uX8Ltxhe+YbXVmNOr2kSVhnqmcWwaTR5dEqPVnsCOAnpLnu2CYBMtDzfoRZNIx
Lrb7KJ0c5152F13bWf8+Zmu3j0tFAEXl3wmMjKonNMuJMp85iC1Cc6wAkv3r8XUC8yfQ7/iXA92G
PZyPTDcNDz5wCqCxpG5LDgVKOchy+l6WafSzABhyotUC50iEOy83K4HRcufxf00dBOHRN/QIdkoa
JyqWaF2IHGYEMD/ZDb4rde+UXqj86oYIOVoAS/foKG9FPdROuWQGlG2m4FL2CSgG2HQFpCEXGJOn
yeQ8qkEP+S2vqir0OOQ8QIqyHPFd7iAsjuPoUMdF/ynLIwrL+d6Rx4T4yxxDmSBZoR6VsuoSvwgG
wWgbuff5rCQskM2RBJJt3IpxWk+gsmdaDjJyuAPtA4Z9WnRxI0fh5xL8HcaQDL8nSIJkT3YRmDsv
IWU/wPprwpUVP9dRnh0EGrSySzuzmjZWJE/ImlQDY8zUg7nl4+3PcMRnKcv8EjNWggRpUqIoMftJ
tHn6eSVkjNoll0mh0rYwJqLL3hfsyIxT3KWK3hsPIx+ydxSpRj4PZ0vwaRCQl/B5tyk6Bp9rAHgy
SRHRRVTCSe63SsithIRpRjBKVFTt7rHuf7O1UEe/mdKVrwuAoPtwnE2LuMNiyOcNtko8rCpxEzLJ
fiHGt3q/kBjyOB72Em8Xm4OZY0ne0KVqiA4Ya2AryP5nbzb/V/DGklT5bIBXyWgCjv7mz/PVx2+f
XZwG9m7IuEsFC7GDC3PuuupdIesM4u3T+DSGqbUmuoUUf+BcSMG8zMXS3OMDjE+4qEsifzCnXk8D
ejU2PVdfVXA5B1xsU6+XHLNO1bRaQBF+m8zeDgauUtKWu2x4wJsIdV0Yne4Y8fx/D//IV59NwnC6
+17cJQjT+JVE9tkaj+jz1RlVtL4q+OXlpHbR/TJLwBgzdibD8KQJs11ep2yKqdfHp26SgPk+AcYY
UNjpPXYqR7EREGDT9qbv4uUYvhuD6SGREArhD2YpQsbfo4OL9VUKCmGPdnzpKxn2w7/U3pJYTjQ/
EZUvNHMcCkPqu42mi3kLHaV1fduZOoVpwxJ/ZxxtdidCIltiruNitBHSDPrym74RWUJbUs6RqD1h
hGo/6Q1JygeRrc+1Y4Azuo5Ml6vqfXqw5L3jxiVQXq4sgKA3Tmj8XTQlA4xDBdglUvUpF5wp+T6b
9W9pSwXfvkjnub7VvQUtcEYDRZhFYCn3r5LlBhFkFcuKEoEcOC/2xa3lWL6o9tDKTOkt/kbNGR0w
zn9Yhd/zs6WFaQKdkMVOlsCEsIHKC7cfxihuGW12aeS0NWga3v3EY5/wwAFwniApTGArvJOpO2AS
JS9b0abkzf424iaADY4UoALPjot8Emi6y/1L46V3FKGi6ownTDaHVObAL/aPzygva1hYhwJxe+Hb
uOorG+BA9+bPvWojkfU9NNNYlqIOib87FLtjZuN//f0ZcxJvNoU5ClE1Q6sqhzqzVBA38gQwIZ+m
lEFGBzwihvJqnCDHerzJRia+AImiGnoYQYLTFwntxQ1IgBgb4c4G4UeCCneKBFzcOgvuhTout3qo
7lhM38H1WJCvPaKkpRjapxk8NG3BlCVoeQhTGTXhnfZsTo8qyOO5Sco2xBnrAHuI4tmkbkKid7DK
HyuOPphaycUA4qSERB3Fcge7O5iffcVdQpJBx6+JqmRVHz+oAI50CFI1Zjum/3PZEBNakRE0pB50
PS79KsJf1mD5WEihXDb+XUuTZbf2dcgzyLZa7ZvC3tGbSo4CSmuNXo6htRrDx74KpvBXazEDQvQI
7CjowIhjBkv9waSA8bNlB38jYCzShLZ7TGL6w8ZYNdootuvSkMtEiX7Q5P6ffi1j9+6zCVZeVD4r
rPtqJoXk0ZAk95jcaQYK0BqZzVRF1oMvIQdGjs9z71CBmQVzGBtv3gPASJ2HMO16OhZNkgXHhweW
EcE4xpaOLxht8RQnXtYkptJEMf765h08f5RNUCEqtKzIqcntAfgbvRjXdTWHCv3TjGV8O/cYC9c/
QtTPuQFOL6Vmim/4kSFmYTQ2UsR7PtJJcYV7xaNJBctlfmEAKucEd3p1MljJDoQUU6moj5tprSlk
jGppIyh2bCmJdAquY7TlSEreUJit1n9dzrbFTUYw6hGudZFNlXem4KbEa67tAt7HkgNfauSk7wJm
Nej1uf/+ynDAaOrCS2sLmWkwPHpNHrog4mdAwmXYIrz3Bu9QQP+zyc8gbLucqIWa3H8eb4JhqzPv
zLFweXZNOR9LWVejKup/Juk6CyQPncyAST4dJe4zWYC4qjuTjiouFtyhb5krUIKPWgEVQ02NaovJ
itM3JTRhYZbtY2qZMh7VQ8H3TMtnAHO+TwukWTm4EViTwkgSwds+c9WFDccn7D5nv979+kV5AMhd
bCl1IzJ4nCaDRPxfaqeJo7T0XRFPhxkxhzkN5w9YGVM6E0uUgq7G4rWEQysevR2Jo3ySu0+JTigt
Wj7+ioBbJ535+gLOqB+vVjJjKZEa5xu5iE2YDtxTsmSUG7Czx+W5qE5yDhDzJKzpM0lwhG60wQGD
t5p7A2162vLi14S21b9ndgQuPk3gVcYMdjb/Cq+03TIRwFUKkkqf2DJi8IpQsKaeiG2i1q0UKDUN
C4Oy2ZkJb7SfXGc+KDNu4FrM92ft5G2gPbVZXur8NYxOMPXBOx/0/RfIg1yq1q+3i+FqwXvPGTfX
0JzSbpo1h0DQPXpOTRXVARYFv9Lmtv9EdmiIukMI+V5yP/+letdUMRMRCENHmKCZTc9dDT3dKXfS
rSdzWUw2JB1oy20MZDOOi/zdFsUiRCfG67ka/ijl6cGv2pR1jSUkSunLGOkdDTlP7nNVzs0R3fqN
Oov4P3Y3uX7G0rQszw81eaNQnyY5+unAenOV/nH8CjPJ4h8sUCFOthv4kOlEc8psrBek9n8qq+Ml
OeXut8CbljQymRYrZq9Ka/FXQrVnL1pWHL4rzoTNrsbpb46glxBbxlbnhRdMRJoqwTH4sWvtSkI2
5NAm1T631U5AzI/uhVIgZEHJkttHHDyM37acF8s30/R/93z7nDhEH/H1yBlmM0hHgCTGCmhOrQJk
JBMf7oI5cl25YQ5nXiLplrUxA3PdafXXFapG/gjF452fJcB51CWm7gbYnAhKL7tcxDJhDx+90Ahx
LwNJLzerNvqZ4ZWhU5BDeJHLgxPCqc/phvVAINc1Lj2UXqh43d539SaXa7Lyw924Mz31S6+eI7s6
eagnnT7ACC/XOW8aMYu0KGCPv6ovc0B/pRvSjBcSFCVLPIYIt1T+lhQT2+xKo4TuHqAyMZ4sYQOC
w1GGeh+b/iittu79DGczgBrWaqgeHhpJOUTHL2d91ZIMFCqIPLCVtBnUO+2i4AmTz4IAWwWZ7Rfc
hD8eJw9TbQqbRxhGczP88m9YGvCPI7Lm3J1iuUbCuTX+Fwt6d1RYCuWI7MIZsPsAiTxR9YRvx2dh
lwswz7qFVummKyQTlnn1ZyuHK94iX6tGzxMq0sD9X/wUVTaENND6D6AOR3i0ItsqADJN+HYLE4F8
+uLo88yY+v7TsMjqFJye8w++7bRPh6MFXE0sVyUDCd9JR2zhp43Y8galcxOawQatMTSmtxnCdRIu
PnaN+c+xQgeKrRqdlMb2rFMMLWb1tjtUYanyAbjCxWM0Kl7l8yZsixZPxGJS8f9YQOieB+Aq2oeY
4iBq3t/ibkhipqSWWq1mKPVHNScoqWsOpS47FUJm71gke89yaqAd5BVuft5F/49+NOTdhHJQE/0/
f/ikSYuK4Y3tbkwSdAYQUeUwXBH9EgB+Bp3gUwp+esLoMWa5Af9Lr+n5A1fZAV+Pzz2wCV8XXSh2
uGw34WcOE6RjKjs+wzKu6wiMsiKJa7WDMsMYvJOHwSI/qdcqKkxxgvfzTdDGMxHbmZuafnrlnpsD
6EWkJz9KP20CRPej84+dLhx+Fn4vm1S3sLR92dN343CUbR+KdK+g+mtKD9Oeb/MwDHuoTK52Y1cU
vvae/17cOY8iE9wE0FYa67CYCTJiSH5SYg2gbPjjfgcj3KAkBnmaN/tk+SL50vzR/o2IliWLJTaf
Ww7IQQqVHWOsKQh33+w09+RJmXaKJET4DpJbEGpHkwRpC/YKpXObsxdmdYiedUcftcSI9LRTl9xR
X6V//RdbPhtFTRkwFaJYsVQEW4IEj8+PbF7IdrQSH1WNpbeYxYizJ3gAqlWeu0nutskV5+vi19rg
nnFsOLkIh5DfK74T/V58TSYcckXsd51rw3X5Axe/pZ485hTm1Qn/hpORdEa1MYhieO8M4Kb5cl48
nYynC9PuqW+sTUCtFAD9sazMEIh3K+ITbNOQ9BYVOaVRr9izP/iyy4Nj11jtxneM1l6jBP2/PM8O
FiuX9HV/07P9YbReYcp2MsjMeGFV/J9L+LZU8EZ8Fw1z698lzP3zgSfMENd1Wuzc5B0wlOhkXFRp
kY9Vf49GcJSqV/PCPo3Tn++/0Vd0tQVwu9KobFHKLdesPu92acygmw3+2QqywA7c8ppT2/1hmebr
x1t6W+jyW61MXrJL7ftT4l1MTpJG6YTtK0Fi5fs42/wowSPFllHcK93X0Re+MzOhB2Wx54a61e/R
VTJWb00QPuxMcofwINoNbrX9MpQy0BEseGgsDQdbPbHlQcA0yy5CRgyrFb/5CTtERqvNT4/E7I2o
xp3fN5APGf+tSUSnVsDQp8OwGqzs3jOT+mL6M90gGbgW6EYb5xZBLYhkI8QaHp3exzgEmNAbdNyy
zxrLfQ0SNHTxzXuHONHJ2rpkoEcqiWrf/18TLlkzogTaCPf148J+EanZ91mKFpJVjuWUju2KBEol
J/L2t75G+N9e+EMbLiqq/ldRv154B/C6T5HHlgPZJ2OhYDnTSXeF52cWxhN45ODssZWjtfNmIz6U
j/CNYupFV8kHxeypMh1XnfnhThGNvRPDG0xEbxfMqE/0/LS7fTn/sZ8r/134C5HzgFI0E/H5FPmG
OqUiPuhn+RavDGzszSF/pSsy5GwucIZOKrkU+/LrGcds5bLMUI6zsRbcAKQKITyShAueYLnkQobX
9H4QqHT1jYOK5VBsnmsjNJxLBPMASiBENJCi/scpY8LcJLqPJ59/UEWHx1LJZIY7y0oCDvVYHoYg
m46kuZzM6LOAsti65kP/2ttos/bIlzcujuqPDMlBvDhYB86fMLd8UYj1DkWU+gJZcj4MGkWj4D4t
SkZwsL/I/7sknX0DANDKXELaeZSmH9MWPe5sHg2YFhiKmBb2CGEB0QsdJX2xl7BZd2bMkKEzJXns
+cldt5uGyuJymaug7XviWaIYeD8lzWspmGcA2kqeEllXj5sSMeSPEFzFT8DZoS6P4sk0hICzp2wJ
vEiX/2lnrU9yjRlNB8h7KBa5X30rEnBlaEveITjSPWtyc4+xezSflY3Qp9nSIKhPo2yw0PMOjdR4
1tS502zc5Hy5XqpLWsmiDz497BJDokHjy5O29OiMheSs9bTRWpWHSMQ6MUO2t6GQuu3zqjqTT3gr
UDE00ygffAH4WEIVgS/CvkqUA9ZleSr0Soyr+PBmeFab4/g9UYNq6DQ4hppAXgguUS58g3Ynpose
5VxnouAowealvEsTEs9jEVik+DHbRCTrcL7Nb7ZZTEW/MBXEULkFpgnc6lvLnC7Wn+b4CBB9wz8Y
6Yca5STM14ZjP7vRBqByu5qfHmfZYhkXto8ro61v9PewF14ZKkBbfs7egMBzmL+ePBVEQDI4r//q
Km0IAp4xCt4lqEar2IonKwLbYCYfLm+wTkRs9CAiC4fqNRiWKoxxKucEfdnKWbAVKDcdClDXAtRx
rM+pBjceTOvqeMdUGqqdGE0Jp2J4FdFy7sXcyUvRiXe8AEkfWxZI5qqOQ2Whr/ZgelpCYeFigXCk
XYOEYhVGqDyRH1aeMMQkKGoaTGSQ2+w0PsJG0bIRHydPj2CCSdMKDKdVyDYvvfVBGGgCbchHcJ/D
jfLR9KJz0mwJHuG9mCmETo5tpPmXCRRsiI78KEl0HL06kNpMv7Wrh1yXAsFXxvIxyH/R2GHL3yUv
TmuFvn7OQFW6fu/V2xZJIuvTfI4oY6e6rRCszxPMffnpgIplPb77q6VmQdlF3uttd0zoeydskiYH
99SaiySE3//sWnqZs/BtgOckpwyiLuxRhi8F2qPgaIuTdpB7RiQ8mQMWxkhRqRWwLHQQOLv/gKiy
kTOFOYJMuDJKzirhywj9uAmywml+IXwv7izwsrwIwBiBaak0JVeJoJDzcOewNe9X2IE6Nstw7YKx
OkVFqHxjLoTA9xb+UULNqA5mf6PPZGq2X2ZIGYGsQ4SHIUIDM4HBmgsXjRnLtDWjwmK1xaoQfauQ
jJxM8U0g9IHbT/rM+SJxdDA/RmpPdTjkRVnvVJpYM8TllvKU4NIxOef721vpsnVfYDeSTtRA2apA
bRltpVE51CrbvTKiHH4U3Nr1pOgg3Z10mNHztFge7Z5OaGmPKZ0PTQr9Zy5XY5ozlGfLq8A4Baqb
tjYcM5JqdFt5A+c1Nf0005W/sD6fTg3uJ+Iu4lEDzrMn9QmSZHs7xA1hczdJL6/6PGkeVRixXQab
rr++RuQII1pt3eJ6JDNgDdbrcxtz6TSuQXap8j/iAUEkQkhWY6Jne6vUO1+3XSI4A7rC373a0AWd
NxOVOTQbj3Z9h90EziRISekrHqsvonQElkw+ghCVhCS3De7+c3Vsi8iIJZ7c/Iyr41RYbLXh6xRr
C/OVLXYzSbiuvgAgSR9wymahz4W57CTVc3iagoGnOb1aevFGpRYhhVmEXsJHeAYzj/JS0VydIBAn
3GyBq8u5yFPOluIKj4qYawLs4y3aH4ZVZWoLf4UYPnWAl0+A8rVgYk4w6mleqEdJVpbh7lLeeu1A
ApN1hiUog143jF6P+ArNpP2iHuwTxTQ4EiphmVkbQa2URlZkk1fwUovilymSJtqfsv7BLDhG0H/8
LmpIBFhu3JpZTJQIlGxIJCw85tl2kuvPZlaHnnf/S6arvUQkhdaJzaEQGYw5K7MCJsCQKvKHmOcF
uDBQD4CTnmqnYK3Qb2jHoJ+Mv8fFJvuLP/4SgFjTbZBvvZeIIUeQ52BRvjjiuluRLPCsCERCoK1k
0Te9LmzLgPL3RbfA4H9Ooj5X0ptAElIwHoj6ZKrTJvPwnX0EkSL26PXO8o5H5/X0de+YujNEbOFP
DgJjLfcQQYCKqOEPl3J4PyVYIMCOWEoD3XU/U26gpdiyNUsQxSlwkKCAa4jkdfL+LEQT0p1eBY+Q
3c5XGci2Wgkk2fm6UtexBfzaRSsBPo93UNBN0fJ9oUcqVCyazI8jo0JR6h6ncR03nbgY2GNden5/
4KZgArQ2/R+YhgjxujdAqIcnIIjPIJCEpoLbleIFzG/b7cio8O9EI6JYN7+bx+qTayZW5hnVGvp7
tYegQ5/vC73pAz6X1KA7xvhepZETqsWK/IYMqbqJOakrMi3sDtjVghNt/iP1FPlZygEq7duj7Giy
UZpp3pZabz50J8+XMGI6SJCAKozm/V3XwAX4VlPgC/NXI859ap0rtxFqTJNA2khi62IcFvLXHGlk
3ofCjGkj5GfUak/XFSQpEJefexp8VzrEblMcH4lhB+TUzNoet+NP+jq1+EDuJcUpPa4XNIon5ZBn
+7lGydVj0VAxJTK4FQYdwXrWliBHLVNs+gRcOB1ioV/sibgZR07ZX2EsTXWkCgUHxkvtgoF4nufo
DJxPgQCE/3tJURJSYRnn6lZrd7ATBo0R661/s/GeB5LAw+6v3K7o8oDrp0hYzuGmLkG84dehDVuU
uHerPIrFDYmp9riUVuGcHFkUbfeVZpCsCEzRVWpN0q57uhTlYdrbETpI0bJEx7wU2YGFmJ5rNef3
hIa9+Pvl7OPImvqXKaiAdkrKqcIeMyKEuZ6PfgSd677hsaOxiDk7K8LExZEsOM6Y1G6oazj7V5sM
WcAuh/LDSOxYdUKu3SREL/WCNRtJAEF0LbPMk61AdUluaBel4wgrg56+/krhiQYQCwem/KF+oJal
PvKLmPpdRDxA9evKNjMHmHhhO7e/JnVy+3HWg4TMHn9wXtxYKXvpQk7aWfNO8xHkjI34xwU1WURv
TbeOey5nW49mFpi+0D6+t6Ir4nAeIJul/kEqfis1Vv1s8mbC2yt5eXxnbGya+1LIk3MRD4IX6gmg
CtSJ6XZNoHPhg5jrWTQV8CZU29arb1S398SsCTE7flvwPLr0s8pAVmM/GlhBJAbLu7YecVCnO7g1
y875dnm8AhF71now4UagUoyRZdmY14oCy6b66kn2sbo2FAD905J4MFyC5AXYXLiKsxV0fM5bVFNu
zhoA9TLeaIfOx3g1bTpYJkWzfUdqdxhOYkFahTlvShAIil9FZcjlb4N2SKiXw3cOtEw5QYkRbIZ0
uomus7MrXjS8xc+39bIQn+8TtQX6rev87tVJ6F3IHBfvfRXU/aItqFV6KoMKm93v2UAipdK/mlJK
TgNXgBEPHU2Dbnlt48nJiieHb+IvqCQMADW3DBh81baL2BmYirYnTmFrkhsCVxKwkL3qP6LZJ7un
fqhTrrs2eF8Bbv2o/5J2WQJKPrdWVts261B3NqtYf6R5oz4LVJ0XKDMRRRrXSK+3nVbo0Iycian0
Bxx02Sk5b/5j5J0RrCNyw/xPVZCK3lBkyS3KcGMq/xenmJ6CMR1MX2jDPn3CiU6tzhukbiuYPpRK
1ohjMsdadqlPVsBuLg9LiPgc4zusPyluKuhfQvZEcWQ4Nw/SlAvDjsyTTE+o3AFv0ZWBcQv+v2+3
v+zciz81U+vjabFIsTxcMP481lV4MJueW54VHxOwUCtRfVcd85xPwBmNxroVK6nUzFttLRP3O6Zh
r/fJxpeEOdmUp/IWfpAujD3V55wODkldlMvk6O92HJAds5rUVj00yMlyEcv972jv+Uln6CeNjWji
Y5orbJyjoxwxJ/XMKv9g4n7VgI3+U5csrW3Dzrzndo2MEciVNN2wuf11BVKiDtIdYX0rAf6bkrLT
ZtHLkEiA2IhYaaJdUBcDCE9fRUyBDy1eDl2IlfTZvaLJsHe/67z8Ir1wLP08s6wfEmYBSouQ7Clf
6nOgSoIDD/0GUY4bvQFMN9GIY5j2YRtXmf2M7WMCwIavdvM3IJWfDmBXMHyrhu4pWY1SL1Vn2M67
SmUMS6hrU3cXPZ5PkNOCzXe7KmvUdGC09c1GauDlYeap0Z/0XuG/cNXyySApCQsgSU0i2/eGL1Mq
f57vtOUtBX/2pHPy64qgeF/DoVjGmE4+nQGiFuv9N49JFQDvVi/2blLYHiRe+11+bGVf89TZa73Y
doKTTsDTV0JjEwWkmusCLVDX498bhHRkPuBYu9GnD4JcrzchZmLQ3VCIQkzpMeEZbDBZw5Va9Hbc
6oX5s+RwXKUBK0kvD6uoVPxe2gYn/5NjH19WPSxAZsD1Ej/AFk6keZuAF7wRlbd6KN+ywgFTpvzw
hn6R9SoAlKOTEjQR7EOzTACh6XDLhPY6X6a1gkLTtcU9NHtxbn0nRj/cH66P2ZpshAulr7D19lcB
mUXU+Kr7bqwOCHap94keRSpsIVCByFxmBPvgJNv80trW9ChsQykvSX/Uuu/VfIdj6vc3UX/+4fu6
S7rXY4Qth+76uon3+s/5CtKjNLAm9JUykooHOOt+Xs58dwuQ78wjZ7wWguvN+nGN/5MisROmmzp8
3G6dzoABxWXFzE/zH30a+JdgAfJh7wH6I3Y4jeh247wq3PqLiE7vYnHNpSHSJM19jQOl60EVZBla
wEAK/debOfKvDJANMIJuIa2xZmS0Cb40tX/Jk/9eQ8QK+5r3SMU7KxXFEbV/xseRBpjpGs2UJEyt
551iEkb0xBikgJ4oWHfnKQoMYA8sWPfVcGhgFC9hBhLX9EhkuuCtjHPeS0/kMRPNo5hGe1OnTi9D
y6ra1sZY+6Iyl6yWHUGCXsOcGGV2fXqGFuh7V/ArFzXMjI3H+tuccLGyFs59jxCo9MmK9YNqIASq
5/PqJeYk1Y7IGpWU7x8l2MV5NcvHZeNaU/kyZBrJIAe++6XsfC3+oAryk1Jp5r0bsgl38ihjT+yx
+ds1ErA1GKp6sBI7+a10I301d94M/3pY9MtnvHAGmaF1q2E8CTA8itRQFwpHU9xfLukt3TLxRPTh
C9hRVbdvcoOH5/x1sfQHSsQUueNSCOesanaUTt6JWBlXkUPzGklBEtlKyVBrXfqf+Zen8adC0vhr
SwXjq/hXCatWqGLRPe8gz9riaiYwyU11AVgFL7DI
%%% protect end_protected
